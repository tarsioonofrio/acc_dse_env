-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use IEEE.std_logic_arith.all;

-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity bram_single is
    generic (
        INPUT_SIZE : integer := 8;
        ADDRESS_SIZE    : integer := 12;
        DEVICE     : string := "7SERIES";
        BRAM_NAME  : string := "default"
        );

    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic;
        DI   : in std_logic_vector(INPUT_SIZE-1 downto 0);
        ADDR : in std_logic_vector(ADDRESS_SIZE-1 downto 0);
        DO   : out std_logic_vector(INPUT_SIZE-1 downto 0)
    );
 end bram_single;

  architecture a1 of bram_single is
    signal bram_wr_en    : std_logic_vector(4-1 downto 0);
    signal bram_addr     : std_logic_vector(9-1 downto 0);

    begin
    bram_wr_en <= (others => '1') when WE = '1' else (others => '0');
    bram_addr <= ADDR(9-1 downto 0);
          

    MEM_IFMAP_LAYER0_ENTITY0 : if BRAM_NAME = "ifmap_layer0_entity0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009e0000009f000000a5000000a6000000a00000009c000000a20000009f",
            INIT_01 => X"0000009e0000009f000000a1000000a0000000a1000000a6000000a9000000aa",
            INIT_02 => X"000000a7000000a2000000a0000000a00000009c000000950000009600000094",
            INIT_03 => X"000000950000008f0000008c0000008d0000008f000000890000007e00000074",
            INIT_04 => X"00000098000000970000009f000000a6000000a2000000a0000000a4000000a2",
            INIT_05 => X"000000a30000009c0000009b0000009f000000a3000000aa000000ab000000ab",
            INIT_06 => X"000000a9000000a00000009a00000097000000910000008b0000008c0000008d",
            INIT_07 => X"0000009500000093000000910000008e0000008f000000880000007d00000077",
            INIT_08 => X"00000097000000970000009e000000a7000000a0000000a3000000a5000000a5",
            INIT_09 => X"000000a3000000a20000009e0000009d000000a1000000a6000000a7000000a9",
            INIT_0A => X"000000aa0000009f00000091000000790000006e000000620000006500000072",
            INIT_0B => X"00000078000000860000008f0000008c0000008e0000008b0000008200000078",
            INIT_0C => X"0000009b0000009b000000a0000000ae000000a7000000a7000000a9000000a9",
            INIT_0D => X"000000a5000000a5000000a7000000bf000000b10000009d000000a2000000a4",
            INIT_0E => X"0000009e000000950000006800000067000000620000005c000000500000004a",
            INIT_0F => X"000000560000005300000071000000840000008c0000008c000000880000007f",
            INIT_10 => X"0000009b0000009c000000a1000000aa000000a9000000a3000000a9000000a6",
            INIT_11 => X"000000a4000000a4000000ad000000f6000000c300000097000000920000008e",
            INIT_12 => X"0000006f0000004e0000005500000071000000700000006a000000610000005d",
            INIT_13 => X"0000004a000000540000005500000069000000800000008a0000008500000081",
            INIT_14 => X"00000094000000850000008200000093000000a1000000a5000000a7000000a7",
            INIT_15 => X"000000a3000000a5000000a3000000b40000009d000000800000006100000042",
            INIT_16 => X"000000450000004200000059000000760000007a00000077000000720000005e",
            INIT_17 => X"000000630000005b0000003a000000430000006c0000008c0000008a00000086",
            INIT_18 => X"0000007f0000006d0000002f0000005800000099000000aa000000a8000000aa",
            INIT_19 => X"000000a9000000a6000000a400000093000000810000007f0000006400000044",
            INIT_1A => X"0000004e000000480000005300000084000000920000007c000000690000006b",
            INIT_1B => X"00000073000000550000003f0000002e0000004f000000840000008d00000086",
            INIT_1C => X"00000083000000630000002a000000460000008f000000a7000000a5000000a8",
            INIT_1D => X"000000ab000000a10000008c0000007800000082000000900000007400000058",
            INIT_1E => X"0000005b000000550000004d0000007c000000a300000088000000660000006a",
            INIT_1F => X"00000064000000550000003600000031000000390000006b0000008a00000088",
            INIT_20 => X"000000aa00000067000000360000007c00000099000000a1000000a3000000a6",
            INIT_21 => X"000000a5000000ae000000710000007d0000009d0000009c0000007900000056",
            INIT_22 => X"000000520000005400000050000000510000008a000000920000007100000057",
            INIT_23 => X"00000053000000560000004700000038000000280000004a0000008500000089",
            INIT_24 => X"000000b4000000860000005e0000009a000000ae0000009e0000009c00000099",
            INIT_25 => X"000000cf000000ed000000cf0000009c000000ae000000940000007d0000005d",
            INIT_26 => X"000000560000004a0000003b0000004c000000890000008f000000850000006a",
            INIT_27 => X"0000005600000057000000540000004b00000032000000280000005f00000084",
            INIT_28 => X"000000b70000006c0000008e000000a5000000b10000009b0000009f0000007a",
            INIT_29 => X"000000d5000000ed000000dc000000a4000000b70000009c0000007d00000078",
            INIT_2A => X"0000004e000000500000002d0000005b000000af0000009d0000009b0000006b",
            INIT_2B => X"0000005700000067000000580000004e0000003b000000290000003b00000068",
            INIT_2C => X"000000bc0000006400000087000000aa000000bb000000a6000000ad00000086",
            INIT_2D => X"00000075000000c2000000c7000000aa000000b9000000bd0000008600000075",
            INIT_2E => X"0000006600000054000000260000007d000000d2000000a0000000920000005d",
            INIT_2F => X"000000530000005e000000680000005500000049000000370000003e0000004c",
            INIT_30 => X"000000bd0000005a0000007f000000af000000ae000000a6000000b20000009f",
            INIT_31 => X"00000061000000a8000000a800000089000000ba000000d8000000a00000007b",
            INIT_32 => X"00000078000000730000003200000096000000c20000009b0000007b0000005b",
            INIT_33 => X"00000054000000540000005f0000005600000054000000490000004f00000049",
            INIT_34 => X"000000bd0000005d00000098000000b90000007700000088000000ad000000a7",
            INIT_35 => X"000000670000009300000091000000a7000000bd000000e2000000b40000008d",
            INIT_36 => X"0000007e00000075000000470000009a000000ba000000950000007200000057",
            INIT_37 => X"00000050000000480000005000000063000000640000005a000000610000005e",
            INIT_38 => X"000000c20000006c000000a8000000ba00000069000000630000009c000000a7",
            INIT_39 => X"00000064000000730000008a000000c6000000be000000ac000000910000009a",
            INIT_3A => X"00000092000000670000004700000098000000b300000089000000820000006e",
            INIT_3B => X"000000550000005b0000005f0000006d00000073000000640000006100000075",
            INIT_3C => X"000000c500000084000000ac000000b8000000820000004e0000008c0000009b",
            INIT_3D => X"00000073000000820000008f000000e6000000f2000000910000008700000083",
            INIT_3E => X"000000790000006c0000005f00000090000000a8000000980000007000000057",
            INIT_3F => X"0000004700000057000000690000007000000078000000670000007900000088",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY0;


    MEM_IFMAP_LAYER0_ENTITY1 : if BRAM_NAME = "ifmap_layer0_entity1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000cb00000092000000a8000000bf000000a80000004e0000007e0000008a",
            INIT_01 => X"0000008a000000600000009a000000ad000000a20000008c0000007100000071",
            INIT_02 => X"000000650000006900000070000000ab0000009c00000094000000870000006d",
            INIT_03 => X"0000004e0000004f0000005e000000650000006b0000007d0000009700000090",
            INIT_04 => X"000000d6000000a3000000a4000000b7000000b00000005e000000600000009c",
            INIT_05 => X"000000940000006a000000810000007600000072000000740000006600000073",
            INIT_06 => X"000000560000006500000090000000760000004400000080000000850000004b",
            INIT_07 => X"0000003c0000003a0000004700000066000000740000008f000000960000008c",
            INIT_08 => X"000000d4000000b2000000a7000000ad000000b00000007c000000560000008d",
            INIT_09 => X"0000009900000087000000680000004d000000860000007c0000008100000093",
            INIT_0A => X"000000550000005c0000009600000084000000750000006b0000004b00000040",
            INIT_0B => X"0000002c0000004100000056000000850000009b000000a00000009a00000097",
            INIT_0C => X"000000c7000000bb000000ab000000ae000000b1000000900000005600000077",
            INIT_0D => X"0000007a000000890000009000000046000000810000006c00000091000000b8",
            INIT_0E => X"0000007400000049000000830000008900000086000000590000003300000034",
            INIT_0F => X"0000002f0000005a00000079000000a3000000ab000000a40000009e00000095",
            INIT_10 => X"000000a5000000c3000000b3000000b1000000b5000000980000006300000083",
            INIT_11 => X"000000ab000000670000005d000000500000005d0000007a000000b2000000bf",
            INIT_12 => X"000000960000006400000059000000570000003c0000002e0000002600000018",
            INIT_13 => X"0000002e0000003c0000006c0000009000000090000000800000007f00000078",
            INIT_14 => X"00000075000000c3000000b1000000b2000000b50000008a0000005300000096",
            INIT_15 => X"000000f5000000db000000850000008600000095000000b0000000be000000c2",
            INIT_16 => X"000000a80000007d0000006e0000003d0000002300000022000000310000003a",
            INIT_17 => X"0000003d0000003a00000045000000480000004e000000450000003b00000037",
            INIT_18 => X"0000004f000000af000000ae000000b0000000b10000008c0000006d000000d3",
            INIT_19 => X"000000fd000000fc000000d00000007c000000720000007c000000740000007a",
            INIT_1A => X"0000006800000044000000440000003c00000034000000320000003300000038",
            INIT_1B => X"00000038000000330000002b000000330000003b000000300000002b0000002a",
            INIT_1C => X"000000290000006000000090000000a8000000b2000000a5000000a5000000f6",
            INIT_1D => X"000000fd000000e30000006e0000003c00000035000000310000003100000030",
            INIT_1E => X"0000002d0000002a0000002e0000002a000000260000002e0000002e0000002b",
            INIT_1F => X"0000002a0000002e0000002e000000320000003700000035000000330000002d",
            INIT_20 => X"0000001d0000001d0000003b00000083000000a600000084000000c2000000fe",
            INIT_21 => X"000000f10000008d0000003d0000003200000032000000330000003100000032",
            INIT_22 => X"0000002f0000002a00000027000000220000002300000027000000260000002a",
            INIT_23 => X"0000002d000000380000003e0000003b00000038000000320000002e00000033",
            INIT_24 => X"000000300000001e00000022000000490000008000000080000000d700000100",
            INIT_25 => X"000000bb00000042000000360000003200000034000000340000002e0000002d",
            INIT_26 => X"0000002b00000029000000240000002700000028000000280000002b0000002e",
            INIT_27 => X"0000003b0000003e000000400000003b00000036000000320000004600000053",
            INIT_28 => X"00000034000000230000001f000000290000004200000080000000e0000000f0",
            INIT_29 => X"0000007c0000003a0000003100000038000000360000002c0000002c0000002f",
            INIT_2A => X"0000002e0000002b0000002b0000002c0000002c0000002d000000360000003a",
            INIT_2B => X"000000360000002e0000002b000000240000003300000049000000550000004c",
            INIT_2C => X"00000032000000230000001d000000230000002c0000004e000000ca000000d3",
            INIT_2D => X"000000610000004100000036000000300000003a00000030000000280000002d",
            INIT_2E => X"0000002f000000300000002f0000002e00000033000000270000002700000030",
            INIT_2F => X"0000002f000000270000001c0000002800000043000000430000002e00000033",
            INIT_30 => X"00000032000000230000002000000021000000290000002e00000068000000aa",
            INIT_31 => X"000000400000003600000034000000350000003d0000003a000000360000002d",
            INIT_32 => X"0000002a000000290000002e000000310000002e0000002a0000002800000027",
            INIT_33 => X"00000025000000280000002c0000003f0000002f0000001f0000000f00000033",
            INIT_34 => X"000000440000002a0000001f00000026000000250000002b0000002a00000047",
            INIT_35 => X"000000310000001f0000001b0000002600000031000000380000003a00000035",
            INIT_36 => X"000000380000003c0000003900000035000000320000002d0000002700000021",
            INIT_37 => X"0000002a0000003e0000004f0000004900000038000000260000000d00000028",
            INIT_38 => X"0000003d00000031000000230000002b000000270000002a0000002c00000028",
            INIT_39 => X"0000002a0000001b000000170000001e0000001b0000001d000000240000002f",
            INIT_3A => X"000000380000003e000000420000004b00000045000000310000002b0000002b",
            INIT_3B => X"0000003c000000550000006d0000005d0000003c0000001a0000001d00000014",
            INIT_3C => X"00000036000000380000002d0000002b00000028000000280000002800000026",
            INIT_3D => X"000000240000001a000000160000001d000000190000001d0000001300000012",
            INIT_3E => X"000000200000002f0000003d0000004a0000004200000035000000340000002d",
            INIT_3F => X"0000004300000059000000690000005900000030000000180000002200000015",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY1;


    MEM_IFMAP_LAYER0_ENTITY2 : if BRAM_NAME = "ifmap_layer0_entity2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000700000006f0000007400000076000000700000006d0000007300000071",
            INIT_01 => X"0000006f00000071000000740000006f0000006f000000750000007500000077",
            INIT_02 => X"00000075000000710000006f000000700000006d0000006b0000006b0000006a",
            INIT_03 => X"0000006b000000650000006200000061000000610000005f0000005b00000055",
            INIT_04 => X"000000700000006e000000720000007400000070000000710000007500000072",
            INIT_05 => X"000000740000006e0000006f0000006e00000071000000770000007500000073",
            INIT_06 => X"000000730000006f00000070000000730000006e000000680000006600000064",
            INIT_07 => X"00000069000000660000006600000061000000620000005f0000005b00000058",
            INIT_08 => X"0000006e0000006d0000006f0000006f0000006a000000730000007500000075",
            INIT_09 => X"0000007300000073000000720000006d0000006f000000730000007200000071",
            INIT_0A => X"00000074000000720000006f000000600000005a0000004e0000004d00000055",
            INIT_0B => X"0000005600000060000000670000006300000063000000620000005f00000059",
            INIT_0C => X"0000006b0000006e0000006d000000700000006e000000750000007800000077",
            INIT_0D => X"00000073000000750000007b00000092000000820000006f0000007300000072",
            INIT_0E => X"000000700000006f00000050000000570000005a0000005a0000004b0000003f",
            INIT_0F => X"000000460000003e00000055000000620000006600000065000000630000005e",
            INIT_10 => X"0000006b00000072000000730000007200000072000000710000007800000074",
            INIT_11 => X"000000710000007400000080000000d60000009c000000720000006f0000006c",
            INIT_12 => X"000000500000003500000045000000670000006e00000072000000660000005e",
            INIT_13 => X"000000480000004e000000490000005300000060000000650000005e0000005d",
            INIT_14 => X"0000006d00000068000000640000007000000073000000710000007400000073",
            INIT_15 => X"0000006f00000074000000760000008a0000007a000000660000004b00000032",
            INIT_16 => X"0000003a000000380000005300000071000000790000007a0000007400000060",
            INIT_17 => X"000000640000005b0000003a0000003a0000005400000069000000620000005f",
            INIT_18 => X"000000640000005f000000250000004a00000075000000760000007300000076",
            INIT_19 => X"0000007500000074000000780000006b000000620000006c0000005700000043",
            INIT_1A => X"000000530000004b00000054000000820000008e000000760000006300000066",
            INIT_1B => X"0000006f00000053000000470000002f0000003d00000062000000630000005d",
            INIT_1C => X"00000073000000600000002b000000400000006f000000750000007200000074",
            INIT_1D => X"00000077000000710000006d0000005e0000006e000000830000006a00000057",
            INIT_1E => X"0000005f000000580000004d00000076000000990000007c0000005d00000062",
            INIT_1F => X"0000005d000000510000003c000000350000002f000000530000006700000061",
            INIT_20 => X"000000a1000000690000003a000000790000007c00000071000000750000007a",
            INIT_21 => X"000000790000008700000059000000690000008d0000008f0000006f00000050",
            INIT_22 => X"00000051000000550000004e000000470000007d00000087000000670000004f",
            INIT_23 => X"0000004d000000520000004900000039000000230000003b0000006a00000067",
            INIT_24 => X"000000b00000008b000000640000009a00000095000000740000007400000076",
            INIT_25 => X"000000b4000000d6000000b40000008300000099000000830000006e00000055",
            INIT_26 => X"000000540000004a00000039000000440000007d000000850000007c00000062",
            INIT_27 => X"0000005100000055000000550000004c000000310000001e0000004b00000067",
            INIT_28 => X"000000b70000007400000097000000a90000009c000000700000007600000059",
            INIT_29 => X"000000c5000000e0000000bf000000870000009f000000890000006c0000006f",
            INIT_2A => X"0000004c000000500000002c00000055000000a5000000930000009300000064",
            INIT_2B => X"0000005300000066000000580000004f0000003b000000240000002e00000051",
            INIT_2C => X"000000bf0000006c00000090000000af000000a7000000780000007b0000005d",
            INIT_2D => X"0000005f000000b6000000ab0000008e000000a1000000ab000000770000006b",
            INIT_2E => X"00000062000000540000002600000079000000c9000000980000008b00000059",
            INIT_2F => X"000000500000005d00000068000000570000004b000000350000003700000038",
            INIT_30 => X"000000c20000006000000086000000b40000009c0000007b0000007b0000006d",
            INIT_31 => X"000000440000009a0000009000000072000000a6000000ca0000009500000071",
            INIT_32 => X"00000072000000720000003200000093000000bb000000950000007600000058",
            INIT_33 => X"00000053000000540000005f0000005700000057000000490000004a00000037",
            INIT_34 => X"000000c00000005f0000009a000000bc0000006e0000006a0000007c00000074",
            INIT_35 => X"00000048000000840000007d00000095000000ae000000d8000000ac00000083",
            INIT_36 => X"00000075000000720000004700000098000000b5000000900000006e00000055",
            INIT_37 => X"0000005000000049000000500000006400000065000000580000005900000049",
            INIT_38 => X"000000c40000006b000000a7000000ba0000006d00000059000000770000007a",
            INIT_39 => X"0000004a0000006a0000007b000000b9000000b4000000a50000008c0000008f",
            INIT_3A => X"00000088000000640000004700000098000000af00000085000000800000006d",
            INIT_3B => X"000000560000005d000000600000006e0000007400000060000000550000005f",
            INIT_3C => X"000000c500000081000000a7000000b20000008900000053000000780000007d",
            INIT_3D => X"0000005e0000007800000083000000dd000000ec0000008a0000008200000079",
            INIT_3E => X"000000700000006800000058000000860000009f000000930000006c00000055",
            INIT_3F => X"0000004800000058000000680000006d0000006e000000560000006000000068",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY2;


    MEM_IFMAP_LAYER0_ENTITY3 : if BRAM_NAME = "ifmap_layer0_entity3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000cb00000092000000a4000000b6000000aa000000560000007d0000007e",
            INIT_01 => X"00000079000000500000008f000000a300000098000000840000006a0000006a",
            INIT_02 => X"00000065000000650000005a0000008f0000008a0000008d0000008200000069",
            INIT_03 => X"0000004c0000004f0000005d0000005b00000053000000580000006c00000068",
            INIT_04 => X"000000d7000000a6000000a7000000b8000000b6000000660000006000000095",
            INIT_05 => X"000000890000005d000000740000006900000066000000690000005b0000006e",
            INIT_06 => X"0000005b00000067000000800000006000000038000000780000007e00000045",
            INIT_07 => X"0000003800000038000000460000005d0000005e00000070000000740000006e",
            INIT_08 => X"000000d3000000b8000000af000000b5000000b800000083000000580000008b",
            INIT_09 => X"00000094000000800000005a00000040000000790000006f000000750000008f",
            INIT_0A => X"0000005c000000600000008b000000750000006d00000063000000440000003b",
            INIT_0B => X"000000290000003e00000045000000690000007700000078000000730000006f",
            INIT_0C => X"000000c0000000bd000000b0000000b3000000b6000000950000005a00000079",
            INIT_0D => X"0000007c00000088000000860000003b000000760000006100000086000000b0",
            INIT_0E => X"000000760000004b000000770000007c00000081000000560000003100000033",
            INIT_0F => X"000000310000005a0000005b0000007600000079000000710000006f0000006b",
            INIT_10 => X"0000009c000000c1000000b2000000ad000000b50000009d0000006700000087",
            INIT_11 => X"000000af000000690000005a0000004d0000005a00000076000000ad000000b6",
            INIT_12 => X"00000094000000640000004e0000004d0000003d000000340000002e00000021",
            INIT_13 => X"0000003900000047000000640000007d0000007b0000006d0000007100000069",
            INIT_14 => X"00000078000000c8000000b2000000a9000000b3000000900000005700000099",
            INIT_15 => X"000000f7000000de0000008c0000008d0000009c000000b6000000c4000000c0",
            INIT_16 => X"000000ac000000850000006d0000003e00000031000000360000004600000051",
            INIT_17 => X"0000005500000054000000630000006500000068000000600000005c0000005a",
            INIT_18 => X"00000069000000c5000000b7000000ac000000b10000009200000070000000d3",
            INIT_19 => X"000000fc000000fd000000e00000008f000000840000008d0000008500000085",
            INIT_1A => X"0000007c0000005d00000057000000520000005400000054000000550000005d",
            INIT_1B => X"0000005e0000005b00000060000000680000006c00000061000000610000005f",
            INIT_1C => X"0000005900000089000000a8000000ae000000b6000000aa000000a6000000f5",
            INIT_1D => X"000000fb000000e70000008800000058000000500000004c0000004b00000048",
            INIT_1E => X"0000004f000000510000005100000052000000560000005a0000005900000057",
            INIT_1F => X"000000590000005d0000005e00000060000000600000005e0000005f0000005a",
            INIT_20 => X"0000005b000000570000006600000099000000b300000088000000bd000000fa",
            INIT_21 => X"000000f50000009f0000005e0000005400000054000000550000005300000054",
            INIT_22 => X"0000005600000054000000520000004f00000053000000560000005500000059",
            INIT_23 => X"0000005c00000067000000670000006500000066000000630000005e00000067",
            INIT_24 => X"0000006f0000005e000000550000006a0000009400000088000000d5000000fd",
            INIT_25 => X"000000c60000005d0000005b000000580000005a0000005a0000005300000052",
            INIT_26 => X"0000005200000051000000500000005300000056000000590000005c0000005f",
            INIT_27 => X"0000006c0000006e0000006d0000006c0000006c000000690000007b00000089",
            INIT_28 => X"000000720000006300000056000000530000005f00000091000000e5000000f5",
            INIT_29 => X"0000008f0000005c000000570000005e0000005c000000520000005200000053",
            INIT_2A => X"000000540000005300000056000000580000005a000000610000006a0000006e",
            INIT_2B => X"00000069000000610000005f0000005b0000006c000000820000008a0000007d",
            INIT_2C => X"0000006e000000620000005900000056000000530000006a000000db000000e4",
            INIT_2D => X"0000007e000000680000005e0000005700000061000000570000005000000052",
            INIT_2E => X"00000054000000570000005900000059000000610000005c0000005d00000066",
            INIT_2F => X"000000650000005d0000005500000065000000810000007e0000006200000060",
            INIT_30 => X"0000006c000000610000005c00000058000000580000005400000085000000c5",
            INIT_31 => X"00000064000000610000005e0000005f00000067000000640000006000000053",
            INIT_32 => X"0000004f00000050000000580000005c0000005c0000005f0000005d0000005c",
            INIT_33 => X"0000005a0000005d000000660000007d0000006e0000005a0000003c0000005d",
            INIT_34 => X"0000007c00000064000000580000005b00000057000000590000004f0000006b",
            INIT_35 => X"000000590000004d00000047000000520000005d00000064000000660000005c",
            INIT_36 => X"0000005e0000006300000063000000610000005f0000005e0000005800000053",
            INIT_37 => X"0000005b00000070000000840000008300000074000000610000004000000055",
            INIT_38 => X"0000007400000066000000550000005b0000005a0000005c0000005800000051",
            INIT_39 => X"0000005500000048000000430000004a00000047000000490000005000000056",
            INIT_3A => X"0000005f000000650000006d00000077000000710000005f0000005800000058",
            INIT_3B => X"00000069000000820000009c0000009100000073000000520000005200000040",
            INIT_3C => X"0000006b000000690000005900000056000000590000005c0000005700000051",
            INIT_3D => X"0000004f00000045000000420000004900000045000000490000003f0000003a",
            INIT_3E => X"000000460000005700000068000000770000006f000000600000005f00000057",
            INIT_3F => X"0000006d000000830000009200000087000000630000004d0000005400000043",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY3;


    MEM_IFMAP_LAYER0_ENTITY4 : if BRAM_NAME = "ifmap_layer0_entity4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000310000002f00000033000000350000002e000000290000002f0000002d",
            INIT_01 => X"0000002c00000029000000290000003400000031000000290000002d0000002c",
            INIT_02 => X"0000002800000026000000270000002b0000002c0000002d0000002d0000002b",
            INIT_03 => X"0000002c000000270000002b0000002900000026000000240000002400000021",
            INIT_04 => X"00000033000000280000002d00000038000000310000002b0000002f0000002d",
            INIT_05 => X"0000002e00000026000000290000003600000034000000290000002800000021",
            INIT_06 => X"0000001e00000021000000290000003200000035000000370000003400000030",
            INIT_07 => X"000000320000002e0000002d00000026000000220000001f0000002000000022",
            INIT_08 => X"0000002f0000002100000024000000300000002a0000002c0000002d0000002d",
            INIT_09 => X"0000002b0000002b000000300000003900000033000000260000002500000023",
            INIT_0A => X"000000270000002f000000360000003100000034000000320000002f00000032",
            INIT_0B => X"0000003000000037000000330000002700000023000000220000002200000021",
            INIT_0C => X"00000028000000200000001f0000002c0000002b0000002e0000003000000030",
            INIT_0D => X"0000002c0000002d000000390000005f0000004b000000290000002f00000036",
            INIT_0E => X"0000003a000000430000002f000000410000004c000000540000004200000032",
            INIT_0F => X"00000034000000270000002d0000002e0000002b000000270000002700000024",
            INIT_10 => X"0000002900000030000000310000002f0000002b000000280000002f0000002c",
            INIT_11 => X"000000290000002a0000003b000000a40000006b000000380000003c00000047",
            INIT_12 => X"000000320000001f00000038000000620000006f00000076000000690000005d",
            INIT_13 => X"00000043000000460000002f0000002d000000300000002e0000002400000024",
            INIT_14 => X"000000360000004000000039000000350000002c000000270000002900000029",
            INIT_15 => X"00000025000000270000002a000000550000004e0000003a0000002b0000001f",
            INIT_16 => X"0000002b0000002d0000004c0000006e000000780000007a0000007400000060",
            INIT_17 => X"00000061000000560000002f00000025000000310000003a0000002c00000028",
            INIT_18 => X"0000003900000050000000110000001c000000300000002b000000280000002b",
            INIT_19 => X"0000002a0000002500000027000000340000003b0000004b0000004600000039",
            INIT_1A => X"00000048000000400000004a00000079000000840000006c0000005a0000005e",
            INIT_1B => X"000000670000004d0000004500000027000000240000003a0000003000000027",
            INIT_1C => X"0000005a0000005c0000002600000029000000380000002a0000002400000027",
            INIT_1D => X"000000310000003300000033000000310000004d0000006b0000005d0000004f",
            INIT_1E => X"0000005800000052000000450000006b0000008c000000700000005100000058",
            INIT_1F => X"000000540000004a0000003a0000003100000020000000320000003300000027",
            INIT_20 => X"00000090000000690000003b00000071000000520000002b0000002900000032",
            INIT_21 => X"000000420000005f0000003b0000004e0000007900000080000000650000004a",
            INIT_22 => X"0000004d00000052000000490000003d000000700000007b0000005d00000046",
            INIT_23 => X"000000450000004c00000043000000350000001b000000230000003b0000002d",
            INIT_24 => X"000000a30000008f000000690000009500000070000000330000002f0000003c",
            INIT_25 => X"00000092000000c6000000a600000077000000910000007d0000006b0000004f",
            INIT_26 => X"0000004f00000047000000350000003a000000700000007a0000007200000059",
            INIT_27 => X"0000004a0000004e0000004e000000470000002b0000000f0000002c00000039",
            INIT_28 => X"000000af0000007a0000009e000000a80000007a00000032000000330000002f",
            INIT_29 => X"000000b3000000e2000000bc000000830000009b000000840000006800000068",
            INIT_2A => X"000000450000004d000000280000004d0000009a000000890000008a0000005c",
            INIT_2B => X"0000004d000000600000004f000000490000003b000000210000001f0000002e",
            INIT_2C => X"000000bd0000007400000099000000b2000000880000003b000000370000002c",
            INIT_2D => X"00000050000000bc000000a400000085000000970000009f0000006a0000005f",
            INIT_2E => X"000000590000004f0000002200000071000000c00000008e0000008200000052",
            INIT_2F => X"0000004b000000580000005e000000510000004e00000037000000300000001a",
            INIT_30 => X"000000c20000006900000090000000b90000008500000044000000350000002f",
            INIT_31 => X"0000002c000000980000007e0000005e00000094000000b70000008100000062",
            INIT_32 => X"000000690000006d0000002f0000008c000000b20000008c0000006f00000053",
            INIT_33 => X"0000004f00000050000000550000005100000059000000490000004000000018",
            INIT_34 => X"000000c100000067000000a3000000c000000062000000420000003a00000032",
            INIT_35 => X"0000002700000078000000670000007f0000009b000000c80000009d00000075",
            INIT_36 => X"0000006b0000006d0000004400000093000000ae000000880000006800000050",
            INIT_37 => X"0000004c00000046000000480000005e00000063000000510000004500000022",
            INIT_38 => X"000000c400000070000000ac000000bc0000006d000000430000003e00000037",
            INIT_39 => X"000000220000005800000067000000a9000000a90000009f0000008c00000086",
            INIT_3A => X"0000007d0000005f0000004600000095000000aa0000007f0000007a00000069",
            INIT_3B => X"000000530000005b0000005a000000680000006f00000050000000350000002f",
            INIT_3C => X"000000c500000088000000ae000000b50000008e0000004d000000580000004d",
            INIT_3D => X"000000340000005d00000074000000d3000000e6000000890000008200000070",
            INIT_3E => X"000000650000005f0000004b00000076000000920000008a0000006500000050",
            INIT_3F => X"000000440000005700000063000000630000005d000000360000003000000030",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY4;


    MEM_IFMAP_LAYER0_ENTITY5 : if BRAM_NAME = "ifmap_layer0_entity5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000cc000000a0000000b2000000bc000000ac0000005a0000007e00000071",
            INIT_01 => X"0000005200000025000000850000009b0000008d00000075000000580000005a",
            INIT_02 => X"0000005c000000570000003a000000680000006d0000007e0000007600000061",
            INIT_03 => X"000000480000004d0000005e00000052000000370000002d000000370000002e",
            INIT_04 => X"000000d7000000b4000000b8000000c2000000ba000000690000006600000091",
            INIT_05 => X"0000006f0000003d000000690000005f00000059000000590000004900000062",
            INIT_06 => X"000000580000005f00000066000000400000002000000069000000730000003d",
            INIT_07 => X"0000003300000035000000410000004e00000040000000440000004000000036",
            INIT_08 => X"000000cd000000c0000000bd000000c1000000bc00000085000000600000008f",
            INIT_09 => X"0000008d0000006f00000050000000370000006c000000600000006400000085",
            INIT_0A => X"0000005d0000005d000000780000005d0000005c000000560000003a00000034",
            INIT_0B => X"000000270000003c000000280000003b0000003e000000360000002d0000002e",
            INIT_0C => X"000000b4000000bb000000b5000000b9000000b8000000980000006300000084",
            INIT_0D => X"00000082000000870000007e000000330000006c000000560000007b000000a8",
            INIT_0E => X"00000076000000490000006700000069000000760000004e0000002c00000032",
            INIT_0F => X"000000340000005d0000003c000000440000004000000034000000320000002e",
            INIT_10 => X"00000092000000bb000000af000000ac000000b4000000a00000006f00000092",
            INIT_11 => X"000000b90000006f00000057000000490000005600000074000000ad000000b1",
            INIT_12 => X"0000009400000065000000420000003f00000039000000360000003300000029",
            INIT_13 => X"00000045000000530000004b000000520000004c0000003d000000450000003f",
            INIT_14 => X"0000007c000000c8000000b0000000a8000000b3000000930000005b0000009f",
            INIT_15 => X"000000fa000000e10000009000000093000000a4000000c0000000d0000000c5",
            INIT_16 => X"000000b50000008f0000006d0000003e0000003a000000440000005700000066",
            INIT_17 => X"0000006e0000006f0000007a0000007700000078000000700000007000000073",
            INIT_18 => X"00000085000000d5000000c0000000b1000000b60000009600000071000000d1",
            INIT_19 => X"000000f7000000fc000000e80000009d00000095000000a20000009c00000098",
            INIT_1A => X"000000940000007700000068000000650000006f0000006e000000730000007d",
            INIT_1B => X"0000008300000082000000870000008d0000008e000000840000008900000084",
            INIT_1C => X"00000087000000a8000000bc000000bc000000c0000000ae000000a4000000ed",
            INIT_1D => X"000000f1000000e4000000990000006f00000069000000690000006b00000065",
            INIT_1E => X"000000730000007800000071000000740000007d0000007d0000007e00000080",
            INIT_1F => X"000000840000008b000000890000008900000087000000860000008b00000085",
            INIT_20 => X"0000008d0000008200000086000000b0000000bf00000089000000b5000000f2",
            INIT_21 => X"000000f5000000af0000007f0000007600000077000000790000007800000074",
            INIT_22 => X"00000075000000750000007300000071000000780000007d0000007d00000082",
            INIT_23 => X"00000086000000910000008e0000008e00000092000000900000008c00000095",
            INIT_24 => X"000000a20000008c0000007c00000088000000a70000008f000000d1000000f9",
            INIT_25 => X"000000cd00000076000000800000007d0000007f0000007f0000007900000073",
            INIT_26 => X"000000710000007000000071000000750000007b00000083000000860000008a",
            INIT_27 => X"000000960000009800000093000000950000009a00000098000000a7000000b6",
            INIT_28 => X"000000a500000093000000820000007a0000007e000000a4000000ea000000f7",
            INIT_29 => X"00000099000000720000007b0000008300000081000000770000007700000077",
            INIT_2A => X"00000077000000770000007b0000007f000000830000008d000000960000009a",
            INIT_2B => X"000000960000008d0000008c0000008a0000009e000000b2000000b6000000a9",
            INIT_2C => X"000000a2000000950000008a000000850000007e0000008a000000e9000000ea",
            INIT_2D => X"0000008c0000007e000000810000007c000000850000007b0000007400000077",
            INIT_2E => X"0000007a0000007e00000082000000840000008c0000008a0000008b00000094",
            INIT_2F => X"000000930000008b0000008500000099000000b6000000b00000008e0000008b",
            INIT_30 => X"000000a1000000930000008f0000008d0000008a0000007d0000009f000000d3",
            INIT_31 => X"000000770000007900000080000000820000008b000000870000008300000078",
            INIT_32 => X"00000076000000780000008200000087000000880000008b0000008a00000088",
            INIT_33 => X"000000870000008a00000097000000b2000000a40000008c0000006700000088",
            INIT_34 => X"000000b10000009400000089000000920000008b000000840000007100000085",
            INIT_35 => X"0000007200000069000000690000007500000080000000870000008900000080",
            INIT_36 => X"00000083000000890000008b0000008a0000008900000088000000830000007d",
            INIT_37 => X"000000850000009a000000b3000000b5000000a8000000920000006c0000007f",
            INIT_38 => X"000000a800000094000000840000008f0000008b000000860000007d00000070",
            INIT_39 => X"0000007300000068000000660000006d0000006a0000006c0000007300000078",
            INIT_3A => X"0000008000000087000000900000009c00000098000000860000007f0000007f",
            INIT_3B => X"00000090000000aa000000c5000000be000000a4000000820000007e0000006b",
            INIT_3C => X"000000a000000095000000840000008600000086000000840000007b00000073",
            INIT_3D => X"0000007200000069000000650000006c000000680000006c0000006200000059",
            INIT_3E => X"000000640000007600000089000000980000009100000083000000820000007b",
            INIT_3F => X"00000091000000a7000000b6000000af000000910000007c000000810000006e",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY5;


    MEM_IFMAP_LAYER0_ENTITY6 : if BRAM_NAME = "ifmap_layer0_entity6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000eb000000e7000000e8000000e8000000e8000000e8000000e8000000e8",
            INIT_01 => X"000000e8000000e8000000e9000000e9000000e9000000e9000000e9000000e9",
            INIT_02 => X"000000e9000000e8000000e7000000e6000000e8000000e8000000e8000000e9",
            INIT_03 => X"000000e8000000e9000000e8000000e8000000e8000000e9000000e9000000e8",
            INIT_04 => X"000000ee000000eb000000eb000000eb000000eb000000eb000000eb000000eb",
            INIT_05 => X"000000eb000000eb000000ec000000ec000000ec000000ec000000ec000000ec",
            INIT_06 => X"000000ed000000ec000000ec000000ea000000ea000000ea000000eb000000ec",
            INIT_07 => X"000000ec000000ec000000eb000000eb000000eb000000ec000000ec000000eb",
            INIT_08 => X"000000ed000000ea000000ea000000ea000000ea000000ea000000ea000000ea",
            INIT_09 => X"000000ea000000ea000000ea000000ea000000ea000000ea000000eb000000eb",
            INIT_0A => X"000000ec000000ec000000eb000000ea000000e3000000e7000000e7000000ea",
            INIT_0B => X"000000ea000000ea000000ea000000ea000000ea000000eb000000eb000000ea",
            INIT_0C => X"000000ee000000eb000000eb000000eb000000eb000000eb000000eb000000eb",
            INIT_0D => X"000000ea000000ea000000ea000000ea000000ea000000ea000000eb000000eb",
            INIT_0E => X"000000e9000000e8000000e4000000df000000ba000000d1000000cf000000e4",
            INIT_0F => X"000000ec000000ea000000ea000000ea000000ea000000eb000000eb000000eb",
            INIT_10 => X"000000ed000000ea000000eb000000eb000000eb000000eb000000eb000000eb",
            INIT_11 => X"000000ea000000ea000000eb000000eb000000ea000000ea000000eb000000eb",
            INIT_12 => X"000000ec000000e9000000db000000cb000000a3000000c3000000d6000000e6",
            INIT_13 => X"000000ed000000eb000000eb000000eb000000eb000000ec000000ec000000ec",
            INIT_14 => X"000000ef000000ec000000ec000000ec000000ec000000ec000000eb000000eb",
            INIT_15 => X"000000ea000000eb000000ed000000ed000000ea000000e8000000eb000000e5",
            INIT_16 => X"000000d0000000c2000000b9000000ae000000a5000000b8000000cf000000e2",
            INIT_17 => X"000000ec000000ec000000ec000000ec000000ec000000ed000000ed000000ed",
            INIT_18 => X"000000e4000000e4000000e8000000e7000000ea000000ed000000ed000000ec",
            INIT_19 => X"000000ed000000ed000000ef000000ef000000e1000000e0000000e9000000dd",
            INIT_1A => X"000000b7000000a10000009f0000009a000000900000008f0000009c000000c6",
            INIT_1B => X"000000e9000000ec000000eb000000eb000000eb000000ec000000ed000000ef",
            INIT_1C => X"000000d4000000e0000000e6000000e3000000e5000000ea000000ed000000ee",
            INIT_1D => X"000000ef000000ef000000ef000000f0000000c9000000db000000e9000000d6",
            INIT_1E => X"000000c1000000b9000000b8000000ad000000a50000009f000000a2000000ba",
            INIT_1F => X"000000e5000000ea000000e9000000e9000000ea000000ec000000ed000000ee",
            INIT_20 => X"000000d8000000dd000000e1000000e1000000e3000000e7000000ec000000ee",
            INIT_21 => X"000000ee000000ee000000ed000000ef000000c5000000dc000000e9000000e6",
            INIT_22 => X"000000d1000000d1000000db000000d0000000d1000000d2000000d9000000da",
            INIT_23 => X"000000e1000000e4000000e4000000e6000000e6000000eb000000ed000000ee",
            INIT_24 => X"00000076000000770000007c00000088000000ac000000e1000000eb000000ed",
            INIT_25 => X"000000ec000000eb000000eb000000e9000000d6000000e2000000e8000000ec",
            INIT_26 => X"000000e4000000e3000000e7000000e1000000e1000000d9000000c9000000b9",
            INIT_27 => X"000000ac000000a7000000a7000000ba000000df000000eb000000ec000000ee",
            INIT_28 => X"0000006d000000670000006c0000006f00000092000000de000000e3000000e5",
            INIT_29 => X"000000ec000000ea000000e7000000e6000000e5000000e7000000e8000000e6",
            INIT_2A => X"000000e7000000e7000000e5000000df000000bf000000a40000009200000089",
            INIT_2B => X"00000086000000800000007900000095000000d8000000ea000000eb000000ed",
            INIT_2C => X"000000c3000000bc000000c7000000c8000000d1000000df000000d5000000d3",
            INIT_2D => X"000000d8000000dc000000db000000d2000000d1000000d3000000d8000000dc",
            INIT_2E => X"000000e1000000e2000000e1000000da000000b7000000af000000b5000000b2",
            INIT_2F => X"000000ba000000aa0000008e000000b9000000db000000e7000000ea000000ec",
            INIT_30 => X"000000c1000000bf000000ca000000d6000000df000000d6000000cb000000ab",
            INIT_31 => X"000000b1000000cf000000ae000000620000005d000000650000006f0000007a",
            INIT_32 => X"0000008900000099000000ca000000df000000da000000dc000000df000000d9",
            INIT_33 => X"000000dd000000d4000000c4000000de000000db000000dd000000e8000000eb",
            INIT_34 => X"000000710000006f000000710000007d0000008a000000aa000000bf000000be",
            INIT_35 => X"000000d0000000d80000009e000000360000002d000000310000003500000042",
            INIT_36 => X"000000660000009f000000dd000000ea000000e9000000e3000000df000000cf",
            INIT_37 => X"000000ca000000d3000000d4000000c7000000b3000000bc000000d3000000dd",
            INIT_38 => X"0000003d000000450000003f000000440000007b0000008b00000097000000c3",
            INIT_39 => X"000000d6000000ce000000a3000000670000005f000000650000008a000000b5",
            INIT_3A => X"000000cf000000dd000000db000000cd000000b70000009e0000009300000083",
            INIT_3B => X"0000007d000000820000008800000085000000800000008a000000b6000000c5",
            INIT_3C => X"000000280000003a000000550000007f000000840000006000000077000000a3",
            INIT_3D => X"000000ad000000b8000000b6000000b5000000b7000000c6000000da000000c8",
            INIT_3E => X"000000ae0000009f000000910000008400000074000000620000005e00000063",
            INIT_3F => X"000000690000006b0000007a0000008a000000960000009d000000bc000000b9",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY6;


    MEM_IFMAP_LAYER0_ENTITY7 : if BRAM_NAME = "ifmap_layer0_entity7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000d0000001a00000086000000ce0000008a000000760000008d000000ac",
            INIT_01 => X"000000b5000000cf000000dc000000e4000000e0000000e6000000e2000000b0",
            INIT_02 => X"000000900000008a0000008e000000910000009a00000095000000950000009a",
            INIT_03 => X"0000009d000000a0000000ad000000bb000000be000000b2000000a50000009d",
            INIT_04 => X"000000050000003a000000c8000000e1000000c5000000c7000000d4000000e2",
            INIT_05 => X"000000e5000000e9000000e8000000e6000000d1000000df000000dd000000d2",
            INIT_06 => X"000000c6000000b4000000c1000000bc000000bd000000c2000000c0000000b8",
            INIT_07 => X"000000ac000000ab000000a1000000900000008800000083000000800000008a",
            INIT_08 => X"0000002700000091000000be000000ba000000b8000000c0000000c2000000c2",
            INIT_09 => X"000000c2000000bf000000c0000000be000000b1000000b40000009a00000093",
            INIT_0A => X"000000910000009c000000920000007100000072000000840000007e0000006f",
            INIT_0B => X"0000005c0000005b0000005d0000005e00000069000000790000008100000081",
            INIT_0C => X"0000007a000000a20000008f0000008900000083000000800000007f00000082",
            INIT_0D => X"00000083000000800000007f00000081000000810000007c0000006800000064",
            INIT_0E => X"0000006600000076000000700000005e0000005e0000005e0000005700000053",
            INIT_0F => X"00000050000000530000005d000000650000006c000000730000007900000082",
            INIT_10 => X"000000490000004c0000004d000000500000005400000057000000570000005a",
            INIT_11 => X"0000005e000000660000006b0000007100000073000000760000007600000078",
            INIT_12 => X"000000730000006e0000006a000000640000005f000000550000004f00000050",
            INIT_13 => X"000000500000004d00000050000000520000005c000000710000007d00000088",
            INIT_14 => X"0000000d00000003000000090000001200000012000000150000001400000016",
            INIT_15 => X"0000001a000000220000002a00000030000000340000003c0000004200000046",
            INIT_16 => X"0000004700000048000000430000003c00000037000000350000003500000039",
            INIT_17 => X"0000003900000039000000480000005700000068000000780000008200000089",
            INIT_18 => X"000000240000000b000000080000002000000024000000160000000800000003",
            INIT_19 => X"0000000100000000000000000000000000000006000000050000000100000003",
            INIT_1A => X"0000000d00000018000000150000001500000015000000160000001e00000027",
            INIT_1B => X"0000003900000055000000710000007b000000740000007a0000008600000099",
            INIT_1C => X"000000230000001a0000000d0000001b0000004700000046000000310000001b",
            INIT_1D => X"0000000f00000005000000020000000000000011000000390000001f0000000a",
            INIT_1E => X"0000000400000004000000070000000e00000019000000290000003e00000056",
            INIT_1F => X"0000007a000000900000008400000072000000750000008400000092000000ac",
            INIT_20 => X"000000100000000d00000004000000030000002d000000410000003600000024",
            INIT_21 => X"000000120000000400000002000000000000000700000076000000a100000083",
            INIT_22 => X"0000007000000069000000690000006d000000760000008a0000009a00000097",
            INIT_23 => X"0000007f000000690000006a00000078000000810000008e000000a4000000b8",
            INIT_24 => X"000000280000000c00000000000000000000000c0000001e0000002000000015",
            INIT_25 => X"000000070000000200000002000000030000000000000044000000b6000000cd",
            INIT_26 => X"000000c4000000c2000000c3000000bb000000ac000000960000007b00000067",
            INIT_27 => X"0000005f000000680000007a000000810000008400000098000000ab000000b9",
            INIT_28 => X"000000450000001a0000000100000001000000040000000c000000120000000c",
            INIT_29 => X"00000004000000020000000200000004000000010000002000000099000000cb",
            INIT_2A => X"000000c3000000bf000000b30000009b000000770000005b000000510000005e",
            INIT_2B => X"000000750000007d0000007d0000008100000090000000a2000000ad000000b8",
            INIT_2C => X"000000530000002f000000010000000200000002000000050000000700000004",
            INIT_2D => X"00000001000000010000000100000003000000010000001b0000008e000000cd",
            INIT_2E => X"000000c6000000a900000079000000550000004a000000550000006600000079",
            INIT_2F => X"000000800000007a000000790000008400000093000000a5000000b0000000ba",
            INIT_30 => X"0000005c00000036000000060000000300000002000000010000000100000001",
            INIT_31 => X"00000001000000010000000100000001000000000000000f000000660000009d",
            INIT_32 => X"000000750000004a000000380000004a00000063000000730000007a0000007c",
            INIT_33 => X"0000007b0000007d000000800000008800000094000000a2000000b1000000bc",
            INIT_34 => X"000000570000002b000000130000000b00000008000000050000000200000002",
            INIT_35 => X"0000000300000003000000030000000200000000000000040000002a00000047",
            INIT_36 => X"0000003500000039000000500000007100000084000000860000007b00000074",
            INIT_37 => X"00000078000000830000008b0000008f0000009c000000a9000000b6000000bc",
            INIT_38 => X"000000520000002e000000240000001f0000001b000000160000001100000010",
            INIT_39 => X"0000001200000013000000140000001300000013000000170000002500000040",
            INIT_3A => X"000000570000006800000074000000800000008b000000830000007500000073",
            INIT_3B => X"0000007b000000830000008b000000940000009f000000ae000000b9000000bb",
            INIT_3C => X"000000550000003e0000003a00000037000000330000002f0000002e00000030",
            INIT_3D => X"000000310000003300000035000000370000003b000000440000005100000068",
            INIT_3E => X"000000740000007f000000850000007f0000007f00000076000000720000007a",
            INIT_3F => X"00000081000000880000008d000000950000009e000000a8000000b4000000ba",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY7;


    MEM_IFMAP_LAYER0_ENTITY8 : if BRAM_NAME = "ifmap_layer0_entity8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000eb000000e7000000e8000000e8000000e8000000e8000000e8000000e8",
            INIT_01 => X"000000e8000000e8000000e9000000e9000000e9000000e9000000e9000000e8",
            INIT_02 => X"000000e7000000e7000000e9000000e9000000e8000000e7000000e8000000e9",
            INIT_03 => X"000000e9000000e9000000e8000000e8000000e8000000e9000000e9000000e8",
            INIT_04 => X"000000ee000000eb000000eb000000eb000000eb000000eb000000eb000000eb",
            INIT_05 => X"000000eb000000eb000000ec000000ec000000ec000000ec000000ec000000ec",
            INIT_06 => X"000000ea000000ea000000ec000000ec000000eb000000ea000000ec000000ec",
            INIT_07 => X"000000ec000000ec000000eb000000eb000000eb000000ec000000ec000000eb",
            INIT_08 => X"000000ed000000ea000000ea000000ea000000ea000000ea000000ea000000ea",
            INIT_09 => X"000000ea000000ea000000ea000000ea000000ea000000ea000000eb000000ea",
            INIT_0A => X"000000e9000000ea000000eb000000eb000000e6000000eb000000e9000000ea",
            INIT_0B => X"000000ea000000ea000000ea000000ea000000ea000000eb000000eb000000ea",
            INIT_0C => X"000000ee000000eb000000eb000000eb000000eb000000eb000000eb000000eb",
            INIT_0D => X"000000ea000000ea000000ea000000ea000000ea000000ea000000eb000000eb",
            INIT_0E => X"000000e9000000e8000000e6000000e2000000c0000000d8000000d2000000e4",
            INIT_0F => X"000000eb000000ea000000ea000000ea000000ea000000eb000000eb000000eb",
            INIT_10 => X"000000ed000000ea000000eb000000eb000000eb000000eb000000eb000000eb",
            INIT_11 => X"000000ea000000ea000000eb000000eb000000ea000000ea000000eb000000eb",
            INIT_12 => X"000000ee000000ed000000e1000000d2000000ac000000cd000000da000000e5",
            INIT_13 => X"000000eb000000eb000000eb000000eb000000ec000000ec000000ec000000ec",
            INIT_14 => X"000000ef000000eb000000eb000000eb000000eb000000eb000000ec000000eb",
            INIT_15 => X"000000ea000000eb000000ec000000ec000000eb000000e9000000ed000000e7",
            INIT_16 => X"000000d8000000cd000000c6000000bc000000b3000000c4000000d7000000e4",
            INIT_17 => X"000000eb000000ec000000ec000000ec000000ec000000ed000000ed000000ed",
            INIT_18 => X"000000e5000000e3000000e6000000e4000000e8000000ec000000ed000000ed",
            INIT_19 => X"000000eb000000eb000000ec000000ed000000e5000000e4000000ed000000e2",
            INIT_1A => X"000000c5000000b4000000b4000000b0000000a30000009f000000a9000000ce",
            INIT_1B => X"000000ee000000ed000000ec000000eb000000ec000000ee000000ed000000ed",
            INIT_1C => X"000000dc000000e6000000ea000000e8000000ea000000ed000000ee000000ed",
            INIT_1D => X"000000ed000000ed000000ec000000ee000000cc000000de000000ec000000da",
            INIT_1E => X"000000cc000000c9000000c9000000bf000000b6000000ae000000b0000000c7",
            INIT_1F => X"000000ef000000ef000000ee000000ee000000ef000000ef000000ef000000ee",
            INIT_20 => X"000000ea000000ec000000ee000000ef000000f0000000ee000000ed000000ec",
            INIT_21 => X"000000ec000000ec000000ed000000ef000000c6000000dd000000ea000000e7",
            INIT_22 => X"000000d5000000d8000000e4000000da000000dd000000e0000000e9000000eb",
            INIT_23 => X"000000f0000000ee000000ef000000f0000000f0000000f0000000f0000000ee",
            INIT_24 => X"0000008c0000008a0000008e0000009b000000bc000000ea000000ec000000ea",
            INIT_25 => X"000000e9000000eb000000ed000000ed000000d8000000e4000000ea000000ed",
            INIT_26 => X"000000e6000000e6000000ec000000e8000000ed000000e9000000db000000cc",
            INIT_27 => X"000000bd000000b3000000b4000000c7000000eb000000f1000000f0000000f0",
            INIT_28 => X"00000082000000790000007d0000007f0000009f000000e5000000e4000000e2",
            INIT_29 => X"000000e8000000ea000000ec000000ed000000ea000000eb000000ed000000eb",
            INIT_2A => X"000000ec000000ed000000ed000000e8000000ce000000b8000000a50000009c",
            INIT_2B => X"000000950000008c00000085000000a2000000e4000000f1000000f0000000f0",
            INIT_2C => X"000000d4000000ca000000d3000000d3000000d9000000e3000000d5000000d1",
            INIT_2D => X"000000d5000000de000000e2000000dd000000db000000dd000000e1000000e5",
            INIT_2E => X"000000ea000000ec000000ed000000e7000000cc000000c6000000c8000000c2",
            INIT_2F => X"000000c5000000b200000097000000c3000000e6000000f0000000f1000000f0",
            INIT_30 => X"000000cf000000ca000000d3000000d9000000e1000000db000000d0000000ae",
            INIT_31 => X"000000b4000000d5000000b8000000700000007200000079000000810000008a",
            INIT_32 => X"00000098000000a7000000d8000000ec000000e8000000e9000000ea000000e2",
            INIT_33 => X"000000e4000000db000000cb000000e6000000e3000000e6000000ef000000f1",
            INIT_34 => X"000000820000007d0000007d0000008300000091000000b6000000c9000000c7",
            INIT_35 => X"000000db000000e6000000ac0000004700000046000000490000004900000054",
            INIT_36 => X"00000072000000a8000000e3000000ef000000ed000000e7000000e4000000d3",
            INIT_37 => X"000000d0000000da000000db000000ce000000ba000000c5000000dd000000e7",
            INIT_38 => X"00000051000000560000004f000000550000008d0000009b0000009d000000c8",
            INIT_39 => X"000000e4000000df000000b400000079000000700000007500000097000000c0",
            INIT_3A => X"000000d4000000de000000db000000cb000000ba000000a60000009a0000008a",
            INIT_3B => X"000000850000008b000000920000008e0000008900000099000000c5000000d4",
            INIT_3C => X"00000035000000460000006200000090000000970000006b000000730000009e",
            INIT_3D => X"000000b4000000c2000000c2000000c1000000c2000000d1000000e4000000d2",
            INIT_3E => X"000000b5000000a500000096000000880000007d0000006f0000006a0000006f",
            INIT_3F => X"00000076000000790000008700000097000000a4000000ae000000ce000000cb",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY8;


    MEM_IFMAP_LAYER0_ENTITY9 : if BRAM_NAME = "ifmap_layer0_entity9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000f0000001d0000008c000000d8000000960000007b00000085000000a2",
            INIT_01 => X"000000b5000000d1000000e0000000ea000000ea000000f1000000ee000000bd",
            INIT_02 => X"0000009f0000009a0000009e000000a3000000ab000000a5000000a5000000ab",
            INIT_03 => X"000000ae000000b1000000be000000cc000000cf000000c4000000b7000000af",
            INIT_04 => X"000000050000003e000000cf000000e8000000cd000000cf000000d4000000e0",
            INIT_05 => X"000000e6000000ec000000ee000000ee000000dd000000ee000000ee000000e4",
            INIT_06 => X"000000d9000000c8000000d8000000d5000000d4000000d6000000d4000000cc",
            INIT_07 => X"000000c1000000bf000000b5000000a50000009c000000920000008f0000009a",
            INIT_08 => X"0000002d0000009b000000cc000000c4000000c5000000d3000000d3000000d0",
            INIT_09 => X"000000ce000000cb000000cf000000cf000000c1000000c6000000b0000000a9",
            INIT_0A => X"000000a1000000ab000000a300000085000000890000009d0000009600000087",
            INIT_0B => X"000000730000007000000072000000740000007d000000850000008d0000008e",
            INIT_0C => X"00000087000000b3000000a00000009a00000098000000980000009600000096",
            INIT_0D => X"0000009600000093000000930000009500000095000000910000007e0000007a",
            INIT_0E => X"0000007800000086000000800000006d00000070000000750000007000000067",
            INIT_0F => X"00000061000000670000006f00000075000000790000007d0000008500000090",
            INIT_10 => X"000000570000005a0000005a0000005d00000062000000660000006600000069",
            INIT_11 => X"0000006f000000770000007c0000008300000089000000880000008400000085",
            INIT_12 => X"00000088000000850000007f000000770000006d00000065000000610000005c",
            INIT_13 => X"0000005e00000064000000640000006200000068000000770000008700000095",
            INIT_14 => X"000000190000000b000000100000001a0000001a00000019000000190000001e",
            INIT_15 => X"000000240000002b000000330000003b000000450000004b0000004d0000004f",
            INIT_16 => X"0000005700000058000000510000004800000043000000440000004500000045",
            INIT_17 => X"000000470000004e0000005900000064000000710000007c0000008800000092",
            INIT_18 => X"0000002e000000100000000d0000002c0000002d000000190000000b00000008",
            INIT_19 => X"000000040000000200000002000000040000000d000000120000001300000017",
            INIT_1A => X"0000001d00000026000000210000001f000000260000002c000000320000003a",
            INIT_1B => X"000000460000005a000000730000007b000000730000007b0000008b000000a0",
            INIT_1C => X"000000290000001b00000013000000290000005100000046000000320000001f",
            INIT_1D => X"0000000f00000005000000020000000000000011000000400000003200000024",
            INIT_1E => X"0000001e0000001e0000001e000000230000002b000000370000004700000061",
            INIT_1F => X"0000007c0000008300000078000000690000006f0000008600000098000000b3",
            INIT_20 => X"0000000f0000000a0000000a0000000c0000002c000000340000002b00000021",
            INIT_21 => X"0000001200000004000000020000000100000008000000750000009e00000080",
            INIT_22 => X"000000700000006900000067000000690000006b000000730000007e0000007e",
            INIT_23 => X"0000006a000000560000005e000000740000008200000093000000ac000000c2",
            INIT_24 => X"000000280000000a0000000300000004000000060000000c0000000c0000000a",
            INIT_25 => X"00000006000000010000000100000002000000000000003a0000008000000082",
            INIT_26 => X"0000007f0000007b00000077000000710000006e000000600000004b00000042",
            INIT_27 => X"000000470000005d00000076000000840000008d000000a2000000b6000000c5",
            INIT_28 => X"0000004d0000001d000000010000000100000001000000020000000300000002",
            INIT_29 => X"00000001000000000000000000000000000000010000000c0000002d0000002f",
            INIT_2A => X"0000002e0000003000000032000000310000002a00000026000000300000004d",
            INIT_2B => X"0000006e0000007e000000800000008700000099000000b0000000bb000000c6",
            INIT_2C => X"0000005e00000034000000010000000100000000000000010000000100000000",
            INIT_2D => X"0000000000000000000000000000000000000002000000030000001900000020",
            INIT_2E => X"0000001900000019000000190000001d00000029000000420000005c00000071",
            INIT_2F => X"0000007c0000007e0000007f0000008b0000009d000000b3000000bf000000c9",
            INIT_30 => X"000000660000003c000000070000000200000002000000030000000300000002",
            INIT_31 => X"000000010000000000000000000000010000000300000001000000130000001f",
            INIT_32 => X"000000110000000d0000001b0000003a0000005a000000730000007e0000007c",
            INIT_33 => X"0000007b0000008200000087000000910000009f000000b0000000c0000000ca",
            INIT_34 => X"0000006300000033000000170000000c0000000a0000000b0000000a00000007",
            INIT_35 => X"0000000400000004000000040000000300000006000000050000000d00000015",
            INIT_36 => X"0000001b000000320000004d00000062000000710000007e0000007e0000007d",
            INIT_37 => X"000000800000008a000000940000009a000000a8000000b8000000c5000000ca",
            INIT_38 => X"00000060000000390000002c000000230000001e0000001c0000001a00000017",
            INIT_39 => X"000000150000001500000016000000170000001b0000001f0000002800000037",
            INIT_3A => X"00000046000000580000006600000070000000790000007a0000007a0000007f",
            INIT_3B => X"000000850000008b00000095000000a0000000ac000000bd000000c8000000ca",
            INIT_3C => X"000000650000004b000000430000003d00000038000000350000003500000037",
            INIT_3D => X"00000037000000380000003a0000003e00000043000000470000005400000060",
            INIT_3E => X"000000670000006d00000074000000790000007f0000007c0000007d00000083",
            INIT_3F => X"000000880000009100000098000000a2000000ab000000b7000000c3000000c8",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY9;


    MEM_IFMAP_LAYER0_ENTITY10 : if BRAM_NAME = "ifmap_layer0_entity10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000eb000000e7000000e8000000e8000000e8000000e8000000e8000000e8",
            INIT_01 => X"000000e8000000e8000000e9000000e9000000e9000000e9000000e9000000e9",
            INIT_02 => X"000000e9000000e9000000e9000000e8000000ea000000ea000000e8000000e6",
            INIT_03 => X"000000e7000000e9000000e8000000e8000000e8000000e9000000e9000000e8",
            INIT_04 => X"000000ee000000eb000000eb000000eb000000eb000000eb000000eb000000eb",
            INIT_05 => X"000000eb000000eb000000ec000000ec000000ec000000ec000000ec000000ec",
            INIT_06 => X"000000e9000000e9000000ea000000ea000000ed000000ee000000ed000000eb",
            INIT_07 => X"000000ea000000ec000000eb000000eb000000eb000000ec000000ec000000eb",
            INIT_08 => X"000000ed000000ea000000ea000000ea000000ea000000ea000000ea000000ea",
            INIT_09 => X"000000ea000000ea000000ea000000ea000000ea000000ea000000eb000000ea",
            INIT_0A => X"000000e7000000e7000000ea000000ec000000e9000000ee000000eb000000ea",
            INIT_0B => X"000000ea000000ea000000ea000000ea000000ea000000eb000000eb000000ea",
            INIT_0C => X"000000ee000000eb000000eb000000eb000000eb000000eb000000eb000000eb",
            INIT_0D => X"000000ea000000ea000000ea000000ea000000ea000000ea000000eb000000ea",
            INIT_0E => X"000000e6000000e7000000e8000000e7000000c5000000db000000d5000000e6",
            INIT_0F => X"000000eb000000ea000000ea000000ea000000ea000000eb000000eb000000eb",
            INIT_10 => X"000000ed000000ea000000eb000000eb000000eb000000eb000000eb000000eb",
            INIT_11 => X"000000ea000000ea000000eb000000eb000000ea000000ea000000eb000000eb",
            INIT_12 => X"000000ec000000ed000000e6000000db000000b3000000d0000000dd000000e8",
            INIT_13 => X"000000ed000000eb000000eb000000eb000000ec000000ec000000ec000000ec",
            INIT_14 => X"000000ee000000eb000000eb000000eb000000eb000000eb000000eb000000eb",
            INIT_15 => X"000000ea000000eb000000ec000000ec000000ec000000ea000000ed000000e8",
            INIT_16 => X"000000da000000d2000000cf000000c8000000bd000000ca000000dc000000e8",
            INIT_17 => X"000000ed000000eb000000eb000000eb000000ec000000ed000000ed000000ed",
            INIT_18 => X"000000e5000000e4000000e7000000e6000000e9000000ec000000eb000000eb",
            INIT_19 => X"000000ec000000ec000000ed000000ee000000e6000000e5000000ee000000e4",
            INIT_1A => X"000000cc000000be000000bf000000be000000b1000000ab000000b1000000d3",
            INIT_1B => X"000000ef000000ea000000e9000000eb000000ec000000ed000000ed000000ee",
            INIT_1C => X"000000de000000e9000000ee000000ea000000ea000000ec000000eb000000ec",
            INIT_1D => X"000000ee000000ee000000ed000000ef000000cb000000dd000000eb000000da",
            INIT_1E => X"000000d2000000d2000000d3000000cb000000c4000000bb000000b9000000cc",
            INIT_1F => X"000000f0000000ee000000ed000000ee000000ee000000ee000000ee000000ee",
            INIT_20 => X"000000f1000000f3000000f6000000f3000000f0000000ed000000eb000000eb",
            INIT_21 => X"000000ed000000ed000000ed000000ef000000c4000000da000000e7000000e5",
            INIT_22 => X"000000d9000000de000000eb000000e3000000ea000000eb000000f0000000f1",
            INIT_23 => X"000000f3000000f0000000f0000000f0000000ef000000ef000000ef000000ee",
            INIT_24 => X"000000950000009400000099000000a1000000bf000000e9000000e9000000e8",
            INIT_25 => X"000000ea000000eb000000ec000000eb000000d6000000e2000000e8000000ec",
            INIT_26 => X"000000e8000000eb000000f1000000ef000000f7000000f3000000e2000000d3",
            INIT_27 => X"000000c3000000ba000000b9000000c9000000eb000000ef000000ef000000ef",
            INIT_28 => X"0000008d000000850000008900000089000000a5000000e7000000e1000000e0",
            INIT_29 => X"000000e9000000ea000000ea000000eb000000eb000000ec000000ee000000ec",
            INIT_2A => X"000000ee000000f0000000f1000000ee000000d5000000bf000000ac000000a3",
            INIT_2B => X"0000009f000000990000008f000000a6000000e5000000ef000000ee000000ef",
            INIT_2C => X"000000e0000000d7000000e0000000df000000e3000000e7000000d3000000ce",
            INIT_2D => X"000000d6000000de000000e1000000db000000df000000e1000000e6000000e9",
            INIT_2E => X"000000ed000000ef000000f1000000ed000000d0000000cb000000cf000000ca",
            INIT_2F => X"000000d3000000c4000000a4000000ca000000e9000000ee000000ef000000ef",
            INIT_30 => X"000000de000000d9000000e0000000ea000000f1000000e3000000d0000000ae",
            INIT_31 => X"000000b7000000d6000000bc000000790000007e000000840000008b00000093",
            INIT_32 => X"000000a1000000ae000000dc000000ed000000eb000000ee000000f0000000e9",
            INIT_33 => X"000000ed000000e5000000d4000000ed000000ea000000e9000000f2000000f2",
            INIT_34 => X"00000098000000930000008d00000097000000a5000000c1000000cd000000cc",
            INIT_35 => X"000000e2000000ea000000b70000005c0000005b0000005b0000005a00000062",
            INIT_36 => X"00000081000000b3000000e9000000f1000000f1000000ed000000e9000000d9",
            INIT_37 => X"000000d4000000dc000000df000000d6000000c4000000cd000000e3000000ea",
            INIT_38 => X"0000006c0000007200000064000000660000009b000000a4000000a4000000cf",
            INIT_39 => X"000000ea000000e4000000be0000008a0000008300000087000000a8000000cf",
            INIT_3A => X"000000df000000e8000000e3000000d4000000c3000000ae000000a300000093",
            INIT_3B => X"0000008c00000090000000980000009700000093000000a0000000cb000000d8",
            INIT_3C => X"0000004d0000005e00000074000000990000009c0000006e00000076000000a1",
            INIT_3D => X"000000b6000000c5000000c6000000c8000000ca000000d9000000ec000000d9",
            INIT_3E => X"000000ba000000ac0000009f000000950000008a0000007b000000760000007b",
            INIT_3F => X"000000800000008200000091000000a1000000ae000000b8000000d5000000d0",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY10;


    MEM_IFMAP_LAYER0_ENTITY11 : if BRAM_NAME = "ifmap_layer0_entity11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000230000002f00000097000000dc000000960000007b00000086000000a2",
            INIT_01 => X"000000b4000000d3000000e1000000e9000000e8000000f0000000ee000000be",
            INIT_02 => X"000000a3000000a2000000aa000000b1000000bb000000b6000000b6000000bb",
            INIT_03 => X"000000bd000000bf000000cc000000d9000000da000000d0000000c1000000b7",
            INIT_04 => X"000000180000004f000000d9000000ef000000d4000000d3000000da000000e5",
            INIT_05 => X"000000ed000000f6000000f5000000ef000000dc000000ef000000f1000000ea",
            INIT_06 => X"000000e4000000d6000000e6000000e5000000e7000000ea000000e8000000e0",
            INIT_07 => X"000000d4000000d1000000c5000000b3000000a9000000a10000009e000000a5",
            INIT_08 => X"00000047000000b3000000de000000d8000000d9000000e5000000e6000000e3",
            INIT_09 => X"000000e3000000e4000000e4000000dd000000cf000000d7000000c1000000bc",
            INIT_0A => X"000000b8000000c3000000ba0000009c000000a1000000b4000000ad0000009e",
            INIT_0B => X"0000008a0000008700000085000000830000008c000000970000009e0000009c",
            INIT_0C => X"000000a1000000cf000000c2000000bd000000bb000000be000000c0000000c1",
            INIT_0D => X"000000c0000000be000000bd000000bd000000bc000000ba000000a30000009a",
            INIT_0E => X"0000009a000000aa000000a30000009100000094000000990000009000000088",
            INIT_0F => X"00000082000000860000008b0000008d0000009000000092000000940000009c",
            INIT_10 => X"0000006d000000710000007a0000007f000000860000008e0000009300000096",
            INIT_11 => X"00000098000000a0000000a5000000ac000000b5000000ba000000b4000000af",
            INIT_12 => X"000000ac000000a8000000a30000009b000000940000008b000000840000007f",
            INIT_13 => X"0000008100000085000000810000007a0000007e0000008a000000920000009c",
            INIT_14 => X"0000002900000019000000230000003000000034000000380000003a0000003d",
            INIT_15 => X"0000003e000000460000004d000000570000006a000000790000007e0000007e",
            INIT_16 => X"0000007f0000007e00000078000000700000006a000000680000006700000066",
            INIT_17 => X"000000690000006e000000730000007700000080000000880000008d00000095",
            INIT_18 => X"000000370000001400000013000000350000003a000000290000001e00000018",
            INIT_19 => X"000000110000000f0000000f000000140000002a000000380000003c0000003e",
            INIT_1A => X"00000047000000510000004d0000004c0000004e0000004f000000530000005a",
            INIT_1B => X"00000065000000760000008a0000008a0000007d00000080000000890000009e",
            INIT_1C => X"0000002d0000001a0000001200000029000000540000004c0000003900000025",
            INIT_1D => X"000000150000000b0000000700000007000000230000005b0000004e0000003e",
            INIT_1E => X"0000003c0000003e0000003f000000450000004a00000053000000630000007b",
            INIT_1F => X"00000092000000950000008700000072000000740000008500000092000000af",
            INIT_20 => X"0000001100000009000000080000000b0000002e000000390000002f00000023",
            INIT_21 => X"000000140000000700000004000000030000000f00000086000000b300000094",
            INIT_22 => X"000000830000007d0000007c0000007f0000007e00000085000000900000008d",
            INIT_23 => X"000000740000005b00000061000000740000008100000090000000a5000000be",
            INIT_24 => X"000000230000000700000003000000040000000700000011000000110000000c",
            INIT_25 => X"0000000700000003000000020000000300000002000000400000009200000094",
            INIT_26 => X"000000900000008d00000089000000810000007a0000006a0000005300000045",
            INIT_27 => X"0000004600000058000000710000007e000000870000009e000000b0000000c2",
            INIT_28 => X"0000004000000015000000010000000200000000000000050000000900000005",
            INIT_29 => X"00000002000000000000000000000001000000010000000b0000003b00000044",
            INIT_2A => X"0000004300000045000000430000003b000000310000002a0000002e00000047",
            INIT_2B => X"0000006600000074000000780000008000000093000000ab000000b7000000c4",
            INIT_2C => X"000000520000002b000000010000000200000000000000020000000500000002",
            INIT_2D => X"0000000000000000000000000000000000000000000000020000002600000036",
            INIT_2E => X"0000002e0000002b000000240000002200000027000000380000005200000069",
            INIT_2F => X"0000007300000073000000760000008300000096000000ae000000bb000000c7",
            INIT_30 => X"0000005d00000032000000030000000100000000000000010000000300000002",
            INIT_31 => X"0000000100000000000000000000000100000002000000000000001c0000002f",
            INIT_32 => X"000000170000000c000000160000003700000051000000630000006f00000070",
            INIT_33 => X"00000071000000770000007e0000008900000097000000ab000000bc000000c9",
            INIT_34 => X"00000059000000250000000b0000000400000002000000040000000400000002",
            INIT_35 => X"0000000100000001000000010000000200000006000000020000000d00000018",
            INIT_36 => X"00000019000000290000003e000000520000006500000071000000700000006f",
            INIT_37 => X"000000730000007e0000008900000091000000a1000000b3000000c1000000c9",
            INIT_38 => X"000000520000002400000016000000110000000f0000000f0000000d0000000c",
            INIT_39 => X"0000000c0000000d0000000e0000000f00000014000000150000001b0000002d",
            INIT_3A => X"00000043000000510000005500000058000000690000006e0000006b00000070",
            INIT_3B => X"000000770000007f0000008a00000097000000a4000000b7000000c4000000c8",
            INIT_3C => X"0000005300000030000000260000002500000023000000210000002200000026",
            INIT_3D => X"00000028000000290000002c0000002e0000002d000000300000003b0000004a",
            INIT_3E => X"000000530000005c00000061000000610000006b0000006a0000006c00000075",
            INIT_3F => X"0000007b000000850000008d00000099000000a3000000b2000000bf000000c7",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY11;


    MEM_IFMAP_LAYER0_ENTITY12 : if BRAM_NAME = "ifmap_layer0_entity12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009e0000009e0000008b00000084000000a6000000b6000000bb000000c1",
            INIT_01 => X"000000c7000000cd000000d1000000ce000000da000000df000000e3000000e6",
            INIT_02 => X"000000d5000000e2000000e7000000eb000000ec000000e8000000ea000000ea",
            INIT_03 => X"000000ec000000e2000000e6000000ee000000e8000000e4000000ed000000ee",
            INIT_04 => X"000000aa000000ac0000009700000089000000ae000000c1000000c5000000c7",
            INIT_05 => X"000000ce000000d7000000d9000000d2000000e1000000e7000000e9000000ed",
            INIT_06 => X"000000db000000e4000000e8000000f2000000f5000000ea000000ec000000f2",
            INIT_07 => X"000000f1000000e4000000eb000000f3000000e9000000e8000000f6000000f6",
            INIT_08 => X"000000ae000000b00000009d0000008e000000b5000000c9000000ce000000c7",
            INIT_09 => X"000000d1000000df000000da000000d4000000e0000000e6000000e6000000ef",
            INIT_0A => X"000000dd000000e4000000e9000000ef000000e8000000d5000000ec000000f3",
            INIT_0B => X"000000f5000000e7000000ee000000f8000000ed000000e6000000fa000000f5",
            INIT_0C => X"000000b4000000b2000000a000000093000000ba000000cb000000d4000000cf",
            INIT_0D => X"000000d6000000e4000000dd000000d6000000dc000000e7000000df000000f0",
            INIT_0E => X"000000e0000000e4000000e9000000e4000000b1000000ac000000e6000000f3",
            INIT_0F => X"000000f8000000e8000000ee000000fa000000ee000000e4000000f9000000f4",
            INIT_10 => X"000000ba000000b9000000a500000093000000bd000000cc000000d9000000cf",
            INIT_11 => X"000000d3000000e7000000de000000d6000000da000000e7000000d3000000eb",
            INIT_12 => X"000000e2000000e0000000e8000000d40000009f000000a8000000e0000000ed",
            INIT_13 => X"000000f7000000e7000000eb000000f6000000e8000000ea000000f8000000f2",
            INIT_14 => X"000000c1000000be000000aa0000008e000000bf000000cb000000db000000d3",
            INIT_15 => X"000000d7000000ea000000dd000000d6000000d6000000e4000000c7000000cd",
            INIT_16 => X"000000cf000000ce000000eb000000c1000000700000009e000000de000000e6",
            INIT_17 => X"000000f5000000e5000000e2000000f1000000e4000000e7000000f3000000eb",
            INIT_18 => X"000000c4000000bf000000ac00000085000000bf000000ca000000de000000d9",
            INIT_19 => X"000000df000000eb000000da000000d6000000d7000000e3000000bc000000b0",
            INIT_1A => X"000000bb000000ba000000cd000000bb0000007800000089000000ac000000b7",
            INIT_1B => X"000000db000000df000000d8000000eb000000e2000000e1000000f0000000eb",
            INIT_1C => X"000000cc000000c5000000ae0000008c000000cb000000da000000e0000000e0",
            INIT_1D => X"000000e8000000ed000000dc000000dc000000dc000000dd000000c9000000cd",
            INIT_1E => X"000000ac0000008a0000006400000053000000470000003e000000410000003c",
            INIT_1F => X"00000068000000b6000000d1000000e4000000da000000d4000000ef000000ec",
            INIT_20 => X"000000af000000aa0000009d00000089000000b0000000ba000000af000000c5",
            INIT_21 => X"000000d1000000d4000000ce000000d2000000d4000000c9000000c1000000c1",
            INIT_22 => X"0000008e00000069000000590000005b00000054000000530000005e00000045",
            INIT_23 => X"0000004e00000079000000a2000000b7000000ae000000a3000000cf000000c3",
            INIT_24 => X"00000072000000730000007100000068000000690000006b0000006f00000080",
            INIT_25 => X"0000008b00000092000000970000009b0000009d000000930000009700000096",
            INIT_26 => X"0000007600000064000000630000006300000055000000560000005600000053",
            INIT_27 => X"0000008b000000800000009a00000099000000760000006d000000840000007b",
            INIT_28 => X"000000420000004c0000004b00000044000000530000005a000000540000005a",
            INIT_29 => X"0000005d0000006a00000066000000670000006a0000006b000000720000006c",
            INIT_2A => X"0000005a0000005a0000005b0000005500000048000000420000005f00000072",
            INIT_2B => X"000000800000006e00000093000000c70000007d000000670000005c0000005e",
            INIT_2C => X"00000035000000410000004b0000004d0000006f0000006a0000005500000046",
            INIT_2D => X"0000005d000000710000005f0000005d0000006c000000730000006b00000061",
            INIT_2E => X"000000620000005f00000062000000610000005a0000005500000095000000bb",
            INIT_2F => X"000000b30000009200000070000000cc0000009a0000005f0000005700000055",
            INIT_30 => X"0000003a000000560000005e0000004a00000064000000640000004d00000055",
            INIT_31 => X"00000078000000850000007f0000006c000000690000006e0000006200000057",
            INIT_32 => X"0000005100000051000000570000005f0000005f00000070000000aa000000c3",
            INIT_33 => X"000000d0000000c10000007f000000ad000000b200000050000000550000004f",
            INIT_34 => X"0000004a00000059000000570000004b00000052000000440000004700000050",
            INIT_35 => X"0000005900000067000000760000006f000000650000006a0000006900000062",
            INIT_36 => X"0000006000000062000000620000006d000000720000008e000000b4000000b8",
            INIT_37 => X"000000bf000000c0000000a000000084000000aa000000500000003c00000043",
            INIT_38 => X"0000004d0000004f000000520000004e0000004f000000480000004600000056",
            INIT_39 => X"0000006d00000079000000810000008500000089000000880000008700000083",
            INIT_3A => X"0000009200000094000000920000009600000094000000a3000000b3000000b5",
            INIT_3B => X"000000b9000000b0000000aa000000650000005a00000049000000370000003b",
            INIT_3C => X"000000600000005e0000006a000000680000006d00000083000000840000008a",
            INIT_3D => X"00000090000000980000009b0000009a0000009b0000009b0000009e00000094",
            INIT_3E => X"000000960000009d0000009c00000092000000770000008200000092000000a9",
            INIT_3F => X"000000b1000000a8000000a70000006900000045000000620000005600000048",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY12;


    MEM_IFMAP_LAYER0_ENTITY13 : if BRAM_NAME = "ifmap_layer0_entity13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000006a0000006500000073000000830000008100000087000000900000008f",
            INIT_01 => X"00000092000000960000009a0000009a0000009a000000990000009700000090",
            INIT_02 => X"00000082000000860000008b0000007f0000005e00000075000000920000009f",
            INIT_03 => X"000000a7000000a3000000a20000008400000090000000c00000009a00000069",
            INIT_04 => X"0000005f0000006c000000760000006d0000005f0000005d0000008100000091",
            INIT_05 => X"00000095000000970000009600000090000000860000007e0000007a0000007b",
            INIT_06 => X"0000007a000000850000009b000000940000008300000093000000a20000009c",
            INIT_07 => X"0000009d0000009700000099000000950000009f000000a40000009d00000094",
            INIT_08 => X"00000066000000590000004900000046000000560000006f0000007b0000008c",
            INIT_09 => X"0000008f000000810000007800000075000000780000007e000000850000008d",
            INIT_0A => X"000000960000008e000000990000009f000000970000009d000000a5000000a1",
            INIT_0B => X"00000099000000980000009a0000009000000083000000790000007d00000095",
            INIT_0C => X"000000560000003d000000470000006e000000800000008a000000820000007b",
            INIT_0D => X"000000760000006c00000076000000840000008f000000980000009c00000099",
            INIT_0E => X"0000009500000089000000910000009a000000990000009a000000a0000000a4",
            INIT_0F => X"00000098000000900000007d000000690000005c0000004b0000005600000084",
            INIT_10 => X"00000068000000670000006b0000007200000073000000740000007b00000076",
            INIT_11 => X"00000074000000860000008d000000900000008f0000008d0000008500000075",
            INIT_12 => X"00000062000000590000008200000096000000970000009a0000009800000091",
            INIT_13 => X"00000075000000600000005a0000005000000041000000470000004900000041",
            INIT_14 => X"000000630000006b0000006f0000006f00000072000000770000007d0000007e",
            INIT_15 => X"000000750000007d0000007d0000008100000083000000820000005b0000003d",
            INIT_16 => X"000000390000003800000073000000940000008b00000082000000720000005f",
            INIT_17 => X"0000005600000053000000490000003a0000003c0000004b000000330000001b",
            INIT_18 => X"0000003e0000006800000074000000720000007400000075000000660000005b",
            INIT_19 => X"00000054000000510000004e000000700000008500000082000000600000004c",
            INIT_1A => X"00000053000000560000006b0000006c00000060000000580000005300000051",
            INIT_1B => X"000000460000003d000000330000002d000000340000002e0000001e00000018",
            INIT_1C => X"00000039000000600000006a000000690000006b000000680000004100000035",
            INIT_1D => X"0000003b00000040000000440000006e00000087000000850000007300000062",
            INIT_1E => X"000000580000004f0000004e0000005000000051000000500000004600000037",
            INIT_1F => X"0000002c000000310000002d00000029000000220000001e0000001b00000018",
            INIT_20 => X"000000410000005a00000068000000690000006d0000006d0000004f00000049",
            INIT_21 => X"0000005500000058000000620000006a00000062000000530000004400000041",
            INIT_22 => X"000000460000004a00000051000000520000004800000033000000290000002c",
            INIT_23 => X"0000003d000000370000002700000023000000200000001e0000001b00000019",
            INIT_24 => X"0000004300000057000000690000006700000066000000630000005800000051",
            INIT_25 => X"0000004c000000450000003b000000390000003a0000003f0000004200000046",
            INIT_26 => X"00000048000000440000003e000000360000002e0000002f000000310000002c",
            INIT_27 => X"000000380000002e0000001e0000001c0000001d00000019000000180000001e",
            INIT_28 => X"000000360000003a000000410000003a00000037000000320000002d0000002c",
            INIT_29 => X"0000002e00000033000000370000003a0000003e000000400000003e0000003a",
            INIT_2A => X"0000003300000026000000250000003000000031000000300000002a00000026",
            INIT_2B => X"00000029000000200000001b0000001c0000001b000000190000001c0000001f",
            INIT_2C => X"0000001e0000001d0000001a0000001b0000001f000000200000002100000027",
            INIT_2D => X"000000310000003400000035000000330000002e000000280000002600000028",
            INIT_2E => X"000000260000002c000000420000003700000029000000250000002400000025",
            INIT_2F => X"0000001f0000001b0000001a0000001b0000001c0000001e0000002100000017",
            INIT_30 => X"000000210000001f0000001b0000001c0000001c0000001e0000001f00000020",
            INIT_31 => X"00000023000000210000001e0000001e0000002200000027000000290000002d",
            INIT_32 => X"0000002a0000003400000049000000310000001e000000230000002600000020",
            INIT_33 => X"0000001b0000001a0000001b0000001d0000001e000000260000001a0000000d",
            INIT_34 => X"0000001f0000001e0000001a0000001a00000019000000190000001a0000001b",
            INIT_35 => X"0000001d0000002000000025000000280000002a00000029000000280000002a",
            INIT_36 => X"000000270000002e00000040000000260000001c000000240000001e0000001d",
            INIT_37 => X"0000001a000000190000001b0000001c00000021000000250000000900000004",
            INIT_38 => X"000000170000001b000000190000001c0000001e000000200000002200000025",
            INIT_39 => X"0000002700000027000000280000002700000026000000230000001e00000021",
            INIT_3A => X"0000001c0000002400000039000000240000001e0000001d0000001d0000001d",
            INIT_3B => X"0000001800000018000000170000001b00000024000000130000000400000005",
            INIT_3C => X"0000001c0000001e000000200000002200000021000000220000002300000025",
            INIT_3D => X"000000260000002600000024000000220000001e000000180000000f0000000c",
            INIT_3E => X"00000008000000130000002d00000020000000190000001b0000001b0000001c",
            INIT_3F => X"0000001800000015000000140000002200000019000000050000000400000007",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY13;


    MEM_IFMAP_LAYER0_ENTITY14 : if BRAM_NAME = "ifmap_layer0_entity14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000be000000bb000000a60000009e000000c1000000d0000000d3000000d8",
            INIT_01 => X"000000db000000dd000000de000000da000000e5000000e8000000eb000000ed",
            INIT_02 => X"000000dc000000e9000000ee000000ef000000f1000000ef000000f1000000f1",
            INIT_03 => X"000000f2000000e7000000eb000000f3000000ed000000e7000000ef000000f1",
            INIT_04 => X"000000c8000000c7000000b0000000a0000000c7000000d9000000da000000da",
            INIT_05 => X"000000df000000e5000000e5000000db000000e9000000ee000000ef000000f3",
            INIT_06 => X"000000e1000000ea000000ee000000f5000000f7000000ed000000ef000000f5",
            INIT_07 => X"000000f5000000e9000000ef000000f8000000ec000000e8000000f6000000f7",
            INIT_08 => X"000000c9000000c8000000b3000000a2000000c9000000dc000000df000000d6",
            INIT_09 => X"000000dd000000e9000000e2000000db000000e5000000ea000000ea000000f4",
            INIT_0A => X"000000e2000000e9000000ee000000f3000000eb000000d6000000ea000000f1",
            INIT_0B => X"000000f7000000e9000000f0000000fa000000ee000000e5000000f9000000f4",
            INIT_0C => X"000000cb000000c7000000b3000000a4000000c9000000d9000000e1000000d9",
            INIT_0D => X"000000df000000eb000000e3000000d9000000dd000000e8000000e2000000f4",
            INIT_0E => X"000000e4000000e7000000ed000000eb000000b8000000af000000e4000000f1",
            INIT_0F => X"000000f8000000e8000000ee000000fa000000ed000000e3000000f7000000f2",
            INIT_10 => X"000000cf000000cc000000b5000000a1000000c9000000d6000000e1000000d5",
            INIT_11 => X"000000d7000000ed000000e2000000d7000000d9000000e5000000d4000000ec",
            INIT_12 => X"000000e3000000e1000000ec000000e1000000aa000000ae000000e0000000ec",
            INIT_13 => X"000000f7000000e7000000eb000000f6000000e7000000e7000000f5000000ef",
            INIT_14 => X"000000d0000000cd000000b70000009a000000c9000000d4000000e2000000d7",
            INIT_15 => X"000000da000000ee000000df000000d7000000d7000000e5000000c7000000cd",
            INIT_16 => X"000000d1000000d0000000ef000000cc0000007c000000a7000000e3000000e9",
            INIT_17 => X"000000f6000000e5000000e1000000ef000000e2000000e6000000f1000000e8",
            INIT_18 => X"000000cc000000c7000000b30000008b000000c2000000cb000000dd000000d5",
            INIT_19 => X"000000db000000e9000000d8000000d4000000d8000000e6000000bc000000b0",
            INIT_1A => X"000000be000000c0000000d4000000c00000008100000097000000b7000000be",
            INIT_1B => X"000000e0000000e0000000d6000000e5000000db000000de000000eb000000e0",
            INIT_1C => X"000000cd000000c6000000af0000008a000000c0000000cb000000ce000000cc",
            INIT_1D => X"000000d4000000df000000d0000000d2000000d5000000d8000000c7000000ce",
            INIT_1E => X"000000b200000095000000710000005d00000055000000500000005000000045",
            INIT_1F => X"0000006c000000b7000000ce000000de000000d0000000c5000000dd000000d4",
            INIT_20 => X"000000ad000000a80000009a00000085000000a5000000ac000000a0000000b3",
            INIT_21 => X"000000be000000c2000000bd000000c3000000c7000000bf000000c1000000c6",
            INIT_22 => X"00000098000000790000006b0000006c00000068000000680000006e0000004f",
            INIT_23 => X"000000520000007a0000009f000000af000000a300000095000000be000000af",
            INIT_24 => X"000000730000007400000072000000690000006d0000006e000000700000007f",
            INIT_25 => X"00000087000000880000008c00000093000000970000008f0000009e000000a1",
            INIT_26 => X"000000860000007700000078000000780000006c0000006c000000660000005c",
            INIT_27 => X"0000008f0000008000000097000000910000006e0000006a0000008200000078",
            INIT_28 => X"0000004e00000057000000560000005200000063000000690000006100000064",
            INIT_29 => X"000000650000006d0000006a0000006f0000007200000076000000840000007f",
            INIT_2A => X"0000006d0000006d0000006e0000006b00000060000000570000006c00000077",
            INIT_2B => X"000000840000006f00000090000000bf000000780000006f0000006600000068",
            INIT_2C => X"0000004a000000550000005f00000062000000800000007a0000006200000051",
            INIT_2D => X"00000068000000810000007100000073000000840000008b000000860000007b",
            INIT_2E => X"0000007800000073000000740000007700000071000000680000009e000000bd",
            INIT_2F => X"000000b7000000940000006d000000c500000095000000670000006300000063",
            INIT_30 => X"000000510000006b000000710000005d00000075000000730000005d00000066",
            INIT_31 => X"0000008900000098000000950000008300000082000000880000007d00000071",
            INIT_32 => X"0000006c0000006c000000720000007b000000760000007f000000af000000c2",
            INIT_33 => X"000000ce000000bd00000076000000a2000000a7000000500000006200000065",
            INIT_34 => X"000000610000006e0000006a0000005d00000062000000540000005900000064",
            INIT_35 => X"0000006e0000007b0000008a000000860000007e00000083000000820000007c",
            INIT_36 => X"0000007b0000007f0000007e000000870000008600000099000000b5000000b4",
            INIT_37 => X"000000b8000000b7000000970000007a000000a00000004d0000004800000059",
            INIT_38 => X"000000660000006500000066000000610000005f00000058000000580000006b",
            INIT_39 => X"000000820000008e000000970000009e000000a3000000a4000000a10000009d",
            INIT_3A => X"000000ab000000ad000000aa000000a9000000a2000000a9000000b1000000ae",
            INIT_3B => X"000000b0000000a8000000a40000006200000057000000460000003f0000004b",
            INIT_3C => X"0000007b000000760000007f0000007c0000007e0000009400000098000000a0",
            INIT_3D => X"000000a7000000af000000b3000000b4000000b7000000b8000000b9000000ae",
            INIT_3E => X"000000ad000000b2000000af000000a000000080000000850000008e000000a1",
            INIT_3F => X"000000a9000000a2000000a60000006c000000460000005f0000005900000052",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY14;


    MEM_IFMAP_LAYER0_ENTITY15 : if BRAM_NAME = "ifmap_layer0_entity15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000850000007d0000008a00000098000000940000009a000000a6000000a7",
            INIT_01 => X"000000aa000000ae000000b3000000b6000000b9000000b9000000b5000000ab",
            INIT_02 => X"00000098000000980000009a0000008b0000006600000078000000900000009b",
            INIT_03 => X"000000a5000000a2000000a30000008800000091000000bb000000990000006c",
            INIT_04 => X"0000007c000000850000008d00000083000000740000007200000098000000aa",
            INIT_05 => X"000000af000000af000000b0000000ad000000a7000000a00000009a00000097",
            INIT_06 => X"0000009000000096000000a8000000a00000008c00000098000000a50000009e",
            INIT_07 => X"000000a30000009b0000009c000000970000009e0000009e0000009800000093",
            INIT_08 => X"0000008100000071000000600000005d0000006e0000008700000094000000a4",
            INIT_09 => X"000000a90000009f000000960000009200000094000000990000009f000000a5",
            INIT_0A => X"000000aa000000a0000000a8000000ac000000a1000000a4000000a8000000a4",
            INIT_0B => X"000000a00000009e0000009e0000009200000084000000790000007d00000096",
            INIT_0C => X"000000700000005500000060000000870000009b000000a50000009c00000093",
            INIT_0D => X"0000008e0000008d00000097000000a0000000a7000000ad000000ae000000ab",
            INIT_0E => X"000000a70000009b000000a2000000a8000000a3000000a1000000a3000000a6",
            INIT_0F => X"0000009e00000097000000820000006f00000062000000520000005c0000008a",
            INIT_10 => X"0000008500000084000000870000008f0000008f0000008f000000960000008e",
            INIT_11 => X"0000008a000000a1000000a9000000ab000000a9000000a50000009700000086",
            INIT_12 => X"000000740000006b00000094000000a4000000a3000000a30000009f00000098",
            INIT_13 => X"000000800000006c000000660000005b0000004b0000004e0000005000000048",
            INIT_14 => X"000000840000008c000000900000008f00000090000000930000009700000096",
            INIT_15 => X"0000008b00000092000000940000009a0000009f0000009c0000006e0000004e",
            INIT_16 => X"0000004b0000004a00000084000000a3000000990000008f0000007e0000006d",
            INIT_17 => X"00000067000000640000005a0000004c0000004b000000520000003900000021",
            INIT_18 => X"0000005e00000089000000940000009200000092000000910000008100000073",
            INIT_19 => X"0000006a0000006600000063000000870000009d0000009a000000720000005d",
            INIT_1A => X"00000065000000680000007d0000007c000000710000006a0000006600000065",
            INIT_1B => X"000000580000004f000000450000003f0000004300000035000000250000001f",
            INIT_1C => X"000000560000007d000000860000008600000089000000850000005c0000004d",
            INIT_1D => X"00000052000000590000005c0000008300000099000000960000008400000073",
            INIT_1E => X"0000006a00000061000000600000006100000063000000650000005f0000004f",
            INIT_1F => X"0000003c000000400000003c000000390000002f00000026000000220000001f",
            INIT_20 => X"0000005a000000740000008100000083000000890000008a0000006a00000061",
            INIT_21 => X"0000006c000000740000007c0000007e000000710000005f0000005400000053",
            INIT_22 => X"000000590000005c00000062000000640000005c0000004a0000004300000045",
            INIT_23 => X"0000004a00000042000000330000002e0000002b000000260000002300000020",
            INIT_24 => X"0000005c00000070000000820000007f0000007c000000780000006e00000066",
            INIT_25 => X"000000610000005a000000500000004c0000004b00000050000000540000005b",
            INIT_26 => X"0000005f0000005900000051000000490000004100000041000000430000003d",
            INIT_27 => X"000000450000003a0000002a000000280000002a000000280000002300000025",
            INIT_28 => X"0000004c0000004f000000560000004e0000004a00000045000000400000003f",
            INIT_29 => X"00000041000000460000004a0000004d00000051000000520000005100000050",
            INIT_2A => X"000000490000003b0000003700000044000000430000003f0000003600000032",
            INIT_2B => X"000000360000002d000000280000002800000029000000280000002700000025",
            INIT_2C => X"0000002d0000002b000000280000002a0000003100000034000000350000003a",
            INIT_2D => X"00000044000000470000004800000046000000410000003b0000003a0000003b",
            INIT_2E => X"000000380000003f000000550000004900000039000000330000002f0000002f",
            INIT_2F => X"0000002c000000280000002700000028000000290000002a0000002a0000001d",
            INIT_30 => X"0000002b0000002800000024000000260000002c000000300000003100000032",
            INIT_31 => X"00000035000000340000003100000031000000350000003b0000003e0000003d",
            INIT_32 => X"00000037000000450000005e000000420000002c0000002e0000002f00000028",
            INIT_33 => X"0000002700000027000000280000002a000000290000002e0000002000000012",
            INIT_34 => X"000000280000002700000023000000240000002700000029000000290000002b",
            INIT_35 => X"0000002e00000033000000380000003a0000003d0000003d0000003c00000037",
            INIT_36 => X"0000002e0000003c0000005500000036000000280000002e0000002500000024",
            INIT_37 => X"0000002600000026000000280000002a0000002b000000280000000d00000007",
            INIT_38 => X"000000220000002600000024000000280000002c0000002f0000003100000033",
            INIT_39 => X"00000036000000390000003b000000390000003900000037000000330000002b",
            INIT_3A => X"0000001f000000300000004e0000003200000029000000250000002300000023",
            INIT_3B => X"000000250000002500000024000000290000002d000000140000000600000007",
            INIT_3C => X"000000290000002b0000002d0000002f00000030000000300000003000000031",
            INIT_3D => X"0000003200000033000000310000002d00000028000000220000001a00000011",
            INIT_3E => X"000000080000001b0000003f0000002c00000021000000220000002200000023",
            INIT_3F => X"0000002300000022000000220000002c0000001f000000060000000500000008",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY15;


    MEM_IFMAP_LAYER0_ENTITY16 : if BRAM_NAME = "ifmap_layer0_entity16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000de000000da000000c2000000ba000000de000000ec000000ee000000f1",
            INIT_01 => X"000000f3000000f5000000f4000000eb000000f0000000f1000000f2000000f5",
            INIT_02 => X"000000e3000000f0000000f5000000f8000000f9000000f3000000f3000000f3",
            INIT_03 => X"000000f5000000eb000000ef000000f7000000f1000000ea000000f3000000f6",
            INIT_04 => X"000000e5000000e2000000c9000000b8000000df000000f0000000f0000000ee",
            INIT_05 => X"000000f3000000f7000000f5000000e8000000f3000000f5000000f5000000f8",
            INIT_06 => X"000000e6000000ef000000f3000000fb000000fb000000ee000000ee000000f4",
            INIT_07 => X"000000f8000000ec000000f3000000fc000000f0000000ec000000fa000000fb",
            INIT_08 => X"000000e1000000de000000c7000000b5000000db000000ee000000ef000000e4",
            INIT_09 => X"000000eb000000f4000000ec000000e4000000eb000000ef000000ee000000f7",
            INIT_0A => X"000000e5000000ec000000f1000000f6000000ec000000d7000000e8000000ef",
            INIT_0B => X"000000f8000000eb000000f2000000fc000000f1000000e8000000fb000000f7",
            INIT_0C => X"000000de000000d8000000c2000000b3000000d6000000e4000000eb000000e1",
            INIT_0D => X"000000e5000000ef000000e6000000dd000000e1000000ec000000e6000000f7",
            INIT_0E => X"000000e6000000ea000000f0000000ee000000ba000000b0000000e5000000f1",
            INIT_0F => X"000000f8000000e9000000ef000000fb000000ee000000e4000000f8000000f3",
            INIT_10 => X"000000df000000d9000000c1000000ac000000d2000000dd000000e7000000d9",
            INIT_11 => X"000000da000000eb000000e1000000d7000000db000000e8000000d6000000ee",
            INIT_12 => X"000000e5000000e3000000ee000000e4000000b0000000b2000000e5000000ef",
            INIT_13 => X"000000f7000000e7000000ea000000f5000000e7000000e8000000f6000000f0",
            INIT_14 => X"000000dc000000d5000000bf000000a4000000ce000000d5000000e1000000d5",
            INIT_15 => X"000000d6000000e6000000da000000d6000000d6000000e3000000c8000000ce",
            INIT_16 => X"000000d0000000ce000000ed000000cf00000082000000ad000000e6000000e9",
            INIT_17 => X"000000f4000000e1000000db000000e8000000dd000000e7000000f2000000e6",
            INIT_18 => X"000000d4000000ca000000b900000096000000c4000000c9000000d9000000d0",
            INIT_19 => X"000000d3000000db000000d0000000d3000000d4000000dd000000b9000000af",
            INIT_1A => X"000000bb000000bd000000d2000000c5000000890000009d000000b8000000bb",
            INIT_1B => X"000000dd000000dc000000ce000000da000000d1000000db000000e7000000d8",
            INIT_1C => X"000000d3000000c9000000b300000093000000c5000000cc000000ce000000cb",
            INIT_1D => X"000000d0000000d2000000c6000000cd000000ce000000ce000000c0000000cb",
            INIT_1E => X"000000b30000009b0000007a0000006a000000640000005e0000005800000049",
            INIT_1F => X"0000006f000000b7000000ca000000d7000000c6000000b9000000ce000000c1",
            INIT_20 => X"000000b3000000ad000000a00000008c000000aa000000af000000a1000000b3",
            INIT_21 => X"000000bb000000b8000000b4000000bd000000c3000000b9000000ba000000c4",
            INIT_22 => X"0000009f0000008900000080000000800000007e0000007e000000800000005a",
            INIT_23 => X"000000580000007c0000009e000000ac0000009c00000089000000b00000009f",
            INIT_24 => X"0000007b0000007e0000007b0000007000000072000000720000007200000080",
            INIT_25 => X"000000860000008600000089000000900000009800000092000000a0000000a7",
            INIT_26 => X"000000930000008b000000900000008c00000082000000830000007800000068",
            INIT_27 => X"0000009500000083000000960000008d0000006a000000690000008000000075",
            INIT_28 => X"000000590000006600000062000000580000006b00000073000000680000006a",
            INIT_29 => X"0000006b0000007600000071000000730000007b000000860000009700000092",
            INIT_2A => X"000000800000007f0000007f000000780000006f000000680000007a00000080",
            INIT_2B => X"000000860000006e0000008b000000b600000072000000750000006d00000070",
            INIT_2C => X"00000058000000680000006e0000006a0000008e00000089000000710000005e",
            INIT_2D => X"00000074000000920000007f0000007d00000094000000a5000000a500000097",
            INIT_2E => X"0000008e000000820000007f0000007f0000007b00000072000000a5000000bf",
            INIT_2F => X"000000b40000008e00000064000000b80000008c0000006d0000006c0000006c",
            INIT_30 => X"0000006400000082000000840000006800000081000000820000006d00000076",
            INIT_31 => X"0000009a000000ab000000a8000000970000009b000000a50000009a0000008b",
            INIT_32 => X"000000820000007d000000810000008c0000008600000089000000b3000000c1",
            INIT_33 => X"000000cb000000b90000007000000098000000a000000054000000690000006d",
            INIT_34 => X"00000078000000860000007e0000006a00000071000000650000006c00000079",
            INIT_35 => X"0000008300000091000000a10000009f00000099000000a10000009e00000095",
            INIT_36 => X"0000009200000093000000910000009b00000096000000a1000000b6000000b1",
            INIT_37 => X"000000b5000000b500000094000000760000009d000000500000004e00000060",
            INIT_38 => X"0000007f000000800000007d0000007200000074000000710000007300000086",
            INIT_39 => X"0000009f000000a8000000b0000000b8000000be000000bf000000be000000b9",
            INIT_3A => X"000000c5000000c4000000be000000b8000000ac000000ad000000af000000a8",
            INIT_3B => X"000000ab000000a5000000a30000006300000057000000470000004300000051",
            INIT_3C => X"00000097000000950000009a0000009100000099000000b3000000b8000000c1",
            INIT_3D => X"000000c9000000cd000000cf000000d0000000d1000000d2000000d4000000c8",
            INIT_3E => X"000000c6000000c9000000c3000000ab00000086000000870000008b0000009b",
            INIT_3F => X"000000a5000000a1000000a800000071000000490000005c0000005a00000056",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY16;


    MEM_IFMAP_LAYER0_ENTITY17 : if BRAM_NAME = "ifmap_layer0_entity17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a50000009f000000a7000000b0000000af000000b9000000c6000000c9",
            INIT_01 => X"000000cd000000d0000000d2000000d2000000d2000000d0000000c9000000be",
            INIT_02 => X"000000aa000000aa000000a9000000940000006c0000007a0000008e00000099",
            INIT_03 => X"000000a7000000a5000000a70000008e00000093000000b5000000980000006f",
            INIT_04 => X"0000009d000000aa000000ae0000009d0000008d0000008f000000b6000000ca",
            INIT_05 => X"000000d0000000d3000000d1000000ca000000bf000000b5000000a7000000a2",
            INIT_06 => X"0000009b000000a0000000b2000000a9000000930000009d000000a7000000a0",
            INIT_07 => X"000000a9000000a2000000a10000009c0000009e000000960000009600000094",
            INIT_08 => X"000000a20000009400000080000000790000008a000000a4000000b1000000c2",
            INIT_09 => X"000000c7000000bc000000b2000000ab000000aa000000ac000000ac000000b0",
            INIT_0A => X"000000b4000000a8000000b0000000b5000000aa000000ad000000af000000ac",
            INIT_0B => X"000000a8000000a5000000a30000009600000085000000760000007d00000099",
            INIT_0C => X"0000008f000000750000007f000000a6000000bc000000c5000000ba000000b0",
            INIT_0D => X"000000a9000000a3000000ab000000b2000000b9000000be000000bf000000ba",
            INIT_0E => X"000000b4000000a5000000ac000000b1000000ad000000ac000000af000000b2",
            INIT_0F => X"000000a40000009c000000880000007400000067000000570000006200000090",
            INIT_10 => X"000000a6000000a5000000a8000000b0000000b0000000ae000000b3000000aa",
            INIT_11 => X"000000a4000000b8000000be000000bd000000b9000000b5000000a800000096",
            INIT_12 => X"00000081000000760000009d000000ad000000ad000000ad000000ab000000a2",
            INIT_13 => X"00000085000000700000006a0000005f0000005000000054000000560000004e",
            INIT_14 => X"000000a5000000ac000000b1000000af000000ae000000b0000000b3000000b0",
            INIT_15 => X"000000a4000000ab000000ab000000ad000000af000000ab0000007e0000005e",
            INIT_16 => X"00000058000000550000008e000000ac000000a2000000980000008800000075",
            INIT_17 => X"0000006c000000680000005e000000500000004f000000580000003f00000027",
            INIT_18 => X"0000007c000000a6000000b2000000af000000af000000ad0000009a0000008b",
            INIT_19 => X"000000820000007e0000007a0000009a000000ae000000a9000000830000006c",
            INIT_1A => X"0000007200000072000000860000008500000079000000710000006d0000006c",
            INIT_1B => X"0000005f000000560000004b00000045000000490000003b0000002b00000026",
            INIT_1C => X"0000006f00000096000000a00000009f000000a30000009e0000007400000064",
            INIT_1D => X"00000068000000700000007300000097000000ac000000a80000009500000083",
            INIT_1E => X"000000770000006b0000006a0000006a0000006a0000006c0000006400000054",
            INIT_1F => X"00000045000000490000004400000041000000370000002c0000002800000025",
            INIT_20 => X"000000710000008a000000970000009a000000a1000000a20000008000000077",
            INIT_21 => X"0000008100000088000000900000009200000084000000720000006500000062",
            INIT_22 => X"00000065000000670000006d0000006c0000006300000050000000480000004b",
            INIT_23 => X"000000550000004d0000003d0000003a000000340000002d0000002900000027",
            INIT_24 => X"00000074000000880000009a00000097000000940000008f000000840000007c",
            INIT_25 => X"00000076000000670000005b00000057000000560000005b0000006300000065",
            INIT_26 => X"00000065000000630000005e0000005200000048000000480000004a00000045",
            INIT_27 => X"0000004e00000044000000340000003200000033000000300000002f00000030",
            INIT_28 => X"00000060000000640000006a000000630000005c000000560000005200000051",
            INIT_29 => X"000000520000004f0000005100000054000000570000005b0000005e00000058",
            INIT_2A => X"0000004d00000044000000440000004c0000004a00000048000000400000003b",
            INIT_2B => X"0000003f00000036000000310000003200000031000000300000003400000030",
            INIT_2C => X"0000003b0000003900000036000000370000003c0000003d0000003e00000044",
            INIT_2D => X"0000004e0000004f0000004f0000004d00000048000000440000004500000042",
            INIT_2E => X"0000003d000000470000006100000052000000410000003c0000003800000039",
            INIT_2F => X"0000003500000031000000300000003100000032000000320000003200000023",
            INIT_30 => X"00000032000000300000002c0000002d00000031000000350000003500000037",
            INIT_31 => X"0000003a0000003b00000038000000380000003c000000420000004700000044",
            INIT_32 => X"0000003b0000004b000000680000004b00000035000000380000003a00000033",
            INIT_33 => X"0000003100000030000000310000003300000032000000350000002500000014",
            INIT_34 => X"0000002d0000002c00000028000000290000002c0000002e0000002e00000030",
            INIT_35 => X"00000033000000390000003f000000410000004400000044000000440000003d",
            INIT_36 => X"00000032000000420000005d0000003f0000003100000038000000300000002f",
            INIT_37 => X"0000002f0000002f0000003100000033000000340000002e0000000e00000005",
            INIT_38 => X"000000270000002b000000290000002d0000003200000036000000380000003b",
            INIT_39 => X"0000003e000000400000004200000040000000400000003d0000003a00000031",
            INIT_3A => X"0000002400000035000000550000003b00000032000000300000002f0000002f",
            INIT_3B => X"0000002e0000002e0000002d0000003200000036000000180000000300000003",
            INIT_3C => X"0000002f0000003200000034000000360000003800000038000000380000003a",
            INIT_3D => X"0000003a0000003700000035000000320000002d000000270000001e00000014",
            INIT_3E => X"0000000b0000002100000048000000360000002c0000002d0000002d0000002e",
            INIT_3F => X"0000002c0000002c0000002b0000003400000025000000080000000300000007",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY17;


    MEM_IFMAP_LAYER0_ENTITY18 : if BRAM_NAME = "ifmap_layer0_entity18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009b000000a7000000b0000000be000000b1000000a6000000a8000000a6",
            INIT_01 => X"000000aa000000b3000000bb000000bb000000bb000000bb000000b8000000b8",
            INIT_02 => X"000000b6000000b4000000b8000000ba000000bb000000bb000000bc000000bd",
            INIT_03 => X"000000bb000000bb000000bc000000c3000000c9000000c9000000ca000000c0",
            INIT_04 => X"00000099000000a3000000ab000000bb000000b30000009b0000009a0000009f",
            INIT_05 => X"0000009f000000a5000000ab000000af000000a9000000ab000000a2000000a5",
            INIT_06 => X"000000aa000000a4000000a6000000a5000000a7000000ad000000a9000000a8",
            INIT_07 => X"000000a9000000ad000000be000000ca000000cc000000ca000000cb000000bd",
            INIT_08 => X"0000009b000000a0000000a8000000b8000000bb000000ae000000b0000000bc",
            INIT_09 => X"000000b6000000b3000000b1000000be000000c0000000c2000000bc000000b9",
            INIT_0A => X"000000c1000000c2000000c1000000c2000000c3000000c5000000c1000000bf",
            INIT_0B => X"000000bf000000c5000000ce000000cf000000d0000000ce000000cc000000bd",
            INIT_0C => X"000000970000009d000000a6000000b1000000b4000000b9000000c7000000c5",
            INIT_0D => X"000000b6000000cc000000cd000000c6000000d2000000c5000000c4000000cb",
            INIT_0E => X"000000cd000000cf000000d2000000cb000000cf000000d2000000c5000000cc",
            INIT_0F => X"000000d0000000c6000000cc000000c9000000d1000000cf000000ce000000c0",
            INIT_10 => X"000000970000009e000000a8000000ae000000b1000000b5000000bf000000c4",
            INIT_11 => X"000000b7000000c2000000bd000000b9000000c4000000b9000000b9000000ca",
            INIT_12 => X"000000c7000000c7000000c8000000c0000000c3000000c7000000be000000bc",
            INIT_13 => X"000000c9000000c7000000c9000000c4000000ce000000cc000000cf000000c4",
            INIT_14 => X"000000940000009c000000a7000000ae000000ab000000ae000000c4000000c3",
            INIT_15 => X"000000c0000000be000000bd000000b8000000bb000000bd000000bd000000bf",
            INIT_16 => X"000000be000000c3000000bb000000c6000000c0000000bc000000c0000000c1",
            INIT_17 => X"000000cd000000ce000000cb000000d1000000d4000000d0000000d1000000c4",
            INIT_18 => X"0000009400000099000000a5000000ae000000a8000000b0000000cb000000c3",
            INIT_19 => X"000000bc000000bc000000bb000000be000000b6000000c2000000c5000000c3",
            INIT_1A => X"000000c4000000c1000000c8000000cd000000c6000000c5000000c5000000c9",
            INIT_1B => X"000000c5000000c8000000c6000000c3000000c5000000cb000000cf000000c3",
            INIT_1C => X"000000990000009b000000a3000000ac000000ac000000bc000000c7000000d1",
            INIT_1D => X"000000c4000000be000000bd000000bf000000c1000000bc000000bb000000c4",
            INIT_1E => X"000000ca000000c2000000c4000000ce000000c2000000c9000000c4000000c8",
            INIT_1F => X"000000b5000000bb000000c8000000c9000000c8000000c4000000c7000000bd",
            INIT_20 => X"000000a00000009f000000a3000000ac000000ae000000b0000000b0000000be",
            INIT_21 => X"000000b4000000af000000b0000000b0000000b5000000aa000000ac000000b6",
            INIT_22 => X"000000bb000000b2000000b5000000bb000000b1000000bc000000b4000000bb",
            INIT_23 => X"000000c7000000c4000000bc000000bc000000c5000000c0000000c2000000b8",
            INIT_24 => X"000000ab000000a7000000a2000000ac000000aa000000ab000000b4000000b0",
            INIT_25 => X"0000009b0000009c000000960000009c0000009600000092000000990000009e",
            INIT_26 => X"000000a6000000a6000000a40000009d0000009d000000a20000009c000000a6",
            INIT_27 => X"000000c8000000c7000000bc000000bd000000c5000000c1000000c2000000b6",
            INIT_28 => X"000000af000000b4000000a8000000b0000000ad000000b1000000b6000000ae",
            INIT_29 => X"0000009c000000a00000009f0000009a0000009f000000a3000000a8000000ad",
            INIT_2A => X"000000aa000000a4000000a0000000a2000000a0000000a8000000a7000000ac",
            INIT_2B => X"000000c2000000c3000000c4000000c4000000c5000000bf000000c1000000b7",
            INIT_2C => X"000000b5000000bb000000b2000000bb000000b7000000aa000000ae000000b6",
            INIT_2D => X"000000b3000000b3000000b4000000b5000000b8000000bb000000c1000000c1",
            INIT_2E => X"000000c1000000c0000000bc000000b9000000b8000000ba000000c0000000c0",
            INIT_2F => X"000000bb000000bc000000c0000000bd000000be000000bf000000c4000000ba",
            INIT_30 => X"000000b9000000be000000ba000000ab000000990000008400000095000000c1",
            INIT_31 => X"000000c6000000bf000000ba000000bc000000bf000000c1000000c3000000c4",
            INIT_32 => X"000000c3000000c0000000be000000bc000000bc000000be000000c0000000bf",
            INIT_33 => X"000000bf000000c1000000c3000000c5000000ca000000ca000000cc000000c1",
            INIT_34 => X"000000ba000000c2000000bc0000009e00000084000000740000005e0000006d",
            INIT_35 => X"00000091000000b1000000c2000000c2000000bf000000c1000000c4000000c7",
            INIT_36 => X"000000c7000000c7000000c8000000c6000000c4000000c4000000c7000000c6",
            INIT_37 => X"000000c5000000c4000000c4000000c4000000c6000000c5000000c6000000b9",
            INIT_38 => X"000000ba000000c5000000c4000000c6000000c2000000b80000008d0000005c",
            INIT_39 => X"00000054000000680000008e000000b3000000c3000000c9000000cc000000cc",
            INIT_3A => X"000000cc000000cc000000cc000000c7000000c2000000c2000000c2000000bf",
            INIT_3B => X"000000bd000000be000000be000000be000000bf000000be000000c0000000b5",
            INIT_3C => X"000000b8000000c7000000c6000000c8000000c5000000c8000000c9000000b1",
            INIT_3D => X"00000075000000540000005d00000080000000ad000000ca000000d0000000cd",
            INIT_3E => X"000000ca000000c8000000c7000000c7000000c3000000c4000000c5000000c3",
            INIT_3F => X"000000c1000000c3000000c2000000bf000000bf000000bd000000be000000b2",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY18;


    MEM_IFMAP_LAYER0_ENTITY19 : if BRAM_NAME = "ifmap_layer0_entity19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b9000000c9000000cb000000d0000000cd000000ce000000d0000000d6",
            INIT_01 => X"000000af0000005c0000004c0000005b000000690000008c000000b5000000cb",
            INIT_02 => X"000000ce000000ca000000c5000000c2000000c1000000c2000000c2000000c2",
            INIT_03 => X"000000c2000000c3000000c1000000bf000000c1000000be000000be000000b4",
            INIT_04 => X"000000bb000000cc000000cf000000d6000000d4000000d4000000d3000000d0",
            INIT_05 => X"000000cb0000007c000000470000005700000054000000540000006300000084",
            INIT_06 => X"000000a7000000be000000cb000000cb000000c3000000c0000000c5000000c4",
            INIT_07 => X"000000c2000000c2000000c0000000bf000000c1000000bf000000c0000000b7",
            INIT_08 => X"000000be000000cf000000cf000000d6000000d4000000d3000000d3000000d0",
            INIT_09 => X"000000d300000089000000480000005700000053000000540000005600000053",
            INIT_0A => X"000000590000006b000000830000009b000000a3000000b6000000cb000000cc",
            INIT_0B => X"000000ca000000c6000000c2000000bf000000c1000000c0000000bf000000b6",
            INIT_0C => X"000000bf000000d2000000d1000000d7000000d5000000d4000000d4000000d5",
            INIT_0D => X"000000cc000000710000002f0000003a0000003f0000004c000000570000005d",
            INIT_0E => X"0000005a00000050000000460000003e0000003a0000004d0000007a0000009f",
            INIT_0F => X"000000b4000000c2000000c9000000c8000000c8000000c4000000c4000000b9",
            INIT_10 => X"000000bf000000d0000000cf000000d3000000d1000000d2000000d1000000d4",
            INIT_11 => X"0000009d00000065000000410000002500000033000000440000004a00000058",
            INIT_12 => X"0000005b000000560000005500000049000000370000002e0000003e00000048",
            INIT_13 => X"0000004e0000006b000000850000009e000000b8000000c3000000c4000000ba",
            INIT_14 => X"000000ba000000ca000000cb000000d1000000cf000000ce000000d1000000c8",
            INIT_15 => X"000000950000008c00000097000000640000002d000000350000003200000060",
            INIT_16 => X"0000009c000000a0000000800000004800000062000000700000005900000042",
            INIT_17 => X"0000004300000083000000a6000000a3000000ad000000b7000000bc000000b2",
            INIT_18 => X"000000b9000000c9000000ca000000d2000000d2000000d0000000d1000000d1",
            INIT_19 => X"000000d2000000d3000000d7000000bd000000900000009200000094000000a8",
            INIT_1A => X"000000ca000000ce000000c00000009a000000a3000000b2000000b10000009f",
            INIT_1B => X"0000009c000000b2000000bf000000c2000000c4000000c1000000bc000000b0",
            INIT_1C => X"000000b0000000bc000000c0000000c4000000c0000000bc000000b9000000b7",
            INIT_1D => X"000000b6000000b2000000b3000000ad000000aa000000aa000000ab000000ad",
            INIT_1E => X"000000a9000000a0000000a1000000a7000000a5000000a1000000a5000000aa",
            INIT_1F => X"000000aa000000a000000098000000960000009d000000a3000000a40000009c",
            INIT_20 => X"00000072000000630000006e0000006b00000066000000610000005e0000005d",
            INIT_21 => X"000000580000005500000058000000500000004d0000004e0000005300000065",
            INIT_22 => X"000000710000006c0000006a0000006b0000006c0000006e0000006f00000071",
            INIT_23 => X"0000007500000077000000780000007700000078000000790000007a0000007c",
            INIT_24 => X"0000007a0000006d000000710000007500000073000000700000007200000071",
            INIT_25 => X"0000006f000000700000006f0000006d0000006e0000006d0000006e0000006c",
            INIT_26 => X"0000007300000070000000690000006b0000006c0000006a0000006500000068",
            INIT_27 => X"0000006a0000006b0000006d0000006d00000067000000660000005e00000065",
            INIT_28 => X"00000078000000610000006b000000700000006d00000068000000620000005e",
            INIT_29 => X"0000005e0000005d0000005800000056000000520000004f000000500000004e",
            INIT_2A => X"000000500000004f000000480000004500000043000000420000004100000041",
            INIT_2B => X"00000040000000410000004200000040000000430000003f000000350000004d",
            INIT_2C => X"0000005b00000037000000410000004500000042000000420000003f0000003d",
            INIT_2D => X"00000042000000400000003c00000039000000390000003c0000003d0000003f",
            INIT_2E => X"0000003f00000042000000400000003a00000038000000390000003b0000003c",
            INIT_2F => X"0000003a00000039000000380000003900000034000000310000004b0000005c",
            INIT_30 => X"0000005d0000003c000000420000004400000043000000430000004000000041",
            INIT_31 => X"00000045000000410000003e0000003b0000003b0000003b0000003c0000003d",
            INIT_32 => X"000000400000003f0000003a0000003800000037000000370000003800000038",
            INIT_33 => X"000000390000003a0000003800000035000000410000005d0000006100000051",
            INIT_34 => X"00000059000000390000003d00000039000000390000003b000000390000003b",
            INIT_35 => X"0000003c0000003a00000038000000360000003c0000003d0000003b0000003d",
            INIT_36 => X"000000410000003d0000003a000000390000003c0000003c0000003d0000003d",
            INIT_37 => X"000000420000003e000000390000004600000061000000590000003b00000043",
            INIT_38 => X"000000590000003c0000003f0000003e0000003e0000003e0000003e0000003f",
            INIT_39 => X"0000003e0000003d000000410000005200000054000000510000004e00000051",
            INIT_3A => X"0000005800000054000000550000005300000050000000430000004200000040",
            INIT_3B => X"000000340000003800000056000000670000004c000000390000003d0000004b",
            INIT_3C => X"0000005c0000003c0000003d0000003c0000003f000000420000004300000041",
            INIT_3D => X"0000004200000043000000410000004800000049000000490000004800000046",
            INIT_3E => X"000000490000004a0000004b0000004b0000004b00000040000000400000003e",
            INIT_3F => X"00000041000000560000005800000040000000390000003c0000004000000049",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY19;


    MEM_IFMAP_LAYER0_ENTITY20 : if BRAM_NAME = "ifmap_layer0_entity20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009c000000b0000000b3000000c0000000b9000000ab000000ad000000ad",
            INIT_01 => X"000000af000000b3000000b6000000b8000000b9000000b8000000b6000000b5",
            INIT_02 => X"000000b3000000b3000000b7000000b9000000ba000000ba000000bb000000bd",
            INIT_03 => X"000000bb000000bb000000bc000000c3000000c5000000c4000000ca000000b7",
            INIT_04 => X"0000009b000000b3000000b8000000c3000000be000000a20000009f000000a4",
            INIT_05 => X"000000a3000000a5000000a9000000b0000000ab000000ae000000a4000000a7",
            INIT_06 => X"000000ac000000a6000000a8000000a6000000a9000000af000000ab000000a9",
            INIT_07 => X"000000aa000000ae000000bf000000cc000000ce000000d0000000d7000000be",
            INIT_08 => X"0000009a000000b2000000b9000000c4000000cb000000c1000000b2000000a8",
            INIT_09 => X"000000a0000000af000000be000000c4000000c3000000c5000000be000000bc",
            INIT_0A => X"000000c4000000c3000000c2000000c3000000c4000000c6000000c1000000bf",
            INIT_0B => X"000000c0000000c4000000cd000000cd000000ce000000d0000000d7000000bf",
            INIT_0C => X"0000009a000000b2000000bc000000c3000000ca000000c5000000bc00000080",
            INIT_0D => X"0000006c000000980000009a0000009b0000009e000000950000009500000094",
            INIT_0E => X"000000a7000000a1000000a3000000ad000000a8000000a3000000ae0000009f",
            INIT_0F => X"000000bc000000d0000000cc000000ce000000cc000000cd000000d4000000bc",
            INIT_10 => X"0000009a000000b1000000bb000000bf000000c6000000c4000000bd0000007e",
            INIT_11 => X"000000800000008b0000006a0000006b00000073000000780000007600000071",
            INIT_12 => X"0000007700000072000000720000007e00000076000000700000008800000070",
            INIT_13 => X"000000a0000000cb000000c9000000ce000000ce000000cd000000d6000000be",
            INIT_14 => X"00000097000000ae000000bb000000bd000000c5000000c8000000b700000093",
            INIT_15 => X"000000a9000000a800000091000000a5000000aa00000092000000950000009d",
            INIT_16 => X"000000b4000000b2000000b0000000bd000000b0000000b3000000bc000000b1",
            INIT_17 => X"000000c4000000d0000000cf000000d0000000d0000000d1000000d8000000be",
            INIT_18 => X"00000098000000ac000000b9000000bd000000c2000000c60000009300000060",
            INIT_19 => X"000000950000009700000090000000980000009800000079000000800000008b",
            INIT_1A => X"0000009c00000097000000aa000000a200000096000000ad00000096000000a4",
            INIT_1B => X"0000009c000000a6000000cc000000d2000000d3000000cf000000d4000000bc",
            INIT_1C => X"0000009b000000ac000000b6000000bb000000c2000000b50000007700000065",
            INIT_1D => X"0000007b0000008300000083000000780000009200000087000000870000007f",
            INIT_1E => X"0000007b0000007b000000830000007b0000006d000000840000007b0000009f",
            INIT_1F => X"0000007b00000084000000bf000000c7000000c9000000c9000000d0000000ba",
            INIT_20 => X"000000a1000000af000000b4000000b9000000c0000000ba000000ab000000af",
            INIT_21 => X"000000a2000000a5000000ac000000a6000000af000000ac000000ad000000aa",
            INIT_22 => X"000000ac000000b2000000b2000000af000000a3000000ac000000b2000000be",
            INIT_23 => X"000000ac000000b0000000c8000000cd000000c8000000c9000000d1000000b9",
            INIT_24 => X"000000ac000000b7000000b4000000ba000000be000000c0000000c2000000b7",
            INIT_25 => X"000000a0000000a5000000a2000000a30000009f0000009e000000a4000000a2",
            INIT_26 => X"000000a7000000ae000000ac000000a2000000a0000000a3000000a5000000b6",
            INIT_27 => X"000000c8000000c6000000ca000000cd000000ca000000ca000000d0000000b8",
            INIT_28 => X"000000b1000000c4000000ba000000be000000c0000000c1000000c1000000b7",
            INIT_29 => X"000000a3000000a7000000a50000009f000000a4000000a6000000aa000000ac",
            INIT_2A => X"000000a8000000a6000000a6000000ab000000a8000000ad000000ab000000b2",
            INIT_2B => X"000000c7000000c6000000c7000000c7000000c8000000c8000000d0000000b8",
            INIT_2C => X"000000b7000000cc000000c3000000c8000000c9000000bb000000be000000c6",
            INIT_2D => X"000000c2000000c1000000c1000000c1000000c1000000c2000000c6000000c6",
            INIT_2E => X"000000c6000000c3000000c3000000c6000000c5000000c4000000c4000000c5",
            INIT_2F => X"000000c9000000cb000000c9000000c9000000ca000000c8000000d1000000bb",
            INIT_30 => X"000000b9000000cd000000c6000000b2000000a60000008d0000009a000000c4",
            INIT_31 => X"000000ca000000ca000000c7000000c5000000c5000000c7000000c9000000ca",
            INIT_32 => X"000000c9000000c7000000c6000000c4000000c4000000c6000000c7000000c6",
            INIT_33 => X"000000c7000000ca000000cb000000ce000000cf000000ce000000d4000000bd",
            INIT_34 => X"000000ba000000d0000000c8000000a5000000900000007c0000005f0000006b",
            INIT_35 => X"0000008f000000b3000000c7000000c7000000c5000000c6000000c9000000cc",
            INIT_36 => X"000000cc000000cd000000ce000000cc000000c9000000c9000000cd000000cd",
            INIT_37 => X"000000cc000000cb000000cb000000cb000000ca000000ca000000cf000000b7",
            INIT_38 => X"000000ba000000d4000000d0000000cc000000ce000000c10000008f0000005b",
            INIT_39 => X"00000051000000650000008e000000b5000000c6000000cc000000cf000000cf",
            INIT_3A => X"000000cf000000cf000000cf000000ca000000c5000000c5000000c6000000c5",
            INIT_3B => X"000000c5000000c5000000c5000000c5000000c4000000c5000000cc000000b5",
            INIT_3C => X"000000b8000000d6000000d2000000ce000000d1000000d4000000cf000000b3",
            INIT_3D => X"00000074000000530000005d00000080000000ae000000cb000000d2000000ce",
            INIT_3E => X"000000cc000000ca000000ca000000c9000000c6000000c7000000c9000000c9",
            INIT_3F => X"000000c8000000ca000000c9000000c7000000c6000000c6000000cb000000b4",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY20;


    MEM_IFMAP_LAYER0_ENTITY21 : if BRAM_NAME = "ifmap_layer0_entity21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ba000000d7000000d6000000d5000000d6000000d6000000d4000000d9",
            INIT_01 => X"000000af0000005b0000004900000056000000650000008a000000b5000000cc",
            INIT_02 => X"000000d0000000cb000000c7000000c6000000c7000000c9000000c9000000c8",
            INIT_03 => X"000000c8000000ca000000c9000000c9000000ca000000c8000000cc000000b6",
            INIT_04 => X"000000bb000000d8000000d8000000d9000000db000000d9000000d6000000d3",
            INIT_05 => X"000000cc0000007b00000044000000520000004f000000510000006100000082",
            INIT_06 => X"000000a5000000bc000000c9000000ca000000c4000000c1000000c7000000c6",
            INIT_07 => X"000000c6000000c7000000c8000000c8000000c9000000c7000000cc000000b6",
            INIT_08 => X"000000bc000000d9000000d5000000d6000000d8000000d8000000d6000000d2",
            INIT_09 => X"000000d40000008800000046000000530000004e00000050000000500000004d",
            INIT_0A => X"00000053000000660000007e000000970000009f000000b2000000c9000000cc",
            INIT_0B => X"000000cb000000c9000000c8000000c6000000c7000000c5000000c9000000b4",
            INIT_0C => X"000000bb000000da000000d6000000d5000000d7000000d8000000d7000000d8",
            INIT_0D => X"000000cc000000700000002d000000370000003a000000450000004d00000051",
            INIT_0E => X"000000500000004d000000460000003e0000003b0000004f0000007c000000a0",
            INIT_0F => X"000000b5000000c4000000cd000000cd000000cb000000c8000000ca000000b4",
            INIT_10 => X"000000bc000000d8000000d2000000d1000000d3000000d6000000d4000000d4",
            INIT_11 => X"0000009a0000005f0000003a00000021000000300000003e000000410000004d",
            INIT_12 => X"00000052000000540000005400000048000000380000002f0000003f00000048",
            INIT_13 => X"0000004e0000006b000000840000009e000000b5000000c1000000ca000000b6",
            INIT_14 => X"000000b8000000d2000000ce000000cf000000d1000000d3000000d4000000c8",
            INIT_15 => X"00000091000000850000008f000000610000002d000000320000002e0000005a",
            INIT_16 => X"000000960000009e0000007f0000004700000061000000700000005800000041",
            INIT_17 => X"0000004300000082000000a5000000a2000000a8000000b5000000c5000000b0",
            INIT_18 => X"000000b7000000d2000000cd000000d0000000d3000000d4000000d5000000d2",
            INIT_19 => X"000000d1000000d1000000d4000000bf000000940000009300000093000000a6",
            INIT_1A => X"000000c8000000d0000000c30000009d000000a6000000b5000000b4000000a2",
            INIT_1B => X"0000009f000000b4000000c1000000c5000000c3000000c1000000c7000000b1",
            INIT_1C => X"000000ae000000c4000000c3000000c2000000c2000000be000000bb000000b9",
            INIT_1D => X"000000b8000000b5000000b7000000b5000000b2000000b0000000ae000000ad",
            INIT_1E => X"000000aa000000a4000000a6000000ac000000aa000000a6000000aa000000b0",
            INIT_1F => X"000000af000000a50000009d0000009b0000009d000000a3000000af0000009e",
            INIT_20 => X"000000700000006c000000700000006900000067000000640000006100000060",
            INIT_21 => X"0000005c0000005a0000005e0000005700000054000000530000005700000067",
            INIT_22 => X"00000073000000700000006f0000007000000071000000730000007400000076",
            INIT_23 => X"0000007a0000007b0000007c0000007b000000790000007a000000840000007c",
            INIT_24 => X"00000075000000730000007100000070000000710000006f0000007100000071",
            INIT_25 => X"0000006f000000700000006f0000006e0000006e0000006d0000006e0000006b",
            INIT_26 => X"00000073000000730000006c0000006e0000006f0000006d000000680000006b",
            INIT_27 => X"0000006d0000006e0000007000000070000000640000005f0000006200000065",
            INIT_28 => X"0000007100000066000000690000006a0000006a00000066000000610000005d",
            INIT_29 => X"0000005f0000005e0000005900000055000000520000004e0000004f0000004e",
            INIT_2A => X"000000500000004f000000470000004400000043000000410000004100000041",
            INIT_2B => X"000000410000004200000042000000410000003c000000370000004700000064",
            INIT_2C => X"000000540000003c000000410000004000000040000000400000003e0000003c",
            INIT_2D => X"00000042000000400000003d00000038000000390000003c0000003d0000003f",
            INIT_2E => X"0000004000000043000000410000003b000000380000003a0000003b0000003c",
            INIT_2F => X"0000003a00000039000000380000003800000038000000480000007500000080",
            INIT_30 => X"000000530000003b0000003f0000003e0000003f000000410000003d0000003f",
            INIT_31 => X"000000430000003e0000003c000000390000003a0000003a0000003c0000003d",
            INIT_32 => X"0000004100000044000000400000003e0000003d0000003c0000003e0000003d",
            INIT_33 => X"0000003a0000003a0000003d000000410000005b000000880000008900000063",
            INIT_34 => X"0000004f000000350000003d00000039000000370000003b0000003a0000003c",
            INIT_35 => X"0000003d0000003c00000039000000370000003c0000003e0000003d0000003f",
            INIT_36 => X"000000430000003f0000003c0000003b0000003e0000003e000000400000003f",
            INIT_37 => X"0000003e0000003c000000470000006e0000008e000000770000004f0000004a",
            INIT_38 => X"000000520000003a00000042000000410000003f0000003e0000003e0000003e",
            INIT_39 => X"0000003f0000003e000000410000004f0000004f0000004c0000004a0000004d",
            INIT_3A => X"0000005400000050000000500000004e0000004c0000003f0000003e00000041",
            INIT_3B => X"00000042000000560000007c0000008d00000066000000420000004000000045",
            INIT_3C => X"0000004e000000340000003a0000003a0000003a0000003a0000003b00000039",
            INIT_3D => X"0000003a0000003b0000003a0000004500000047000000470000004600000045",
            INIT_3E => X"0000004800000048000000490000004a000000490000003f0000003f00000044",
            INIT_3F => X"0000005a000000800000008000000058000000420000003f0000004100000044",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY21;


    MEM_IFMAP_LAYER0_ENTITY22 : if BRAM_NAME = "ifmap_layer0_entity22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000095000000bb000000c1000000cd000000ca000000b7000000b5000000b4",
            INIT_01 => X"000000b6000000bd000000c1000000c0000000c0000000c0000000bd000000bd",
            INIT_02 => X"000000ba000000b9000000bd000000c0000000c1000000c1000000c0000000be",
            INIT_03 => X"000000bb000000bb000000bc000000c3000000ca000000d1000000d4000000ab",
            INIT_04 => X"0000009d000000cc000000d7000000e3000000e0000000be000000b3000000b3",
            INIT_05 => X"000000b3000000bb000000c3000000c3000000bb000000be000000b4000000b7",
            INIT_06 => X"000000bc000000b7000000b8000000b7000000b9000000bf000000bc000000bc",
            INIT_07 => X"000000be000000c2000000d3000000e0000000df000000de000000e3000000b7",
            INIT_08 => X"00000099000000c9000000d5000000db000000df000000d5000000c4000000b8",
            INIT_09 => X"000000b1000000c3000000d3000000d4000000d0000000d2000000cc000000ca",
            INIT_0A => X"000000d1000000d1000000d0000000d1000000d2000000d4000000d0000000d0",
            INIT_0B => X"000000d0000000d5000000de000000df000000da000000d7000000e0000000b8",
            INIT_0C => X"000000a6000000cf000000d3000000de000000e2000000dc000000c900000083",
            INIT_0D => X"000000770000009e000000a6000000b1000000b2000000a7000000a6000000ab",
            INIT_0E => X"000000b7000000b2000000b2000000ba000000b9000000ba000000b4000000a5",
            INIT_0F => X"000000cf000000e4000000dc000000dd000000e0000000df000000e6000000ba",
            INIT_10 => X"000000a7000000cb000000ca000000da000000e0000000e1000000d60000008e",
            INIT_11 => X"00000099000000980000007800000081000000810000007e0000007c00000083",
            INIT_12 => X"0000008600000084000000820000008a00000088000000880000008d0000007b",
            INIT_13 => X"000000ba000000e3000000da000000d9000000de000000dc000000e3000000b9",
            INIT_14 => X"000000a4000000c9000000cb000000d9000000dc000000da000000d1000000a5",
            INIT_15 => X"000000c4000000b50000009c000000b4000000b3000000a0000000a3000000ac",
            INIT_16 => X"000000bf000000c1000000be000000c9000000bf000000c0000000c6000000be",
            INIT_17 => X"000000d4000000e1000000e1000000e1000000df000000e1000000e8000000bc",
            INIT_18 => X"000000a4000000c6000000c8000000d9000000d9000000d6000000ac00000068",
            INIT_19 => X"0000009e000000a5000000a6000000af000000a50000009000000097000000a0",
            INIT_1A => X"000000b2000000ad000000bd000000b6000000aa000000b7000000ad000000b9",
            INIT_1B => X"000000a6000000b2000000dc000000e2000000dd000000e0000000e7000000bc",
            INIT_1C => X"000000a9000000c9000000c7000000d8000000da000000cb000000920000006f",
            INIT_1D => X"00000086000000950000009d000000900000009b0000008f0000008f00000090",
            INIT_1E => X"000000930000008e000000940000008e0000007f0000008d0000008e000000b0",
            INIT_1F => X"0000008900000095000000d1000000dc000000d9000000dc000000e4000000ba",
            INIT_20 => X"000000b1000000ce000000c7000000d9000000db000000cd000000c1000000c5",
            INIT_21 => X"000000b8000000b7000000bb000000b8000000c0000000ba000000bb000000bd",
            INIT_22 => X"000000c0000000c2000000c2000000bf000000b2000000ba000000bc000000c8",
            INIT_23 => X"000000c1000000c6000000d6000000db000000db000000dd000000e4000000b9",
            INIT_24 => X"000000ba000000d4000000c5000000d6000000d7000000d6000000dc000000d2",
            INIT_25 => X"000000b9000000bb000000b6000000ba000000b6000000b4000000b9000000ba",
            INIT_26 => X"000000c1000000c6000000c3000000b8000000b5000000b6000000b6000000c6",
            INIT_27 => X"000000de000000de000000dd000000df000000df000000de000000e3000000b7",
            INIT_28 => X"000000bc000000de000000c8000000d8000000d7000000d4000000d6000000cc",
            INIT_29 => X"000000b5000000b8000000b6000000b0000000b5000000b8000000bc000000bf",
            INIT_2A => X"000000bd000000ba000000b8000000b9000000b6000000b8000000ba000000c9",
            INIT_2B => X"000000df000000dd000000dc000000db000000db000000dc000000e3000000b8",
            INIT_2C => X"000000bf000000e2000000cf000000e0000000dc000000d1000000d7000000de",
            INIT_2D => X"000000d9000000d7000000d6000000d7000000d9000000db000000df000000df",
            INIT_2E => X"000000df000000dd000000db000000da000000d8000000d6000000d9000000db",
            INIT_2F => X"000000db000000db000000d9000000d6000000d7000000db000000e3000000ba",
            INIT_30 => X"000000bc000000dc000000d4000000ce000000b500000099000000ac000000d9",
            INIT_31 => X"000000e2000000e1000000dd000000dc000000de000000df000000e1000000e2",
            INIT_32 => X"000000e1000000dd000000dc000000da000000d9000000db000000dc000000da",
            INIT_33 => X"000000d9000000dc000000de000000e0000000e0000000e0000000e6000000bb",
            INIT_34 => X"000000bd000000df000000d6000000c10000009d0000007e0000006300000073",
            INIT_35 => X"0000009d000000c6000000dd000000dd000000da000000dc000000df000000e2",
            INIT_36 => X"000000e2000000e0000000e1000000df000000dc000000dd000000e0000000e0",
            INIT_37 => X"000000df000000de000000de000000de000000dd000000dd000000e2000000b7",
            INIT_38 => X"000000bd000000e2000000de000000e9000000dc000000c4000000920000005a",
            INIT_39 => X"0000005400000071000000a1000000ca000000da000000e0000000e3000000e4",
            INIT_3A => X"000000e2000000e1000000e0000000dc000000d7000000d7000000d8000000d9",
            INIT_3B => X"000000d8000000d8000000d8000000d8000000d7000000da000000e1000000b6",
            INIT_3C => X"000000bb000000e5000000e0000000ea000000e1000000e1000000da000000b3",
            INIT_3D => X"00000073000000580000006a00000091000000c0000000dd000000e4000000e1",
            INIT_3E => X"000000df000000db000000da000000d9000000d6000000d6000000d9000000db",
            INIT_3F => X"000000db000000dd000000dc000000da000000d9000000dc000000e2000000b7",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY22;


    MEM_IFMAP_LAYER0_ENTITY23 : if BRAM_NAME = "ifmap_layer0_entity23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000be000000e9000000de000000e9000000e4000000e2000000e0000000e1",
            INIT_01 => X"000000b500000062000000500000005b0000006a00000092000000c0000000d9",
            INIT_02 => X"000000e0000000e1000000dd000000da000000d9000000da000000da000000d9",
            INIT_03 => X"000000da000000dd000000dd000000dd000000dd000000dc000000e3000000bc",
            INIT_04 => X"000000bf000000ea000000dd000000e9000000e7000000e3000000e2000000dd",
            INIT_05 => X"000000d500000082000000490000004f0000004b000000500000006400000088",
            INIT_06 => X"000000ad000000c8000000d7000000dc000000d9000000d9000000df000000de",
            INIT_07 => X"000000dd000000dd000000db000000db000000da000000db000000e3000000bd",
            INIT_08 => X"000000bd000000e8000000d9000000e4000000e3000000e1000000e2000000dc",
            INIT_09 => X"000000dd000000900000004a000000500000004a0000004c0000004e0000004c",
            INIT_0A => X"000000530000006400000081000000a1000000b0000000c9000000e1000000e2",
            INIT_0B => X"000000df000000dc000000d9000000d7000000d7000000d9000000e1000000bb",
            INIT_0C => X"000000bb000000e8000000d7000000e1000000e0000000e1000000e3000000e2",
            INIT_0D => X"000000d50000007700000032000000380000003b000000450000004d00000052",
            INIT_0E => X"0000005000000048000000420000003f000000410000005b00000085000000a2",
            INIT_0F => X"000000b8000000cc000000da000000df000000dd000000dd000000e3000000bc",
            INIT_10 => X"000000b7000000e7000000de000000df000000df000000e6000000e4000000e1",
            INIT_11 => X"000000a2000000620000003c000000270000003500000043000000440000004e",
            INIT_12 => X"0000005100000052000000530000004800000039000000310000003f00000043",
            INIT_13 => X"0000004b0000006d0000008b000000a8000000c6000000d7000000df000000c3",
            INIT_14 => X"000000b0000000e2000000e2000000de000000de000000e2000000e2000000d4",
            INIT_15 => X"0000009b0000008b000000960000006a0000003500000039000000330000005e",
            INIT_16 => X"0000009a000000a1000000820000004900000063000000720000005a00000043",
            INIT_17 => X"0000004500000086000000ab000000a9000000b7000000c5000000d0000000be",
            INIT_18 => X"000000af000000e1000000e1000000df000000df000000de000000de000000de",
            INIT_19 => X"000000de000000e0000000e4000000cc0000009f0000009f000000a0000000b3",
            INIT_1A => X"000000d6000000dc000000cf000000a9000000b2000000c1000000c0000000ad",
            INIT_1B => X"000000ab000000c3000000d2000000d6000000d8000000d1000000d2000000bd",
            INIT_1C => X"000000a6000000d4000000d7000000d1000000ce000000cc000000c9000000c7",
            INIT_1D => X"000000c7000000c3000000c5000000c2000000c0000000c1000000c2000000c4",
            INIT_1E => X"000000c4000000c2000000c4000000ca000000c8000000c4000000c8000000cd",
            INIT_1F => X"000000ce000000c5000000c0000000bf000000c5000000c5000000c9000000b5",
            INIT_20 => X"0000006500000078000000820000007800000076000000700000006b0000006a",
            INIT_21 => X"0000006500000062000000660000006300000062000000650000006c00000080",
            INIT_22 => X"000000900000009200000092000000930000009400000096000000980000009e",
            INIT_23 => X"000000a4000000a6000000a8000000a8000000a8000000a5000000a700000092",
            INIT_24 => X"0000006f0000008200000086000000860000008a000000880000008900000088",
            INIT_25 => X"0000008400000086000000830000007e0000007f000000800000008300000083",
            INIT_26 => X"0000008a000000860000007f0000008100000081000000800000007c0000007e",
            INIT_27 => X"0000008100000082000000840000008400000077000000730000007300000060",
            INIT_28 => X"000000680000007100000078000000780000007a000000760000006c00000064",
            INIT_29 => X"000000600000005b000000550000005900000058000000550000005700000056",
            INIT_2A => X"000000560000004f000000460000004300000042000000410000003f0000003c",
            INIT_2B => X"0000003b0000003c0000003c0000003b00000036000000320000003f0000004b",
            INIT_2C => X"0000003d000000370000003d000000390000003a0000003f0000003b00000036",
            INIT_2D => X"00000038000000330000002f0000002f00000030000000320000003100000032",
            INIT_2E => X"0000003300000037000000350000002f0000002d0000002e0000003200000037",
            INIT_2F => X"00000036000000340000003400000034000000300000003a0000006800000068",
            INIT_30 => X"000000440000003d000000410000003c0000003e0000003d0000003700000039",
            INIT_31 => X"0000003d00000038000000370000003a0000003b000000380000003800000036",
            INIT_32 => X"000000390000003b000000370000003400000033000000330000003400000034",
            INIT_33 => X"000000330000003500000037000000390000004b00000071000000780000004b",
            INIT_34 => X"0000003e000000340000003b0000003500000039000000390000003400000036",
            INIT_35 => X"0000003600000032000000300000003200000039000000380000003400000035",
            INIT_36 => X"0000003900000036000000340000003300000036000000370000003500000030",
            INIT_37 => X"00000032000000340000003d0000005f0000007c000000650000003e00000032",
            INIT_38 => X"0000003e000000350000003a000000370000003b0000003d0000003c0000003c",
            INIT_39 => X"00000039000000370000003a0000004b0000004c000000480000004400000045",
            INIT_3A => X"0000004b0000004a0000004b00000049000000460000003a0000003700000035",
            INIT_3B => X"00000033000000450000006b0000007f0000005b0000003a0000003600000033",
            INIT_3C => X"0000004000000033000000330000002e00000033000000380000003900000035",
            INIT_3D => X"0000003400000033000000320000003e000000400000003e0000003c00000039",
            INIT_3E => X"0000003c0000003e000000400000004000000040000000350000003400000037",
            INIT_3F => X"0000004600000067000000690000004800000035000000320000003400000032",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY23;


    MEM_IFMAP_LAYER0_ENTITY24 : if BRAM_NAME = "ifmap_layer0_entity24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004100000046000000300000001e00000017000000280000002c0000002d",
            INIT_01 => X"0000002d000000280000000a0000000f0000002c000000350000003300000030",
            INIT_02 => X"000000410000005a0000005d0000005b0000005f000000510000003c00000037",
            INIT_03 => X"000000700000006f00000029000000440000004d000000330000003600000043",
            INIT_04 => X"000000450000004f0000003c0000001e00000029000000410000003100000031",
            INIT_05 => X"0000003100000023000000070000001900000041000000450000003700000031",
            INIT_06 => X"0000004d0000005500000053000000500000005700000051000000370000003b",
            INIT_07 => X"00000083000000790000001f0000002f0000003800000036000000410000003d",
            INIT_08 => X"00000049000000540000004800000029000000400000004a0000003200000036",
            INIT_09 => X"00000036000000200000000b000000240000003c000000430000002f00000027",
            INIT_0A => X"0000004b0000004d0000003b0000003e0000005300000055000000300000003f",
            INIT_0B => X"0000008b000000800000001700000029000000460000004e0000004900000030",
            INIT_0C => X"000000580000004b00000050000000360000005000000044000000370000003f",
            INIT_0D => X"0000003a0000001c00000011000000250000002b000000330000002800000027",
            INIT_0E => X"00000055000000620000004b0000004600000056000000540000003200000044",
            INIT_0F => X"0000008e000000890000002f0000004b000000640000005d0000004100000026",
            INIT_10 => X"0000005f000000590000006f00000042000000510000003d0000003d00000044",
            INIT_11 => X"0000003e000000160000000f000000160000001f00000023000000330000003f",
            INIT_12 => X"000000480000004b00000048000000470000004d00000053000000330000004e",
            INIT_13 => X"000000950000009c0000005700000057000000630000005f0000004b00000058",
            INIT_14 => X"0000005200000053000000520000004d000000470000003a0000004000000039",
            INIT_15 => X"0000003b00000014000000110000001c000000320000003d0000004700000047",
            INIT_16 => X"000000450000004300000044000000380000002900000053000000460000004e",
            INIT_17 => X"0000009c000000ac00000062000000590000005e0000006f0000007000000063",
            INIT_18 => X"0000004500000040000000200000003b000000480000004a0000004900000031",
            INIT_19 => X"00000031000000120000001d0000003e0000005200000055000000560000003f",
            INIT_1A => X"00000022000000340000005f0000002b000000190000005e000000550000004e",
            INIT_1B => X"000000a6000000b40000006d0000006b0000006c00000083000000560000002f",
            INIT_1C => X"0000003b000000350000001900000046000000510000004e000000500000003d",
            INIT_1D => X"000000280000000a000000350000005e00000057000000580000004b00000019",
            INIT_1E => X"0000000d0000002d0000005c0000003900000032000000650000005900000062",
            INIT_1F => X"00000090000000b3000000780000007c0000007c000000800000003400000018",
            INIT_20 => X"000000440000002f000000310000006600000077000000590000003f0000004f",
            INIT_21 => X"00000042000000220000005100000060000000590000005a000000290000000e",
            INIT_22 => X"000000340000005c00000043000000470000006f000000710000006e00000073",
            INIT_23 => X"000000880000009c000000790000007f0000007c000000730000001f00000016",
            INIT_24 => X"0000004d000000350000003700000072000000800000007b0000004100000037",
            INIT_25 => X"0000004f000000520000006f0000006e0000006a000000450000001400000025",
            INIT_26 => X"0000005c0000006900000053000000610000007600000078000000730000005c",
            INIT_27 => X"00000090000000930000007d0000007f000000770000005f0000000e00000017",
            INIT_28 => X"000000550000003a000000360000007000000081000000840000006400000031",
            INIT_29 => X"0000002700000054000000680000006d0000007d0000005d0000003f00000053",
            INIT_2A => X"000000610000005e000000680000006e0000006d0000007f0000005500000039",
            INIT_2B => X"00000098000000960000007b0000007c000000720000005d0000000c00000015",
            INIT_2C => X"0000006c00000035000000320000006b0000007e00000083000000800000004b",
            INIT_2D => X"000000330000005b000000550000006b0000008a0000006e0000008100000093",
            INIT_2E => X"0000008400000078000000710000007700000075000000730000005a0000005d",
            INIT_2F => X"000000a00000008d000000710000007d00000079000000650000000e00000009",
            INIT_30 => X"000000600000002a0000002b0000005c0000006a000000800000008200000077",
            INIT_31 => X"000000780000007b0000007200000089000000940000006e0000006900000084",
            INIT_32 => X"000000920000008700000080000000860000008c000000780000007e00000077",
            INIT_33 => X"0000009800000091000000630000006a00000082000000630000001200000028",
            INIT_34 => X"00000061000000420000003b00000059000000640000006f0000008500000088",
            INIT_35 => X"000000930000008c00000096000000910000008e00000088000000830000007f",
            INIT_36 => X"0000007d0000007b0000008800000093000000970000008e0000009c00000088",
            INIT_37 => X"00000092000000900000006d00000070000000820000005c0000003200000053",
            INIT_38 => X"00000069000000480000004b0000005f000000680000005e0000008500000085",
            INIT_39 => X"0000008f0000008700000080000000850000009300000096000000a000000098",
            INIT_3A => X"000000910000009000000084000000870000008a0000008a000000a2000000a5",
            INIT_3B => X"000000a30000007f0000007e00000077000000760000005f0000003b0000004d",
            INIT_3C => X"0000005e00000044000000440000005b00000065000000620000007b00000083",
            INIT_3D => X"00000093000000c10000008a0000004f0000007c0000009300000093000000a2",
            INIT_3E => X"000000b4000000ab0000009800000090000000900000007900000094000000b3",
            INIT_3F => X"000000b4000000a0000000800000007b000000700000003f0000001a00000054",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY24;


    MEM_IFMAP_LAYER0_ENTITY25 : if BRAM_NAME = "ifmap_layer0_entity25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000580000004f0000004a000000590000006e000000780000007800000081",
            INIT_01 => X"00000078000000b8000000c000000057000000720000009c000000a4000000a6",
            INIT_02 => X"0000009a000000a1000000b7000000b6000000bb000000ad000000940000008f",
            INIT_03 => X"000000b5000000c30000008e0000007c0000006b0000002c0000002900000076",
            INIT_04 => X"0000005b00000059000000670000006000000074000000640000006f0000006a",
            INIT_05 => X"0000007200000080000000bb000000a80000008c00000099000000ac000000ac",
            INIT_06 => X"000000a7000000a40000009d000000a3000000a1000000a5000000ab0000009c",
            INIT_07 => X"000000a100000091000000a7000000720000006a0000004a0000002a0000005e",
            INIT_08 => X"0000006500000061000000780000007a000000720000004e0000005f0000005b",
            INIT_09 => X"000000730000006e00000081000000cc000000a700000089000000a000000099",
            INIT_0A => X"000000b3000000ba000000aa000000b2000000b30000009c000000a2000000a5",
            INIT_0B => X"0000009c0000008c000000680000004800000054000000590000004600000072",
            INIT_0C => X"0000006e0000006b0000007a000000600000005a0000004c0000004800000064",
            INIT_0D => X"0000006d0000007f000000570000008c000000bd0000009f000000a6000000b4",
            INIT_0E => X"000000ae000000ad000000be000000bc000000a200000099000000a2000000a1",
            INIT_0F => X"00000099000000950000004b0000004a000000420000003e000000700000008a",
            INIT_10 => X"000000770000006a000000590000004e00000059000000470000003c00000067",
            INIT_11 => X"0000004b0000005f00000072000000420000007f000000b5000000ae000000be",
            INIT_12 => X"000000ba000000ab000000b8000000c1000000a4000000a0000000ab000000a5",
            INIT_13 => X"000000920000008b000000680000005c0000004d0000005e0000007000000073",
            INIT_14 => X"0000007e0000005e0000003a000000670000006a0000004c000000480000005f",
            INIT_15 => X"0000005e0000004100000078000000630000005b000000a1000000c4000000bc",
            INIT_16 => X"000000b6000000c1000000a7000000a7000000aa000000a00000009a000000a1",
            INIT_17 => X"000000910000008a0000006e0000005100000069000000880000006d00000064",
            INIT_18 => X"0000006f000000520000004600000068000000710000005e0000004500000054",
            INIT_19 => X"000000740000006d000000550000007d0000007f0000009b000000ba000000c8",
            INIT_1A => X"000000bb000000bb000000b10000009d00000094000000a2000000a4000000a6",
            INIT_1B => X"000000a200000095000000790000006100000078000000730000006100000061",
            INIT_1C => X"000000650000005c0000008c000000b4000000970000007b000000550000004c",
            INIT_1D => X"000000670000007c0000005a0000005400000092000000af000000ad000000c8",
            INIT_1E => X"000000bc000000ad000000ad0000009f0000009f000000ac000000a3000000ad",
            INIT_1F => X"000000a40000008b0000008300000083000000700000005f0000006400000060",
            INIT_20 => X"0000007700000090000000c0000000d1000000c20000009d0000007f0000006c",
            INIT_21 => X"0000006a0000005e0000006a0000006f0000007c000000af000000b0000000c5",
            INIT_22 => X"000000b8000000aa000000b0000000a50000009c000000c5000000af000000a3",
            INIT_23 => X"00000093000000830000007a0000006500000064000000600000006b00000066",
            INIT_24 => X"0000006e000000740000008a000000a9000000c5000000c4000000a000000088",
            INIT_25 => X"00000081000000630000005c0000008a000000920000009f000000b4000000a9",
            INIT_26 => X"0000008e0000008d000000af000000b2000000a6000000bc000000b300000097",
            INIT_27 => X"0000008f0000009a000000700000003a0000005b000000650000006600000049",
            INIT_28 => X"0000005b000000570000004a0000006b000000a5000000b9000000bf000000a3",
            INIT_29 => X"00000086000000800000006a0000006600000076000000840000009200000074",
            INIT_2A => X"0000004d00000063000000a1000000b6000000b70000009f000000ad000000a7",
            INIT_2B => X"0000009c000000870000005e0000002b0000005b0000005c000000440000004d",
            INIT_2C => X"000000510000005f000000320000002c0000005f00000094000000a6000000bb",
            INIT_2D => X"000000ae000000900000007e000000720000006800000072000000770000006b",
            INIT_2E => X"00000051000000520000009d000000b6000000a9000000b2000000a900000096",
            INIT_2F => X"000000980000006c0000002c0000003f00000061000000450000005000000056",
            INIT_30 => X"0000005a0000005f00000034000000150000001c0000006d00000092000000b0",
            INIT_31 => X"000000ca000000b50000008e0000007f00000078000000770000007200000082",
            INIT_32 => X"000000810000007600000090000000a90000009f000000ad000000b400000098",
            INIT_33 => X"00000077000000440000002c000000550000003300000072000000a70000006a",
            INIT_34 => X"0000005f0000005b00000039000000340000001800000031000000770000009c",
            INIT_35 => X"000000bb000000cb000000ba0000009b0000008d000000850000007400000075",
            INIT_36 => X"0000006d000000770000008b000000990000009f000000a70000009c0000007d",
            INIT_37 => X"000000650000004100000044000000400000003700000090000000aa0000007a",
            INIT_38 => X"0000005e0000004b00000020000000490000002e000000210000003600000073",
            INIT_39 => X"00000096000000b0000000c3000000c2000000b10000009b0000008800000092",
            INIT_3A => X"0000008b000000650000005e00000077000000650000005f0000006000000069",
            INIT_3B => X"00000083000000760000006b0000006d000000800000008f0000009a0000006a",
            INIT_3C => X"0000004e00000023000000180000004c00000041000000280000001b0000003b",
            INIT_3D => X"000000780000008800000096000000b0000000c0000000b7000000a5000000ba",
            INIT_3E => X"000000cf000000aa0000006b000000560000004200000055000000700000008c",
            INIT_3F => X"000000a9000000950000008900000089000000960000008f0000009a00000080",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY25;


    MEM_IFMAP_LAYER0_ENTITY26 : if BRAM_NAME = "ifmap_layer0_entity26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004400000051000000400000002e00000021000000390000004b00000050",
            INIT_01 => X"00000053000000460000001400000022000000470000004b0000004600000042",
            INIT_02 => X"00000057000000780000007c000000790000007e0000006c0000005400000052",
            INIT_03 => X"00000088000000810000003b0000005b00000060000000430000004c00000057",
            INIT_04 => X"00000050000000660000004a0000002f000000380000005c0000005400000054",
            INIT_05 => X"000000580000003e00000012000000300000005d0000005c0000004d00000049",
            INIT_06 => X"0000006b000000750000006f0000006a000000750000006c0000004d00000053",
            INIT_07 => X"000000970000008b0000002d0000004100000047000000420000005a00000051",
            INIT_08 => X"0000005f0000006d00000058000000380000005400000069000000560000005a",
            INIT_09 => X"0000005c00000035000000140000003c0000005900000058000000420000003c",
            INIT_0A => X"00000067000000660000004e0000005400000072000000720000004200000056",
            INIT_0B => X"0000009e0000008f00000023000000370000005400000062000000620000003b",
            INIT_0C => X"000000740000006400000064000000490000006d000000660000005800000060",
            INIT_0D => X"0000005e0000002d0000001a0000003800000041000000430000003600000037",
            INIT_0E => X"0000006a0000007500000061000000620000007600000072000000450000005b",
            INIT_0F => X"000000a000000096000000400000005d000000780000007e0000005e00000032",
            INIT_10 => X"0000007800000068000000800000005d000000720000005e0000005a0000005e",
            INIT_11 => X"0000005d000000270000001a000000240000002f000000370000004900000056",
            INIT_12 => X"00000069000000710000006b00000065000000670000006d0000004a00000067",
            INIT_13 => X"000000a2000000ac00000070000000740000008100000084000000670000006c",
            INIT_14 => X"000000690000006600000062000000620000005f000000590000005b0000004e",
            INIT_15 => X"00000058000000230000001b0000002b0000004d0000005d0000006a0000006c",
            INIT_16 => X"0000006700000065000000640000004e000000390000006e0000006200000066",
            INIT_17 => X"000000a7000000ba000000820000007f00000081000000900000008400000078",
            INIT_18 => X"0000005e00000060000000300000004f0000005a000000640000005d0000003f",
            INIT_19 => X"0000004a0000001d000000260000005a0000007e000000810000008200000063",
            INIT_1A => X"0000003a000000470000007300000039000000250000007b000000710000006a",
            INIT_1B => X"000000b7000000c10000008d0000008c00000089000000a0000000650000003b",
            INIT_1C => X"00000056000000540000002f0000006900000067000000610000005e00000047",
            INIT_1D => X"0000003800000014000000490000008b0000008a0000008c0000007200000029",
            INIT_1E => X"0000001a00000041000000730000004f0000003b0000007d000000780000008c",
            INIT_1F => X"000000b0000000c30000009600000094000000900000009b0000003f00000018",
            INIT_20 => X"000000620000004e0000004a0000008c0000009500000072000000500000005c",
            INIT_21 => X"000000470000002c000000710000009000000088000000860000003f00000017",
            INIT_22 => X"000000450000007c0000005e00000056000000700000008b0000009b000000a5",
            INIT_23 => X"000000aa000000b10000009600000096000000920000008e0000002900000016",
            INIT_24 => X"00000074000000510000004e00000094000000a30000009b0000005400000045",
            INIT_25 => X"000000510000005a000000890000008e0000008a0000005d0000002100000038",
            INIT_26 => X"0000007c0000008f0000007300000080000000970000009c0000009c00000081",
            INIT_27 => X"000000a7000000ad000000980000009a00000094000000790000001600000018",
            INIT_28 => X"000000780000004f0000004900000091000000a5000000a60000007f00000041",
            INIT_29 => X"00000036000000720000008e0000007f0000007e0000005d000000470000006c",
            INIT_2A => X"000000870000008500000092000000a10000009c000000a50000007500000057",
            INIT_2B => X"000000a9000000af000000970000009c00000091000000740000001300000017",
            INIT_2C => X"0000007b00000045000000420000008a000000a1000000a8000000a50000005f",
            INIT_2D => X"0000004b0000008c0000008a000000700000006d0000006600000088000000a2",
            INIT_2E => X"000000990000009a00000097000000870000007c000000850000007600000088",
            INIT_2F => X"000000bd000000aa000000920000009d0000009400000077000000140000000b",
            INIT_30 => X"0000006a000000390000003c0000007900000087000000a4000000ad00000098",
            INIT_31 => X"00000090000000930000007f00000076000000730000005c000000660000008b",
            INIT_32 => X"0000008d0000008a0000008500000074000000780000006b0000007700000088",
            INIT_33 => X"000000b0000000ae0000008700000091000000a1000000720000001a0000002b",
            INIT_34 => X"00000074000000550000004e000000740000007f0000008c000000ac000000ab",
            INIT_35 => X"000000990000007c00000082000000780000007700000076000000710000006e",
            INIT_36 => X"000000690000006c000000770000007d000000830000007a0000008100000075",
            INIT_37 => X"00000090000000a20000008d0000009a000000a600000070000000410000005f",
            INIT_38 => X"000000840000006000000063000000780000008200000072000000a5000000a8",
            INIT_39 => X"0000008b0000006b00000068000000700000007c000000810000008e00000084",
            INIT_3A => X"0000007a000000770000006b0000006f00000073000000760000008d00000090",
            INIT_3B => X"0000008e0000007b000000920000009f0000009d00000070000000480000005e",
            INIT_3C => X"000000790000005a0000005d000000760000007f0000007c00000097000000a6",
            INIT_3D => X"00000099000000ab00000079000000450000006b0000007c0000007b0000008b",
            INIT_3E => X"0000009b0000009000000080000000770000007a0000006700000083000000a7",
            INIT_3F => X"0000009f0000008c00000080000000a0000000950000004b0000002200000068",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY26;


    MEM_IFMAP_LAYER0_ENTITY27 : if BRAM_NAME = "ifmap_layer0_entity27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007000000064000000640000007e0000008d0000009800000095000000a3",
            INIT_01 => X"0000008a000000a3000000a60000004700000064000000850000008b0000008d",
            INIT_02 => X"0000008100000088000000a00000009e000000a3000000970000007d0000007e",
            INIT_03 => X"000000a9000000b10000007a0000008f0000008f0000003d000000330000008b",
            INIT_04 => X"00000070000000700000008300000081000000930000007c0000009000000089",
            INIT_05 => X"0000008f00000079000000a8000000990000007a0000007f0000009200000093",
            INIT_06 => X"0000008d0000008b000000840000008a000000860000008f0000009900000086",
            INIT_07 => X"0000009100000082000000920000007a00000086000000640000003a0000006f",
            INIT_08 => X"0000007900000076000000950000008e0000008d000000610000007b00000076",
            INIT_09 => X"0000008f0000007e00000079000000bb000000910000006e0000008800000082",
            INIT_0A => X"0000009a000000a1000000940000009a00000097000000860000009600000091",
            INIT_0B => X"000000860000007b000000610000005700000067000000770000006100000086",
            INIT_0C => X"0000008800000087000000970000006f0000007a000000650000005d0000007d",
            INIT_0D => X"0000008600000099000000600000007d000000a90000008800000092000000a0",
            INIT_0E => X"0000009600000094000000a6000000a70000008d000000800000009000000091",
            INIT_0F => X"00000084000000820000004b0000005e000000530000005700000095000000a9",
            INIT_10 => X"000000940000008c000000700000005e00000079000000680000005400000082",
            INIT_11 => X"00000066000000740000008d0000004a00000076000000a30000009b000000aa",
            INIT_12 => X"000000a5000000950000009d000000a700000092000000890000009300000091",
            INIT_13 => X"0000007f0000007c0000006d0000007100000060000000770000009c000000a1",
            INIT_14 => X"0000009800000077000000480000007d00000081000000650000006300000079",
            INIT_15 => X"000000780000005b0000009a0000007d0000005d00000096000000b5000000a9",
            INIT_16 => X"000000a2000000ad000000910000008f0000008f00000087000000810000008b",
            INIT_17 => X"0000007d00000078000000750000006600000081000000ab0000009a00000099",
            INIT_18 => X"0000008800000068000000520000007b00000088000000760000006200000073",
            INIT_19 => X"000000960000008d00000075000000940000008100000095000000ad000000b3",
            INIT_1A => X"000000a5000000a80000009f0000008f0000007e0000008b0000008c0000008d",
            INIT_1B => X"00000088000000850000007a0000006d00000098000000a40000009600000095",
            INIT_1C => X"0000007d0000006f00000096000000bf000000ac0000009e000000790000006f",
            INIT_1D => X"0000009100000099000000730000006900000094000000a10000009a000000ac",
            INIT_1E => X"000000a10000009b0000009c0000008d0000008900000093000000880000008f",
            INIT_1F => X"000000890000008c0000007b000000860000009c000000950000009e00000095",
            INIT_20 => X"00000095000000a2000000c8000000dc000000d1000000bd000000aa00000093",
            INIT_21 => X"000000910000007a0000007d000000880000008b0000009f00000096000000a4",
            INIT_22 => X"0000009b0000009b0000009f0000008e00000085000000a90000009300000088",
            INIT_23 => X"0000007f0000007e0000006b000000720000009a0000008f000000a00000009c",
            INIT_24 => X"0000008b000000890000009d000000be000000d5000000d7000000bf000000b0",
            INIT_25 => X"000000a90000008400000075000000a3000000ad000000970000009a0000008f",
            INIT_26 => X"0000007c00000081000000990000009800000091000000a3000000950000007c",
            INIT_27 => X"0000007700000083000000600000004a00000091000000950000009700000078",
            INIT_28 => X"000000730000006f0000006100000086000000bf000000cf000000d3000000c1",
            INIT_29 => X"000000b1000000ad000000910000007f000000900000008f0000008600000068",
            INIT_2A => X"000000490000005c0000008b0000009b000000a10000008a000000940000008e",
            INIT_2B => X"0000008300000075000000550000003c00000092000000910000006f0000006d",
            INIT_2C => X"0000006a00000072000000410000004000000078000000b2000000c3000000d5",
            INIT_2D => X"000000ca000000b9000000ad000000990000008e000000960000008d0000007d",
            INIT_2E => X"0000006c000000600000008e0000009a00000090000000a1000000950000007f",
            INIT_2F => X"00000083000000620000003100000061000000930000006c0000007600000075",
            INIT_30 => X"00000074000000700000003e000000260000002900000087000000b4000000c7",
            INIT_31 => X"000000d4000000cc000000b7000000b2000000ab000000a40000009e000000a1",
            INIT_32 => X"0000009d0000008b000000870000008d00000087000000990000009c0000007e",
            INIT_33 => X"00000067000000420000003b0000007c0000005400000088000000c500000083",
            INIT_34 => X"0000007f0000007b0000004f0000004e000000250000004200000095000000bf",
            INIT_35 => X"000000d0000000db000000d6000000c2000000b8000000b4000000a50000009f",
            INIT_36 => X"000000870000007d0000007b000000830000008a000000930000008700000072",
            INIT_37 => X"0000006c0000004f000000550000005b0000004e000000ac000000c90000008f",
            INIT_38 => X"0000007d00000068000000340000006b00000043000000300000004e00000097",
            INIT_39 => X"000000bd000000cb000000d9000000da000000cd000000c3000000b4000000b6",
            INIT_3A => X"000000a5000000740000005e0000007a0000006100000059000000590000006f",
            INIT_3B => X"000000960000008a00000082000000860000009f000000b5000000bc00000081",
            INIT_3C => X"00000066000000330000002800000073000000600000003a000000290000004e",
            INIT_3D => X"000000a0000000b5000000b9000000cf000000da000000d2000000c4000000ce",
            INIT_3E => X"000000d6000000b40000007c00000071000000560000006600000084000000a0",
            INIT_3F => X"000000ba000000a7000000a7000000a7000000b4000000b3000000b90000009c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY27;


    MEM_IFMAP_LAYER0_ENTITY28 : if BRAM_NAME = "ifmap_layer0_entity28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000032000000400000002e0000001e00000016000000240000003700000039",
            INIT_01 => X"0000003b000000360000000c000000120000002b0000002c0000003100000032",
            INIT_02 => X"0000003a0000004d000000510000004d000000530000004e0000003800000039",
            INIT_03 => X"000000610000005d0000001f0000003a00000041000000290000003500000042",
            INIT_04 => X"0000003a00000051000000390000001d000000230000003d0000003b0000003c",
            INIT_05 => X"000000400000002f000000070000001b000000380000003e0000003b0000002f",
            INIT_06 => X"000000440000004a0000004a000000440000004e00000051000000330000003c",
            INIT_07 => X"0000006f0000006000000015000000270000002d0000002c0000004500000042",
            INIT_08 => X"0000004800000057000000460000002300000035000000480000003c00000041",
            INIT_09 => X"0000004500000026000000070000002300000034000000410000003000000021",
            INIT_0A => X"000000430000004200000032000000370000004d000000520000002d0000003e",
            INIT_0B => X"000000740000006300000010000000260000003f0000004b0000004d00000033",
            INIT_0C => X"0000005e0000004c000000500000002f0000004700000048000000410000004a",
            INIT_0D => X"000000480000001e0000000c000000220000002800000034000000230000001e",
            INIT_0E => X"0000004b000000570000004400000045000000510000004d0000002e00000043",
            INIT_0F => X"000000770000006b0000002a000000490000005f000000600000004400000022",
            INIT_10 => X"000000610000004f0000006a0000003c0000004b00000044000000480000004c",
            INIT_11 => X"00000049000000180000000c000000110000001c00000025000000330000003b",
            INIT_12 => X"000000480000004f0000004b0000004700000047000000490000002d0000004d",
            INIT_13 => X"000000800000008100000052000000550000005e000000610000004900000050",
            INIT_14 => X"000000520000004d0000004b000000430000003d000000450000004d0000003d",
            INIT_15 => X"00000043000000130000000d000000160000002c0000003b0000004700000049",
            INIT_16 => X"0000004800000048000000490000003500000022000000490000003e0000004d",
            INIT_17 => X"0000008800000093000000600000005b0000005c0000006e000000680000005c",
            INIT_18 => X"000000480000004600000019000000330000003e0000004f0000004f00000032",
            INIT_19 => X"000000380000000f0000001800000036000000490000004b0000004d0000003e",
            INIT_1A => X"0000002200000033000000600000002a0000001600000058000000480000004a",
            INIT_1B => X"00000095000000a1000000680000006c0000006b00000083000000510000002b",
            INIT_1C => X"0000003f0000003b00000015000000460000004d000000480000004b0000003a",
            INIT_1D => X"00000029000000080000002f000000510000004b0000004b0000003e00000012",
            INIT_1E => X"000000060000002700000059000000400000002a0000005e0000004800000053",
            INIT_1F => X"00000083000000a2000000720000007800000076000000850000003400000015",
            INIT_20 => X"0000004900000035000000310000006800000079000000580000003900000046",
            INIT_21 => X"000000330000001700000047000000530000004e0000004f0000002200000007",
            INIT_22 => X"00000028000000510000003c0000003e00000050000000630000005b0000005d",
            INIT_23 => X"000000730000008d0000007800000079000000790000007c0000002100000014",
            INIT_24 => X"000000560000003a0000003800000076000000830000007f0000004000000033",
            INIT_25 => X"0000003b0000004000000061000000630000005e0000003a0000000d0000001c",
            INIT_26 => X"000000530000005d000000490000005000000062000000690000005f0000004a",
            INIT_27 => X"0000007400000084000000770000007e0000007f000000650000000d00000017",
            INIT_28 => X"0000005b0000003b000000350000007400000084000000870000006700000030",
            INIT_29 => X"000000200000004b0000006000000061000000660000004a0000003200000049",
            INIT_2A => X"0000005a000000520000005900000061000000620000006c0000004700000031",
            INIT_2B => X"000000770000007c000000770000008a0000007b0000005b0000000a00000014",
            INIT_2C => X"00000065000000330000002f0000006e00000081000000870000008700000048",
            INIT_2D => X"0000002e00000054000000520000004f0000005e000000560000007500000087",
            INIT_2E => X"00000078000000660000005d0000005e0000005c000000580000004a00000058",
            INIT_2F => X"0000008400000073000000760000008d000000770000005b0000000b00000007",
            INIT_30 => X"000000580000002800000028000000600000006b000000830000008b00000077",
            INIT_31 => X"0000006b0000006600000057000000590000005f0000004a000000510000006c",
            INIT_32 => X"000000760000006e000000640000005d0000006600000055000000570000005f",
            INIT_33 => X"0000007c0000007800000065000000710000007b000000590000000f00000020",
            INIT_34 => X"0000005f0000003f000000370000005c000000640000006e0000008b00000089",
            INIT_35 => X"0000007b00000061000000650000005c0000005a000000580000005600000056",
            INIT_36 => X"0000005500000058000000640000006c000000720000006c0000006e0000005f",
            INIT_37 => X"0000006d000000750000006b000000730000008000000058000000310000004c",
            INIT_38 => X"0000006a00000045000000470000006000000068000000560000008600000087",
            INIT_39 => X"0000007400000057000000510000005800000060000000600000006e0000006a",
            INIT_3A => X"000000620000005f000000570000005c000000610000006b0000007f00000080",
            INIT_3B => X"0000007a0000005e00000074000000770000007a0000005c0000003500000046",
            INIT_3C => X"0000006000000040000000400000005c000000670000005f0000007900000085",
            INIT_3D => X"0000008100000096000000640000003300000058000000650000006200000071",
            INIT_3E => X"0000008300000077000000650000005f00000060000000530000007100000098",
            INIT_3F => X"0000009400000078000000620000007c00000076000000390000000d00000048",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY28;


    MEM_IFMAP_LAYER0_ENTITY29 : if BRAM_NAME = "ifmap_layer0_entity29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000570000004c000000470000005a000000730000007c0000007800000082",
            INIT_01 => X"0000006e0000008e000000960000003a00000054000000740000007700000078",
            INIT_02 => X"0000006c000000710000008500000086000000890000007e000000670000006e",
            INIT_03 => X"0000009f000000a30000006300000072000000750000002a000000210000006b",
            INIT_04 => X"0000005600000058000000640000005d00000075000000630000007500000069",
            INIT_05 => X"0000006e000000660000009b0000008b0000006b0000006f0000008100000081",
            INIT_06 => X"0000007c000000770000006d0000007600000071000000760000007c00000071",
            INIT_07 => X"0000008300000075000000830000006300000069000000480000002700000057",
            INIT_08 => X"0000005f0000006000000078000000730000006d000000470000006300000056",
            INIT_09 => X"0000006c000000630000006a000000b0000000820000005e0000007b00000075",
            INIT_0A => X"000000890000008d0000008100000088000000830000006f0000007800000079",
            INIT_0B => X"000000750000006b00000050000000430000004800000051000000430000006e",
            INIT_0C => X"0000006d000000700000007d000000570000005800000048000000470000005e",
            INIT_0D => X"0000006400000079000000490000007300000098000000760000008700000094",
            INIT_0E => X"000000850000008200000094000000950000007d00000071000000790000007a",
            INIT_0F => X"00000072000000710000003a0000004e0000003d00000038000000730000008a",
            INIT_10 => X"0000007700000074000000590000004300000058000000480000003c00000066",
            INIT_11 => X"00000048000000570000006d0000003700000065000000920000008d0000009c",
            INIT_12 => X"00000098000000880000008c00000098000000860000007b0000007f0000007c",
            INIT_13 => X"0000006d000000690000005d000000620000004d000000620000007a00000077",
            INIT_14 => X"0000007e00000061000000320000005d00000060000000460000004b00000060",
            INIT_15 => X"0000005a0000003b00000076000000610000004900000083000000a200000097",
            INIT_16 => X"00000096000000a3000000840000007f0000007d000000760000006e00000075",
            INIT_17 => X"00000069000000660000005e0000004f0000006b0000008e000000700000006a",
            INIT_18 => X"000000700000005100000037000000590000005c0000004e0000004500000059",
            INIT_19 => X"000000770000006b00000053000000760000006b0000007d000000970000009c",
            INIT_1A => X"000000940000009b000000940000007e0000006c0000007b0000007800000075",
            INIT_1B => X"0000007200000066000000540000005600000081000000790000006300000069",
            INIT_1C => X"0000006200000056000000780000009a000000770000005f000000450000004e",
            INIT_1D => X"000000730000007e000000570000004e0000007d0000008b0000008400000096",
            INIT_1E => X"0000008d0000008e000000920000007e0000007900000084000000760000007b",
            INIT_1F => X"0000007300000058000000520000006f00000079000000650000006a00000067",
            INIT_20 => X"0000007400000088000000a7000000b60000009f00000077000000600000005c",
            INIT_21 => X"000000660000005a000000660000006f0000007000000088000000830000008f",
            INIT_22 => X"000000860000008e0000009600000080000000750000009c0000008400000077",
            INIT_23 => X"00000066000000590000004e000000530000006a00000060000000710000006c",
            INIT_24 => X"0000006c0000006d0000007100000092000000a60000009e0000007b00000069",
            INIT_25 => X"0000006600000052000000550000008c000000910000007e000000860000007b",
            INIT_26 => X"00000068000000730000008a0000008900000083000000960000008a0000006a",
            INIT_27 => X"000000610000006f0000004a0000002d0000006000000065000000690000004b",
            INIT_28 => X"000000580000005500000037000000560000008b00000097000000970000007e",
            INIT_29 => X"000000680000006800000057000000570000006f0000006e0000006e00000052",
            INIT_2A => X"000000350000004b000000790000008c0000009100000078000000810000007a",
            INIT_2B => X"00000074000000620000003e0000002000000061000000620000004100000040",
            INIT_2C => X"000000520000005c00000022000000200000004b00000075000000860000009c",
            INIT_2D => X"0000008d0000006d0000006200000057000000520000005a0000005b0000005f",
            INIT_2E => X"0000005200000046000000790000008b000000810000008f000000800000006b",
            INIT_2F => X"000000710000004e0000001d0000003f00000063000000470000004700000042",
            INIT_30 => X"0000005a00000056000000230000000d0000000f0000004e0000007200000094",
            INIT_31 => X"000000a20000008b0000006f00000062000000610000005b0000005600000071",
            INIT_32 => X"000000780000006a000000730000007e0000007600000087000000870000006a",
            INIT_33 => X"0000004f0000002a000000260000005b0000002c000000600000009900000053",
            INIT_34 => X"0000005c000000560000002d000000250000000d0000001f000000570000007a",
            INIT_35 => X"00000096000000ad0000009e0000007a00000075000000720000005d0000005c",
            INIT_36 => X"0000004d0000005500000067000000710000007e00000085000000730000005b",
            INIT_37 => X"0000004e000000320000003b0000003c0000002a0000006c0000008600000062",
            INIT_38 => X"0000005200000047000000180000003800000024000000170000002300000054",
            INIT_39 => X"0000007600000092000000a5000000a500000096000000820000006f00000079",
            INIT_3A => X"0000006c000000420000003f000000620000004e000000450000004600000056",
            INIT_3B => X"000000750000006c000000600000006200000078000000740000007b00000059",
            INIT_3C => X"000000410000001b0000001100000040000000340000001d0000000f00000025",
            INIT_3D => X"00000059000000640000007400000096000000aa00000098000000880000009c",
            INIT_3E => X"000000a600000079000000450000004a0000002f00000047000000660000007f",
            INIT_3F => X"0000009c0000008b000000830000008200000093000000880000009200000075",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY29;


    MEM_IFMAP_LAYER0_ENTITY30 : if BRAM_NAME = "ifmap_layer0_entity30" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b30000008b0000004d000000580000008d0000009d0000009c00000097",
            INIT_01 => X"0000009c0000009e000000900000009700000097000000880000007900000076",
            INIT_02 => X"0000007e0000006c000000540000005400000062000000620000005e00000053",
            INIT_03 => X"0000005a00000056000000540000006000000075000000570000004c0000004d",
            INIT_04 => X"000000b80000008500000080000000920000009f0000009f0000009e000000a7",
            INIT_05 => X"000000a5000000a2000000990000009a0000009600000096000000880000007d",
            INIT_06 => X"000000810000006d0000005a000000520000005d000000620000005e00000058",
            INIT_07 => X"0000004e0000004c0000005b0000006a00000076000000620000005b0000005a",
            INIT_08 => X"000000b400000098000000b0000000aa000000a4000000980000009b000000a4",
            INIT_09 => X"000000a2000000aa000000a20000009f0000009c00000097000000920000008c",
            INIT_0A => X"000000920000007c00000058000000470000005500000062000000670000006b",
            INIT_0B => X"000000650000006d0000006f0000006f0000006f000000650000005d0000005f",
            INIT_0C => X"000000af000000ae000000b8000000b5000000a800000098000000a4000000a3",
            INIT_0D => X"000000a6000000b3000000a7000000a8000000ae000000a20000009f000000a4",
            INIT_0E => X"0000009700000089000000590000003a000000480000005a000000630000006b",
            INIT_0F => X"00000075000000800000007d0000007900000069000000610000006d0000006f",
            INIT_10 => X"000000af000000ae000000a7000000ac000000a2000000a1000000b0000000af",
            INIT_11 => X"000000b2000000b2000000b3000000b4000000b0000000a8000000a0000000a4",
            INIT_12 => X"000000ad0000009c0000007800000045000000420000005a000000630000005e",
            INIT_13 => X"000000690000007c0000007f0000007b00000070000000680000007100000074",
            INIT_14 => X"000000b5000000ae00000090000000aa000000a9000000a6000000b0000000b3",
            INIT_15 => X"000000b4000000b4000000b4000000b5000000b0000000ae0000009f00000096",
            INIT_16 => X"000000b5000000af0000009b00000074000000600000007d0000008300000070",
            INIT_17 => X"00000075000000780000007a000000790000007900000078000000760000007c",
            INIT_18 => X"000000c00000009c0000008a000000b2000000af000000ae000000b0000000af",
            INIT_19 => X"000000b8000000b4000000ba000000b8000000bb000000bb000000ad00000099",
            INIT_1A => X"000000a6000000ad000000ad000000a700000096000000950000009400000079",
            INIT_1B => X"00000073000000750000006d0000006f000000780000007a0000007b00000080",
            INIT_1C => X"000000b90000007d0000009c000000ab000000ad000000af000000af000000b8",
            INIT_1D => X"000000bc000000b7000000c1000000c2000000bd000000b9000000b8000000a6",
            INIT_1E => X"000000a4000000ac000000b1000000b0000000aa000000890000008f0000007a",
            INIT_1F => X"0000006b0000006e000000600000006700000075000000760000007b0000007d",
            INIT_20 => X"0000009b000000950000009f000000a0000000ac000000ad000000b2000000b4",
            INIT_21 => X"000000bb000000ba000000ba000000bf000000bb000000af000000ac000000a0",
            INIT_22 => X"0000009a00000097000000a6000000b0000000b70000009b000000a600000085",
            INIT_23 => X"00000068000000680000007000000077000000760000007a0000007a0000007d",
            INIT_24 => X"0000009a0000009800000093000000a9000000b2000000b2000000b7000000aa",
            INIT_25 => X"000000b0000000bc000000c6000000c1000000ae000000a7000000a5000000a9",
            INIT_26 => X"0000009d0000008c00000092000000a9000000b3000000a0000000ab0000008d",
            INIT_27 => X"0000005f000000680000007500000077000000740000007b000000760000007d",
            INIT_28 => X"00000086000000700000009f000000b1000000ae000000b8000000b8000000ba",
            INIT_29 => X"000000ba000000c2000000bf000000b00000009b0000009e000000a7000000bb",
            INIT_2A => X"000000ae000000930000008600000097000000a00000009c0000009b0000007c",
            INIT_2B => X"0000004a0000006600000069000000660000006b000000750000007b0000007f",
            INIT_2C => X"000000410000005b000000ae0000009d00000093000000b1000000bf000000be",
            INIT_2D => X"000000bc000000b0000000ac000000b0000000b8000000ae00000094000000a3",
            INIT_2E => X"000000b00000009a000000850000009500000098000000950000008300000050",
            INIT_2F => X"000000420000006100000067000000660000006700000071000000780000007d",
            INIT_30 => X"000000150000005c000000bf000000b1000000bc000000ca000000bd000000b6",
            INIT_31 => X"000000b30000009c000000a5000000bc000000c8000000ae0000009800000072",
            INIT_32 => X"0000005f0000007f00000078000000890000009700000088000000720000004e",
            INIT_33 => X"0000004000000049000000590000006200000062000000710000007500000076",
            INIT_34 => X"0000002c00000063000000a8000000ad000000c8000000c3000000bc000000bb",
            INIT_35 => X"000000a500000095000000b4000000c2000000b9000000a8000000a80000009a",
            INIT_36 => X"0000006b00000092000000910000008a0000009c0000007f0000006400000048",
            INIT_37 => X"00000039000000400000005300000060000000620000006a0000006c0000006f",
            INIT_38 => X"0000006900000076000000750000009f000000c4000000be000000b4000000bb",
            INIT_39 => X"000000ad000000ad000000c6000000c1000000ab000000a5000000b4000000bc",
            INIT_3A => X"000000ae000000bb000000ad000000b3000000a0000000800000006900000048",
            INIT_3B => X"0000004300000045000000570000006c00000063000000640000006100000066",
            INIT_3C => X"0000008a00000071000000680000009d000000c6000000c4000000b4000000a8",
            INIT_3D => X"000000b4000000bf000000cb000000cd000000d2000000bf000000c4000000c8",
            INIT_3E => X"000000c0000000bb000000bc000000be000000a8000000990000007100000050",
            INIT_3F => X"00000046000000400000006000000087000000780000005a0000005a00000062",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY30;


    MEM_IFMAP_LAYER0_ENTITY31 : if BRAM_NAME = "ifmap_layer0_entity31" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000960000008a0000007300000093000000be000000bb000000b000000096",
            INIT_01 => X"000000ab000000c7000000d3000000c6000000d3000000c2000000be000000cb",
            INIT_02 => X"000000bf000000ba000000b8000000bd000000be000000a60000006400000046",
            INIT_03 => X"0000002f000000380000006a0000008f000000950000005c0000004a0000005e",
            INIT_04 => X"0000009b0000009b00000092000000a5000000bd000000c0000000bf00000091",
            INIT_05 => X"0000009c000000d2000000a900000095000000c0000000c2000000b2000000a8",
            INIT_06 => X"000000a9000000b5000000aa000000a70000009a00000075000000430000002b",
            INIT_07 => X"0000002200000031000000680000008f0000009c0000006a0000003f00000050",
            INIT_08 => X"000000a5000000a20000008a000000a6000000c4000000be000000ba00000089",
            INIT_09 => X"00000074000000c90000009d000000a9000000d2000000b6000000800000008f",
            INIT_0A => X"0000007c000000930000007f0000006100000052000000380000002f00000033",
            INIT_0B => X"0000002b00000040000000690000009d0000009d0000007b0000003900000041",
            INIT_0C => X"000000a900000096000000780000009e000000be000000be000000be00000098",
            INIT_0D => X"0000003c00000099000000bc000000b9000000c3000000a500000090000000ce",
            INIT_0E => X"000000b100000089000000650000003d00000037000000330000004700000050",
            INIT_0F => X"000000370000004a0000006e000000a0000000b00000008e0000003600000032",
            INIT_10 => X"000000aa000000a000000096000000a6000000ba000000bc000000ba0000009a",
            INIT_11 => X"00000020000000310000007e000000920000009b0000008c0000008c000000c0",
            INIT_12 => X"000000cc0000009c000000610000003e00000049000000490000005200000057",
            INIT_13 => X"0000003a0000003e0000006b000000a6000000bc000000a70000004800000033",
            INIT_14 => X"000000b2000000ab000000970000009c000000b5000000b2000000a30000007c",
            INIT_15 => X"000000240000001d00000028000000370000004e000000630000006500000082",
            INIT_16 => X"000000900000007b0000005f0000003700000034000000330000003c00000055",
            INIT_17 => X"0000004e0000004d0000006600000099000000bb000000b10000005900000037",
            INIT_18 => X"000000b5000000ab0000009200000098000000a9000000a70000009500000069",
            INIT_19 => X"0000004f0000005e000000420000002e0000002f000000470000005c00000078",
            INIT_1A => X"0000005a00000037000000380000002900000023000000220000001e00000037",
            INIT_1B => X"00000052000000560000006100000077000000ad000000ae0000006a0000003c",
            INIT_1C => X"000000b10000009c0000009e000000a30000009c000000a00000009400000089",
            INIT_1D => X"0000008f00000076000000660000006b0000006e0000006d0000007d00000067",
            INIT_1E => X"0000002f000000110000001000000013000000180000001c0000000e00000013",
            INIT_1F => X"0000002b0000004100000060000000630000008c000000ad0000008500000043",
            INIT_20 => X"0000009e0000008b000000a7000000b6000000970000008c000000ab000000c0",
            INIT_21 => X"000000ac000000740000008500000088000000920000008d0000007f00000065",
            INIT_22 => X"0000004100000025000000200000001900000018000000110000000a0000000f",
            INIT_23 => X"0000001400000042000000610000004e00000062000000940000009c00000069",
            INIT_24 => X"000000a0000000a4000000ae000000ab0000009e0000008800000094000000b1",
            INIT_25 => X"000000b800000093000000a9000000970000007f0000008b0000008e0000007d",
            INIT_26 => X"000000670000004d0000003f0000002b0000002100000018000000110000001a",
            INIT_27 => X"0000001f0000003e0000004800000032000000480000005a0000007800000088",
            INIT_28 => X"000000a0000000a3000000a7000000a7000000b1000000a80000008c00000078",
            INIT_29 => X"000000ab0000008f00000076000000820000007b0000009c000000a600000091",
            INIT_2A => X"0000007c000000690000005b0000004e0000004c000000420000003800000043",
            INIT_2B => X"00000046000000410000004100000049000000640000007b000000510000006a",
            INIT_2C => X"0000009c0000009f0000008c00000093000000b4000000aa000000990000007b",
            INIT_2D => X"0000008b0000009c000000730000007e000000830000009e000000a8000000a2",
            INIT_2E => X"0000007f000000770000007b0000007800000070000000680000006900000077",
            INIT_2F => X"0000007400000069000000680000006d0000007a000000860000005c00000068",
            INIT_30 => X"000000a40000009e0000007b0000008b000000ad0000009c0000008d0000008c",
            INIT_31 => X"0000008d0000007900000082000000a1000000970000009d000000a6000000a8",
            INIT_32 => X"000000900000008a0000008f0000008400000081000000850000008a00000094",
            INIT_33 => X"0000008f00000089000000860000008400000078000000640000007300000093",
            INIT_34 => X"0000008e0000009500000090000000a8000000a7000000a10000009e0000009e",
            INIT_35 => X"000000a50000009000000097000000a9000000a1000000a00000009e000000a2",
            INIT_36 => X"0000009900000091000000890000007f0000008d00000095000000960000009e",
            INIT_37 => X"0000009f00000096000000940000008f0000007b000000770000008b0000009f",
            INIT_38 => X"00000098000000a6000000b3000000b9000000a7000000a7000000aa000000a8",
            INIT_39 => X"000000a7000000a4000000ad000000b2000000a90000009d0000008900000085",
            INIT_3A => X"000000920000008f0000008c000000880000008c00000097000000980000009d",
            INIT_3B => X"000000a60000009c000000990000009000000085000000830000009000000099",
            INIT_3C => X"0000009f000000b2000000b7000000ab0000008b0000007d000000910000009f",
            INIT_3D => X"000000a20000008b000000950000009c0000009e000000980000008300000073",
            INIT_3E => X"000000840000008e000000940000008f000000900000009d0000009c000000a1",
            INIT_3F => X"000000a70000009f000000940000009c0000009c000000960000009900000098",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY31;


    MEM_IFMAP_LAYER0_ENTITY32 : if BRAM_NAME = "ifmap_layer0_entity32" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007600000060000000310000003b000000600000005f0000005400000053",
            INIT_01 => X"0000005f00000061000000530000005a0000005c000000520000004b0000004f",
            INIT_02 => X"0000005b000000500000003b0000003200000037000000380000003800000033",
            INIT_03 => X"0000003c00000038000000330000003a0000004c000000350000002f0000002f",
            INIT_04 => X"000000820000005800000059000000690000006c000000600000005d00000068",
            INIT_05 => X"00000065000000620000005a0000005b00000054000000570000004f00000048",
            INIT_06 => X"00000052000000480000003d0000003200000037000000380000003700000033",
            INIT_07 => X"0000002b0000002800000035000000410000004b0000003d0000003a00000039",
            INIT_08 => X"0000008400000068000000810000007a0000006c000000590000005f0000006a",
            INIT_09 => X"0000006200000069000000620000005e00000055000000500000004f0000004c",
            INIT_0A => X"000000550000004c000000360000002a000000330000003a0000003f00000042",
            INIT_0B => X"0000003c000000420000004300000042000000430000003e0000003800000039",
            INIT_0C => X"000000810000007f0000008800000084000000700000005a0000006800000069",
            INIT_0D => X"00000065000000710000006500000066000000670000005a000000570000005d",
            INIT_0E => X"0000004f0000004e000000330000001f0000002a00000033000000390000003e",
            INIT_0F => X"000000460000004d0000004b0000004a0000003c000000370000004300000045",
            INIT_10 => X"000000800000007f000000790000007f0000006d000000630000007200000072",
            INIT_11 => X"0000006f0000006f00000070000000710000006c00000063000000590000005c",
            INIT_12 => X"0000005e000000590000004e0000002c0000002700000034000000380000002e",
            INIT_13 => X"00000035000000430000004700000049000000420000003b0000004500000047",
            INIT_14 => X"0000008900000083000000680000007f000000760000006a0000007100000074",
            INIT_15 => X"000000730000007500000074000000710000006d000000690000005a00000054",
            INIT_16 => X"0000006a00000068000000670000004f0000003a0000004d000000520000003d",
            INIT_17 => X"0000003e0000003f00000043000000460000004900000048000000460000004b",
            INIT_18 => X"000000980000007700000066000000870000007a00000075000000730000006f",
            INIT_19 => X"000000790000007b0000007c000000700000007300000071000000660000005c",
            INIT_1A => X"00000064000000650000006d0000006e0000005c000000570000005b00000043",
            INIT_1B => X"0000003e00000040000000380000003b00000045000000480000004a0000004e",
            INIT_1C => X"0000009300000059000000780000007e00000078000000760000007200000079",
            INIT_1D => X"000000800000007a0000007c00000073000000730000006d0000006c00000064",
            INIT_1E => X"00000065000000680000006d0000006a000000660000004b0000005700000048",
            INIT_1F => X"0000003b0000003c0000002e000000350000004200000044000000490000004b",
            INIT_20 => X"000000760000006f000000780000007200000077000000740000007500000077",
            INIT_21 => X"000000800000007a0000006f0000006d0000007300000067000000610000005e",
            INIT_22 => X"0000005e0000005900000061000000640000006d0000005f0000007200000059",
            INIT_23 => X"0000003e0000003a00000040000000470000004600000048000000480000004b",
            INIT_24 => X"000000770000007100000069000000780000007c0000007a0000007b0000006f",
            INIT_25 => X"000000760000007b0000007d00000079000000760000006d000000650000006f",
            INIT_26 => X"000000690000005500000052000000600000006a000000640000007a00000067",
            INIT_27 => X"0000003d0000003e0000004700000049000000470000004b000000440000004b",
            INIT_28 => X"0000006400000048000000720000007e000000780000007f0000007c0000007e",
            INIT_29 => X"0000007f00000081000000800000007b00000079000000770000007800000090",
            INIT_2A => X"00000083000000630000004f000000580000005f000000610000006c0000005b",
            INIT_2B => X"0000002e0000003e0000003d0000003b0000004000000046000000490000004c",
            INIT_2C => X"00000022000000340000007f000000690000005d0000007a0000008400000083",
            INIT_2D => X"0000008100000073000000780000008c000000a6000000970000007400000085",
            INIT_2E => X"0000008d0000006e0000005600000061000000600000005c0000005600000031",
            INIT_2F => X"0000002a0000003c0000003e0000003c0000003e00000042000000450000004a",
            INIT_30 => X"00000004000000400000008e0000007d0000008c0000009a0000008c00000084",
            INIT_31 => X"0000007f0000006b0000007b0000009c000000b2000000930000007700000053",
            INIT_32 => X"000000400000005b00000053000000640000006f0000005c0000004d00000031",
            INIT_33 => X"000000290000002f00000037000000390000003b000000430000004200000044",
            INIT_34 => X"00000018000000480000007a0000007b0000009c000000960000008f0000008d",
            INIT_35 => X"000000770000006a0000008f000000a000000097000000810000008000000077",
            INIT_36 => X"0000004d00000074000000730000006d0000007b0000005a000000440000002d",
            INIT_37 => X"000000230000002b00000033000000370000003b0000003e0000003a0000003e",
            INIT_38 => X"00000045000000520000004a000000700000009600000091000000860000008f",
            INIT_39 => X"0000008300000084000000a10000009c0000007d000000720000008500000097",
            INIT_3A => X"00000091000000a00000009200000098000000810000005d0000004b0000002f",
            INIT_3B => X"0000002f0000003000000038000000440000003c0000003c0000003600000039",
            INIT_3C => X"00000057000000410000003b000000700000009800000096000000860000007d",
            INIT_3D => X"0000008f0000009b000000a7000000a50000009b000000840000008f000000a0",
            INIT_3E => X"000000a20000009e0000009f000000a100000089000000780000005400000039",
            INIT_3F => X"000000330000002b000000400000005f00000051000000370000003600000039",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY32;


    MEM_IFMAP_LAYER0_ENTITY33 : if BRAM_NAME = "ifmap_layer0_entity33" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000580000004e0000004000000066000000900000008d000000810000006c",
            INIT_01 => X"0000008b000000a5000000af0000009d0000009e00000086000000860000009f",
            INIT_02 => X"0000009a0000009400000093000000980000009a000000870000004900000031",
            INIT_03 => X"0000001e000000230000004b000000670000006f0000003d0000002c00000039",
            INIT_04 => X"000000560000005700000057000000740000008f000000930000009100000069",
            INIT_05 => X"00000080000000b3000000850000006c000000910000008b0000007a00000079",
            INIT_06 => X"0000007d000000870000007c0000007900000072000000580000002a00000018",
            INIT_07 => X"000000130000001d00000049000000660000007500000050000000270000002e",
            INIT_08 => X"0000005c0000005c0000004d000000760000009c000000990000009100000062",
            INIT_09 => X"0000005c000000aa000000740000007a000000a5000000830000004b00000062",
            INIT_0A => X"0000004c000000610000005500000040000000360000001b000000110000001b",
            INIT_0B => X"0000001a0000002800000045000000750000007f000000640000002400000028",
            INIT_0C => X"0000005e000000540000003c0000006e0000009c000000a30000009b00000073",
            INIT_0D => X"000000270000007c00000094000000890000009500000071000000570000009c",
            INIT_0E => X"00000078000000500000003d000000270000002700000018000000220000002e",
            INIT_0F => X"0000001f0000002d0000004500000078000000990000007b0000002200000020",
            INIT_10 => X"000000610000005d000000590000007200000096000000a20000009800000075",
            INIT_11 => X"0000000d0000001d00000064000000740000007300000056000000490000007c",
            INIT_12 => X"000000860000005b0000002f0000001b00000031000000320000003100000032",
            INIT_13 => X"000000190000001e000000420000007d000000a2000000960000003800000020",
            INIT_14 => X"0000006a0000006800000057000000630000008d000000960000008100000057",
            INIT_15 => X"0000000f0000000b00000016000000250000003600000039000000290000003e",
            INIT_16 => X"0000005300000048000000360000001a00000020000000230000002200000033",
            INIT_17 => X"000000280000002b0000003e000000700000009b0000009e0000004a0000001f",
            INIT_18 => X"00000070000000680000004f0000005a0000007b000000890000007300000042",
            INIT_19 => X"0000002f0000004200000028000000170000001b000000260000002c00000045",
            INIT_1A => X"000000360000001f000000260000001d00000019000000160000000f0000001f",
            INIT_1B => X"00000031000000330000003a0000004e0000008600000094000000570000001f",
            INIT_1C => X"0000006d0000005800000059000000600000006900000081000000730000005e",
            INIT_1D => X"0000006100000047000000360000003c000000420000003e0000004b0000003c",
            INIT_1E => X"0000001a0000000a000000090000000e00000011000000130000000b0000000c",
            INIT_1F => X"000000170000001f0000003a0000003b0000005e000000880000006900000023",
            INIT_20 => X"0000005b00000046000000600000007000000060000000680000008900000093",
            INIT_21 => X"000000750000003a00000045000000430000004a000000450000003f00000035",
            INIT_22 => X"0000002900000019000000130000000d0000000c000000090000000d00000012",
            INIT_23 => X"0000000c000000240000003e0000002700000034000000680000007900000047",
            INIT_24 => X"0000005b0000005c000000620000006200000061000000560000006900000086",
            INIT_25 => X"0000008e0000006b0000007c0000006100000044000000490000004e00000049",
            INIT_26 => X"0000003e0000002b000000260000001c000000160000000e0000000b00000014",
            INIT_27 => X"000000140000002a000000300000001400000025000000380000005800000064",
            INIT_28 => X"0000005b0000005e0000006100000062000000710000006f0000005b0000004c",
            INIT_29 => X"000000840000006e0000005000000051000000470000005f0000006300000054",
            INIT_2A => X"000000480000003d0000003800000033000000350000002b000000200000002b",
            INIT_2B => X"0000002e000000280000002500000028000000400000005a0000003000000042",
            INIT_2C => X"00000057000000600000005000000052000000710000006d0000006200000048",
            INIT_2D => X"0000005c0000007300000045000000460000004a0000005e0000006000000058",
            INIT_2E => X"00000045000000470000004c0000004a000000420000003c0000003d0000004b",
            INIT_2F => X"00000049000000400000003f000000410000004c0000005e000000360000003a",
            INIT_30 => X"0000006000000061000000430000004c000000690000005a0000004e00000050",
            INIT_31 => X"00000057000000480000004c00000062000000570000005c0000005d0000005a",
            INIT_32 => X"0000004f00000054000000550000004600000042000000480000004d00000057",
            INIT_33 => X"0000005300000052000000500000004f0000004300000035000000460000005e",
            INIT_34 => X"00000049000000540000005100000065000000610000005b000000580000005b",
            INIT_35 => X"00000069000000590000005b00000063000000590000005d0000005d0000005a",
            INIT_36 => X"0000005800000055000000490000003c0000004900000052000000540000005b",
            INIT_37 => X"0000005d00000056000000570000005500000043000000440000005700000064",
            INIT_38 => X"00000053000000600000006a00000071000000600000005f000000600000005f",
            INIT_39 => X"00000066000000690000006d000000680000005b0000005a000000520000004a",
            INIT_3A => X"000000520000004e0000004d0000004a0000004d00000055000000570000005c",
            INIT_3B => X"00000064000000590000005a000000540000004e0000004d000000570000005a",
            INIT_3C => X"0000005c0000006b000000710000006800000052000000420000004d0000005c",
            INIT_3D => X"0000005f000000510000005b0000005a000000580000005b0000004d0000003d",
            INIT_3E => X"000000460000004d0000005600000052000000530000005c0000005b00000060",
            INIT_3F => X"000000650000005c000000570000005b0000005c0000005a0000005b00000057",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY33;


    MEM_IFMAP_LAYER0_ENTITY34 : if BRAM_NAME = "ifmap_layer0_entity34" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000530000003d0000001a0000002400000041000000430000003a00000036",
            INIT_01 => X"0000003f00000041000000340000003b0000003e000000350000002e00000034",
            INIT_02 => X"00000047000000410000002b000000270000002f0000002f0000002d00000026",
            INIT_03 => X"0000002f0000002d0000002a00000032000000450000002e0000002900000029",
            INIT_04 => X"00000061000000350000003a000000460000004600000043000000440000004d",
            INIT_05 => X"000000440000004100000038000000390000003400000039000000320000002e",
            INIT_06 => X"0000003c000000340000002b000000260000002f0000002f0000002c00000028",
            INIT_07 => X"000000200000001e0000002b0000003800000043000000350000003300000031",
            INIT_08 => X"00000064000000470000005c000000510000004400000039000000440000004e",
            INIT_09 => X"00000040000000470000003f0000003b00000034000000300000003100000030",
            INIT_0A => X"0000003b00000032000000210000001e0000002b000000300000003500000038",
            INIT_0B => X"0000003300000038000000390000003800000039000000350000002f00000031",
            INIT_0C => X"000000600000005f000000610000005900000049000000370000004900000048",
            INIT_0D => X"000000410000004e00000042000000420000004300000037000000360000003f",
            INIT_0E => X"0000002f0000002e0000001a0000001200000022000000290000002f00000035",
            INIT_0F => X"0000003d00000044000000400000003e000000300000002d0000003a0000003c",
            INIT_10 => X"0000005c000000610000005400000057000000490000003f0000004c0000004b",
            INIT_11 => X"0000004a0000004a0000004b0000004b000000430000003b000000350000003b",
            INIT_12 => X"0000003b00000034000000330000001e0000001f000000290000002e00000027",
            INIT_13 => X"0000002e0000003b0000003d0000003d00000034000000300000003a0000003c",
            INIT_14 => X"0000006500000066000000470000005900000051000000460000004c0000004c",
            INIT_15 => X"0000004c000000510000004e0000004700000044000000430000003500000031",
            INIT_16 => X"000000430000004100000048000000390000002b0000003e0000004200000032",
            INIT_17 => X"0000003800000036000000380000003a0000003c0000003d0000003c00000041",
            INIT_18 => X"000000780000005900000049000000630000005300000050000000510000004b",
            INIT_19 => X"000000510000005700000055000000420000004c0000004f0000004300000035",
            INIT_1A => X"0000003c000000400000004a0000004d0000004100000040000000410000002f",
            INIT_1B => X"00000035000000360000002d000000300000003a0000003d0000003f00000042",
            INIT_1C => X"000000750000003b0000005b0000005b00000051000000510000004f00000054",
            INIT_1D => X"000000570000005600000056000000480000004d0000004c0000004a0000003f",
            INIT_1E => X"00000042000000490000004c00000049000000470000002f000000380000002f",
            INIT_1F => X"0000002c00000031000000230000002a00000037000000390000003e00000040",
            INIT_20 => X"0000005c000000540000005b00000051000000530000004f0000005000000050",
            INIT_21 => X"000000580000005300000049000000460000005100000048000000430000003d",
            INIT_22 => X"000000430000004100000046000000460000004f000000400000004f0000003c",
            INIT_23 => X"0000002c0000002d000000340000003b0000003a0000003d0000003d00000040",
            INIT_24 => X"00000061000000580000004c0000005a0000005b000000560000005300000047",
            INIT_25 => X"0000004f00000052000000540000005300000058000000530000004d00000055",
            INIT_26 => X"000000510000003e00000039000000460000005000000048000000590000004b",
            INIT_27 => X"0000002b000000310000003a0000003c0000003a0000003f0000003900000040",
            INIT_28 => X"00000051000000300000005600000062000000590000005b0000005200000054",
            INIT_29 => X"0000005b0000005400000050000000500000005e00000065000000670000007e",
            INIT_2A => X"0000006b0000004900000037000000430000004b0000004c0000005100000044",
            INIT_2B => X"00000020000000310000002f0000002d000000330000003a0000003e00000041",
            INIT_2C => X"000000140000001f000000630000004d00000040000000560000005a0000005a",
            INIT_2D => X"0000005f00000045000000450000005f0000008f000000880000006700000079",
            INIT_2E => X"00000076000000520000003f00000050000000520000004d0000004200000021",
            INIT_2F => X"0000002100000030000000300000002e00000030000000360000003b0000003f",
            INIT_30 => X"0000000000000032000000700000005c0000006e0000007a0000006900000062",
            INIT_31 => X"000000600000004800000054000000770000009d0000007d0000005f00000049",
            INIT_32 => X"00000034000000470000004100000054000000600000004f000000410000002a",
            INIT_33 => X"000000250000002500000029000000290000002d00000038000000390000003a",
            INIT_34 => X"000000140000003c000000610000005c0000007d00000078000000700000006f",
            INIT_35 => X"000000590000004c0000006e000000800000007f00000064000000620000006c",
            INIT_36 => X"0000004400000063000000620000005b0000006a0000004c0000003a00000029",
            INIT_37 => X"000000210000002300000025000000260000002e000000340000003200000035",
            INIT_38 => X"0000003b000000460000003a000000580000007b000000750000006a00000073",
            INIT_39 => X"0000006600000067000000820000007d0000005f000000500000006600000089",
            INIT_3A => X"000000830000008c0000007e000000840000006f0000004e000000400000002a",
            INIT_3B => X"0000002b000000280000002a000000320000002f000000320000002e00000031",
            INIT_3C => X"0000004900000035000000320000005e0000007e0000007c0000006c00000062",
            INIT_3D => X"000000720000007d0000008a000000880000007b00000062000000710000008c",
            INIT_3E => X"0000008f000000890000008a0000008c00000075000000690000004900000033",
            INIT_3F => X"0000002f00000023000000320000004d000000430000002d0000002d00000032",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY34;


    MEM_IFMAP_LAYER0_ENTITY35 : if BRAM_NAME = "ifmap_layer0_entity35" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000048000000410000003a0000005600000077000000750000006900000053",
            INIT_01 => X"0000006e000000890000009300000082000000820000006b0000006d00000087",
            INIT_02 => X"000000840000007f0000007e0000008300000087000000770000003d0000002a",
            INIT_03 => X"0000001a0000001b0000003c0000005500000061000000330000002400000033",
            INIT_04 => X"00000047000000480000005100000066000000780000007c0000007a00000050",
            INIT_05 => X"00000063000000970000006a000000540000007c00000079000000650000005c",
            INIT_06 => X"000000630000007300000068000000650000005e000000480000001f00000011",
            INIT_07 => X"0000000e000000150000003a0000005500000068000000460000001f00000029",
            INIT_08 => X"0000004f0000004e000000440000006400000086000000880000007d0000004b",
            INIT_09 => X"00000047000000930000005b000000610000008e000000710000003700000048",
            INIT_0A => X"000000350000004f00000045000000320000002a000000140000000d00000016",
            INIT_0B => X"000000140000002300000037000000600000006f0000005b0000001e00000023",
            INIT_0C => X"0000005100000048000000320000005800000087000000990000008a0000005d",
            INIT_0D => X"0000001f0000006f0000007f000000710000007c0000005c000000470000008d",
            INIT_0E => X"000000670000004100000033000000210000002400000019000000240000002c",
            INIT_0F => X"0000001a0000002b000000360000006000000089000000730000001e0000001a",
            INIT_10 => X"00000053000000520000004f0000005f00000082000000960000008600000062",
            INIT_11 => X"0000000a000000170000005600000063000000650000004c0000004200000074",
            INIT_12 => X"0000007a0000004e00000027000000170000002e0000002f0000002f0000002e",
            INIT_13 => X"000000140000001b000000340000006700000092000000890000002f00000019",
            INIT_14 => X"0000005c0000005c0000004e000000530000007b000000870000006e00000046",
            INIT_15 => X"0000000c00000008000000100000001d0000002f000000340000002500000038",
            INIT_16 => X"00000046000000390000002b00000012000000190000001c0000001d0000002c",
            INIT_17 => X"0000002100000026000000310000005e0000008c0000008d0000003d00000018",
            INIT_18 => X"000000610000005d000000460000004e0000006b000000760000006000000030",
            INIT_19 => X"000000250000003a0000002200000013000000130000001f000000260000003b",
            INIT_1A => X"00000027000000130000001b0000001200000011000000110000000a00000018",
            INIT_1B => X"0000002a0000002c000000300000004000000078000000800000004600000018",
            INIT_1C => X"0000005e0000004d00000052000000580000005b0000006b0000005f0000004b",
            INIT_1D => X"0000004a0000003700000030000000390000003a000000350000004300000033",
            INIT_1E => X"000000100000000400000003000000080000000e000000130000000700000006",
            INIT_1F => X"0000001100000017000000300000002f0000005100000073000000570000001b",
            INIT_20 => X"0000004b0000003b00000057000000690000005300000052000000750000007e",
            INIT_21 => X"0000005500000022000000390000003e000000420000003d000000390000002e",
            INIT_22 => X"0000002400000017000000120000000d0000000f0000000e0000000c0000000e",
            INIT_23 => X"000000070000001c000000360000001e0000002800000055000000680000003e",
            INIT_24 => X"0000004d0000004d000000510000005600000055000000450000005700000070",
            INIT_25 => X"0000006f0000004f000000640000004f0000003b00000043000000450000003a",
            INIT_26 => X"00000033000000260000002000000015000000110000000c000000060000000e",
            INIT_27 => X"0000000f00000022000000290000000f0000001f0000002e0000004c0000005a",
            INIT_28 => X"0000004f00000051000000520000005500000065000000600000004a00000039",
            INIT_29 => X"0000006d000000570000003a0000003e0000003d000000580000005a00000044",
            INIT_2A => X"0000003b000000350000002f0000002a0000002c000000230000001800000023",
            INIT_2B => X"000000260000001d0000001b0000001f00000039000000520000002700000038",
            INIT_2C => X"0000004c000000570000004a0000004a000000660000005f0000005300000039",
            INIT_2D => X"0000004d00000063000000370000003a0000003f00000054000000570000004d",
            INIT_2E => X"000000390000003c00000043000000440000003b00000031000000310000003f",
            INIT_2F => X"0000003c0000003100000030000000330000003f000000540000002d0000002f",
            INIT_30 => X"000000550000005a00000040000000450000005e0000004e0000004100000044",
            INIT_31 => X"0000004c0000003c000000420000005a0000004a0000004e0000005300000051",
            INIT_32 => X"00000043000000470000004c000000400000003b000000390000003e00000048",
            INIT_33 => X"0000004400000042000000400000003e00000032000000290000003d00000053",
            INIT_34 => X"0000003d0000004b000000490000005c00000057000000510000004e00000050",
            INIT_35 => X"0000005d0000004c00000050000000590000004a0000004c0000004e00000050",
            INIT_36 => X"0000004a000000450000003e000000350000004000000042000000440000004b",
            INIT_37 => X"0000004d00000048000000480000004400000032000000380000004e00000059",
            INIT_38 => X"00000046000000510000005a0000006400000056000000550000005700000055",
            INIT_39 => X"00000056000000570000005d0000005a0000004a000000460000003f0000003c",
            INIT_3A => X"000000420000003c0000003e0000003e0000004100000046000000470000004c",
            INIT_3B => X"000000550000004d0000004e000000470000003e000000410000004d0000004f",
            INIT_3C => X"0000004f0000005d0000005f0000005900000046000000390000004600000051",
            INIT_3D => X"000000530000004000000047000000470000004a0000004c0000003d0000002f",
            INIT_3E => X"000000380000003f0000004800000046000000450000004c0000004b00000050",
            INIT_3F => X"000000560000004f000000490000004e0000004f0000004c0000004f00000049",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY35;


    MEM_IFMAP_LAYER0_ENTITY36 : if BRAM_NAME = "ifmap_layer0_entity36" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a0000000b9000000d1000000d9000000e6000000f6000000f9000000f6",
            INIT_01 => X"000000f8000000f3000000e6000000dd000000da000000dd000000d8000000c7",
            INIT_02 => X"000000bc000000bb000000b8000000b4000000a600000090000000790000008b",
            INIT_03 => X"0000006a00000066000000660000004f0000005e000000650000005b0000005e",
            INIT_04 => X"000000e1000000ef000000f2000000e6000000e8000000f5000000f3000000eb",
            INIT_05 => X"000000ed000000e6000000d8000000cd000000c9000000cb000000c8000000ba",
            INIT_06 => X"000000af000000ab000000a10000007f0000008e0000008d0000007a00000087",
            INIT_07 => X"000000760000005200000025000000340000005f0000006b0000006100000064",
            INIT_08 => X"000000fc000000f9000000f1000000dc000000d9000000e2000000df000000d6",
            INIT_09 => X"000000d5000000cf000000c3000000b8000000b3000000b6000000b3000000a7",
            INIT_0A => X"0000009f000000980000009400000081000000800000008c0000008000000072",
            INIT_0B => X"0000005700000028000000040000002600000063000000730000006900000069",
            INIT_0C => X"000000e9000000e1000000de000000d3000000d3000000cb000000c8000000c0",
            INIT_0D => X"000000bb000000b7000000ae000000a4000000a0000000a5000000a000000099",
            INIT_0E => X"000000910000008d0000008c0000008a0000007d0000007d0000007f00000069",
            INIT_0F => X"0000003b000000250000001a000000370000007000000078000000700000006d",
            INIT_10 => X"000000cf000000c3000000cf000000c9000000be000000b4000000b3000000ab",
            INIT_11 => X"000000a30000009f00000099000000920000009100000097000000930000008d",
            INIT_12 => X"00000087000000880000008300000087000000810000007a000000840000005a",
            INIT_13 => X"0000003a0000003d00000030000000560000007500000078000000720000006d",
            INIT_14 => X"000000b6000000ab000000aa000000a2000000990000009c0000009f00000097",
            INIT_15 => X"000000900000008d0000008c0000008a0000008b0000008d0000008a0000008a",
            INIT_16 => X"000000870000008c000000860000008a0000008c000000890000006600000045",
            INIT_17 => X"0000004b0000003e00000043000000740000008100000080000000700000006e",
            INIT_18 => X"0000008d00000088000000880000008600000088000000860000008c00000085",
            INIT_19 => X"00000087000000890000008b0000008d0000008f000000920000008e00000091",
            INIT_1A => X"00000091000000910000008a0000008f0000008e0000006b0000002f00000021",
            INIT_1B => X"000000480000004b0000006c0000007f00000084000000840000006f00000070",
            INIT_1C => X"000000760000007d000000800000008100000088000000830000008a00000084",
            INIT_1D => X"000000880000008c0000009000000093000000960000009e0000009a00000099",
            INIT_1E => X"0000009200000095000000930000009400000080000000420000000d00000011",
            INIT_1F => X"0000005000000075000000800000007a0000007b000000800000007200000070",
            INIT_20 => X"000000730000007e00000084000000850000008b000000870000008f00000089",
            INIT_21 => X"0000008b000000910000009500000098000000940000009a000000a3000000aa",
            INIT_22 => X"0000009e000000a20000009d00000094000000730000002c0000000e0000001e",
            INIT_23 => X"000000690000008b000000880000007e000000770000007a000000740000006f",
            INIT_24 => X"000000760000008000000088000000880000008d00000088000000910000008d",
            INIT_25 => X"0000008d000000930000009a000000a50000009d0000009a000000a2000000a7",
            INIT_26 => X"0000009b00000093000000910000008a00000063000000380000002e00000037",
            INIT_27 => X"0000006d0000007c0000007a0000007e0000007300000074000000750000006e",
            INIT_28 => X"0000007d000000840000008b000000890000008e00000088000000900000008c",
            INIT_29 => X"0000008b000000900000009600000099000000830000008b0000009000000098",
            INIT_2A => X"000000a6000000ba000000d3000000d6000000800000005c000000450000002a",
            INIT_2B => X"000000550000005f0000006300000073000000700000006f000000710000006b",
            INIT_2C => X"00000085000000890000008e0000008a0000008d000000880000008e0000008a",
            INIT_2D => X"000000890000008f00000088000000840000008e000000b6000000c9000000cb",
            INIT_2E => X"000000d2000000ce000000cf000000c0000000a2000000bd000000920000002a",
            INIT_2F => X"0000001b0000002800000067000000720000006d0000006a0000006c00000068",
            INIT_30 => X"0000008c0000008b0000008f0000008b0000008f0000008c0000008a00000089",
            INIT_31 => X"000000870000008500000090000000a4000000ab000000a00000008900000073",
            INIT_32 => X"0000006a0000005d0000004b0000003b0000006f000000dc000000c90000005f",
            INIT_33 => X"0000000d000000070000003e0000007400000063000000650000006900000064",
            INIT_34 => X"000000900000008a0000008f0000008c00000092000000920000008200000087",
            INIT_35 => X"00000082000000910000008c0000006e0000005e0000005c0000003100000013",
            INIT_36 => X"0000001d00000032000000190000001200000078000000d1000000d20000009d",
            INIT_37 => X"000000260000000600000013000000440000004500000052000000630000005f",
            INIT_38 => X"000000910000008b000000920000008e000000900000008e0000007900000080",
            INIT_39 => X"000000850000007f000000540000004400000056000000520000002e00000016",
            INIT_3A => X"00000013000000320000001e00000041000000af000000c9000000cd000000cb",
            INIT_3B => X"0000006600000010000000120000001600000023000000380000004f00000058",
            INIT_3C => X"0000008f0000008b00000094000000900000008a000000840000008b00000083",
            INIT_3D => X"000000750000004200000048000000560000006a0000004e0000002800000022",
            INIT_3E => X"000000240000004600000073000000b6000000cb000000c5000000cd000000c3",
            INIT_3F => X"0000006c0000003d0000002500000012000000180000004f0000006400000053",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY36;


    MEM_IFMAP_LAYER0_ENTITY37 : if BRAM_NAME = "ifmap_layer0_entity37" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000008e0000008b000000930000009000000085000000720000008400000079",
            INIT_01 => X"00000051000000590000003c000000450000005500000044000000530000009b",
            INIT_02 => X"000000c0000000db000000ed000000eb000000d7000000d7000000d300000072",
            INIT_03 => X"000000300000005d0000003500000014000000410000008b0000008f00000054",
            INIT_04 => X"0000008f0000008d0000008e0000008900000074000000450000003a00000043",
            INIT_05 => X"000000510000004b0000001d0000001c00000024000000190000008c000000f2",
            INIT_06 => X"000000ec000000eb000000e3000000dc000000db000000df000000950000003a",
            INIT_07 => X"00000039000000540000004e0000004e00000085000000a1000000a70000005b",
            INIT_08 => X"0000008f0000008c00000088000000860000008d000000470000002d00000034",
            INIT_09 => X"000000430000002100000017000000160000002f000000290000009b000000d9",
            INIT_0A => X"000000c7000000be000000bf000000d0000000dc000000df000000ad00000067",
            INIT_0B => X"0000005d0000007300000087000000950000009800000094000000a500000059",
            INIT_0C => X"0000008f0000008c0000007e000000b5000000bd0000004c000000210000002b",
            INIT_0D => X"0000003900000015000000100000001700000039000000420000009e000000c2",
            INIT_0E => X"000000b6000000b3000000c4000000c9000000c2000000ce000000de000000b3",
            INIT_0F => X"000000970000009c000000950000009700000096000000920000008800000042",
            INIT_10 => X"0000008c000000850000009a000000ea000000b50000005a000000260000002a",
            INIT_11 => X"000000340000000b0000000b0000000b0000001400000031000000a0000000ba",
            INIT_12 => X"000000b0000000b9000000b900000073000000450000005a000000a1000000c4",
            INIT_13 => X"000000b7000000aa000000a00000009900000093000000880000004d00000026",
            INIT_14 => X"0000008200000080000000a3000000a30000008b0000006a0000002d0000002e",
            INIT_15 => X"0000001c00000003000000090000000f0000001e00000036000000a2000000b4",
            INIT_16 => X"000000ac000000be000000710000001500000014000000150000003000000095",
            INIT_17 => X"000000bb000000ab0000008e0000008500000080000000430000001500000027",
            INIT_18 => X"0000007c00000084000000670000001a000000480000006c0000003400000030",
            INIT_19 => X"00000012000000070000000b0000003b0000005a00000063000000a5000000b0",
            INIT_1A => X"000000b1000000a90000002a0000001d0000002f000000260000000e00000046",
            INIT_1B => X"000000950000008800000075000000750000003c0000000e0000001500000030",
            INIT_1C => X"000000790000007c000000490000001e0000003b00000072000000440000001f",
            INIT_1D => X"0000000d0000000e00000018000000480000004f0000006c000000bb000000bb",
            INIT_1E => X"000000bf0000008b0000001b0000002b0000001e0000001b0000001c0000001b",
            INIT_1F => X"0000006c000000840000007b0000005900000016000000150000002a0000003b",
            INIT_20 => X"0000006d00000066000000470000003f0000003c000000710000004d0000001c",
            INIT_21 => X"000000100000001f00000030000000470000004600000088000000bd000000b3",
            INIT_22 => X"000000b4000000740000001f0000003600000035000000290000001b0000000e",
            INIT_23 => X"00000048000000850000007c0000003c0000001200000022000000320000003b",
            INIT_24 => X"00000057000000510000003d0000003c0000003a000000690000004b00000015",
            INIT_25 => X"000000140000002e0000004c000000600000006100000091000000a4000000a3",
            INIT_26 => X"000000aa00000071000000200000003900000047000000310000002500000011",
            INIT_27 => X"000000290000006c00000060000000210000000c0000001d0000002800000032",
            INIT_28 => X"0000004900000049000000400000003c000000390000005f000000570000002f",
            INIT_29 => X"0000003d0000006200000089000000a5000000a9000000b0000000b7000000b6",
            INIT_2A => X"000000b60000007c0000002200000036000000600000005c000000330000001b",
            INIT_2B => X"00000011000000460000003b0000000c00000006000000120000001d00000028",
            INIT_2C => X"0000004900000049000000450000004e0000004100000059000000450000002f",
            INIT_2D => X"000000340000003c0000004a000000560000005b000000600000006200000060",
            INIT_2E => X"0000006200000053000000200000003c0000003b0000003e0000001d00000014",
            INIT_2F => X"00000004000000110000000a00000003000000070000000a0000001100000021",
            INIT_30 => X"0000004b0000005300000048000000360000002d000000270000000f00000004",
            INIT_31 => X"0000000300000002000000050000000700000007000000080000000a0000000b",
            INIT_32 => X"0000000b0000000d0000000800000042000000430000002f000000380000000f",
            INIT_33 => X"00000002000000020000000100000003000000060000000a0000000f00000020",
            INIT_34 => X"0000005000000059000000510000002f000000150000000a0000001000000019",
            INIT_35 => X"0000000e0000000a0000000e0000000e0000000e0000000e0000000e0000000c",
            INIT_36 => X"0000000a0000000900000006000000170000003e000000480000002a00000007",
            INIT_37 => X"00000003000000040000000500000005000000070000000b0000001500000021",
            INIT_38 => X"000000490000004f00000049000000370000002e0000002f0000003b0000003a",
            INIT_39 => X"0000001a00000011000000190000001c0000001f000000200000001d0000001c",
            INIT_3A => X"0000001800000015000000100000000c00000014000000160000000800000006",
            INIT_3B => X"000000080000000700000008000000080000000b0000000f0000001b0000001f",
            INIT_3C => X"00000045000000480000004c0000004e00000058000000530000004800000038",
            INIT_3D => X"00000020000000260000002b0000002a0000002f000000330000003200000031",
            INIT_3E => X"0000002c000000260000001e0000001c0000002200000022000000130000000c",
            INIT_3F => X"0000000e000000100000000f0000000d000000120000001a0000001e0000001d",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY37;


    MEM_IFMAP_LAYER0_ENTITY38 : if BRAM_NAME = "ifmap_layer0_entity38" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002500000031000000390000003a000000420000004e0000005000000051",
            INIT_01 => X"0000005600000052000000490000004200000041000000430000004300000038",
            INIT_02 => X"0000003200000032000000400000007300000034000000380000003200000027",
            INIT_03 => X"00000016000000220000002e000000240000001d000000120000001500000013",
            INIT_04 => X"00000043000000480000004d00000044000000430000004a0000004800000042",
            INIT_05 => X"000000440000004000000039000000340000003200000036000000370000002e",
            INIT_06 => X"000000290000002a000000270000002900000028000000230000001e00000021",
            INIT_07 => X"000000220000002e0000001e0000001b0000001c000000150000001600000012",
            INIT_08 => X"0000004800000044000000480000003e0000003a0000003d0000003800000031",
            INIT_09 => X"000000300000002d0000002b00000028000000260000002a0000002b00000026",
            INIT_0A => X"00000022000000230000001e0000001c00000023000000210000001f00000022",
            INIT_0B => X"00000030000000220000000d0000000e00000015000000140000001300000011",
            INIT_0C => X"00000038000000360000003d0000003c0000003e000000300000002b00000024",
            INIT_0D => X"000000230000002300000022000000200000001f000000210000002200000020",
            INIT_0E => X"0000001d0000001e0000001b0000001d000000200000001c0000001d00000025",
            INIT_0F => X"0000002a000000120000000b0000000f00000016000000130000001000000011",
            INIT_10 => X"0000003900000039000000420000003b0000003400000024000000200000001b",
            INIT_11 => X"0000001c0000001d0000001c0000001a0000001a0000001a0000001c0000001e",
            INIT_12 => X"0000001c0000001c0000001c0000001c0000001c00000030000000430000002a",
            INIT_13 => X"00000019000000120000000d000000190000001b0000001f0000001300000011",
            INIT_14 => X"0000003b0000003a0000002f000000210000001a0000001a0000001900000016",
            INIT_15 => X"00000017000000190000001a0000001900000018000000180000001b0000001f",
            INIT_16 => X"0000001d0000001e000000210000001e000000210000005d0000005e0000003c",
            INIT_17 => X"000000290000001b0000001e0000002c0000002b0000002d0000001800000013",
            INIT_18 => X"000000220000001c000000170000001400000016000000170000001600000015",
            INIT_19 => X"0000001600000016000000190000001a00000018000000190000001d00000023",
            INIT_1A => X"000000200000001f000000230000001e00000033000000590000003700000025",
            INIT_1B => X"00000038000000280000002b0000002d000000240000001e0000001700000015",
            INIT_1C => X"0000001100000011000000100000001200000016000000170000001600000016",
            INIT_1D => X"00000018000000170000001a0000001b000000190000001b0000001d00000027",
            INIT_1E => X"000000280000002d00000033000000300000004100000040000000120000000b",
            INIT_1F => X"00000022000000250000001f0000002000000019000000160000001600000015",
            INIT_20 => X"0000001100000012000000120000001200000015000000160000001700000017",
            INIT_21 => X"00000019000000180000001c0000001e0000002500000038000000330000003b",
            INIT_22 => X"0000003b0000003a00000037000000360000003d000000280000001100000010",
            INIT_23 => X"0000001a00000019000000180000001b0000001a000000170000001500000014",
            INIT_24 => X"0000001300000012000000120000001200000015000000140000001600000018",
            INIT_25 => X"000000180000001900000020000000310000003e0000004c0000003900000034",
            INIT_26 => X"000000310000002e000000320000003a0000003800000031000000300000002c",
            INIT_27 => X"0000002900000023000000190000001900000019000000180000001400000014",
            INIT_28 => X"0000001400000012000000130000001200000015000000150000001500000017",
            INIT_29 => X"0000001900000019000000240000003500000031000000420000003e0000004a",
            INIT_2A => X"0000006800000089000000a6000000b80000007c000000680000004b00000021",
            INIT_2B => X"000000380000003d000000260000001900000018000000190000001200000013",
            INIT_2C => X"0000001500000012000000140000001300000018000000180000001600000018",
            INIT_2D => X"000000190000001d0000001f000000300000005500000097000000b2000000be",
            INIT_2E => X"000000cd000000cd000000ca000000c5000000b2000000d00000009800000016",
            INIT_2F => X"0000001800000025000000460000002800000015000000160000001100000011",
            INIT_30 => X"000000140000001400000016000000150000001800000018000000190000001a",
            INIT_31 => X"00000019000000200000004200000070000000900000009b0000008c00000075",
            INIT_32 => X"0000006400000058000000470000003d00000075000000e8000000d50000004e",
            INIT_33 => X"0000000f0000000a00000032000000460000001a000000150000001100000010",
            INIT_34 => X"000000140000001600000019000000160000001700000017000000190000001a",
            INIT_35 => X"0000001a00000048000000670000005b00000050000000560000003400000012",
            INIT_36 => X"00000011000000220000000f000000100000007c000000dd000000e00000009b",
            INIT_37 => X"0000002400000007000000160000003b00000021000000130000001200000010",
            INIT_38 => X"00000018000000170000001b0000001600000018000000190000001300000015",
            INIT_39 => X"00000037000000550000003a000000290000003d0000004e0000003200000018",
            INIT_3A => X"0000000b0000002b0000001e00000049000000bf000000d8000000d1000000cd",
            INIT_3B => X"000000670000000e00000010000000170000001b000000160000001400000012",
            INIT_3C => X"0000001a000000160000001a0000001700000019000000250000003c00000034",
            INIT_3D => X"0000004c00000034000000380000003b000000500000004d0000002e00000026",
            INIT_3E => X"00000023000000490000007c000000c4000000df000000d8000000d9000000d2",
            INIT_3F => X"0000007600000039000000150000000e0000001f000000470000003e00000011",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY38;


    MEM_IFMAP_LAYER0_ENTITY39 : if BRAM_NAME = "ifmap_layer0_entity39" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000190000001400000019000000170000002100000035000000600000005c",
            INIT_01 => X"000000490000005d0000003e0000004200000051000000470000005a000000a2",
            INIT_02 => X"000000c4000000df000000f5000000f5000000e3000000e4000000de00000079",
            INIT_03 => X"000000250000003b0000001100000009000000480000008c0000007500000013",
            INIT_04 => X"0000001900000015000000180000001a000000280000002c0000003500000045",
            INIT_05 => X"00000058000000520000002500000029000000310000002000000094000000fb",
            INIT_06 => X"000000f6000000f2000000e9000000e2000000e1000000e20000008b0000001f",
            INIT_07 => X"0000000b00000019000000280000004300000085000000a20000009700000022",
            INIT_08 => X"000000160000001300000016000000260000005d000000460000002e00000036",
            INIT_09 => X"0000004b00000026000000180000001b0000003800000031000000a3000000e3",
            INIT_0A => X"000000d6000000cd000000cb000000da000000e5000000e4000000a30000004a",
            INIT_0B => X"000000390000005a00000080000000950000009700000096000000a000000033",
            INIT_0C => X"000000130000000f000000260000007c000000af0000005a000000240000002a",
            INIT_0D => X"0000003f000000170000000b00000015000000400000004f000000aa000000d0",
            INIT_0E => X"000000c7000000c5000000d3000000d6000000ce000000d9000000e3000000b1",
            INIT_0F => X"00000098000000a8000000a7000000a20000009a00000097000000880000002a",
            INIT_10 => X"000000120000000a00000065000000dc000000be0000006f0000002f0000002e",
            INIT_11 => X"000000390000000a000000090000000e0000001f00000042000000b1000000cc",
            INIT_12 => X"000000c2000000ca000000c60000007c0000004f00000066000000ac000000d3",
            INIT_13 => X"000000c8000000b8000000b1000000a90000009c0000008c0000004a00000011",
            INIT_14 => X"0000000e0000001400000084000000a500000096000000800000003700000034",
            INIT_15 => X"0000001e000000030000000a000000160000002d00000048000000b4000000c6",
            INIT_16 => X"000000be000000cd0000007b000000190000001a0000001e00000038000000a3",
            INIT_17 => X"000000ca000000b80000009e0000009300000088000000440000000d00000011",
            INIT_18 => X"0000000a00000023000000530000002100000053000000820000003e00000035",
            INIT_19 => X"000000130000000700000010000000480000006c00000075000000b7000000c2",
            INIT_1A => X"000000c3000000b70000002f0000001e000000310000002b000000140000004f",
            INIT_1B => X"000000a1000000940000008400000081000000400000000a0000000900000018",
            INIT_1C => X"0000000a00000021000000370000002300000046000000880000004e00000024",
            INIT_1D => X"0000000f000000110000002200000058000000610000007e000000cd000000cd",
            INIT_1E => X"000000d000000098000000200000002b000000200000001f000000200000001f",
            INIT_1F => X"00000075000000910000008a00000063000000170000000c0000001900000021",
            INIT_20 => X"0000000a00000015000000360000004100000047000000880000005700000021",
            INIT_21 => X"00000015000000270000003f00000057000000560000009a000000cf000000c5",
            INIT_22 => X"000000c6000000810000002500000038000000370000002c0000001c0000000f",
            INIT_23 => X"0000004d000000930000008b000000430000000e000000140000001c0000001f",
            INIT_24 => X"000000070000000e0000002f0000003e0000004500000080000000560000001c",
            INIT_25 => X"0000001e0000003c0000005e0000006f0000006f000000a2000000b6000000b4",
            INIT_26 => X"000000bc0000007f000000290000003c0000004b00000035000000230000000f",
            INIT_27 => X"0000002c0000007a0000006f00000026000000070000000d0000001000000016",
            INIT_28 => X"0000000b00000011000000270000003b0000004600000075000000680000003d",
            INIT_29 => X"00000051000000790000009f000000b7000000b9000000c3000000c9000000c7",
            INIT_2A => X"000000c6000000880000002a0000003c0000006600000062000000340000001c",
            INIT_2B => X"000000150000004f000000450000001000000003000000070000000c00000016",
            INIT_2C => X"00000013000000140000001d000000430000004900000067000000550000003c",
            INIT_2D => X"00000045000000500000005b000000640000006800000071000000710000006d",
            INIT_2E => X"0000006d00000059000000250000004100000040000000420000001f00000017",
            INIT_2F => X"00000008000000140000000e0000000500000006000000060000000b00000018",
            INIT_30 => X"000000170000001c0000001d000000250000002c0000002c0000001600000007",
            INIT_31 => X"0000000a0000000a0000000c0000000c0000000d000000100000001100000010",
            INIT_32 => X"0000000f0000000f000000090000004300000044000000300000003800000010",
            INIT_33 => X"0000000400000003000000030000000400000006000000090000000e00000019",
            INIT_34 => X"0000002100000025000000270000002000000017000000120000001900000020",
            INIT_35 => X"000000170000001500000017000000170000001700000015000000130000000f",
            INIT_36 => X"0000000b0000000a00000007000000180000003e000000470000002900000008",
            INIT_37 => X"00000004000000050000000500000006000000090000000e000000180000001d",
            INIT_38 => X"000000230000002500000029000000320000003c00000043000000510000004d",
            INIT_39 => X"0000002c000000240000002d00000030000000310000002c0000002700000023",
            INIT_3A => X"0000001d0000001b000000150000001000000017000000190000000a00000009",
            INIT_3B => X"0000000b000000090000000a0000000b0000000e000000140000001f0000001e",
            INIT_3C => X"0000002a0000002a0000003b000000570000006d0000006f0000006600000052",
            INIT_3D => X"000000370000003e00000045000000470000004a000000480000004600000043",
            INIT_3E => X"0000003b000000330000002b000000290000002f0000002c0000001800000012",
            INIT_3F => X"00000014000000160000001500000013000000160000001c000000200000001e",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY39;


    MEM_IFMAP_LAYER0_ENTITY40 : if BRAM_NAME = "ifmap_layer0_entity40" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000d0000000b0000000e0000000a000000090000000a0000000500000002",
            INIT_01 => X"0000000300000003000000010000000200000004000000060000000500000000",
            INIT_02 => X"0000000100000000000000230000005600000016000000170000001d00000008",
            INIT_03 => X"0000000d0000001b000000270000001d00000013000000080000000600000005",
            INIT_04 => X"0000000d0000000c0000000a0000000400000007000000080000000300000000",
            INIT_05 => X"0000000400000002000000010000000100000002000000040000000400000001",
            INIT_06 => X"0000000100000001000000100000001300000007000000060000000600000007",
            INIT_07 => X"000000210000002e000000170000001600000013000000080000000400000006",
            INIT_08 => X"0000000700000004000000030000000000000004000000040000000100000000",
            INIT_09 => X"0000000400000004000000040000000400000004000000060000000500000003",
            INIT_0A => X"00000004000000030000000c000000090000000400000007000000060000000a",
            INIT_0B => X"00000028000000230000000d0000000c0000000f000000060000000300000006",
            INIT_0C => X"0000000100000003000000080000000b00000012000000040000000300000003",
            INIT_0D => X"0000000500000006000000080000000700000008000000090000000600000006",
            INIT_0E => X"00000007000000050000000a00000009000000040000000a0000001000000017",
            INIT_0F => X"0000001e00000016000000110000000e0000000f000000060000000500000008",
            INIT_10 => X"0000000c000000130000001d0000001a00000017000000060000000700000008",
            INIT_11 => X"00000007000000080000000900000008000000090000000a0000000700000008",
            INIT_12 => X"0000000900000007000000080000000700000008000000250000004000000027",
            INIT_13 => X"00000010000000100000000e000000150000000e0000000f0000000d00000009",
            INIT_14 => X"000000180000001e000000160000000c00000009000000060000000900000008",
            INIT_15 => X"0000000500000005000000090000000a0000000b0000000a0000000700000009",
            INIT_16 => X"0000000a0000000b0000000b0000000700000014000000550000005d0000003b",
            INIT_17 => X"000000220000000e0000001300000020000000170000001b0000001000000009",
            INIT_18 => X"0000000c0000000b0000000a0000000700000008000000080000000a00000007",
            INIT_19 => X"00000006000000050000000a0000000e0000000d0000000c0000000a0000000c",
            INIT_1A => X"000000090000000e0000000e0000000700000025000000560000003c00000028",
            INIT_1B => X"000000350000001c0000001c0000001c00000014000000100000000600000007",
            INIT_1C => X"000000030000000600000006000000070000000b0000000a0000000c00000009",
            INIT_1D => X"00000009000000080000000c0000000e0000000e000000120000001000000013",
            INIT_1E => X"00000010000000150000001a00000016000000310000003e000000140000000a",
            INIT_1F => X"0000001e0000001a000000100000000d00000009000000080000000400000007",
            INIT_20 => X"000000070000000a00000009000000080000000b0000000a0000000e0000000b",
            INIT_21 => X"0000000d0000000c0000000e0000000f00000013000000240000002200000028",
            INIT_22 => X"00000024000000200000002200000022000000330000002b0000000f00000009",
            INIT_23 => X"000000140000000c000000090000000a00000008000000080000000800000008",
            INIT_24 => X"0000000c0000000c0000000b000000080000000c0000000a0000000e0000000d",
            INIT_25 => X"0000000e0000000e000000140000002200000027000000310000002800000026",
            INIT_26 => X"000000200000001b0000002700000032000000360000003b0000003400000026",
            INIT_27 => X"00000023000000150000000b0000000c00000006000000090000000b0000000a",
            INIT_28 => X"0000000c0000000b0000000b000000090000000c0000000a0000000d0000000d",
            INIT_29 => X"0000000d000000100000001b000000280000002000000032000000320000003f",
            INIT_2A => X"0000005800000077000000a1000000b400000079000000710000005400000022",
            INIT_2B => X"00000032000000310000001d00000011000000090000000a0000000c0000000a",
            INIT_2C => X"000000090000000a0000000e0000000b0000000e0000000c0000000d0000000c",
            INIT_2D => X"0000000c0000001200000018000000270000004d00000093000000af000000ba",
            INIT_2E => X"000000c8000000c8000000d2000000ca000000b1000000d50000009e0000001c",
            INIT_2F => X"000000130000002200000046000000250000000a000000090000000b00000009",
            INIT_30 => X"000000080000000a0000000f0000000d000000100000000e0000000d0000000e",
            INIT_31 => X"0000000c000000180000003e0000006c0000008e000000a2000000930000007d",
            INIT_32 => X"0000006e0000005e000000540000004a0000007e000000f1000000d700000054",
            INIT_33 => X"0000000c000000090000003400000049000000190000000d0000000900000008",
            INIT_34 => X"0000000b0000000b0000000f0000000e00000011000000100000000c0000000e",
            INIT_35 => X"0000001400000044000000670000005d000000560000005f0000003d00000019",
            INIT_36 => X"0000001600000023000000110000001700000089000000eb000000eb000000a7",
            INIT_37 => X"0000002a00000007000000170000004200000028000000110000000900000007",
            INIT_38 => X"0000000f0000000d000000120000000e00000010000000120000000b00000012",
            INIT_39 => X"00000036000000530000003b0000002e0000004400000053000000370000001b",
            INIT_3A => X"0000000c000000270000001c0000004c000000c8000000e8000000e7000000e0",
            INIT_3B => X"0000007300000016000000130000001a0000001f000000160000000d00000008",
            INIT_3C => X"000000100000000d000000130000000e0000000e0000001e0000003900000037",
            INIT_3D => X"0000004f00000035000000390000003c000000520000004e0000003200000029",
            INIT_3E => X"00000023000000470000007c000000c8000000e7000000e6000000ec000000dd",
            INIT_3F => X"0000007e000000440000001a0000000e00000020000000490000003f00000009",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY40;


    MEM_IFMAP_LAYER0_ENTITY41 : if BRAM_NAME = "ifmap_layer0_entity41" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000110000000e0000001300000011000000180000002f0000005d0000005c",
            INIT_01 => X"0000004f000000620000003c0000003d0000004c000000470000005e000000a6",
            INIT_02 => X"000000c6000000e2000000fa000000fc000000ed000000f0000000e70000007c",
            INIT_03 => X"0000002a0000004a0000001c0000000c0000004c000000950000007e00000011",
            INIT_04 => X"00000012000000100000001200000015000000240000002a0000003800000048",
            INIT_05 => X"000000600000005800000024000000240000002d000000220000009a00000100",
            INIT_06 => X"000000fa000000f9000000f4000000ed000000ed000000ee0000009600000027",
            INIT_07 => X"000000150000002e0000003b0000004d0000008e000000ae000000a300000026",
            INIT_08 => X"000000110000001000000010000000220000005c000000490000003c00000042",
            INIT_09 => X"000000540000002c0000001c000000210000003e00000037000000ae000000f0",
            INIT_0A => X"000000e1000000d9000000d9000000e7000000ef000000ee000000b100000056",
            INIT_0B => X"000000450000006a00000092000000a4000000a4000000a1000000a900000037",
            INIT_0C => X"0000000d0000000a000000200000007d000000b4000000620000003500000038",
            INIT_0D => X"000000480000001c0000000e0000001b0000004900000059000000b9000000e0",
            INIT_0E => X"000000d5000000d5000000e4000000e3000000d7000000e1000000f2000000c0",
            INIT_0F => X"000000a5000000b4000000b5000000b0000000a60000009f0000008d0000002a",
            INIT_10 => X"0000000c0000000700000065000000e5000000c90000007b0000003e00000039",
            INIT_11 => X"000000410000000f000000090000000f000000260000004f000000bf000000da",
            INIT_12 => X"000000d0000000db000000d80000008a000000580000006d000000b8000000e4",
            INIT_13 => X"000000da000000c9000000bf000000b5000000a6000000930000004d0000000e",
            INIT_14 => X"0000000d000000180000008b000000b3000000a20000008d000000450000003d",
            INIT_15 => X"00000023000000040000000b0000001b0000003600000056000000c2000000d4",
            INIT_16 => X"000000cc000000db0000008800000024000000200000002200000040000000b1",
            INIT_17 => X"000000dd000000cc000000ad0000009f00000090000000490000000f0000000d",
            INIT_18 => X"00000009000000270000005b00000031000000600000008f0000004c0000003e",
            INIT_19 => X"000000150000000700000015000000510000007900000083000000c5000000d0",
            INIT_1A => X"000000d1000000c10000003800000026000000370000002e0000001900000059",
            INIT_1B => X"000000b2000000a9000000950000008d000000480000000e0000000800000014",
            INIT_1C => X"00000005000000220000003b0000003000000053000000950000005c0000002d",
            INIT_1D => X"0000000f000000130000002a000000640000006f0000008c000000db000000db",
            INIT_1E => X"000000de000000a0000000260000003300000025000000230000002400000027",
            INIT_1F => X"00000082000000a40000009b0000006e0000001d0000000c000000160000001e",
            INIT_20 => X"00000007000000170000003a0000004d0000005400000094000000650000002a",
            INIT_21 => X"000000160000002b0000004a0000006500000064000000a8000000dd000000d3",
            INIT_22 => X"000000d4000000890000002b000000400000003f000000340000002300000015",
            INIT_23 => X"00000056000000a20000009a0000004e0000001300000012000000180000001c",
            INIT_24 => X"0000000900000015000000370000004c000000520000008c0000006500000025",
            INIT_25 => X"00000021000000430000006c0000007f0000007e000000b0000000c3000000c2",
            INIT_26 => X"000000c900000087000000300000004600000056000000410000002e00000015",
            INIT_27 => X"00000032000000830000007b000000310000000b0000000a0000000b00000014",
            INIT_28 => X"0000000b0000001700000031000000490000005700000084000000780000004b",
            INIT_29 => X"0000005d00000086000000b1000000c8000000c8000000cf000000d4000000d5",
            INIT_2A => X"000000d6000000940000003500000048000000710000006e0000004000000022",
            INIT_2B => X"00000018000000550000004c0000001600000007000000090000000d00000016",
            INIT_2C => X"0000000f00000016000000250000004e00000057000000730000006000000048",
            INIT_2D => X"000000520000005d0000006900000072000000770000007d0000007e0000007b",
            INIT_2E => X"0000007c00000066000000300000004c0000004b0000004e000000290000001b",
            INIT_2F => X"00000009000000180000001000000006000000080000000a0000000f00000019",
            INIT_30 => X"000000150000001f000000230000002b0000003200000030000000190000000c",
            INIT_31 => X"0000000e0000000e000000110000001100000014000000180000001a00000019",
            INIT_32 => X"00000018000000140000000d0000004a0000004e0000003b0000004100000012",
            INIT_33 => X"0000000300000005000000040000000300000005000000090000000d0000001a",
            INIT_34 => X"00000021000000280000002c000000250000001e000000170000001e00000025",
            INIT_35 => X"0000001c000000190000001c0000001c0000001b000000180000001700000013",
            INIT_36 => X"0000000f00000009000000060000001c00000047000000530000002f00000008",
            INIT_37 => X"00000002000000050000000500000004000000060000000b000000150000001c",
            INIT_38 => X"0000002500000029000000300000003b000000490000004f0000005c00000059",
            INIT_39 => X"000000380000002f000000380000003b00000039000000300000002b00000028",
            INIT_3A => X"000000230000001b000000150000001500000021000000250000001000000008",
            INIT_3B => X"00000008000000090000000a0000000a0000000d000000120000001d0000001c",
            INIT_3C => X"0000002c00000031000000460000006500000080000000800000007600000063",
            INIT_3D => X"000000470000004e00000054000000550000005700000053000000510000004f",
            INIT_3E => X"000000470000003c00000031000000310000003a000000380000002000000013",
            INIT_3F => X"00000013000000180000001800000015000000190000001f000000220000001c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY41;


    MEM_IFMAP_LAYER0_ENTITY42 : if BRAM_NAME = "ifmap_layer0_entity42" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005300000052000000510000004d00000051000000550000005b0000005c",
            INIT_01 => X"0000005c0000005f000000650000005c0000005700000052000000500000004c",
            INIT_02 => X"00000044000000410000003f0000003e0000003c00000038000000340000002f",
            INIT_03 => X"0000002a000000250000002300000022000000240000001d0000001900000015",
            INIT_04 => X"0000005400000053000000530000004d00000050000000540000005a0000005d",
            INIT_05 => X"0000005a000000580000005f0000006100000058000000520000004e0000004c",
            INIT_06 => X"000000470000004400000040000000420000003d00000036000000340000002e",
            INIT_07 => X"0000002a000000260000002400000023000000240000001e0000001d0000001f",
            INIT_08 => X"0000005200000051000000500000004b0000004b00000054000000580000004c",
            INIT_09 => X"0000005200000056000000570000006300000065000000580000004d0000004c",
            INIT_0A => X"000000490000004400000040000000400000003a00000037000000340000002d",
            INIT_0B => X"0000002b00000028000000290000002c00000031000000300000003100000035",
            INIT_0C => X"0000005300000051000000500000004e0000004a000000570000005000000032",
            INIT_0D => X"0000005500000061000000570000005b00000068000000660000005800000050",
            INIT_0E => X"00000049000000400000003f0000003f0000003b00000038000000390000003a",
            INIT_0F => X"0000003d0000003f000000440000004700000049000000470000004500000045",
            INIT_10 => X"0000004f0000004f0000004f0000004f0000004a000000530000004c00000037",
            INIT_11 => X"00000053000000540000004b0000004b0000004e000000590000005a00000057",
            INIT_12 => X"000000530000004200000043000000460000004e000000500000005400000057",
            INIT_13 => X"0000005700000056000000590000005900000058000000540000004f00000049",
            INIT_14 => X"0000004c0000004a0000004b0000004d00000049000000490000004600000046",
            INIT_15 => X"000000460000004500000047000000490000004b0000004e0000004e00000051",
            INIT_16 => X"0000005a00000059000000600000006200000064000000680000006600000068",
            INIT_17 => X"000000630000005f000000610000005e00000057000000500000004900000042",
            INIT_18 => X"0000004a0000004800000047000000490000004a0000003e0000002b00000033",
            INIT_19 => X"000000440000004000000044000000470000004b0000004a000000510000005e",
            INIT_1A => X"00000060000000620000006e000000720000006600000064000000680000006d",
            INIT_1B => X"000000630000005b00000055000000500000004c000000490000004600000043",
            INIT_1C => X"00000047000000480000004700000048000000470000003a0000002a00000029",
            INIT_1D => X"00000039000000360000003a0000003f00000041000000470000005200000060",
            INIT_1E => X"000000690000005e0000005d00000067000000670000006a0000006c00000061",
            INIT_1F => X"0000005d0000005b000000540000005000000050000000500000004f0000004d",
            INIT_20 => X"00000049000000490000004b000000520000005800000067000000570000002e",
            INIT_21 => X"0000003800000038000000450000005200000051000000570000005a00000057",
            INIT_22 => X"00000062000000630000005e0000005b00000061000000660000006a00000066",
            INIT_23 => X"0000005e00000063000000610000005c00000059000000590000005b0000005f",
            INIT_24 => X"000000560000005f0000006d0000007b00000088000000990000006800000033",
            INIT_25 => X"0000003c0000003b0000004900000061000000650000006c000000660000005a",
            INIT_26 => X"0000005f00000061000000610000005d0000005d00000063000000690000006e",
            INIT_27 => X"00000067000000690000006c0000006c0000006d0000006e0000006e0000006e",
            INIT_28 => X"0000007f0000008b000000960000009d000000a0000000a20000005700000032",
            INIT_29 => X"0000004300000038000000350000005800000065000000700000006b0000005a",
            INIT_2A => X"0000005e000000600000005e00000060000000600000005f0000006000000065",
            INIT_2B => X"00000068000000710000007d0000007e0000007b000000770000007400000070",
            INIT_2C => X"000000980000009d0000009f000000a2000000a00000009f0000005a0000002c",
            INIT_2D => X"00000048000000450000003a00000056000000670000005a000000610000005c",
            INIT_2E => X"0000005a000000600000005f0000005e0000006300000062000000570000005c",
            INIT_2F => X"000000610000007000000083000000830000007f00000079000000740000006c",
            INIT_30 => X"0000009b0000009e000000a00000009d00000098000000940000007200000030",
            INIT_31 => X"00000044000000580000005e000000670000007300000060000000580000005d",
            INIT_32 => X"0000005900000065000000620000005e00000063000000650000005400000055",
            INIT_33 => X"000000690000006e0000007d000000840000007f000000760000006b0000005f",
            INIT_34 => X"00000094000000940000009500000092000000900000008e0000008800000050",
            INIT_35 => X"0000002f000000480000005e0000006800000072000000710000005c0000005e",
            INIT_36 => X"0000005d00000067000000610000005d00000060000000610000005500000052",
            INIT_37 => X"0000006b0000006b0000006f000000790000007000000064000000570000004d",
            INIT_38 => X"00000086000000870000008a0000008c0000008e000000930000009700000089",
            INIT_39 => X"0000005d00000049000000320000003e000000590000005e0000005a00000062",
            INIT_3A => X"000000660000006900000067000000610000005e0000005e0000005600000053",
            INIT_3B => X"0000005f000000650000005c000000660000005f000000520000004a0000004b",
            INIT_3C => X"00000083000000860000008b00000090000000980000009f0000009a00000098",
            INIT_3D => X"0000009e00000076000000350000003900000067000000640000005f00000066",
            INIT_3E => X"0000006e000000740000006f0000006a000000610000005b0000005700000055",
            INIT_3F => X"0000005400000062000000550000005300000053000000550000005a0000005f",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY42;


    MEM_IFMAP_LAYER0_ENTITY43 : if BRAM_NAME = "ifmap_layer0_entity43" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000870000009000000098000000a0000000a4000000a10000008900000073",
            INIT_01 => X"0000009d00000091000000800000006e0000007b0000007a0000006800000067",
            INIT_02 => X"000000690000006d0000006c00000068000000610000005a0000005800000057",
            INIT_03 => X"0000004f0000005c00000057000000550000006500000069000000690000005e",
            INIT_04 => X"000000940000009a0000009f000000a4000000aa000000b3000000b00000007f",
            INIT_05 => X"000000b0000000c50000009d0000009800000071000000910000008000000067",
            INIT_06 => X"00000067000000650000006800000066000000610000005f0000005b00000059",
            INIT_07 => X"0000004f000000560000005b0000005b0000006d000000680000005600000046",
            INIT_08 => X"0000009b000000a4000000b2000000c5000000dd000000ee000000f8000000c4",
            INIT_09 => X"0000009c000000c8000000b0000000b80000006c0000008e000000890000006a",
            INIT_0A => X"0000006400000063000000640000006500000065000000630000005f00000059",
            INIT_0B => X"00000050000000510000005c0000005300000058000000520000004900000047",
            INIT_0C => X"000000bf000000d6000000eb000000f9000000fd000000f6000000fb000000f4",
            INIT_0D => X"000000a00000009e000000ac000000c300000071000000720000008b0000006e",
            INIT_0E => X"000000620000006200000061000000630000006700000068000000660000005c",
            INIT_0F => X"000000530000004e00000055000000490000004b000000500000004a00000048",
            INIT_10 => X"000000f5000000fc000000fd000000fe000000f3000000bb000000ba000000c9",
            INIT_11 => X"0000009100000080000000970000009c000000740000006a0000008000000072",
            INIT_12 => X"000000680000006700000065000000670000006c0000006e000000690000005c",
            INIT_13 => X"000000520000004c00000054000000550000004e000000530000004d00000049",
            INIT_14 => X"000000fb000000fc000000fc00000100000000e90000007e0000006b00000072",
            INIT_15 => X"0000006900000073000000780000006e00000063000000630000006800000067",
            INIT_16 => X"0000006d0000006e0000006b0000006b000000700000006e0000006000000056",
            INIT_17 => X"0000004e0000004c0000005a000000680000005b00000052000000520000004f",
            INIT_18 => X"000000f8000000f8000000f6000000eb000000c80000007c0000007200000076",
            INIT_19 => X"0000005d00000057000000530000004f00000050000000560000004b00000044",
            INIT_1A => X"0000005f00000064000000620000006100000062000000610000006100000061",
            INIT_1B => X"0000005b000000570000005b0000006f0000006e000000550000005200000052",
            INIT_1C => X"000000eb000000d6000000b5000000960000008a000000880000008500000084",
            INIT_1D => X"000000640000003d000000390000003c0000004300000059000000600000003a",
            INIT_1E => X"000000330000004500000047000000500000005e000000650000006800000065",
            INIT_1F => X"0000005d000000570000005e0000006d00000077000000620000005100000051",
            INIT_20 => X"00000099000000820000007a000000780000007c0000007a0000006f00000067",
            INIT_21 => X"0000006a0000005a000000390000003400000045000000660000006a00000053",
            INIT_22 => X"00000040000000470000004d000000550000006400000067000000660000006d",
            INIT_23 => X"0000006a000000570000005d0000006300000071000000730000005c00000050",
            INIT_24 => X"0000006d0000006f000000720000006d0000006500000061000000660000006d",
            INIT_25 => X"000000750000007800000067000000550000005d000000650000005f00000059",
            INIT_26 => X"0000004a0000004b000000520000005a00000072000000770000006900000066",
            INIT_27 => X"0000006f0000006b0000005e0000006200000065000000750000006b0000004f",
            INIT_28 => X"00000069000000620000005d0000005b000000630000006a0000006f00000071",
            INIT_29 => X"0000007000000068000000610000005f000000500000004c000000540000005c",
            INIT_2A => X"00000051000000480000004f00000059000000750000007b000000690000005e",
            INIT_2B => X"0000006000000067000000670000006500000060000000690000006f0000005a",
            INIT_2C => X"00000057000000570000005e000000650000006c0000006e0000006b00000064",
            INIT_2D => X"0000005b0000005100000056000000680000005d000000490000004c0000005c",
            INIT_2E => X"000000580000004d0000004f0000004f0000005b000000640000005d00000056",
            INIT_2F => X"000000570000005c000000610000006000000060000000600000006600000065",
            INIT_30 => X"0000005a000000600000006700000069000000650000005f0000005600000050",
            INIT_31 => X"0000005100000055000000600000006a0000006200000055000000600000005d",
            INIT_32 => X"00000058000000510000004f0000004c000000470000004c000000540000005b",
            INIT_33 => X"0000005c00000056000000530000005a00000062000000600000005b00000060",
            INIT_34 => X"00000064000000630000005f00000056000000500000004f0000004f0000004f",
            INIT_35 => X"0000005200000053000000620000006c00000063000000600000006100000059",
            INIT_36 => X"0000005c000000540000004f000000510000004c0000004a0000005200000059",
            INIT_37 => X"0000005a0000005500000052000000560000005d0000005c0000005300000053",
            INIT_38 => X"000000570000004e00000049000000470000004d000000570000005900000053",
            INIT_39 => X"000000510000004f000000610000006a0000006400000067000000590000005c",
            INIT_3A => X"00000060000000570000005800000059000000520000004f0000005400000053",
            INIT_3B => X"000000560000005a000000560000005300000056000000560000004f00000049",
            INIT_3C => X"0000003e0000003f000000460000004900000054000000560000005300000051",
            INIT_3D => X"0000004e0000004a0000005e0000006b0000005f000000680000005b00000058",
            INIT_3E => X"0000005b00000058000000580000005900000055000000500000005500000053",
            INIT_3F => X"000000540000005900000056000000500000004c0000004d0000004c00000048",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY43;


    MEM_IFMAP_LAYER0_ENTITY44 : if BRAM_NAME = "ifmap_layer0_entity44" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005e0000005e0000005d000000590000005a0000005a0000006000000060",
            INIT_01 => X"00000061000000660000006e000000650000005e000000580000005500000052",
            INIT_02 => X"0000004e0000004b000000490000004800000045000000410000003d00000038",
            INIT_03 => X"000000330000002e000000290000002700000028000000220000001d00000019",
            INIT_04 => X"000000600000005f0000005f0000005900000059000000590000005f00000062",
            INIT_05 => X"00000061000000600000006a0000006b00000060000000590000005500000052",
            INIT_06 => X"0000004f0000004b0000004700000049000000440000003d0000003b00000035",
            INIT_07 => X"000000310000002c000000270000002500000026000000200000001f0000001f",
            INIT_08 => X"0000005e0000005c0000005c00000057000000540000005a0000005d00000051",
            INIT_09 => X"0000005900000060000000630000006e00000070000000620000005600000054",
            INIT_0A => X"0000004f0000004900000044000000460000003f0000003a0000003600000030",
            INIT_0B => X"0000002e0000002b000000290000002b0000002f0000002e0000003000000031",
            INIT_0C => X"0000005f0000005d0000005c0000005a000000530000005d0000005600000039",
            INIT_0D => X"0000005d0000006b00000063000000680000007400000072000000650000005a",
            INIT_0E => X"0000004e0000004300000042000000420000003e000000380000003800000039",
            INIT_0F => X"0000003c0000003e000000410000004200000043000000410000003f0000003d",
            INIT_10 => X"0000005c0000005b0000005b0000005b0000005300000059000000520000003e",
            INIT_11 => X"0000005c0000005f00000058000000580000005c000000680000006900000064",
            INIT_12 => X"0000005b000000460000004500000048000000500000004d0000005000000053",
            INIT_13 => X"000000530000005100000051000000500000004f0000004b000000460000003f",
            INIT_14 => X"00000058000000560000005700000059000000520000004f0000004c0000004d",
            INIT_15 => X"000000500000005200000055000000570000005a0000005e0000005e0000005f",
            INIT_16 => X"000000630000005e000000620000006300000064000000640000006000000062",
            INIT_17 => X"0000005d0000005800000058000000530000004c000000450000003e00000037",
            INIT_18 => X"00000055000000540000005200000054000000510000003d0000002a00000037",
            INIT_19 => X"000000530000005700000058000000590000005b000000570000005d00000065",
            INIT_1A => X"0000006200000064000000700000007300000069000000670000006700000067",
            INIT_1B => X"0000005b000000500000004e0000004a000000440000003f0000003900000036",
            INIT_1C => X"000000520000005300000052000000540000004c00000037000000260000002c",
            INIT_1D => X"0000004c00000055000000520000005100000050000000530000005b00000063",
            INIT_1E => X"0000006700000060000000610000006c0000006d00000072000000710000005e",
            INIT_1F => X"000000520000004d0000004d0000004b0000004700000044000000400000003b",
            INIT_20 => X"0000005100000052000000540000005b0000005e000000680000005500000031",
            INIT_21 => X"00000049000000540000005b000000630000006100000064000000650000005e",
            INIT_22 => X"000000650000006800000065000000620000006a0000006f0000007200000067",
            INIT_23 => X"0000005700000055000000520000004e0000004a000000460000004700000048",
            INIT_24 => X"0000005c0000006500000073000000800000008e0000009d0000006800000036",
            INIT_25 => X"0000004b000000540000005d00000071000000750000007c0000007500000065",
            INIT_26 => X"000000670000006a0000006b00000067000000680000006e0000007400000076",
            INIT_27 => X"000000640000005a000000550000005400000055000000550000005500000052",
            INIT_28 => X"000000820000008e00000099000000a0000000a6000000aa0000005900000035",
            INIT_29 => X"000000500000004d000000460000006800000077000000820000007f0000006b",
            INIT_2A => X"0000006a0000006c000000690000006a0000006a000000690000006e00000072",
            INIT_2B => X"000000690000006200000062000000600000005e0000005b0000005900000055",
            INIT_2C => X"0000009a0000009f000000a2000000a4000000a7000000a90000005d0000002e",
            INIT_2D => X"00000051000000560000004a000000670000007b000000700000007a00000072",
            INIT_2E => X"0000006a0000006d0000006a000000670000006b00000069000000670000006e",
            INIT_2F => X"00000066000000610000006500000063000000600000005e0000005a00000055",
            INIT_30 => X"0000009d0000009f000000a10000009e0000009e0000009f0000007500000030",
            INIT_31 => X"00000049000000650000006c0000007800000087000000780000007400000075",
            INIT_32 => X"0000006b000000730000006c00000066000000690000006a0000006400000069",
            INIT_33 => X"00000070000000600000006000000065000000620000005d000000550000004c",
            INIT_34 => X"000000990000009800000097000000930000009300000093000000870000004c",
            INIT_35 => X"0000002c00000049000000670000007500000083000000850000007300000071",
            INIT_36 => X"0000006c00000077000000710000006b0000006a0000006a0000006500000064",
            INIT_37 => X"00000075000000690000005d000000620000005d000000550000004a00000040",
            INIT_38 => X"0000008f0000008e0000008e0000008e0000008f000000940000009500000083",
            INIT_39 => X"00000054000000410000003500000046000000630000006b000000680000006d",
            INIT_3A => X"000000720000007c0000007d000000750000006e0000006c0000006500000062",
            INIT_3B => X"0000006c0000006f000000580000005a0000005500000048000000410000003f",
            INIT_3C => X"0000008c0000008d0000008e0000009100000099000000a00000009900000093",
            INIT_3D => X"000000970000006f000000340000003a0000006a00000068000000650000006e",
            INIT_3E => X"0000007b000000890000008700000080000000730000006c0000006800000065",
            INIT_3F => X"000000630000006f000000590000004e0000004a000000480000004a0000004d",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY44;


    MEM_IFMAP_LAYER0_ENTITY45 : if BRAM_NAME = "ifmap_layer0_entity45" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000008f000000950000009b0000009f000000a4000000a00000008800000072",
            INIT_01 => X"0000009b0000008f0000007a000000680000007600000077000000660000006c",
            INIT_02 => X"00000078000000840000008500000080000000750000006d0000006b0000006a",
            INIT_03 => X"000000610000006c00000062000000560000005a000000540000004f00000044",
            INIT_04 => X"0000009a0000009d0000009f000000a1000000a7000000b1000000b000000081",
            INIT_05 => X"000000b3000000c7000000970000008e00000068000000890000007b0000006c",
            INIT_06 => X"000000790000007e00000083000000800000007700000073000000700000006e",
            INIT_07 => X"00000063000000690000006a0000005e0000005c0000004a0000003400000027",
            INIT_08 => X"0000009d000000a4000000b0000000c1000000da000000ec000000f7000000c7",
            INIT_09 => X"000000a3000000ce000000ad000000b100000065000000880000008600000071",
            INIT_0A => X"000000770000007e00000082000000810000007d0000007a0000007600000071",
            INIT_0B => X"00000068000000670000006a000000500000003e0000002c0000002500000027",
            INIT_0C => X"000000c0000000d4000000e8000000f6000000fa000000f2000000fa000000f7",
            INIT_0D => X"000000a9000000aa000000ae000000c10000006e000000700000008b00000078",
            INIT_0E => X"000000760000007e0000008000000080000000800000007f0000007e00000074",
            INIT_0F => X"0000006c00000066000000600000003e0000002a00000025000000270000002b",
            INIT_10 => X"000000f5000000fb000000fa000000fb000000f1000000ba000000be000000d2",
            INIT_11 => X"000000a1000000920000009c000000a00000007d00000073000000870000007a",
            INIT_12 => X"000000780000007f00000081000000800000007f0000007f0000007d00000074",
            INIT_13 => X"0000006a0000006200000057000000420000002d0000002a0000002900000029",
            INIT_14 => X"000000fb000000fb000000fb000000fe000000ea000000830000007400000082",
            INIT_15 => X"0000007f0000008a000000820000007c0000007a00000077000000720000006b",
            INIT_16 => X"0000007600000080000000820000007f0000007d000000770000006f0000006c",
            INIT_17 => X"000000630000005a00000052000000500000003d0000002f0000002c00000029",
            INIT_18 => X"000000fc000000fc000000f9000000ef000000cb000000800000007b00000083",
            INIT_19 => X"0000006f0000006c00000066000000670000006a000000690000005100000044",
            INIT_1A => X"000000660000007500000078000000740000006e0000006b0000007000000073",
            INIT_1B => X"00000068000000590000004b0000005400000051000000340000002d0000002d",
            INIT_1C => X"000000f5000000df000000bf000000a00000009000000089000000890000008a",
            INIT_1D => X"0000006d0000004b00000051000000570000005a00000066000000630000003a",
            INIT_1E => X"0000003a000000560000005f000000650000006d000000740000007a00000074",
            INIT_1F => X"000000610000004d000000460000005000000059000000420000002f0000002f",
            INIT_20 => X"000000a50000008d0000008600000084000000820000007b0000007000000069",
            INIT_21 => X"0000006b0000005e0000004a00000047000000530000006e0000006f00000056",
            INIT_22 => X"000000480000005a000000660000006c000000760000007b0000007b0000007c",
            INIT_23 => X"0000006c00000049000000420000004400000052000000540000003d00000030",
            INIT_24 => X"00000075000000780000007a000000750000006a00000061000000650000006a",
            INIT_25 => X"00000070000000730000006a000000570000005c000000680000006800000061",
            INIT_26 => X"000000540000005f0000006c00000072000000860000008e000000820000007a",
            INIT_27 => X"0000007700000064000000450000004000000045000000570000004f00000032",
            INIT_28 => X"0000006c00000066000000600000005e000000650000006b0000006e0000006b",
            INIT_29 => X"000000670000005d000000560000005100000042000000480000005d00000068",
            INIT_2A => X"0000005e0000005f0000006b000000710000008900000094000000850000007a",
            INIT_2B => X"000000720000006b0000005100000042000000400000004b000000550000003f",
            INIT_2C => X"00000058000000570000005d000000630000006b0000006c0000006500000057",
            INIT_2D => X"000000490000003c00000041000000530000004a0000003f0000004e0000005e",
            INIT_2E => X"00000059000000570000005f0000005d000000690000007b0000007a00000072",
            INIT_2F => X"0000006d000000680000004e0000003b0000003c0000003f0000004a0000004b",
            INIT_30 => X"0000005d0000005f000000610000005f0000005b000000540000004500000038",
            INIT_31 => X"0000003200000031000000420000005500000053000000490000005500000048",
            INIT_32 => X"0000003e0000003e000000430000004400000045000000580000006400000068",
            INIT_33 => X"000000650000005a000000400000003300000035000000360000003a00000045",
            INIT_34 => X"000000600000005b00000051000000440000003b000000370000003400000030",
            INIT_35 => X"0000002f0000002e0000004000000052000000520000004f0000004d00000039",
            INIT_36 => X"0000003500000032000000340000003a0000003a0000003f000000470000004a",
            INIT_37 => X"0000004800000041000000340000002e00000030000000310000003000000036",
            INIT_38 => X"000000490000003c000000310000002b0000002c000000300000003400000030",
            INIT_39 => X"000000300000002c0000003a000000490000004b0000004f0000003e00000035",
            INIT_3A => X"000000320000002e0000003400000039000000340000002f000000330000002f",
            INIT_3B => X"0000002f000000310000002e0000002a0000002b0000002d0000002b0000002a",
            INIT_3C => X"000000290000002500000027000000250000002a00000029000000290000002d",
            INIT_3D => X"0000002f0000002b0000003600000047000000430000004c0000003b0000002e",
            INIT_3E => X"0000002b0000002a0000002d000000300000002f0000002d000000310000002d",
            INIT_3F => X"0000002b0000002d0000002a0000002700000025000000280000002800000026",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY45;


    MEM_IFMAP_LAYER0_ENTITY46 : if BRAM_NAME = "ifmap_layer0_entity46" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005500000054000000530000004f00000050000000520000005d0000005f",
            INIT_01 => X"0000005a000000550000004f000000480000004b0000004e000000540000004f",
            INIT_02 => X"000000440000003e0000003c0000003d0000003c0000003b0000003800000033",
            INIT_03 => X"0000002e000000290000002500000023000000240000001e0000001900000015",
            INIT_04 => X"0000005600000055000000550000004f0000004e000000500000005a0000005d",
            INIT_05 => X"0000005400000049000000460000004700000044000000450000004700000048",
            INIT_06 => X"00000046000000430000003e0000003e0000003800000035000000340000002e",
            INIT_07 => X"00000029000000250000002200000020000000210000001b0000001a0000001b",
            INIT_08 => X"0000005400000053000000520000004e00000049000000500000005600000048",
            INIT_09 => X"00000046000000410000003800000043000000480000003f000000360000003c",
            INIT_0A => X"00000042000000410000003d0000003a000000300000002f0000002d00000026",
            INIT_0B => X"000000240000002100000022000000250000002a000000290000002a0000002c",
            INIT_0C => X"0000005500000053000000520000005000000048000000520000004d0000002b",
            INIT_0D => X"00000043000000450000003200000034000000410000003f000000320000002f",
            INIT_0E => X"000000320000003400000039000000360000002d0000002b0000002b0000002c",
            INIT_0F => X"0000002f00000032000000380000003b0000003c0000003b0000003800000037",
            INIT_10 => X"00000052000000510000005100000051000000480000004c000000460000002c",
            INIT_11 => X"0000003d00000033000000220000001d0000001f000000270000002600000023",
            INIT_12 => X"000000290000002b000000390000003b0000003d0000003d0000004100000044",
            INIT_13 => X"0000004400000042000000470000004800000047000000430000003e00000038",
            INIT_14 => X"0000004d0000004c0000004c0000004f00000047000000420000003e00000038",
            INIT_15 => X"0000002c000000210000001a0000001700000016000000140000000f0000000e",
            INIT_16 => X"0000001f000000350000004f0000005400000053000000520000004e00000050",
            INIT_17 => X"0000004c000000480000004d0000004b000000440000003c000000350000002e",
            INIT_18 => X"0000004900000047000000460000004800000047000000370000002000000020",
            INIT_19 => X"00000026000000180000001400000013000000120000000b0000000e00000015",
            INIT_1A => X"0000001800000029000000460000005900000056000000500000004f00000052",
            INIT_1B => X"0000004b0000004800000048000000430000003b000000340000002d0000002a",
            INIT_1C => X"0000004400000045000000440000004500000043000000330000001c00000011",
            INIT_1D => X"000000170000000c0000000a0000000b000000090000000b0000001100000018",
            INIT_1E => X"0000001c00000016000000210000003f0000004d0000004f0000004d00000040",
            INIT_1F => X"000000410000004900000048000000420000003c000000360000002f0000002b",
            INIT_20 => X"0000004400000045000000470000004e000000520000005d0000004600000013",
            INIT_21 => X"000000120000000c000000190000002500000020000000210000002100000014",
            INIT_22 => X"0000001600000018000000190000002100000031000000380000003c0000003b",
            INIT_23 => X"0000003b0000004b000000490000003f00000039000000340000003400000035",
            INIT_24 => X"00000050000000590000006700000075000000800000008d0000005500000016",
            INIT_25 => X"000000150000000f0000002100000038000000390000003d000000350000001c",
            INIT_26 => X"0000001500000016000000160000001400000018000000230000002d0000003a",
            INIT_27 => X"0000003d00000048000000460000004100000041000000400000003f0000003d",
            INIT_28 => X"00000077000000830000008e0000009500000098000000980000004700000018",
            INIT_29 => X"0000001e0000001100000015000000310000003c000000440000003f00000021",
            INIT_2A => X"000000190000001b00000015000000110000000f000000140000001c0000002b",
            INIT_2B => X"00000037000000460000004d0000004a00000049000000470000004400000041",
            INIT_2C => X"0000008f00000094000000960000009900000099000000990000004f00000017",
            INIT_2D => X"0000002800000022000000190000002e0000003d000000300000003700000027",
            INIT_2E => X"0000001d000000240000001f000000150000001300000015000000120000001f",
            INIT_2F => X"0000002a0000003b0000004c0000004d0000004d0000004c0000004a00000045",
            INIT_30 => X"0000009200000095000000970000009400000092000000920000006b00000020",
            INIT_31 => X"0000002b00000037000000340000003b00000047000000340000002c00000029",
            INIT_32 => X"00000022000000320000002c0000001e0000001a0000001c0000001200000019",
            INIT_33 => X"0000002e000000320000004500000051000000510000004f0000004900000042",
            INIT_34 => X"000000900000008f0000008f0000008b0000008a000000890000007e00000040",
            INIT_35 => X"0000001a0000002e0000003d0000004100000046000000400000002800000024",
            INIT_36 => X"00000024000000360000003300000028000000210000001d0000001200000013",
            INIT_37 => X"0000002f000000330000003c0000004e0000004f0000004a0000004000000037",
            INIT_38 => X"0000008500000084000000860000008600000086000000880000008900000077",
            INIT_39 => X"00000047000000310000001b000000210000002e0000002a0000002000000022",
            INIT_3A => X"00000028000000390000003d00000032000000270000001c0000001100000011",
            INIT_3B => X"00000024000000330000003000000041000000460000003e0000003600000032",
            INIT_3C => X"0000007d0000007f00000081000000850000008c000000910000008800000081",
            INIT_3D => X"000000840000005a0000001e0000001e00000040000000330000002700000027",
            INIT_3E => X"0000003100000045000000450000003d0000002c0000001c0000001400000013",
            INIT_3F => X"0000001900000030000000290000002d00000035000000390000003c0000003d",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY46;


    MEM_IFMAP_LAYER0_ENTITY47 : if BRAM_NAME = "ifmap_layer0_entity47" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007d000000840000008b000000910000009500000091000000750000005a",
            INIT_01 => X"00000080000000720000006200000050000000570000004d0000003100000028",
            INIT_02 => X"0000002e0000003f000000440000003c0000002d0000001f0000001900000017",
            INIT_03 => X"000000150000002a0000002b0000002d00000040000000420000003e00000032",
            INIT_04 => X"000000880000008c00000090000000930000009a000000a40000009e00000068",
            INIT_05 => X"00000095000000a60000007a0000007700000050000000670000004b00000029",
            INIT_06 => X"0000002d00000038000000410000003c00000030000000280000001f0000001b",
            INIT_07 => X"00000015000000230000002f0000003200000041000000390000002300000014",
            INIT_08 => X"0000009000000097000000a4000000b6000000d2000000e6000000eb000000b2",
            INIT_09 => X"00000085000000ab0000008a000000950000004d00000067000000550000002d",
            INIT_0A => X"0000002b000000380000003f0000003c0000003500000030000000270000001d",
            INIT_0B => X"000000170000001d0000002f00000027000000270000001f0000001600000015",
            INIT_0C => X"000000b7000000cd000000e1000000f0000000f8000000f2000000f2000000e6",
            INIT_0D => X"0000008d00000084000000840000009f000000530000004d0000005600000031",
            INIT_0E => X"0000002a000000370000003c0000003a00000039000000370000002f00000021",
            INIT_0F => X"000000190000001a000000270000001c000000190000001d0000001c0000001b",
            INIT_10 => X"000000f1000000f8000000f7000000f9000000ec000000b0000000ab000000b5",
            INIT_11 => X"000000780000006200000072000000760000004d0000003c0000004700000034",
            INIT_12 => X"0000002e00000036000000390000003a0000003b000000390000003000000020",
            INIT_13 => X"000000180000001700000025000000250000001c000000200000001f0000001a",
            INIT_14 => X"000000f8000000f9000000f9000000fd000000e00000006a0000005300000055",
            INIT_15 => X"000000470000004e0000005100000041000000300000002e0000003400000031",
            INIT_16 => X"000000330000003700000036000000390000003d00000033000000240000001b",
            INIT_17 => X"00000015000000160000002700000036000000280000001f0000001f0000001c",
            INIT_18 => X"000000f7000000f8000000f5000000eb000000c20000006d000000600000005e",
            INIT_19 => X"000000410000003500000023000000190000001c0000002b0000002d00000020",
            INIT_1A => X"0000002e000000330000002f0000002f000000300000002d0000002b00000029",
            INIT_1B => X"000000220000001e000000240000003a00000039000000210000001d0000001e",
            INIT_1C => X"000000ec000000d7000000b60000009800000088000000810000007a00000074",
            INIT_1D => X"00000051000000230000000d0000000900000014000000340000004900000022",
            INIT_1E => X"000000110000001c0000001a000000200000002f0000003b0000003b00000031",
            INIT_1F => X"000000230000001a00000022000000340000003f0000002c0000001c0000001d",
            INIT_20 => X"0000009a000000820000007a000000780000007b00000076000000680000005c",
            INIT_21 => X"0000005a000000460000001f000000120000001d0000003d0000004500000034",
            INIT_22 => X"000000220000002400000024000000280000003a00000047000000410000003d",
            INIT_23 => X"00000030000000170000001f00000028000000380000003c000000270000001c",
            INIT_24 => X"000000690000006b0000006d000000680000005f000000580000005b0000005d",
            INIT_25 => X"0000006000000062000000560000003e00000038000000380000002f00000031",
            INIT_26 => X"00000028000000250000002a000000300000004c0000005b0000004800000039",
            INIT_27 => X"000000360000002c0000001d000000230000002a0000003d000000370000001d",
            INIT_28 => X"0000005f00000059000000530000005100000056000000580000005b00000058",
            INIT_29 => X"0000005300000049000000440000003e00000028000000230000002c00000034",
            INIT_2A => X"000000280000001e0000002700000031000000510000005f0000004700000032",
            INIT_2B => X"000000290000002a000000250000002300000022000000300000003a00000028",
            INIT_2C => X"0000004b000000490000004f0000005500000057000000530000004c00000040",
            INIT_2D => X"00000033000000270000002a0000003b00000032000000220000002900000031",
            INIT_2E => X"000000260000001e000000240000002700000037000000450000003c0000002d",
            INIT_2F => X"0000002600000026000000220000001d00000020000000240000003000000033",
            INIT_30 => X"0000004c0000004e0000004f0000004d00000044000000390000002c00000021",
            INIT_31 => X"0000001d0000001e0000002e0000003d00000037000000290000003200000026",
            INIT_32 => X"0000001d0000001a0000001d0000001e0000001d000000250000002e00000030",
            INIT_33 => X"0000002e0000002500000019000000180000001e00000020000000240000002f",
            INIT_34 => X"000000500000004a000000400000003200000026000000200000001e0000001b",
            INIT_35 => X"0000001b0000001b0000002d0000003c000000350000002f0000002c0000001d",
            INIT_36 => X"0000001c00000017000000170000001c00000019000000180000002000000025",
            INIT_37 => X"000000230000001d00000015000000150000001a0000001e0000001c00000022",
            INIT_38 => X"0000003a0000002d000000210000001a0000001a0000001d000000210000001c",
            INIT_39 => X"0000001b0000001800000027000000330000003100000032000000210000001c",
            INIT_3A => X"0000001b00000015000000190000001d00000018000000150000001900000017",
            INIT_3B => X"000000170000001a0000001600000012000000150000001a0000001900000017",
            INIT_3C => X"0000001b0000001700000018000000150000001a000000190000001800000019",
            INIT_3D => X"0000001a0000001600000021000000300000002a000000330000002300000018",
            INIT_3E => X"0000001500000014000000150000001800000017000000170000001d00000019",
            INIT_3F => X"000000180000001b000000160000001200000011000000160000001800000016",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY47;


    MEM_IFMAP_LAYER0_ENTITY48 : if BRAM_NAME = "ifmap_layer0_entity48" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000017000000130000001500000041000000a4000000bc000000b7000000b2",
            INIT_01 => X"000000aa000000ac000000ba000000ba000000b8000000b7000000b6000000b7",
            INIT_02 => X"000000b4000000a40000007f0000005c0000006b0000006e00000099000000c2",
            INIT_03 => X"000000c3000000c9000000c5000000c6000000c9000000c8000000c7000000c5",
            INIT_04 => X"0000001700000013000000150000002e00000099000000ca000000bf000000b2",
            INIT_05 => X"000000a40000009e000000a9000000b7000000ba000000b8000000b4000000b2",
            INIT_06 => X"000000b4000000ad0000008a000000560000004a0000006a000000b4000000ce",
            INIT_07 => X"000000cf000000d5000000d0000000ce000000cf000000cd000000cc000000ca",
            INIT_08 => X"0000001700000014000000170000001f0000007f000000c8000000b9000000a8",
            INIT_09 => X"0000009f0000009e0000009a000000a2000000b2000000b2000000b3000000b2",
            INIT_0A => X"000000b5000000be000000b60000007d0000004700000072000000c5000000d1",
            INIT_0B => X"000000d5000000d8000000d5000000d3000000d4000000d3000000d0000000ce",
            INIT_0C => X"0000001700000015000000180000001700000063000000bd000000af000000a0",
            INIT_0D => X"000000a8000000a8000000a600000095000000aa000000ba000000bf000000c3",
            INIT_0E => X"000000c3000000c8000000bc0000008d0000006300000092000000d2000000d6",
            INIT_0F => X"000000d5000000d4000000d4000000d5000000d9000000d9000000d7000000d6",
            INIT_10 => X"0000001900000017000000170000001500000048000000aa000000a500000097",
            INIT_11 => X"000000af000000b7000000b90000009b000000920000009d000000a9000000bc",
            INIT_12 => X"000000c5000000c4000000b20000008d00000079000000ac000000d3000000db",
            INIT_13 => X"000000dd000000d9000000d9000000d9000000d6000000d4000000d1000000ce",
            INIT_14 => X"0000001a0000001b0000001a00000017000000310000008f000000a40000009a",
            INIT_15 => X"000000a9000000c2000000c8000000a6000000820000007d0000008000000097",
            INIT_16 => X"000000a5000000a5000000940000008f00000093000000b6000000bc000000c9",
            INIT_17 => X"000000d4000000d9000000d5000000db000000dc000000d7000000d7000000d3",
            INIT_18 => X"0000001e0000001a0000001b00000019000000250000007d000000b4000000ab",
            INIT_19 => X"000000a9000000c5000000ca000000b30000008b000000710000007a00000082",
            INIT_1A => X"00000077000000850000007a0000008c000000b9000000cb000000bf000000c9",
            INIT_1B => X"000000d7000000da000000d7000000db000000dc000000da000000dc000000e0",
            INIT_1C => X"0000005e000000300000001f0000002400000064000000af000000c1000000a8",
            INIT_1D => X"000000a3000000c0000000c6000000c3000000ae000000910000008e00000084",
            INIT_1E => X"0000006a000000790000007a0000008b000000c0000000d1000000bd000000d5",
            INIT_1F => X"000000f2000000ed000000ef000000e8000000d0000000d5000000de000000e5",
            INIT_20 => X"000000b40000009e000000720000007a000000b1000000be000000be000000a0",
            INIT_21 => X"00000085000000ad000000c5000000c8000000c2000000b9000000a700000092",
            INIT_22 => X"0000008100000081000000850000008d000000b1000000c9000000bd000000dc",
            INIT_23 => X"000000f1000000eb000000e8000000d5000000bd000000c7000000e1000000ea",
            INIT_24 => X"000000c5000000c0000000b2000000ba000000c1000000c3000000c50000009d",
            INIT_25 => X"00000080000000a3000000b9000000bf000000c1000000c3000000b200000097",
            INIT_26 => X"00000072000000810000008300000086000000aa000000c2000000d0000000ea",
            INIT_27 => X"000000ec000000f0000000eb000000c9000000b9000000bb000000d0000000eb",
            INIT_28 => X"000000ca000000c4000000bb000000c0000000c8000000cd000000c500000097",
            INIT_29 => X"00000095000000af000000b8000000bd000000c1000000bb000000a800000088",
            INIT_2A => X"00000075000000800000008000000081000000a7000000b5000000cd000000f0",
            INIT_2B => X"000000f3000000f3000000ee000000ce000000ba000000bb000000c1000000dd",
            INIT_2C => X"000000cd000000cd000000c5000000c0000000cb000000d0000000c2000000a0",
            INIT_2D => X"000000a8000000bf000000c1000000bf000000c1000000ac0000009200000077",
            INIT_2E => X"0000007c0000008e0000008500000087000000a7000000b0000000bf000000ea",
            INIT_2F => X"000000f3000000f1000000ec000000d7000000ba000000b8000000b9000000c4",
            INIT_30 => X"000000ce000000cc000000c8000000c1000000c5000000c7000000bf000000b4",
            INIT_31 => X"000000ac000000b3000000b7000000ad000000ae000000ae0000009800000083",
            INIT_32 => X"0000008d000000a60000008e0000009a000000a9000000ac000000bf000000e6",
            INIT_33 => X"000000f0000000f1000000ef000000e4000000c8000000ba000000b8000000c0",
            INIT_34 => X"000000d2000000ca000000c6000000bf000000c9000000b4000000b1000000ca",
            INIT_35 => X"000000ab0000009a0000008e0000008e000000a8000000a8000000930000009c",
            INIT_36 => X"000000af000000a900000096000000a40000009e000000a0000000c5000000e6",
            INIT_37 => X"000000f1000000f1000000f4000000f2000000e2000000bf000000c3000000d7",
            INIT_38 => X"000000d3000000c9000000c7000000c0000000cf000000aa000000a1000000d7",
            INIT_39 => X"000000bd000000ba000000ad000000ac000000be000000b1000000890000007f",
            INIT_3A => X"000000b4000000ae00000096000000a0000000af000000b0000000c1000000ec",
            INIT_3B => X"000000f5000000f2000000f3000000fb000000ef000000c9000000d4000000e1",
            INIT_3C => X"000000d3000000c4000000c5000000c1000000d1000000b50000009a000000d9",
            INIT_3D => X"000000ce000000c5000000c3000000b9000000aa000000ad000000a600000098",
            INIT_3E => X"000000a3000000b8000000a600000098000000c0000000b5000000af000000cc",
            INIT_3F => X"000000ee000000f3000000f4000000f7000000df000000d5000000e2000000e2",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY48;


    MEM_IFMAP_LAYER0_ENTITY49 : if BRAM_NAME = "ifmap_layer0_entity49" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d6000000c2000000b4000000b5000000c5000000c40000009b000000c6",
            INIT_01 => X"000000d6000000c0000000ae000000b7000000ad000000a1000000ae000000b2",
            INIT_02 => X"00000080000000a4000000bd00000093000000a7000000b40000009c00000076",
            INIT_03 => X"0000009d000000d7000000ef000000eb000000ce000000d6000000ea000000e4",
            INIT_04 => X"000000d7000000c6000000a6000000a3000000b4000000ca000000be000000b9",
            INIT_05 => X"000000cf000000d2000000cd000000d6000000c1000000ae000000b0000000ad",
            INIT_06 => X"0000008100000089000000bf00000099000000a3000000c8000000ab00000087",
            INIT_07 => X"0000007400000090000000b8000000c1000000bb000000d2000000ef000000eb",
            INIT_08 => X"000000d8000000cd000000ae000000a4000000b9000000cb000000d2000000c2",
            INIT_09 => X"000000bf000000d3000000da000000e2000000e1000000cb000000be000000b3",
            INIT_0A => X"0000009700000079000000a80000009e000000a7000000c2000000aa000000ac",
            INIT_0B => X"0000009a0000008300000099000000a9000000a2000000b8000000de000000ec",
            INIT_0C => X"000000d8000000d0000000c0000000b4000000c5000000ca000000d1000000d2",
            INIT_0D => X"000000ba000000bd000000c5000000cc000000d1000000d5000000cf000000b5",
            INIT_0E => X"000000b20000009500000092000000af000000b7000000ae0000009c000000ab",
            INIT_0F => X"000000a300000094000000a9000000b4000000a6000000a0000000ac000000cc",
            INIT_10 => X"000000da000000d5000000ca000000b6000000bf000000cb000000c9000000ca",
            INIT_11 => X"000000ca000000c3000000c1000000c0000000b2000000c6000000cf000000c7",
            INIT_12 => X"000000d3000000cb000000a6000000bb000000b10000009b00000093000000a6",
            INIT_13 => X"000000a7000000ab000000b6000000af0000009c0000009c0000009f000000a7",
            INIT_14 => X"000000d9000000d7000000d1000000ba000000b3000000c8000000d0000000c8",
            INIT_15 => X"000000d1000000d7000000d2000000ba000000a1000000b6000000c4000000c2",
            INIT_16 => X"000000cb000000cf000000be000000b90000009b0000008e0000009b000000a6",
            INIT_17 => X"000000ac000000b3000000ad0000009f000000960000009e0000009e0000008f",
            INIT_18 => X"000000d6000000d5000000d6000000c0000000a9000000c5000000da000000d9",
            INIT_19 => X"000000d7000000d9000000d4000000c3000000aa000000b3000000c3000000bf",
            INIT_1A => X"000000be000000c0000000c0000000aa000000840000008e000000a7000000aa",
            INIT_1B => X"000000aa000000b3000000ad0000009d0000009d00000093000000860000007d",
            INIT_1C => X"000000d5000000d1000000d3000000ca000000a8000000c1000000d8000000de",
            INIT_1D => X"000000df000000de000000d3000000cd000000c2000000c2000000c9000000c6",
            INIT_1E => X"000000c6000000c4000000bc00000099000000860000009b000000ab000000a7",
            INIT_1F => X"000000a6000000bd000000b2000000a5000000a30000008e0000008500000089",
            INIT_20 => X"000000d3000000ce000000ce000000ca000000af000000bf000000d3000000d5",
            INIT_21 => X"000000d6000000d8000000c6000000ab000000c2000000ce000000c9000000c9",
            INIT_22 => X"000000c8000000c5000000b100000096000000900000009e000000a70000009d",
            INIT_23 => X"0000009f000000b5000000b0000000a800000098000000960000009500000090",
            INIT_24 => X"000000d2000000cc000000c9000000c1000000b5000000bc000000d0000000d2",
            INIT_25 => X"000000cd000000ce000000a00000007a000000b1000000d0000000c6000000c2",
            INIT_26 => X"000000c1000000b8000000a6000000960000008b0000009c000000a000000099",
            INIT_27 => X"0000009b000000a00000009f0000009b00000098000000980000008c00000083",
            INIT_28 => X"000000d2000000ca000000c6000000bb000000ae000000b2000000cd000000d6",
            INIT_29 => X"000000d1000000cb000000a400000083000000b4000000ca000000bb000000b6",
            INIT_2A => X"000000b6000000a90000009d0000008b00000086000000990000009a00000090",
            INIT_2B => X"000000970000008d000000830000008d0000009d0000009b0000009600000093",
            INIT_2C => X"000000d2000000c8000000c2000000b5000000a8000000a8000000c4000000d7",
            INIT_2D => X"000000d4000000c7000000bd000000b8000000cb000000b9000000ad000000ac",
            INIT_2E => X"000000a30000009b00000093000000760000008300000094000000910000008d",
            INIT_2F => X"00000090000000840000007f0000008500000095000000a3000000a20000009c",
            INIT_30 => X"000000d0000000c2000000bd000000b4000000a20000009e000000bd000000d3",
            INIT_31 => X"000000d3000000c5000000c2000000c7000000bf000000ac000000a3000000a4",
            INIT_32 => X"0000009e00000093000000820000006d00000089000000900000009000000091",
            INIT_33 => X"00000090000000840000007c0000008600000097000000a20000009f00000093",
            INIT_34 => X"000000c2000000b1000000b0000000b50000009f0000008f000000b3000000cd",
            INIT_35 => X"000000d0000000c7000000c2000000be000000b5000000a50000009c000000a1",
            INIT_36 => X"0000009500000088000000700000007200000089000000850000008a00000092",
            INIT_37 => X"000000920000008300000083000000900000009600000095000000940000008d",
            INIT_38 => X"000000ac0000009d000000a5000000b2000000a7000000850000009c000000c7",
            INIT_39 => X"000000ce000000c7000000c7000000c2000000a000000085000000840000008b",
            INIT_3A => X"0000008c0000007e0000006b0000007e00000082000000810000008a00000095",
            INIT_3B => X"0000008d0000008c000000910000008e000000880000008c0000009500000098",
            INIT_3C => X"0000009700000086000000900000009b0000009e0000007d00000082000000b7",
            INIT_3D => X"000000c5000000bf000000b7000000a500000080000000670000005e00000069",
            INIT_3E => X"0000007700000070000000750000007c000000790000007d0000008b0000008f",
            INIT_3F => X"0000008b0000008c000000810000007d00000084000000950000009b00000096",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY49;


    MEM_IFMAP_LAYER0_ENTITY50 : if BRAM_NAME = "ifmap_layer0_entity50" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001300000015000000100000002f0000008300000093000000930000008e",
            INIT_01 => X"0000008700000089000000900000008e0000008d0000008c0000008c0000008f",
            INIT_02 => X"0000008c0000007e00000060000000490000005f0000005d00000082000000a4",
            INIT_03 => X"0000009b0000009c0000009b0000009d0000009e0000009b0000009800000097",
            INIT_04 => X"0000001400000014000000110000001f0000007a000000a10000009b00000092",
            INIT_05 => X"0000008a000000880000008b0000009500000098000000960000009200000097",
            INIT_06 => X"0000009f00000096000000750000004900000041000000580000009c000000af",
            INIT_07 => X"000000a8000000a9000000ab000000ad000000ac000000a8000000a4000000a3",
            INIT_08 => X"0000001400000014000000140000001500000066000000a2000000970000008c",
            INIT_09 => X"0000008d00000095000000880000008b0000009a00000099000000980000009f",
            INIT_0A => X"000000a6000000ab000000a10000006d0000003a00000061000000b1000000b7",
            INIT_0B => X"000000b3000000b2000000b1000000b2000000b1000000ad000000a9000000a6",
            INIT_0C => X"000000140000001400000015000000110000004f000000990000008c00000082",
            INIT_0D => X"00000097000000a40000009d0000008700000099000000a6000000a9000000b0",
            INIT_0E => X"000000b0000000af000000a1000000760000005200000085000000c4000000c3",
            INIT_0F => X"000000bd000000b7000000b4000000b3000000b3000000b1000000ad000000ab",
            INIT_10 => X"0000001500000014000000150000001300000038000000890000008200000077",
            INIT_11 => X"0000009c000000b2000000b300000092000000840000008b00000094000000a7",
            INIT_12 => X"000000af000000a900000098000000780000006d000000a7000000ce000000d2",
            INIT_13 => X"000000d1000000c9000000c3000000bf000000ba000000b6000000b1000000ac",
            INIT_14 => X"0000001600000016000000170000001600000026000000730000008200000078",
            INIT_15 => X"00000092000000b9000000c30000009e000000760000006c0000006b00000084",
            INIT_16 => X"000000920000008f00000081000000840000008f000000b7000000be000000c7",
            INIT_17 => X"000000cf000000d1000000cc000000d1000000d1000000ca000000c7000000c2",
            INIT_18 => X"000000180000001300000015000000140000001e00000071000000a100000094",
            INIT_19 => X"00000097000000ba000000c2000000aa00000080000000620000006900000071",
            INIT_1A => X"00000068000000740000006b00000080000000b2000000ca000000c0000000c5",
            INIT_1B => X"000000ce000000cf000000d1000000d7000000d8000000d6000000d7000000da",
            INIT_1C => X"0000005800000029000000180000001d00000060000000ae000000ba0000009c",
            INIT_1D => X"00000095000000b5000000bd000000ba000000a4000000840000008100000076",
            INIT_1E => X"0000005c0000006b0000006c0000007c000000b4000000cc000000bb000000ce",
            INIT_1F => X"000000e6000000e0000000e7000000e4000000cd000000d3000000dc000000e2",
            INIT_20 => X"000000b1000000990000006d00000075000000af000000bd000000b700000093",
            INIT_21 => X"00000078000000a1000000bc000000c0000000b8000000ad0000009a00000083",
            INIT_22 => X"0000007300000073000000770000007f000000a6000000c5000000bc000000d8",
            INIT_23 => X"000000e9000000e2000000e3000000d3000000bc000000c6000000e0000000e8",
            INIT_24 => X"000000c2000000bc000000af000000b6000000bf000000c2000000be00000090",
            INIT_25 => X"0000007300000098000000b1000000b6000000b7000000b6000000a40000008a",
            INIT_26 => X"0000006600000076000000770000007b000000a0000000bd000000d0000000e9",
            INIT_27 => X"000000e8000000eb000000ea000000cb000000bb000000bd000000d1000000eb",
            INIT_28 => X"000000c7000000c0000000b7000000bb000000c6000000cd000000bf0000008a",
            INIT_29 => X"00000088000000a5000000b0000000b5000000b8000000af0000009a0000007c",
            INIT_2A => X"0000006b0000007600000077000000780000009e000000b0000000cd000000f0",
            INIT_2B => X"000000f3000000f4000000f2000000d4000000c0000000c0000000c6000000e0",
            INIT_2C => X"000000c9000000c9000000c1000000bb000000c9000000d1000000bc00000092",
            INIT_2D => X"0000009b000000b6000000b9000000b7000000b70000009f000000840000006b",
            INIT_2E => X"00000073000000850000007c0000007e0000009e000000aa000000bd000000eb",
            INIT_2F => X"000000f6000000f6000000f2000000de000000c2000000c0000000c0000000ca",
            INIT_30 => X"000000cb000000c9000000c5000000bd000000c4000000c6000000b7000000a5",
            INIT_31 => X"0000009f000000aa000000b0000000a5000000a4000000a20000008a00000078",
            INIT_32 => X"000000850000009f0000008700000092000000a1000000a5000000bd000000e7",
            INIT_33 => X"000000f4000000f8000000f7000000ea000000d0000000c3000000c1000000c7",
            INIT_34 => X"000000d0000000ca000000c4000000b9000000c1000000a70000009c000000b9",
            INIT_35 => X"000000a1000000910000008700000087000000a10000009e000000890000008f",
            INIT_36 => X"000000a4000000a400000095000000a2000000990000009d000000c3000000e4",
            INIT_37 => X"000000f2000000f7000000f9000000f5000000e8000000c7000000cc000000de",
            INIT_38 => X"000000d2000000cc000000c5000000b6000000bf0000008e0000007d000000c1",
            INIT_39 => X"000000b5000000b1000000a6000000a7000000b8000000aa0000008200000072",
            INIT_3A => X"000000a5000000aa000000980000009e000000ab000000ae000000bd000000e7",
            INIT_3B => X"000000f2000000f4000000f5000000fb000000f2000000cf000000dd000000e9",
            INIT_3C => X"000000d4000000c8000000c5000000b9000000bd0000009100000070000000c0",
            INIT_3D => X"000000c7000000be000000bd000000b4000000a4000000a7000000a000000089",
            INIT_3E => X"00000092000000b0000000a200000091000000b8000000b1000000a8000000c3",
            INIT_3F => X"000000e8000000f1000000f5000000f9000000e4000000dd000000ec000000eb",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY50;


    MEM_IFMAP_LAYER0_ENTITY51 : if BRAM_NAME = "ifmap_layer0_entity51" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d8000000c7000000b6000000ae000000b00000009b0000006e000000ad",
            INIT_01 => X"000000d0000000ba000000a8000000b2000000a80000009b000000a7000000a4",
            INIT_02 => X"0000006e00000096000000b1000000860000009a000000ab0000009000000068",
            INIT_03 => X"00000091000000d1000000ee000000ed000000d2000000dd000000f3000000ed",
            INIT_04 => X"000000db000000ce000000a90000009e000000a3000000a700000095000000a2",
            INIT_05 => X"000000ca000000cd000000c8000000d1000000bc000000a8000000aa000000a1",
            INIT_06 => X"0000007000000078000000ad0000008700000093000000ba0000009b00000073",
            INIT_07 => X"0000006200000084000000b2000000bc000000b9000000d4000000f3000000ef",
            INIT_08 => X"000000dd000000d6000000b3000000a1000000af000000b5000000b3000000b1",
            INIT_09 => X"000000bd000000cf000000d4000000dd000000dc000000c5000000b8000000ab",
            INIT_0A => X"0000008b00000067000000950000008c00000097000000b10000009400000093",
            INIT_0B => X"00000083000000700000008a0000009c00000097000000b1000000d9000000ea",
            INIT_0C => X"000000df000000da000000c6000000b2000000c2000000c2000000be000000c8",
            INIT_0D => X"000000ba000000b8000000bf000000c7000000cb000000d0000000c8000000b1",
            INIT_0E => X"000000ab000000870000007f0000009e000000a80000009b000000830000008f",
            INIT_0F => X"000000890000007e000000940000009f00000093000000900000009e000000c5",
            INIT_10 => X"000000e1000000dd000000d0000000b7000000bf000000c7000000be000000c2",
            INIT_11 => X"000000c6000000bc000000be000000ba000000ab000000c1000000c6000000bf",
            INIT_12 => X"000000cf000000bf00000094000000a9000000a0000000870000007b0000008d",
            INIT_13 => X"0000008e000000950000009f0000009800000087000000880000008c0000009a",
            INIT_14 => X"000000de000000dd000000d6000000be000000b3000000c3000000c8000000be",
            INIT_15 => X"000000c6000000cd000000d1000000b200000097000000b3000000b6000000b5",
            INIT_16 => X"000000c5000000c4000000ae000000a5000000860000007c0000008900000093",
            INIT_17 => X"00000099000000a1000000990000008b000000830000008b0000008b0000007d",
            INIT_18 => X"000000db000000da000000db000000c6000000aa000000bf000000d2000000cf",
            INIT_19 => X"000000cb000000ce000000cf000000b40000009c000000ae000000b4000000b0",
            INIT_1A => X"000000b6000000b5000000b0000000960000006f0000007d0000009600000098",
            INIT_1B => X"00000098000000a10000009a0000008a0000008a00000080000000730000006a",
            INIT_1C => X"000000da000000d6000000d9000000cf000000aa000000bc000000d2000000d5",
            INIT_1D => X"000000d4000000d3000000c7000000b6000000ae000000ba000000ba000000b5",
            INIT_1E => X"000000ba000000b6000000ab0000008500000072000000890000009a00000095",
            INIT_1F => X"00000094000000ab0000009f00000092000000900000007b0000007300000076",
            INIT_20 => X"000000d8000000d4000000d4000000d1000000b3000000bd000000cf000000cd",
            INIT_21 => X"000000cd000000cd000000b10000008a000000a7000000c3000000bb000000b6",
            INIT_22 => X"000000b9000000b50000009e000000820000007d0000008d000000960000008c",
            INIT_23 => X"0000008d000000a30000009d000000950000008500000083000000820000007c",
            INIT_24 => X"000000d7000000d2000000d0000000c8000000bb000000be000000ce000000cc",
            INIT_25 => X"000000c6000000c4000000830000005000000091000000c2000000b8000000ae",
            INIT_26 => X"000000ae000000a50000009300000083000000780000008b0000008f00000088",
            INIT_27 => X"000000890000008e0000008c0000008800000085000000850000007900000070",
            INIT_28 => X"000000d7000000d0000000cd000000c2000000b5000000b7000000cd000000d1",
            INIT_29 => X"000000cc000000c200000081000000510000008e000000ba000000ab000000a1",
            INIT_2A => X"000000a10000009500000089000000780000007300000087000000890000007e",
            INIT_2B => X"000000850000007b000000700000007a0000008a000000880000008300000080",
            INIT_2C => X"000000d6000000cd000000c8000000bc000000b0000000af000000c6000000d4",
            INIT_2D => X"000000d0000000c0000000a00000008e000000aa000000a80000009b00000095",
            INIT_2E => X"0000008d000000850000007f000000640000007100000083000000800000007b",
            INIT_2F => X"0000007e000000720000006c0000007200000082000000900000009000000089",
            INIT_30 => X"000000d2000000c4000000c0000000b7000000a9000000a6000000c0000000d2",
            INIT_31 => X"000000d1000000c0000000b6000000b4000000ab000000990000008d0000008c",
            INIT_32 => X"000000860000007d0000006f0000005c000000780000007e0000007e0000007f",
            INIT_33 => X"0000007e00000072000000690000007400000085000000900000008d00000081",
            INIT_34 => X"000000c4000000b3000000b3000000b9000000a600000097000000b5000000cc",
            INIT_35 => X"000000cd000000c2000000ba000000b3000000a6000000920000008500000088",
            INIT_36 => X"0000007e000000720000005d0000006100000078000000730000007800000080",
            INIT_37 => X"0000008000000071000000710000007e0000008400000083000000820000007b",
            INIT_38 => X"000000b1000000a1000000aa000000b8000000ae0000008c0000009c000000c3",
            INIT_39 => X"000000c9000000c1000000bf000000b600000091000000710000006c00000073",
            INIT_3A => X"000000760000006a000000590000006e00000072000000700000007800000083",
            INIT_3B => X"0000007b0000007a0000007f0000007c000000750000007a0000008200000086",
            INIT_3C => X"0000009d0000008c00000097000000a1000000a60000008200000080000000b1",
            INIT_3D => X"000000bf000000b7000000af0000009a00000070000000530000004700000053",
            INIT_3E => X"000000630000005e000000650000006e0000006c0000006c000000790000007e",
            INIT_3F => X"000000790000007a0000006f0000006b00000073000000840000008900000084",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY51;


    MEM_IFMAP_LAYER0_ENTITY52 : if BRAM_NAME = "ifmap_layer0_entity52" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000170000001c000000130000002800000071000000730000006d00000074",
            INIT_01 => X"00000071000000670000006a000000690000006900000069000000690000006b",
            INIT_02 => X"0000006a000000630000004c0000003a00000054000000560000007200000089",
            INIT_03 => X"0000007c0000007d0000007c0000007d0000007f0000007d0000007a00000078",
            INIT_04 => X"000000180000001b000000140000001a0000006a00000082000000760000007c",
            INIT_05 => X"0000007d000000720000006d0000007500000078000000760000007200000079",
            INIT_06 => X"00000085000000830000006a000000440000003e000000510000008c00000096",
            INIT_07 => X"0000008a0000008c000000890000008800000088000000850000008100000080",
            INIT_08 => X"000000180000001a00000017000000120000005800000083000000740000007b",
            INIT_09 => X"0000008b0000008d0000007400000074000000810000007f0000007d00000084",
            INIT_0A => X"0000008e0000009a000000980000006900000037000000590000009f0000009e",
            INIT_0B => X"0000009700000097000000920000008e0000008e0000008b0000008800000084",
            INIT_0C => X"00000018000000190000001900000012000000450000007c0000006a00000073",
            INIT_0D => X"0000009c000000a6000000920000007800000089000000940000009500000097",
            INIT_0E => X"000000960000009c000000940000006d0000004a0000007a000000b1000000a9",
            INIT_0F => X"000000a10000009d00000098000000950000009600000094000000910000008e",
            INIT_10 => X"00000019000000180000001900000017000000330000006d0000006000000068",
            INIT_11 => X"000000a1000000b8000000b20000008d0000007c000000800000008600000093",
            INIT_12 => X"0000009700000096000000890000006c0000006000000098000000b7000000b5",
            INIT_13 => X"000000b3000000ae000000a8000000a4000000a00000009c0000009800000093",
            INIT_14 => X"0000001a0000001a0000001b0000001c00000023000000590000005f00000066",
            INIT_15 => X"00000096000000c1000000c70000009f00000074000000660000006200000076",
            INIT_16 => X"0000008200000083000000770000007a00000084000000a7000000a6000000aa",
            INIT_17 => X"000000b2000000b7000000b3000000b7000000b7000000b1000000af000000a9",
            INIT_18 => X"0000001a00000016000000190000001a0000001d0000005c000000800000007b",
            INIT_19 => X"00000093000000c3000000c7000000ab0000007e0000005e000000630000006a",
            INIT_1A => X"000000600000006d000000650000007a000000ac000000c0000000aa000000b0",
            INIT_1B => X"000000c3000000c4000000c5000000ca000000c5000000bf000000bf000000c2",
            INIT_1C => X"0000004d000000210000001100000019000000580000009a0000009b0000007e",
            INIT_1D => X"0000008c000000be000000c1000000b9000000a3000000810000007b00000071",
            INIT_1E => X"00000058000000670000006800000079000000b1000000c6000000a5000000bd",
            INIT_1F => X"000000e4000000db000000e0000000da000000ba000000bb000000c4000000cd",
            INIT_20 => X"000000950000008000000056000000600000009b000000a70000009900000077",
            INIT_21 => X"0000006f000000a8000000bf000000bf000000b7000000aa000000940000007f",
            INIT_22 => X"0000007000000070000000740000007c000000a3000000bb000000a2000000c1",
            INIT_23 => X"000000df000000d5000000cf000000bb0000009d000000a6000000c4000000d2",
            INIT_24 => X"000000a10000009e000000920000009b000000a7000000a90000009f00000075",
            INIT_25 => X"000000680000009b000000b3000000b5000000b6000000b40000009f00000087",
            INIT_26 => X"000000640000007400000075000000790000009e000000b2000000b2000000cc",
            INIT_27 => X"000000d8000000d6000000cb000000a70000009300000096000000b0000000cf",
            INIT_28 => X"000000aa000000a50000009e000000a5000000af000000b0000000a000000070",
            INIT_29 => X"0000007b000000a4000000b1000000b4000000b6000000ac0000009500000079",
            INIT_2A => X"0000006a0000007400000075000000760000009c000000a6000000af000000d1",
            INIT_2B => X"000000de000000d8000000cd000000a900000091000000930000009f000000ba",
            INIT_2C => X"000000ac000000ae000000a9000000a6000000b0000000b00000009d0000007a",
            INIT_2D => X"0000008d000000b1000000b9000000b6000000b60000009d0000007f00000068",
            INIT_2E => X"00000073000000840000007b0000007d0000009f000000a4000000a3000000ce",
            INIT_2F => X"000000e0000000d9000000cd000000b5000000920000008e000000930000009c",
            INIT_30 => X"000000a7000000a7000000a5000000a0000000a5000000a4000000990000008f",
            INIT_31 => X"00000091000000a3000000ae000000a4000000a30000009f0000008500000076",
            INIT_32 => X"000000860000009f0000008700000092000000a3000000a3000000a8000000cd",
            INIT_33 => X"000000df000000dc000000d6000000c7000000a3000000900000009000000098",
            INIT_34 => X"000000a9000000a2000000a00000009b000000a30000008800000083000000a4",
            INIT_35 => X"000000920000008800000084000000850000009f0000009e0000008700000092",
            INIT_36 => X"000000a7000000a2000000900000009e0000009800000098000000b0000000cb",
            INIT_37 => X"000000d7000000d8000000dd000000da000000c50000009f000000a2000000b6",
            INIT_38 => X"000000ae000000a4000000a20000009d000000a8000000780000006d000000b2",
            INIT_39 => X"000000a6000000a7000000a1000000a3000000b6000000ab0000008400000078",
            INIT_3A => X"000000a9000000a30000008c00000095000000a6000000a4000000aa000000cc",
            INIT_3B => X"000000d3000000d5000000da000000e4000000d6000000b0000000bb000000c7",
            INIT_3C => X"000000af000000a0000000a10000009f000000aa0000008400000068000000b7",
            INIT_3D => X"000000bc000000b6000000b8000000b0000000a2000000a8000000a30000008d",
            INIT_3E => X"00000091000000a50000009200000085000000af000000a500000096000000a9",
            INIT_3F => X"000000ca000000d4000000d9000000dd000000c4000000ba000000c7000000c7",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY52;


    MEM_IFMAP_LAYER0_ENTITY53 : if BRAM_NAME = "ifmap_layer0_entity53" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b30000009f0000009200000094000000a1000000970000006d000000a8",
            INIT_01 => X"000000c7000000b5000000a4000000ae000000a50000009c000000aa000000a6",
            INIT_02 => X"00000069000000880000009f000000770000008f0000009e0000007e00000050",
            INIT_03 => X"00000076000000b7000000d1000000cd000000af000000b7000000c9000000c5",
            INIT_04 => X"000000b5000000a4000000850000008300000095000000a5000000970000009f",
            INIT_05 => X"000000c2000000c7000000c4000000cd000000b9000000a8000000ac000000a2",
            INIT_06 => X"00000068000000690000009b0000007700000086000000ad000000880000005c",
            INIT_07 => X"0000004b0000006f000000980000009e00000098000000b0000000cb000000c8",
            INIT_08 => X"000000b7000000ac0000008e000000850000009f000000b0000000b1000000aa",
            INIT_09 => X"000000b1000000c5000000cf000000d9000000d9000000c6000000bb000000aa",
            INIT_0A => X"000000830000005a000000850000007e0000008b000000a2000000820000007e",
            INIT_0B => X"0000006f0000006000000076000000840000007c00000092000000b8000000c7",
            INIT_0C => X"000000b9000000b0000000a100000095000000af000000b7000000b6000000bc",
            INIT_0D => X"000000aa000000aa000000b9000000c2000000c9000000d0000000ca000000af",
            INIT_0E => X"000000a40000007b00000071000000910000009d0000008c000000710000007b",
            INIT_0F => X"0000007700000070000000860000008e0000007f0000007900000084000000a6",
            INIT_10 => X"000000bd000000b7000000ad0000009b000000ab000000ba000000b1000000b2",
            INIT_11 => X"000000b4000000ac000000b2000000b1000000a4000000bc000000c3000000bd",
            INIT_12 => X"000000c9000000b6000000880000009d00000093000000780000006a0000007c",
            INIT_13 => X"000000800000008a000000940000008a00000078000000770000007a00000082",
            INIT_14 => X"000000bd000000bc000000b7000000a10000009e000000b7000000bb000000b0",
            INIT_15 => X"000000b8000000bf000000c0000000a40000008b000000a6000000ad000000b1",
            INIT_16 => X"000000c0000000bc000000a200000096000000760000006b0000007900000085",
            INIT_17 => X"0000008e000000960000008d0000007d000000750000007c0000007d0000006c",
            INIT_18 => X"000000ba000000ba000000bb000000a600000094000000b4000000c7000000c5",
            INIT_19 => X"000000c1000000c3000000c0000000a8000000910000009f000000a9000000aa",
            INIT_1A => X"000000af000000ac000000a3000000860000005d0000006c000000860000008b",
            INIT_1B => X"0000008d000000970000008e0000007c0000007c00000072000000650000005b",
            INIT_1C => X"000000ba000000b5000000b7000000ac0000008f000000b0000000c9000000cf",
            INIT_1D => X"000000ce000000cb000000bd000000af000000a5000000ab000000ae000000ac",
            INIT_1E => X"000000b2000000ab0000009e0000007500000061000000780000008a00000088",
            INIT_1F => X"0000008a000000a10000009200000084000000820000006d0000006400000068",
            INIT_20 => X"000000b8000000b2000000af000000a900000092000000aa000000c6000000ca",
            INIT_21 => X"000000c8000000c5000000ab00000088000000a1000000b4000000ab000000aa",
            INIT_22 => X"000000ad000000a800000090000000730000006c0000007c000000860000007e",
            INIT_23 => X"000000820000009900000091000000870000007700000075000000740000006f",
            INIT_24 => X"000000b8000000b0000000a80000009d00000093000000a2000000c0000000c8",
            INIT_25 => X"000000bf000000b900000081000000520000008d000000b3000000a60000009f",
            INIT_26 => X"0000009f000000960000008400000074000000690000007a0000007f0000007a",
            INIT_27 => X"0000007f00000084000000800000007a00000077000000770000006b00000062",
            INIT_28 => X"000000b8000000ac000000a3000000940000008600000092000000ba000000ca",
            INIT_29 => X"000000c0000000b200000082000000580000008c000000ac0000009800000090",
            INIT_2A => X"00000091000000840000007a0000006900000064000000770000007900000070",
            INIT_2B => X"0000007a00000071000000640000006c0000007c0000007a0000007500000072",
            INIT_2C => X"000000b7000000a90000009e0000008e0000007e00000084000000b2000000cc",
            INIT_2D => X"000000c3000000af0000009d00000090000000a4000000980000008700000083",
            INIT_2E => X"0000007c000000740000006f000000540000006100000073000000710000006d",
            INIT_2F => X"00000072000000660000005f000000640000007400000082000000820000007b",
            INIT_30 => X"000000b1000000a1000000990000008e000000770000007a000000b2000000cc",
            INIT_31 => X"000000c5000000b4000000aa000000a80000009d000000870000007a0000007b",
            INIT_32 => X"000000770000006d0000005e0000004b000000680000006f0000007000000071",
            INIT_33 => X"00000070000000640000005c0000006600000077000000820000007e00000073",
            INIT_34 => X"000000a3000000900000008d00000091000000740000006b000000a9000000c8",
            INIT_35 => X"000000c2000000b7000000ac000000a300000096000000810000007300000079",
            INIT_36 => X"00000070000000640000004e0000005100000068000000650000006a00000072",
            INIT_37 => X"000000720000006300000063000000700000007600000075000000740000006e",
            INIT_38 => X"0000008e0000007e000000830000008f0000007c0000005f00000091000000c0",
            INIT_39 => X"000000be000000b7000000b2000000a800000082000000620000005c00000065",
            INIT_3A => X"000000680000005c0000004b0000005f00000063000000610000006a00000074",
            INIT_3B => X"0000006d0000006c000000710000006e000000670000006c0000007400000077",
            INIT_3C => X"0000007b000000680000007000000078000000740000005700000076000000ae",
            INIT_3D => X"000000b5000000ae000000a40000008d00000063000000450000003900000046",
            INIT_3E => X"000000570000005100000058000000600000005d0000005e0000006b00000070",
            INIT_3F => X"0000006b0000006c000000610000005d00000065000000760000007b00000076",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY53;


    MEM_IFMAP_LAYER0_ENTITY54 : if BRAM_NAME = "ifmap_layer0_entity54" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d9000000d2000000cd000000c7000000da000000d6000000cf000000bd",
            INIT_01 => X"000000bb000000ae000000a6000000a9000000960000009a0000008c0000008f",
            INIT_02 => X"000000a7000000bf000000db000000df000000db000000d7000000e2000000e1",
            INIT_03 => X"000000db000000be000000af000000bb000000c8000000aa000000a1000000a2",
            INIT_04 => X"000000de000000dd000000dc000000d7000000d8000000e1000000d3000000b3",
            INIT_05 => X"000000b4000000c0000000be000000bc000000c7000000ce000000d1000000db",
            INIT_06 => X"000000e5000000eb000000ec000000ec000000e9000000e2000000e1000000e5",
            INIT_07 => X"000000e7000000d4000000d0000000cd000000d8000000b7000000ba000000c8",
            INIT_08 => X"000000ea000000e9000000e7000000e8000000e9000000ef000000d9000000ad",
            INIT_09 => X"000000a4000000b4000000ad000000b7000000be000000bc000000d4000000e0",
            INIT_0A => X"000000da000000eb000000e3000000e1000000e5000000df000000d6000000e1",
            INIT_0B => X"000000ea000000e8000000e6000000d8000000d1000000ca000000d0000000d3",
            INIT_0C => X"000000f5000000f4000000f4000000f2000000f4000000f3000000e40000009e",
            INIT_0D => X"000000920000009d000000830000009f0000009100000088000000a20000009f",
            INIT_0E => X"000000a9000000cb000000c3000000d3000000d1000000cb000000d0000000e2",
            INIT_0F => X"000000e6000000e9000000e4000000d5000000c7000000db000000e0000000d4",
            INIT_10 => X"000000f5000000f3000000f4000000f4000000f5000000f1000000cf00000075",
            INIT_11 => X"000000630000006c000000590000006b000000640000005b000000640000005c",
            INIT_12 => X"000000660000007c0000007c00000095000000b6000000b9000000ca000000e9",
            INIT_13 => X"000000e1000000e2000000e3000000cd000000c2000000d5000000e2000000de",
            INIT_14 => X"000000f5000000f4000000f4000000f3000000f5000000ed000000d80000007e",
            INIT_15 => X"000000480000005a0000005b0000006600000065000000670000006b00000063",
            INIT_16 => X"00000059000000590000005b0000005d0000007e000000be000000d8000000eb",
            INIT_17 => X"000000e7000000df000000d8000000c4000000ae000000bd000000d9000000ec",
            INIT_18 => X"000000f5000000f3000000f3000000f4000000f1000000db000000d90000009e",
            INIT_19 => X"000000500000007200000084000000970000008c000000840000008f0000008a",
            INIT_1A => X"000000820000007a00000072000000780000006e0000009b000000dd000000e9",
            INIT_1B => X"000000eb000000e0000000c6000000c0000000a7000000ab000000cc000000eb",
            INIT_1C => X"000000f4000000f3000000f3000000f6000000e3000000c7000000d700000099",
            INIT_1D => X"0000005100000092000000bb000000ca000000cf0000009e0000008300000083",
            INIT_1E => X"000000810000008d00000083000000840000009f000000840000009f000000d7",
            INIT_1F => X"000000e5000000d7000000d4000000d1000000c5000000ab000000b2000000dd",
            INIT_20 => X"000000f4000000f3000000f4000000f5000000e3000000ce000000da00000082",
            INIT_21 => X"00000051000000820000008000000081000000b800000091000000740000007d",
            INIT_22 => X"0000007c000000890000008e0000007d000000990000009300000090000000c6",
            INIT_23 => X"000000d6000000db000000e9000000dc000000b8000000a4000000a9000000c9",
            INIT_24 => X"000000f3000000f3000000f4000000f2000000e4000000be000000a80000006e",
            INIT_25 => X"0000005300000086000000770000006e0000008f000000800000007300000078",
            INIT_26 => X"0000007d00000083000000920000007d000000950000009b0000008c000000c4",
            INIT_27 => X"000000e9000000f0000000f0000000e9000000c8000000c8000000d7000000dc",
            INIT_28 => X"000000ef000000f1000000f4000000f5000000dc00000085000000820000005f",
            INIT_29 => X"0000004e00000074000000740000006c0000006d0000006b0000006d0000006c",
            INIT_2A => X"0000007300000078000000780000007300000088000000960000008f000000a7",
            INIT_2B => X"000000d0000000e4000000f5000000f3000000f4000000f5000000f5000000f4",
            INIT_2C => X"000000de000000e9000000f2000000f4000000d8000000a9000000a500000059",
            INIT_2D => X"0000003d000000430000005b000000640000005f0000005f0000006200000060",
            INIT_2E => X"000000600000005f0000005a000000610000006900000079000000810000007e",
            INIT_2F => X"0000009b000000d8000000f8000000f3000000f4000000f4000000f4000000f4",
            INIT_30 => X"000000d0000000df000000ec000000e3000000bf000000b7000000b500000064",
            INIT_31 => X"000000370000003800000058000000650000006f000000630000005600000054",
            INIT_32 => X"00000052000000540000005d000000710000006d000000620000007000000081",
            INIT_33 => X"000000ae000000e2000000f5000000f4000000f4000000f4000000f4000000f4",
            INIT_34 => X"000000c8000000cc000000db000000c3000000aa0000009a0000009c00000066",
            INIT_35 => X"00000068000000630000006c0000006600000073000000750000005e00000055",
            INIT_36 => X"0000005a0000006a0000007a0000008c00000080000000680000006c0000007c",
            INIT_37 => X"00000096000000b3000000c3000000d4000000ef000000f5000000f4000000f4",
            INIT_38 => X"000000c8000000d2000000cf000000a9000000a400000094000000930000008a",
            INIT_39 => X"000000810000005c0000006a0000005d000000590000005d000000540000004d",
            INIT_3A => X"0000004c0000005100000051000000510000004f0000004a0000004b00000052",
            INIT_3B => X"000000650000007b0000008c0000008f000000bf000000f4000000f4000000f4",
            INIT_3C => X"000000d2000000e2000000c4000000770000007000000096000000ba000000c0",
            INIT_3D => X"0000006c0000004d0000004d000000370000002d0000002f0000003c0000003f",
            INIT_3E => X"0000003b0000003f0000003b0000003600000031000000320000003d00000040",
            INIT_3F => X"000000470000004b0000005b0000006700000087000000e1000000f6000000f4",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY54;


    MEM_IFMAP_LAYER0_ENTITY55 : if BRAM_NAME = "ifmap_layer0_entity55" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000c7000000c1000000b4000000600000005d00000091000000c0000000a1",
            INIT_01 => X"00000056000000490000005c00000062000000680000004f0000004f00000047",
            INIT_02 => X"000000250000001c0000001e0000001b0000003400000032000000160000001c",
            INIT_03 => X"00000018000000350000005b0000006800000080000000ce000000f7000000f3",
            INIT_04 => X"000000d3000000c7000000c200000071000000780000009d0000009f00000047",
            INIT_05 => X"000000440000005a000000740000007c00000095000000790000008000000066",
            INIT_06 => X"0000004e00000062000000700000006400000094000000930000005c00000063",
            INIT_07 => X"0000005e0000006c000000870000008e0000009c000000b7000000f2000000f5",
            INIT_08 => X"000000dc000000ca000000b7000000660000006e000000a5000000840000001e",
            INIT_09 => X"00000039000000620000006b0000005300000052000000650000008100000064",
            INIT_0A => X"00000099000000ae0000009e0000009f000000ac000000a8000000a2000000a3",
            INIT_0B => X"000000a0000000af0000009c000000770000007200000087000000e4000000f7",
            INIT_0C => X"000000db000000cf000000bc00000062000000530000008d0000006f0000002a",
            INIT_0D => X"0000003a000000480000004c0000003e0000003500000038000000400000005d",
            INIT_0E => X"000000a00000007c0000005b00000065000000740000006b0000006700000067",
            INIT_0F => X"000000630000009b0000007e000000430000005100000076000000d9000000f8",
            INIT_10 => X"000000d9000000d2000000c70000006500000038000000580000005d0000003c",
            INIT_11 => X"000000380000002e0000003f000000460000003c000000360000004000000041",
            INIT_12 => X"0000006300000072000000690000006700000064000000600000005d00000061",
            INIT_13 => X"000000660000006f00000064000000490000005200000072000000d4000000f9",
            INIT_14 => X"000000d1000000cd000000ca0000007500000053000000460000005100000044",
            INIT_15 => X"00000032000000230000002b00000033000000440000004d000000570000003f",
            INIT_16 => X"0000003400000047000000520000004800000040000000430000003e0000005d",
            INIT_17 => X"000000580000003c000000530000006c000000700000006c000000cc000000fa",
            INIT_18 => X"000000cd000000ca000000c5000000680000005d0000006f0000004700000049",
            INIT_19 => X"0000003f0000002900000026000000220000004b000000630000008e0000004f",
            INIT_1A => X"0000001e00000056000000930000007600000063000000720000006600000099",
            INIT_1B => X"000000b20000003f0000004a0000008d000000770000005a000000c3000000f6",
            INIT_1C => X"000000c6000000c2000000b900000057000000310000006c0000006100000063",
            INIT_1D => X"0000005f00000033000000270000002400000028000000320000005700000037",
            INIT_1E => X"000000200000004f000000970000007f0000007a00000088000000740000009c",
            INIT_1F => X"0000009f00000037000000350000004a0000003e0000004e000000c2000000f0",
            INIT_20 => X"000000b6000000b4000000a90000004d000000250000003b0000006c00000090",
            INIT_21 => X"0000006a0000003c0000002b000000200000001d0000001c0000001e00000021",
            INIT_22 => X"000000270000002a0000003a000000580000006a000000790000007a00000075",
            INIT_23 => X"000000430000002f00000033000000320000003300000050000000ba000000e1",
            INIT_24 => X"000000a8000000a5000000a40000007d0000005b000000600000006f0000008d",
            INIT_25 => X"000000600000004a00000037000000240000001e0000001e0000001d0000001f",
            INIT_26 => X"000000230000001800000040000000ae000000cd000000cb000000b3000000b5",
            INIT_27 => X"00000057000000260000002b00000030000000420000005b000000ae000000d3",
            INIT_28 => X"000000a2000000a3000000af000000b400000098000000760000006c0000008d",
            INIT_29 => X"0000005b000000530000004e000000300000001900000018000000190000001d",
            INIT_2A => X"000000270000002600000047000000a4000000b8000000b1000000a9000000a6",
            INIT_2B => X"000000510000001e0000001e000000310000004e0000005f000000a9000000ce",
            INIT_2C => X"0000009a000000ac000000b3000000a600000092000000750000006700000092",
            INIT_2D => X"00000057000000550000005200000036000000200000001e0000002100000025",
            INIT_2E => X"000000360000004d00000056000000650000006b000000790000008e00000089",
            INIT_2F => X"0000003c0000001e00000021000000360000004e0000005b000000a5000000c7",
            INIT_30 => X"000000a6000000a90000009e000000940000008f000000850000006700000071",
            INIT_31 => X"0000004f000000510000004b0000003c0000002a000000270000002a0000002c",
            INIT_32 => X"0000003000000036000000410000004d0000005a0000006e000000830000008b",
            INIT_33 => X"000000350000001d0000002600000036000000460000005b000000a9000000c4",
            INIT_34 => X"000000a200000097000000930000008d00000089000000850000006b0000004e",
            INIT_35 => X"000000480000004e000000460000003c000000320000002a0000002e00000030",
            INIT_36 => X"00000031000000330000003b000000420000004c000000590000006500000071",
            INIT_37 => X"000000450000001d00000023000000340000003f00000062000000ae000000ba",
            INIT_38 => X"000000940000008d0000008e0000008c0000008f0000008c0000006a0000003c",
            INIT_39 => X"000000420000004a00000042000000370000003900000034000000360000003a",
            INIT_3A => X"0000003a0000003a00000041000000460000004900000050000000570000005d",
            INIT_3B => X"0000004d0000002500000026000000370000004a00000083000000b3000000b4",
            INIT_3C => X"0000009000000095000000a0000000a20000009e000000920000007e0000003d",
            INIT_3D => X"00000039000000390000003a0000004300000046000000450000004900000048",
            INIT_3E => X"000000440000004900000059000000620000005e000000610000006300000061",
            INIT_3F => X"0000005200000045000000400000004700000077000000a4000000b6000000ba",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY55;


    MEM_IFMAP_LAYER0_ENTITY56 : if BRAM_NAME = "ifmap_layer0_entity56" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d7000000d0000000d0000000ca000000d7000000d1000000ca000000b9",
            INIT_01 => X"000000b8000000a800000098000000a00000009d000000a70000009a0000009d",
            INIT_02 => X"000000b5000000cb000000e1000000e1000000de000000db000000e5000000e4",
            INIT_03 => X"000000dd000000c5000000b8000000c4000000d0000000b8000000b0000000a5",
            INIT_04 => X"000000e2000000e0000000e1000000d9000000d5000000dd000000cc000000ab",
            INIT_05 => X"000000b4000000bd000000b2000000b1000000c4000000cd000000d0000000e0",
            INIT_06 => X"000000ec000000f0000000f2000000f3000000ee000000e5000000e4000000e7",
            INIT_07 => X"000000e7000000d6000000d4000000d2000000de000000be000000bf000000c5",
            INIT_08 => X"000000eb000000ea000000ea000000eb000000ea000000ef000000d6000000a6",
            INIT_09 => X"000000a6000000b1000000a8000000b1000000b8000000b7000000ce000000df",
            INIT_0A => X"000000dc000000ec000000e3000000e8000000eb000000e4000000d9000000e0",
            INIT_0B => X"000000e9000000e9000000e6000000dd000000d9000000ce000000d1000000d2",
            INIT_0C => X"000000f5000000f4000000f4000000f3000000f4000000f4000000e300000099",
            INIT_0D => X"000000920000009b000000820000009f000000900000008a000000a2000000a0",
            INIT_0E => X"000000ac000000cd000000c2000000dc000000de000000d3000000d3000000e0",
            INIT_0F => X"000000e6000000e9000000e5000000db000000cf000000df000000e2000000d4",
            INIT_10 => X"000000f5000000f4000000f4000000f4000000f5000000f0000000cd00000070",
            INIT_11 => X"000000620000006d0000005b0000006d000000650000005c000000640000005c",
            INIT_12 => X"000000680000007d0000007c0000009a000000c2000000c2000000c9000000e3",
            INIT_13 => X"000000dc000000de000000e3000000d3000000cb000000dc000000e8000000e1",
            INIT_14 => X"000000f5000000f4000000f4000000f3000000f6000000eb000000d40000007b",
            INIT_15 => X"000000470000005d0000005f00000069000000670000006a0000006e00000066",
            INIT_16 => X"0000005b000000590000005b0000005d00000081000000c5000000d9000000e6",
            INIT_17 => X"000000dd000000da000000d6000000c6000000b4000000c5000000e2000000ed",
            INIT_18 => X"000000f5000000f3000000f3000000f4000000f0000000d6000000d50000009c",
            INIT_19 => X"0000004f00000077000000890000009a000000900000008b0000009b00000096",
            INIT_1A => X"0000008e00000080000000790000007e00000072000000a0000000e1000000e9",
            INIT_1B => X"000000e9000000da000000c0000000ba000000a5000000b0000000d4000000ec",
            INIT_1C => X"000000f4000000f3000000f3000000f7000000e2000000c1000000d300000096",
            INIT_1D => X"0000005100000098000000bc000000c8000000cd000000a50000008d00000090",
            INIT_1E => X"0000008e000000960000008d0000008f000000a70000008c000000a3000000d6",
            INIT_1F => X"000000e0000000d1000000d3000000d2000000c7000000ae000000af000000dc",
            INIT_20 => X"000000f4000000f3000000f4000000f5000000e1000000ca000000d80000007f",
            INIT_21 => X"00000051000000860000008400000087000000b9000000970000007c00000087",
            INIT_22 => X"00000086000000910000009600000088000000a40000009e0000008e000000c0",
            INIT_23 => X"000000cf000000d8000000e7000000d7000000b10000009e0000009c000000c4",
            INIT_24 => X"000000f2000000f2000000f4000000f2000000e3000000bd000000a80000006e",
            INIT_25 => X"000000530000008c000000800000007600000093000000870000007c00000081",
            INIT_26 => X"000000850000008b00000097000000860000009e000000a400000091000000c1",
            INIT_27 => X"000000e5000000ef000000ef000000e6000000c1000000be000000cc000000d7",
            INIT_28 => X"000000e8000000ef000000f3000000f4000000da00000081000000800000005e",
            INIT_29 => X"0000004f0000007a0000007a0000007000000071000000700000007300000073",
            INIT_2A => X"0000007c000000800000007f0000007e000000900000009e00000099000000aa",
            INIT_2B => X"000000ce000000e3000000f6000000f4000000f3000000f3000000f5000000f4",
            INIT_2C => X"000000cd000000e3000000f2000000f2000000d3000000a10000009f00000058",
            INIT_2D => X"0000003c000000450000005e0000006600000062000000610000006700000066",
            INIT_2E => X"00000068000000640000005f00000067000000710000007f0000008900000080",
            INIT_2F => X"00000099000000d7000000f8000000f3000000f4000000f4000000f4000000f4",
            INIT_30 => X"000000bc000000d5000000e4000000dc000000b4000000aa000000ad00000063",
            INIT_31 => X"00000037000000390000005a0000006600000072000000670000005800000055",
            INIT_32 => X"00000055000000550000005d0000007300000070000000650000007600000086",
            INIT_33 => X"000000b0000000e1000000f5000000f4000000f4000000f4000000f4000000f4",
            INIT_34 => X"000000b8000000bc000000ca000000b500000098000000860000008d00000063",
            INIT_35 => X"00000067000000660000006f0000006700000076000000780000006000000056",
            INIT_36 => X"0000005c0000006b0000007d00000092000000840000006a0000006e0000007f",
            INIT_37 => X"00000098000000b3000000c3000000d2000000ee000000f5000000f4000000f4",
            INIT_38 => X"000000b6000000c2000000bd00000098000000920000007b0000007f0000007e",
            INIT_39 => X"0000007c0000005d000000690000005e0000005a0000005d000000550000004f",
            INIT_3A => X"0000004e000000530000005400000055000000510000004b0000004c00000053",
            INIT_3B => X"000000650000007a0000008a0000008a000000bc000000f4000000f4000000f4",
            INIT_3C => X"000000bd000000cc000000a700000065000000650000007d000000a9000000ae",
            INIT_3D => X"000000670000004d0000004f000000360000002b0000002f0000003b0000003e",
            INIT_3E => X"0000003b0000003e00000039000000340000002f000000300000003d00000040",
            INIT_3F => X"000000460000004a0000005a0000006100000080000000df000000f6000000f4",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY56;


    MEM_IFMAP_LAYER0_ENTITY57 : if BRAM_NAME = "ifmap_layer0_entity57" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ae000000a40000009700000054000000520000007c000000ac00000092",
            INIT_01 => X"0000005300000049000000570000005a000000640000004b0000004c00000044",
            INIT_02 => X"00000021000000170000001a00000017000000300000002f0000001400000019",
            INIT_03 => X"0000001500000032000000560000006400000078000000ca000000f7000000f3",
            INIT_04 => X"000000c0000000b4000000b30000006800000068000000870000008e00000040",
            INIT_05 => X"00000041000000570000006c0000007800000095000000760000007d00000062",
            INIT_06 => X"00000046000000590000006a0000006000000090000000900000005900000060",
            INIT_07 => X"0000005a00000067000000820000008b00000097000000b2000000f1000000f4",
            INIT_08 => X"000000d1000000bd000000ab0000005e0000006200000092000000760000001c",
            INIT_09 => X"000000360000005f000000670000004f0000005300000064000000800000005f",
            INIT_0A => X"00000092000000aa0000009b0000009e000000ab000000a8000000a0000000a1",
            INIT_0B => X"0000009e000000ac0000009b000000770000006f00000080000000e2000000f7",
            INIT_0C => X"000000d0000000c1000000b00000005b0000004c0000007f0000006400000028",
            INIT_0D => X"0000003500000044000000490000003900000032000000350000003d00000059",
            INIT_0E => X"0000009c00000077000000570000006200000071000000680000006300000064",
            INIT_0F => X"00000060000000980000007a0000003f0000004d00000070000000d6000000f8",
            INIT_10 => X"000000ca000000c3000000be0000005f000000330000004e0000005300000038",
            INIT_11 => X"00000033000000270000003c0000004400000039000000330000003b0000003d",
            INIT_12 => X"0000005f0000006e0000006600000065000000630000005f0000005c00000060",
            INIT_13 => X"000000640000006c00000060000000460000004f0000006c000000d0000000f9",
            INIT_14 => X"000000c2000000c0000000c00000006e0000004c0000003e000000490000003f",
            INIT_15 => X"0000002e0000001d00000028000000300000004100000048000000530000003b",
            INIT_16 => X"00000030000000430000004d000000430000003c000000400000003b00000058",
            INIT_17 => X"00000052000000360000004e000000690000006b00000065000000c9000000f9",
            INIT_18 => X"000000c3000000be000000bb0000006100000055000000630000004100000043",
            INIT_19 => X"0000003a00000026000000230000002000000048000000600000008d0000004c",
            INIT_1A => X"000000190000004f0000008c000000710000005e0000006d0000006100000092",
            INIT_1B => X"000000ab0000003a000000450000008a0000007400000053000000c0000000f4",
            INIT_1C => X"000000bd000000b7000000b0000000520000002c00000063000000590000005e",
            INIT_1D => X"0000005a000000300000002400000021000000260000002f0000005500000034",
            INIT_1E => X"0000001c0000004a000000910000007b00000077000000860000007100000097",
            INIT_1F => X"0000009c0000003300000032000000470000003b00000047000000c0000000ee",
            INIT_20 => X"000000ae000000ad000000a3000000480000002200000036000000650000008b",
            INIT_21 => X"000000660000003a000000280000001e0000001a000000190000001a0000001e",
            INIT_22 => X"0000002500000026000000350000005600000068000000750000007600000072",
            INIT_23 => X"0000003e0000002b000000300000002e0000002f0000004b000000b8000000df",
            INIT_24 => X"000000a2000000a00000009e0000007800000057000000590000006700000088",
            INIT_25 => X"0000005c0000004800000034000000220000001c0000001b0000001b0000001d",
            INIT_26 => X"00000020000000150000003d000000af000000cf000000ca000000b1000000b4",
            INIT_27 => X"0000005400000022000000280000002c0000003e00000057000000ab000000d1",
            INIT_28 => X"0000009c0000009c000000a8000000b000000093000000700000006600000088",
            INIT_29 => X"00000056000000510000004b0000002d0000001600000016000000170000001a",
            INIT_2A => X"000000230000002200000045000000a4000000b9000000b1000000a9000000a5",
            INIT_2B => X"0000004e000000190000001a0000002d0000004b0000005c000000a7000000cc",
            INIT_2C => X"00000095000000a7000000ad000000a10000008d00000071000000630000008e",
            INIT_2D => X"00000053000000530000004f000000330000001d0000001c0000001f00000022",
            INIT_2E => X"0000003200000048000000510000006100000066000000740000008a00000085",
            INIT_2F => X"000000370000001b0000001d000000320000004c00000059000000a4000000c6",
            INIT_30 => X"000000a4000000a60000009b000000900000008b00000082000000630000006c",
            INIT_31 => X"0000004c00000050000000480000003800000026000000240000002700000029",
            INIT_32 => X"0000002d000000330000003d0000004800000054000000670000007c00000083",
            INIT_33 => X"000000310000001a00000021000000320000004500000059000000a9000000c3",
            INIT_34 => X"000000a000000094000000920000008d00000087000000820000006600000049",
            INIT_35 => X"000000450000004d00000042000000380000002f000000280000002b0000002d",
            INIT_36 => X"0000002e00000030000000360000003d00000046000000540000005e0000006a",
            INIT_37 => X"000000400000001a0000001f000000300000003d00000062000000af000000ba",
            INIT_38 => X"000000930000008d0000008e0000008c0000008f0000008b0000006800000039",
            INIT_39 => X"000000400000004a0000003f0000003400000037000000310000003300000036",
            INIT_3A => X"00000036000000360000003d00000042000000440000004a0000005100000057",
            INIT_3B => X"000000480000002100000023000000340000004800000084000000b6000000b5",
            INIT_3C => X"0000009200000096000000a1000000a30000009d000000910000007c0000003a",
            INIT_3D => X"0000003700000038000000390000004100000043000000420000004600000045",
            INIT_3E => X"0000004300000048000000570000005f0000005c0000005f000000600000005e",
            INIT_3F => X"00000051000000440000003e0000004600000076000000a3000000b6000000b9",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY57;


    MEM_IFMAP_LAYER0_ENTITY58 : if BRAM_NAME = "ifmap_layer0_entity58" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d1000000ca000000bf000000b6000000d1000000d1000000c6000000af",
            INIT_01 => X"000000ab000000a50000009d000000a0000000950000009a0000008d0000008f",
            INIT_02 => X"000000a4000000bc000000d6000000db000000d1000000ca000000d9000000d6",
            INIT_03 => X"000000d0000000b1000000a1000000ad000000b70000009d0000009500000095",
            INIT_04 => X"000000d4000000d4000000d2000000cd000000cf000000db000000c8000000a3",
            INIT_05 => X"000000a5000000b6000000b8000000b6000000c2000000c9000000cd000000d7",
            INIT_06 => X"000000df000000e3000000e3000000e4000000dd000000d4000000d3000000d7",
            INIT_07 => X"000000df000000cd000000c3000000bb000000c6000000aa000000ad000000ba",
            INIT_08 => X"000000e6000000e5000000e3000000e2000000e3000000ec000000d3000000a4",
            INIT_09 => X"0000009f000000ad000000b7000000b8000000bc000000bf000000cf000000e0",
            INIT_0A => X"000000db000000e5000000e0000000d6000000d6000000d0000000c8000000d3",
            INIT_0B => X"000000de000000e0000000db000000c5000000b9000000bc000000c5000000c6",
            INIT_0C => X"000000f5000000f4000000f4000000f1000000f2000000f1000000e3000000af",
            INIT_0D => X"000000a8000000b0000000a1000000bb000000ae000000a0000000b8000000b6",
            INIT_0E => X"000000b9000000d5000000d0000000ca000000b9000000ba000000c4000000d4",
            INIT_0F => X"000000d7000000dc000000d5000000bb000000a9000000c5000000d4000000c8",
            INIT_10 => X"000000f5000000f3000000f4000000f4000000f5000000f1000000cd00000084",
            INIT_11 => X"0000008b000000a10000008a000000a70000009f0000008b0000009b0000008d",
            INIT_12 => X"0000008e000000a600000099000000a4000000a9000000a9000000c4000000e0",
            INIT_13 => X"000000d1000000d1000000d4000000b1000000a0000000b8000000cc000000d2",
            INIT_14 => X"000000f5000000f4000000f4000000f3000000f6000000ee000000d700000081",
            INIT_15 => X"000000710000009c000000a0000000aa000000aa000000aa000000b1000000a7",
            INIT_16 => X"0000009d0000009d000000980000008f00000094000000b3000000cd000000e4",
            INIT_17 => X"000000da000000ce000000c1000000aa00000093000000a0000000c0000000df",
            INIT_18 => X"000000f5000000f3000000f3000000f4000000f1000000dd000000dd000000b4",
            INIT_19 => X"00000083000000b4000000c4000000cf000000c8000000cb000000d9000000d3",
            INIT_1A => X"000000cc000000c3000000c0000000bf000000a3000000a6000000cd000000e1",
            INIT_1B => X"000000e3000000d5000000b1000000a90000009100000092000000b2000000da",
            INIT_1C => X"000000f4000000f2000000f2000000f7000000e6000000ca000000d9000000c0",
            INIT_1D => X"00000086000000c2000000e0000000e8000000ea000000d7000000ce000000d1",
            INIT_1E => X"000000cf000000d0000000ca000000cf000000e0000000b40000009a000000cc",
            INIT_1F => X"000000dc000000c9000000c4000000bc000000ab000000920000009a000000c7",
            INIT_20 => X"000000f5000000f3000000f3000000f5000000e3000000d1000000df000000ae",
            INIT_21 => X"00000087000000ba000000c1000000c1000000dd000000cc000000c1000000c9",
            INIT_22 => X"000000ca000000cd000000cd000000c6000000dc000000d0000000a3000000bc",
            INIT_23 => X"000000cb000000d1000000df000000cb000000a10000008b00000094000000b2",
            INIT_24 => X"000000f2000000f1000000f3000000f2000000e5000000cd000000c2000000a4",
            INIT_25 => X"0000008c000000c1000000bd000000b8000000ca000000c4000000c0000000c4",
            INIT_26 => X"000000c7000000ca000000d0000000c6000000d7000000e0000000bc000000c8",
            INIT_27 => X"000000e6000000ee000000ed000000e3000000bc000000ba000000ca000000d3",
            INIT_28 => X"000000ea000000ee000000f3000000f4000000df000000a0000000a90000009c",
            INIT_29 => X"00000086000000b1000000b3000000ac000000ae000000ae000000b4000000b7",
            INIT_2A => X"000000bb000000be000000bc000000be000000cd000000dc000000d0000000c4",
            INIT_2B => X"000000d9000000e6000000f6000000f4000000f4000000f4000000f4000000f4",
            INIT_2C => X"000000d3000000e6000000f2000000f2000000d8000000b6000000be00000097",
            INIT_2D => X"0000006a0000006e00000093000000a00000009e0000009f000000a6000000aa",
            INIT_2E => X"000000a9000000a30000009e000000a6000000ad000000bd000000c6000000af",
            INIT_2F => X"000000b7000000e0000000f8000000f3000000f4000000f4000000f4000000f4",
            INIT_30 => X"000000c4000000da000000e9000000e1000000bd000000b4000000c30000009f",
            INIT_31 => X"0000005d0000005c0000008d000000a0000000ba000000a80000008f0000008c",
            INIT_32 => X"0000008b0000008900000092000000a700000098000000830000008f00000096",
            INIT_33 => X"000000bc000000e3000000f3000000f4000000f4000000f4000000f4000000f4",
            INIT_34 => X"000000c3000000c7000000d3000000c1000000a400000095000000a200000089",
            INIT_35 => X"00000096000000aa000000b2000000a6000000bd000000cd000000a600000092",
            INIT_36 => X"00000099000000ac000000c0000000d3000000af00000080000000800000008a",
            INIT_37 => X"000000a0000000b1000000bf000000d3000000ef000000f5000000f3000000f3",
            INIT_38 => X"000000c2000000cf000000c8000000a20000009c000000880000008e00000089",
            INIT_39 => X"000000a2000000b2000000b10000009f00000096000000a3000000950000008b",
            INIT_3A => X"0000008d000000920000009200000093000000860000007c0000007f00000085",
            INIT_3B => X"00000095000000a3000000ad000000a6000000cc000000f5000000f3000000f4",
            INIT_3C => X"000000c3000000d0000000ad0000006e000000710000008b000000b4000000b9",
            INIT_3D => X"000000850000009a0000007f00000057000000490000004c000000590000005f",
            INIT_3E => X"0000005c000000600000005e0000005800000056000000560000006300000067",
            INIT_3F => X"0000006d000000740000008f0000009b000000af000000e8000000f5000000f5",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY58;


    MEM_IFMAP_LAYER0_ENTITY59 : if BRAM_NAME = "ifmap_layer0_entity59" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b7000000aa000000a1000000650000006000000088000000b5000000a1",
            INIT_01 => X"000000800000008400000081000000870000008c0000007d0000007d0000006a",
            INIT_02 => X"000000350000002b0000002c000000270000004d000000470000002300000028",
            INIT_03 => X"00000020000000500000009100000097000000a7000000db000000f6000000f3",
            INIT_04 => X"000000ca000000c1000000c20000007c00000078000000920000009900000049",
            INIT_05 => X"00000069000000870000008300000094000000b80000009f000000a900000083",
            INIT_06 => X"0000006600000076000000840000007a000000af000000aa0000006f00000073",
            INIT_07 => X"0000006f00000091000000b2000000b5000000bb000000c5000000f2000000f4",
            INIT_08 => X"000000d8000000c8000000b800000072000000730000009d0000008200000024",
            INIT_09 => X"0000004f0000009500000081000000630000006f000000810000009d00000084",
            INIT_0A => X"000000b1000000c1000000b7000000b9000000c8000000c1000000ba000000bd",
            INIT_0B => X"000000b5000000c7000000b60000009700000094000000a2000000e8000000f6",
            INIT_0C => X"000000d9000000cc000000bb00000071000000600000008b000000710000003d",
            INIT_0D => X"0000004e00000070000000730000005d00000055000000530000005e0000007d",
            INIT_0E => X"000000bf0000009f0000007f0000008a000000a0000000950000008c0000008f",
            INIT_0F => X"0000008a000000bd0000009f00000063000000730000009a000000e2000000f7",
            INIT_10 => X"000000d5000000d0000000c700000075000000490000005c0000006300000054",
            INIT_11 => X"0000004b0000004100000061000000690000005f00000057000000670000005f",
            INIT_12 => X"00000086000000a200000099000000970000009600000090000000890000008f",
            INIT_13 => X"00000093000000990000008f0000006f0000007300000092000000de000000f7",
            INIT_14 => X"000000cc000000ce000000cc0000008300000065000000510000005c0000005a",
            INIT_15 => X"000000460000002d0000003900000045000000620000006f0000007d00000057",
            INIT_16 => X"0000004a00000066000000700000006700000062000000650000005e0000007d",
            INIT_17 => X"000000730000005200000071000000950000009a00000089000000d4000000f8",
            INIT_18 => X"000000d1000000d0000000ce00000075000000690000007a000000560000005e",
            INIT_19 => X"0000005600000036000000330000002f0000006600000083000000ad00000063",
            INIT_1A => X"0000002d000000640000009e00000082000000790000008a0000007c000000ab",
            INIT_1B => X"000000bb0000004b0000005f000000ab0000009800000075000000cf000000fa",
            INIT_1C => X"000000dd000000d6000000cc000000680000003b000000740000007200000080",
            INIT_1D => X"0000007c00000041000000340000003000000038000000460000006c0000004b",
            INIT_1E => X"000000300000005f000000a60000008f00000091000000a70000008f000000af",
            INIT_1F => X"000000af0000004a00000048000000620000005400000068000000d6000000fb",
            INIT_20 => X"000000d7000000d4000000c9000000630000002f0000004400000080000000b0",
            INIT_21 => X"0000008700000050000000380000002d00000028000000270000002b0000002f",
            INIT_22 => X"000000370000003c000000500000006e0000007d00000093000000900000008b",
            INIT_23 => X"0000005c000000430000004600000043000000450000006d000000d9000000fb",
            INIT_24 => X"000000cf000000cf000000cb0000009d000000730000007500000085000000aa",
            INIT_25 => X"0000007e0000006500000048000000300000002800000029000000290000002d",
            INIT_26 => X"000000320000002700000053000000c0000000da000000dc000000c7000000c9",
            INIT_27 => X"0000006b00000034000000380000003f0000005a0000007e000000d2000000f7",
            INIT_28 => X"000000bc000000c0000000ce000000d8000000bf0000009a00000086000000a1",
            INIT_29 => X"0000007900000073000000680000003e00000021000000220000002300000029",
            INIT_2A => X"000000330000003100000055000000b3000000c7000000c0000000be000000bb",
            INIT_2B => X"000000600000002700000026000000420000006f00000085000000d1000000f5",
            INIT_2C => X"000000bf000000c6000000cd000000c6000000b50000009e00000084000000a0",
            INIT_2D => X"00000072000000760000006f0000004600000027000000260000002c00000031",
            INIT_2E => X"000000440000005d000000690000007e0000008700000096000000ad000000a6",
            INIT_2F => X"00000048000000280000002a000000470000007100000082000000cf000000f2",
            INIT_30 => X"000000ce000000d1000000c6000000b8000000ab000000a30000008200000085",
            INIT_31 => X"0000006b0000006f000000680000004d000000320000002f0000003500000039",
            INIT_32 => X"0000003f0000004800000057000000680000007800000091000000a8000000b0",
            INIT_33 => X"00000045000000280000003000000047000000660000007e000000d4000000ee",
            INIT_34 => X"000000c7000000c2000000c2000000bd000000b2000000a60000008600000065",
            INIT_35 => X"0000006300000069000000600000004f0000003e000000360000003b0000003e",
            INIT_36 => X"00000041000000450000004e000000570000006400000074000000810000008f",
            INIT_37 => X"00000057000000270000002c000000470000005900000085000000df000000e8",
            INIT_38 => X"000000c1000000bc000000be000000bc000000bd000000bc0000009000000050",
            INIT_39 => X"0000005a00000063000000580000004600000049000000450000004a0000004e",
            INIT_3A => X"0000004e0000004e000000560000005d00000061000000660000006d00000072",
            INIT_3B => X"0000005e00000030000000300000004a00000064000000ad000000e8000000e7",
            INIT_3C => X"000000c4000000c7000000d0000000cd000000c8000000bb000000a500000055",
            INIT_3D => X"0000004c0000004c0000004e0000005400000054000000590000006200000063",
            INIT_3E => X"0000005e00000063000000720000007c0000007d00000081000000800000007f",
            INIT_3F => X"000000700000005b000000540000006000000094000000cc000000e1000000df",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY59;


    MEM_GOLD_LAYER0_ENTITY0 : if BRAM_NAME = "gold_layer0_entity0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a000000012000000400000010400000051000000bc0000010100000000",
            INIT_01 => X"0000000000000047000000000000001c0000000000000000000000ba00000000",
            INIT_02 => X"0000000000000000000000000000003100000000000000000000009200000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000104000000000000000000000002",
            INIT_05 => X"0000000000000000000000000000000000000000000000a80000000000000038",
            INIT_06 => X"0000000000000000000000000000000000000000000000020000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000530000003700000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_0A => X"00000000000000a80000017a00000134000000370000011300000082000000b7",
            INIT_0B => X"0000003500000000000000000000002d00000079000000000000014d00000062",
            INIT_0C => X"00000000000000000000000000000000000000000000007e0000001000000035",
            INIT_0D => X"000000000000006a00000000000000d100000000000000000000000000000000",
            INIT_0E => X"000000b0000000b000000000000000a00000003300000077000000d200000081",
            INIT_0F => X"000000c6000000000000000000000008000000a9000000570000000000000065",
            INIT_10 => X"000000c800000000000000a10000003c00000000000000580000007a00000000",
            INIT_11 => X"000000000000000000000006000000000000005c000000000000000000000000",
            INIT_12 => X"000000000000002c000000e600000000000000770000004800000000000000ff",
            INIT_13 => X"0000002400000000000000000000001900000000000000360000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"00000000000000000000005d0000004d000000b50000006c000000aa00000000",
            INIT_17 => X"000000000000000000000000000000000000003f000000000000001b00000030",
            INIT_18 => X"0000001500000000000000000000000000000119000000b30000000000000012",
            INIT_19 => X"00000000000000aa00000000000000bd000000b6000000260000000000000000",
            INIT_1A => X"0000002800000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"00000000000000c000000124000001440000014f000000d00000006800000017",
            INIT_1D => X"0000000000000040000000000000000000000009000000570000001600000000",
            INIT_1E => X"000000cf0000005d000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000a800000001000000b8",
            INIT_21 => X"0000001e00000028000000960000009000000015000000630000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000011b0000009e",
            INIT_24 => X"00000000000000000000006c0000000000000000000000000000000000000079",
            INIT_25 => X"000000f80000004300000004000000ff00000067000000120000001100000000",
            INIT_26 => X"000000000000001c00000000000000690000004100000000000000860000004e",
            INIT_27 => X"000000310000000000000000000000910000006c000000510000001700000026",
            INIT_28 => X"0000004600000000000000b0000000fd000000e0000000000000007800000000",
            INIT_29 => X"00000010000000000000000000000000000000000000000000000059000000ab",
            INIT_2A => X"000000c1000000fb000000ef0000006a0000008f000000db0000003b00000053",
            INIT_2B => X"000000140000001000000000000000000000007b00000046000000ab00000062",
            INIT_2C => X"0000005a0000013c000000a20000006d0000008c0000007a0000012300000051",
            INIT_2D => X"00000097000000a1000000000000000000000000000000000000003c00000000",
            INIT_2E => X"0000000700000000000000000000000000000000000000000000000000000104",
            INIT_2F => X"000000000000000000000000000000000000001e0000004f000000a20000012f",
            INIT_30 => X"0000008c00000000000000000000015b0000013a0000016100000083000000a1",
            INIT_31 => X"00000072000001380000001200000000000000000000008800000070000000dc",
            INIT_32 => X"000000e0000000ad0000013e000000cd000000ae000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000000000000000000000000000c80000001f",
            INIT_34 => X"000000bf000000460000004b0000004e0000001b00000026000000000000001e",
            INIT_35 => X"000000730000013b0000009f000000360000001e00000006000000aa000000a5",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"000000000000000000000000000000000000006a000000430000007600000101",
            INIT_3B => X"000000660000007c000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000059",
            INIT_3D => X"000000690000000000000031000000000000000000000000000000000000003d",
            INIT_3E => X"0000000000000000000000100000003100000072000000ed0000000000000000",
            INIT_3F => X"000000000000000000000000000000000000000000000000000000700000012c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY0;


    MEM_GOLD_LAYER0_ENTITY1 : if BRAM_NAME = "gold_layer0_entity1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000017f000000d0000000000000000000000000000000000000003200000000",
            INIT_01 => X"00000067000000080000003900000021000000de0000006d0000004400000076",
            INIT_02 => X"0000008400000141000000eb0000000000000000000000000000000000000000",
            INIT_03 => X"00000000000000000000000000000000000000b2000000780000006e0000003f",
            INIT_04 => X"0000007f0000009200000000000000000000000000000000000000000000001c",
            INIT_05 => X"00000191000000000000001e0000003400000087000001480000000000000000",
            INIT_06 => X"000000000000000000000000000000000000000000000000000000580000004a",
            INIT_07 => X"0000004600000000000000000000000000000000000000f3000000d7000000c5",
            INIT_08 => X"000000000000000000000000000000000000000000000000000001180000006b",
            INIT_09 => X"00000000000000000000003100000000000000fe0000003a00000071000001a4",
            INIT_0A => X"00000130000000b6000000000000000000000000000000000000000000000000",
            INIT_0B => X"000000e300000000000000f30000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000001690000004d000000c7",
            INIT_0E => X"000000f5000000aa0000002a0000000000000100000000780000005200000000",
            INIT_0F => X"00000000000000000000000000000076000001c0000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000007d00000000",
            INIT_12 => X"0000000000000000000000110000000000000000000000000000000000000074",
            INIT_13 => X"00000000000000c80000013900000006000000b9000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"000000000000000000000000000000000000000000000000000000000000005c",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"00000000000000000000000000000000000000450000000000000000000000c3",
            INIT_19 => X"000000eb0000016c000001a1000001d5000000d4000001b4000001db00000149",
            INIT_1A => X"0000000000000000000000000000007c000000830000005c0000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000007900000176000000d1000000a0000000d40000004d0000020300000255",
            INIT_1E => X"000002180000022a00000270000001b600000129000000000000006300000000",
            INIT_1F => X"0000000000000000000000000000005900000000000000000000000000000000",
            INIT_20 => X"00000000000000000000003d000000da00000000000000000000000000000000",
            INIT_21 => X"000000a80000004a000000dd0000005f00000148000001d60000002200000000",
            INIT_22 => X"0000000000000000000000af00000000000000000000000e000000900000018a",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000f9000000d40000009000000042000001370000013d",
            INIT_26 => X"00000138000000b7000000160000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000001450000019b000000b8",
            INIT_29 => X"000001150000014f00000106000000000000002c000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"000000000000000000000000000000b90000016d0000019d000000000000029f",
            INIT_2C => X"000000000000000000000000000000000000000000000000000000fb00000121",
            INIT_2D => X"000000fa00000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"000000d30000000000000000000000d0000000830000009f0000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"000000000000000000000000000000000000000000000000000000000000003d",
            INIT_32 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000000000006f000000380000000000000000",
            INIT_34 => X"000000340000003400000000000000000000008b00000000000000790000007a",
            INIT_35 => X"0000018e00000143000000a00000005400000000000000000000000000000000",
            INIT_36 => X"0000000000000090000000e4000001240000009a000000a4000000c200000000",
            INIT_37 => X"00000028000000a6000000000000000800000000000000000000000000000000",
            INIT_38 => X"0000006f0000000b00000000000000e4000000db000000ec0000016e0000009d",
            INIT_39 => X"0000005f000001d9000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000008b0000001f",
            INIT_3C => X"0000001c00000000000000000000000000000033000000000000000000000000",
            INIT_3D => X"00000000000000000000000000000000000000000000000e0000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000011b00000000",
            INIT_3F => X"00000000000000000000000000000000000000000000000000000000000000c1",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY1;


    MEM_GOLD_LAYER0_ENTITY2 : if BRAM_NAME = "gold_layer0_entity2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009f00000093000000000000000000000000000000000000000000000000",
            INIT_01 => X"000000f500000000000000dc0000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000c5000000f50000006f",
            INIT_04 => X"0000009e0000003c000000d60000000000000000000000210000000000000000",
            INIT_05 => X"000000000000000000000000000000480000026000000161000000d30000018f",
            INIT_06 => X"00000002000000c1000001a3000000d1000000790000008f000001a40000002f",
            INIT_07 => X"00000000000000000000000000000000000000520000005b00000071000000b2",
            INIT_08 => X"000000000000002d00000062000000b700000096000000e9000000dc00000000",
            INIT_09 => X"0000010500000008000000470000006f000000b0000001c5000001ed000001db",
            INIT_0A => X"000001b6000002dc000001dc0000000000000000000000000000000000000000",
            INIT_0B => X"00000000000000fd000000c00000005300000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000037000000000000000000000000",
            INIT_0D => X"000000000000000000000000000000000000000000000000000001a7000000c7",
            INIT_0E => X"000000c0000000b3000000610000010400000000000000000000007000000000",
            INIT_0F => X"00000045000000c700000167000001c1000001ac00000111000000e3000000d2",
            INIT_10 => X"0000000000000031000000000000000000000000000000000000000000000000",
            INIT_11 => X"00000000000000fe0000009f0000004a000000000000000000000000000000ec",
            INIT_12 => X"000000b300000025000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"000000000000000000000000000000000000000000000084000000000000002b",
            INIT_16 => X"000000c2000001040000008b000000c20000009d0000007400000131000000e1",
            INIT_17 => X"000000b9000000000000000000000000000000f1000000f70000010c00000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000089000000000000002700000061",
            INIT_1C => X"000000000000000700000000000000000000000000000000000000720000006b",
            INIT_1D => X"0000009000000000000000000000000000000000000000000000000000000007",
            INIT_1E => X"000000000000000000000000000000000000001f000000000000000000000030",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"000000030000004300000000000000000000000000000000000000000000018b",
            INIT_21 => X"000000de0000017900000038000000a000000053000001130000010d0000009d",
            INIT_22 => X"0000000000000000000000000000004e00000017000000d70000002500000000",
            INIT_23 => X"000000dc00000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000140000002a0000000d000000000000000000000000",
            INIT_25 => X"00000000000000000000000000000099000000e50000007c000000a0000000df",
            INIT_26 => X"000000a6000000c600000073000000a000000023000000150000000000000023",
            INIT_27 => X"000000000000000000000000000000180000001a000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000003600000000000000820000007300000057",
            INIT_29 => X"0000015800000018000000450000001e000000660000009c0000008c00000000",
            INIT_2A => X"00000000000000000000000000000067000000000000001c0000005100000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_2D => X"000000000000000000000181000000cf000000d000000000000000c5000000d5",
            INIT_2E => X"000000b1000000cf000000620000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000a2000000b400000029",
            INIT_31 => X"0000009f0000005800000053000000940000006c0000006a0000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"000000500000002c0000007e00000000000000000000006300000000000000c0",
            INIT_34 => X"0000000000000000000000000000008500000000000000000000000000000000",
            INIT_35 => X"0000002200000000000000000000000000000067000000b00000001800000012",
            INIT_36 => X"0000004900000030000000000000000000000000000000000000000000000000",
            INIT_37 => X"000000000000001d000000590000003800000028000000000000000000000000",
            INIT_38 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"000000d60000007700000071000000000000000b000000100000000000000011",
            INIT_3B => X"000000000000000900000000000000000000000000000000000000080000001f",
            INIT_3C => X"000000000000009200000053000000a2000000830000000000000090000000eb",
            INIT_3D => X"00000054000000cc000000000000000b00000000000000000000000000000000",
            INIT_3E => X"0000000000000093000000db00000090000000b7000000b7000000a900000032",
            INIT_3F => X"0000004d000000200000000c0000001b00000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY2;


    MEM_GOLD_LAYER0_ENTITY3 : if BRAM_NAME = "gold_layer0_entity3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000010000000840000000900000150000001230000011e0000000000000000",
            INIT_01 => X"000000300000006c000000bb0000008900000000000000000000000000000018",
            INIT_02 => X"000000000000004a000000000000000000000000000000000000000000000000",
            INIT_03 => X"000000000000000000000000000000000000000000000000000000a0000000a7",
            INIT_04 => X"0000005100000012000000670000000000000028000000a90000009c00000000",
            INIT_05 => X"000000000000000000000000000000000000000000000000000000000000002e",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000500000000000000000000000000000000",
            INIT_09 => X"0000004800000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"000000000000000000000000000000000000000000000071000000bc00000000",
            INIT_0C => X"000000a5000000c9000000000000005d00000025000000000000000000000000",
            INIT_0D => X"0000002f00000000000000000000000000000075000000310000004900000197",
            INIT_0E => X"000000910000013c0000005b000000470000007f0000001f0000004200000000",
            INIT_0F => X"00000041000000000000004e0000013c0000000e00000000000000ae0000006d",
            INIT_10 => X"0000007d000000b40000000000000116000000a100000001000000000000003e",
            INIT_11 => X"000000000000000e000000fc0000007d000000d9000000fa000000bb00000182",
            INIT_12 => X"00000102000001050000014d0000000000000000000000000000000000000000",
            INIT_13 => X"000000000000003e0000004f0000000a00000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"000000000000001a0000005c0000000000000000000000000000019f000000fc",
            INIT_16 => X"000000c2000000e1000000940000008000000106000000b20000007a000000eb",
            INIT_17 => X"0000010700000011000000a50000008e00000000000000f50000008e00000074",
            INIT_18 => X"000000370000002600000000000000000000000000000000000000a80000014c",
            INIT_19 => X"000000880000000000000000000000000000000000000305000002120000002c",
            INIT_1A => X"000000000000006d0000000000000000000000750000000000000101000000a9",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000012000000c90000005400000000",
            INIT_1D => X"00000000000000000000000000000000000000000000006a0000000000000000",
            INIT_1E => X"000000a0000001aa0000016a0000000000000054000000610000000000000000",
            INIT_1F => X"00000002000000000000000000000000000000a8000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"000000000000000000000000000000e1000000260000001b0000000000000000",
            INIT_23 => X"00000097000000b400000044000000000000002c000000000000000000000083",
            INIT_24 => X"000000000000000000000000000000560000004a000000240000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"00000000000000000000005f0000001300000000000000000000000a00000000",
            INIT_27 => X"00000044000000910000000a0000000000000048000000a30000000000000000",
            INIT_28 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000a900000167000000ac000000bd00000155000001ba",
            INIT_2A => X"0000000c0000009a0000007900000083000000140000000200000000000000a2",
            INIT_2B => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"00000000000000000000000000000000000000000000000e000000800000000a",
            INIT_2D => X"00000027000000000000006e0000004500000107000000ca00000009000000f9",
            INIT_2E => X"000000cd00000266000002bc0000035e000000770000004d00000000000000b5",
            INIT_2F => X"0000005f00000119000000000000000000000000000000000000002500000000",
            INIT_30 => X"0000000000000000000000000000000600000117000000c50000000000000000",
            INIT_31 => X"00000000000000880000005f000000000000008f0000013c0000012500000000",
            INIT_32 => X"000000000000000000000042000000000000001f000000ff0000008a000000b8",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000a40000006b00000000000000000000000000000000",
            INIT_35 => X"00000000000000000000009f000000600000009a000000d90000003400000028",
            INIT_36 => X"0000016800000164000001780000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000c90000011b00000115",
            INIT_39 => X"0000004000000077000001730000007e0000000c000000230000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"000000be000000a2000000000000000000000000000001370000021c0000028e",
            INIT_3C => X"000000000000003e000000490000000000000000000000000000000000000073",
            INIT_3D => X"0000008a000000930000005a00000053000000ff000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"00000000000000000000000000000081000000a700000181000000430000005b",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY3;


    MEM_GOLD_LAYER0_ENTITY4 : if BRAM_NAME = "gold_layer0_entity4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009c00000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000f00000071",
            INIT_02 => X"00000000000000000000000000000000000000000000002d0000000000000000",
            INIT_03 => X"0000000a0000002b0000000000000000000000720000004f00000032000000c7",
            INIT_04 => X"0000003a00000000000000530000000000000000000001db0000017600000128",
            INIT_05 => X"00000083000000cc0000009e0000002c0000003f000001040000008c00000000",
            INIT_06 => X"000000000000012900000064000000000000007b000000000000008a0000007e",
            INIT_07 => X"0000005c0000000a000000000000000000000000000000430000000000000051",
            INIT_08 => X"000000000000000000000000000000210000002b000000000000000000000178",
            INIT_09 => X"000000f100000001000000240000008d00000079000000420000005800000060",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000300000044",
            INIT_0C => X"0000000e00000000000000960000002b00000000000000100000000800000000",
            INIT_0D => X"00000000000000000000001f0000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"000000000000000000000000000000000000000000000000000000000000003b",
            INIT_10 => X"00000000000000000000000000000000000000500000005a000000f800000062",
            INIT_11 => X"0000000000000000000000e20000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"00000000000000000000000000000000000000000000005100000087000000ae",
            INIT_14 => X"0000000000000090000000cf0000011a000000e30000010d0000000000000000",
            INIT_15 => X"00000000000000000000009100000000000000000000005200000138000000ae",
            INIT_16 => X"000000470000005000000000000001970000007c0000006a0000007f000000f9",
            INIT_17 => X"0000002b000000bc00000101000000ef00000000000000000000000000000098",
            INIT_18 => X"000000e3000000000000003d00000021000000000000017b0000010a00000033",
            INIT_19 => X"000001c3000001620000013b00000089000000590000013b000000e700000030",
            INIT_1A => X"00000115000001130000017f0000000000000000000000000000000000000000",
            INIT_1B => X"00000000000000630000009b0000013200000000000000000000000000000000",
            INIT_1C => X"000000a5000000000000000f0000002700000008000001aa000000ca00000000",
            INIT_1D => X"0000016200000000000000000000000000000000000000000000013800000164",
            INIT_1E => X"00000158000000000000009500000192000000320000002d0000015400000042",
            INIT_1F => X"000001140000007c000000490000015e000000da0000012e000002120000026d",
            INIT_20 => X"0000003f00000000000000000000001400000000000000000000000000000076",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"000000000000000b000000000000000900000055000000000000003600000049",
            INIT_23 => X"00000000000000000000009c0000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000002b0000001c000000000000000000000000000000aa0000010d00000000",
            INIT_26 => X"000000e0000000cf000000740000010e000000b10000004e0000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000007100000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"00000000000000340000006100000059000000000000006e0000017c00000032",
            INIT_2B => X"0000000000000100000000c5000000a0000001d3000000ee0000009c000000e8",
            INIT_2C => X"000001900000014e00000075000000ed00000069000000ff000000fc000000e6",
            INIT_2D => X"0000002e00000055000000de00000000000000d4000000650000012600000084",
            INIT_2E => X"000000940000007b000000520000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000005400000000",
            INIT_30 => X"0000000000000000000000000000003e00000000000000000000000800000083",
            INIT_31 => X"0000004f0000000300000000000000000000004c000000730000000000000000",
            INIT_32 => X"0000000000000016000000000000000000000083000000800000003200000000",
            INIT_33 => X"000000000000006900000000000000f500000077000000bf000000ad00000078",
            INIT_34 => X"0000005a0000007900000000000000fb0000001100000000000000a900000076",
            INIT_35 => X"000000370000000000000000000000000000001a000000000000000000000000",
            INIT_36 => X"0000000000000008000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000005a0000002a000000080000000700000000",
            INIT_38 => X"0000001a00000000000000000000001b0000000000000000000000440000008d",
            INIT_39 => X"000000000000003e000000000000000000000000000000600000000000000000",
            INIT_3A => X"0000001000000000000000000000001f0000001b000000660000001000000048",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000097000000370000003d000000590000014a000000be00000086",
            INIT_3D => X"00000073000000e100000000000000000000000000000000000000000000001c",
            INIT_3E => X"00000000000000000000002e0000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY4;


    MEM_GOLD_LAYER0_ENTITY5 : if BRAM_NAME = "gold_layer0_entity5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000000000000000000000000002c0000002a00000089",
            INIT_01 => X"0000004800000037000000810000003900000001000000f80000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000003700000000000000000000003e00000000000000300000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"00000000000000ee000000d1000000b200000152000000d9000000ec0000001b",
            INIT_06 => X"0000008e0000009b000000a6000000de0000006f000000680000000000000042",
            INIT_07 => X"000000000000000000000000000000000000000000000000000000000000000d",
            INIT_08 => X"000000be000000000000003b000000d300000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000dd000001510000015c",
            INIT_0A => X"00000156000000e6000000a9000001150000009c000000000000000000000000",
            INIT_0B => X"000000000000000000000000000000420000000000000000000000120000010e",
            INIT_0C => X"00000052000000780000010f0000000000000000000000af000000080000002b",
            INIT_0D => X"0000000700000000000000000000000000000000000000170000000000000055",
            INIT_0E => X"000000b800000000000000370000000000000000000000470000000000000039",
            INIT_0F => X"000000540000000000000000000000000000000e0000003f0000000000000000",
            INIT_10 => X"0000000000000000000000190000000000000000000000000000000000000000",
            INIT_11 => X"000000000000000000000000000000390000004700000000000000ad00000075",
            INIT_12 => X"000000000000000c0000003f000000f000000000000000000000000000000000",
            INIT_13 => X"000000000000000000000000000000000000000000000000000000f40000010e",
            INIT_14 => X"00000191000001530000000000000000000001a20000016600000000000000d1",
            INIT_15 => X"00000000000000170000003b0000000000000000000000040000001500000039",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000066000000000000000000000085",
            INIT_1B => X"0000003f0000000000000005000000a300000000000000000000004500000000",
            INIT_1C => X"0000000000000000000000600000003c00000000000000000000002800000005",
            INIT_1D => X"0000000000000000000000000000009200000000000000000000006d00000000",
            INIT_1E => X"0000000000000022000000950000003e000000000000004a000000a200000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"000000000000000000000111000000000000003c000000ab00000016000000ce",
            INIT_21 => X"0000000000000000000000c70000007f0000002b00000096000000a500000043",
            INIT_22 => X"000000ba000000dd0000001e000000260000015b000000ab000000d70000003f",
            INIT_23 => X"00000000000000f4000000da00000000000001610000015a00000139000000f2",
            INIT_24 => X"000000b20000011b000001900000007b00000114000000000000000000000000",
            INIT_25 => X"0000009800000000000000000000000000000044000000000000000000000000",
            INIT_26 => X"0000000000000000000000370000000000000023000000a60000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"00000070000000a50000010e000000c600000000000000e0000000de00000089",
            INIT_29 => X"00000083000000190000008600000078000000a0000000510000005400000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000031",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"00000000000000000000000000000000000000e400000118000000cd0000002d",
            INIT_2D => X"000000c4000000000000003b00000091000000960000007d0000000000000000",
            INIT_2E => X"0000007600000026000000000000000000000000000000000000000000000000",
            INIT_2F => X"000000560000000000000000000000d40000003d000000000000002c00000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000480000008a000000be0000005d0000009700000000",
            INIT_33 => X"000000560000004e0000004d000000030000005c0000000000000001000000dd",
            INIT_34 => X"0000001a000000000000002a0000002000000000000000000000005500000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000004100000000",
            INIT_36 => X"0000000000000000000000be0000002f0000002b000000000000000000000000",
            INIT_37 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"000000000000002600000000000000550000000000000049000000b000000000",
            INIT_39 => X"0000000000000000000000000000001e000000220000003e0000009300000025",
            INIT_3A => X"00000034000000540000003d0000004c000000be000000000000000000000029",
            INIT_3B => X"000000000000006d000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"000000000000000000000000000000000000002b0000000000000000000000df",
            INIT_3E => X"00000000000000000000005a00000000000000cf00000086000000000000006d",
            INIT_3F => X"0000001e00000000000000000000003200000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY5;


    MEM_GOLD_LAYER0_ENTITY6 : if BRAM_NAME = "gold_layer0_entity6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000022",
            INIT_01 => X"0000004100000000000000820000002d00000044000000ea0000010e00000000",
            INIT_02 => X"0000000000000000000000270000002f00000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"00000000000000cf00000087000000a4000000de000000c2000000bf000000c3",
            INIT_05 => X"000000cc000000e4000000000000000000000000000000000000000300000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000820000007000000000",
            INIT_09 => X"000000e40000009d00000000000000ae00000073000000100000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"000000000000000000000000000000000000001b000000000000005400000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000031",
            INIT_0D => X"0000007d000000ed0000007e00000072000001090000000000000000000000d3",
            INIT_0E => X"0000002300000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"000000000000000000000000000000ca000000b80000009e000000a600000000",
            INIT_10 => X"0000003a00000066000000000000004e000000920000008f000000830000004e",
            INIT_11 => X"000000060000007c000000db000000b500000136000000000000000000000000",
            INIT_12 => X"00000000000000000000000000000000000000000000004d0000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000004000000000",
            INIT_15 => X"000000bc000000f800000015000000e400000031000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"00000000000000000000000000000000000000000000000000000049000000a5",
            INIT_18 => X"0000006500000000000000000000000000000000000000000000005c00000034",
            INIT_19 => X"000000c40000000000000000000000000000002d000000690000007000000000",
            INIT_1A => X"0000000000000064000000b5000000840000006f000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"000000000000000000000000000000000000000000000000000000000000003b",
            INIT_1D => X"000000000000005c000000c300000000000000bc000000ae0000002a00000078",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000004b00000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"00000000000000000000000000000000000000940000006e000000ae000000b9",
            INIT_23 => X"000000770000012c0000006e000000bc00000077000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000004700000000000000000000001900000000",
            INIT_25 => X"0000005d000000820000007e0000007000000082000000aa000000e300000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000070",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"000000000000000000000115000000ae000000e0000000fe0000014500000116",
            INIT_2A => X"000000590000011c000000f50000000000000000000000000000000000000000",
            INIT_2B => X"000000000000000000000000000000000000005a0000005700000034000000bc",
            INIT_2C => X"000000ac00000096000000640000006600000034000000320000000000000000",
            INIT_2D => X"0000000000000000000000000000004e00000080000000a70000005e0000000b",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"000000250000000000000000000000c100000000000000000000004000000060",
            INIT_30 => X"0000004b00000040000001080000012000000009000000e2000000d300000057",
            INIT_31 => X"000001690000016d0000021500000004000001b9000000000000000000000000",
            INIT_32 => X"000001b7000001da000000000000000000000000000000730000004100000000",
            INIT_33 => X"0000008f000000af000000000000000000000000000000000000000000000000",
            INIT_34 => X"000000000000000000000000000000000000037c000002790000012000000149",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000016000000000",
            INIT_37 => X"000000000000004b000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000080000009e0000013b000001bf000000eb0000003b",
            INIT_3B => X"00000000000000be000000000000000000000000000000000000000000000134",
            INIT_3C => X"0000001e00000142000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000e300000000000000000000000000000069000000d1",
            INIT_3F => X"000000fe000000eb0000000e0000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY6;


    MEM_GOLD_LAYER0_ENTITY7 : if BRAM_NAME = "gold_layer0_entity7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000163000000cc0000016c000000d0000000ca000000b4",
            INIT_01 => X"0000007300000000000000000000000000000065000000260000009400000156",
            INIT_02 => X"00000000000000000000006c0000000000000000000000860000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"000000000000000000000000000001ec0000022f00000042000000db00000262",
            INIT_06 => X"0000005f0000009e0000008c00000000000000c60000017a0000003100000027",
            INIT_07 => X"0000000d00000000000000000000006a0000000000000011000001b700000000",
            INIT_08 => X"000001700000012000000000000000000000000000000000000000510000008c",
            INIT_09 => X"0000014800000082000000c4000000a4000000a1000000970000013900000000",
            INIT_0A => X"0000000000000000000000000000000000000100000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000006200000029000000e60000011c00000109",
            INIT_0D => X"0000009f00000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000002360000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"000000000000000000000000000000000000000000000084000000aa00000033",
            INIT_11 => X"0000004000000000000000000000000000000046000000f50000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"000000c80000000000000194000001f90000008a000000000000000000000000",
            INIT_14 => X"0000028f0000026b0000016a000001d200000356000000000000012700000000",
            INIT_15 => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000008e00000200000000d8000001350000002a000000000000000000000000",
            INIT_18 => X"000000000000000800000000000000000000000000000000000000fb00000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000087000001cf0000003f00000124000000000000001100000000",
            INIT_1B => X"00000000000000f400000112000000000000012d000000000000005900000000",
            INIT_1C => X"0000004f000000880000008400000000000000bc0000000000000000000000c7",
            INIT_1D => X"00000115000001c900000082000001bf0000009a000000000000000000000046",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000008900000000",
            INIT_1F => X"0000017900000000000000000000000000000000000000000000000000000028",
            INIT_20 => X"000000d7000001ba0000019b000000a6000002a2000001a800000374000000b3",
            INIT_21 => X"000001c7000000260000027b00000231000000640000005e0000007a00000053",
            INIT_22 => X"0000005a000000d7000000ca0000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000001a0000009c",
            INIT_25 => X"00000000000000000000002b000000780000005100000000000000b10000009d",
            INIT_26 => X"000000bb00000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000078",
            INIT_28 => X"0000000000000050000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"00000000000000000000000000000000000000ce000000590000012700000017",
            INIT_2B => X"00000000000000b3000000000000000000000037000000000000000000000000",
            INIT_2C => X"000000000000000000000000000000000000000000000000000002240000007f",
            INIT_2D => X"00000040000000f3000000720000000000000175000001680000019800000000",
            INIT_2E => X"0000001100000000000000000000011e00000000000000450000010300000000",
            INIT_2F => X"00000000000000000000000000000000000000b5000000000000000000000078",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000002c8000001de000001340000012c0000026700000182",
            INIT_32 => X"0000015400000138000001650000000000000000000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000ad00000000000000000000000000000010",
            INIT_34 => X"0000000000000000000000590000000000000000000000c30000000000000000",
            INIT_35 => X"0000000000000000000000c10000000000000000000000100000001a00000153",
            INIT_36 => X"00000000000000200000000000000000000000000000000000000000000001a5",
            INIT_37 => X"000001d100000089000001a00000009600000004000000af0000013400000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000330000007500000000000000000000006f00000000",
            INIT_3B => X"000000000000002e000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"000000000000001e00000000000000290000002a0000017e000001b500000155",
            INIT_3E => X"000000bd00000168000001ea000000810000018f000001e8000000000000006f",
            INIT_3F => X"00000000000000000000001600000091000000f1000000d30000003d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY7;


    MEM_GOLD_LAYER0_ENTITY8 : if BRAM_NAME = "gold_layer0_entity8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"00000000000000e700000000000000000000010c0000011400000000000000e3",
            INIT_03 => X"000000b900000000000000fe000000f200000092000000f60000018200000143",
            INIT_04 => X"00000081000001040000013a0000000000000001000000cb0000000000000000",
            INIT_05 => X"0000005c0000000000000000000000210000001a000000360000006900000064",
            INIT_06 => X"00000093000000000000012e000000b300000036000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"00000066000000000000003800000166000000b5000000000000011900000000",
            INIT_0B => X"000000000000004f000000be000000720000001c000001340000009000000000",
            INIT_0C => X"000000890000004e000000240000001100000000000000000000000100000000",
            INIT_0D => X"0000000c000000940000002e000000000000000f0000008a0000000000000000",
            INIT_0E => X"00000000000000a400000000000000000000005e00000060000000000000009f",
            INIT_0F => X"00000000000000810000000000000000000000ae000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"000000000000000000000000000000000000002b000000000000000000000010",
            INIT_12 => X"00000000000000cd0000013d0000002900000000000000600000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"00000000000000000000000000000000000000b100000000000000000000001f",
            INIT_15 => X"000000000000000000000000000000000000002e000000000000000000000000",
            INIT_16 => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000a30000005e00000000",
            INIT_19 => X"00000096000000980000000000000063000000c3000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000018000000000000000000000000000000870000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"00000000000000cd000000db00000146000000d6000000890000010b00000000",
            INIT_1E => X"0000007200000104000000410000000000000000000000000000007100000000",
            INIT_1F => X"000000a7000000d20000001b000000a200000075000000090000005000000130",
            INIT_20 => X"000000c500000000000001150000009400000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000820000000000000045",
            INIT_22 => X"000000fd00000046000000000000000d00000000000000000000000000000000",
            INIT_23 => X"0000003c00000000000000000000001900000000000000000000000000000145",
            INIT_24 => X"0000008800000020000001e6000000660000000e000001720000003900000000",
            INIT_25 => X"00000021000000e60000006900000000000000240000014c0000000000000000",
            INIT_26 => X"0000012200000000000000000000000000000000000000000000006200000000",
            INIT_27 => X"000000000000008b000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000050000003100000000000000000000000000000007",
            INIT_29 => X"000000000000000000000000000000000000000000000050000000b500000055",
            INIT_2A => X"00000000000000d100000000000000000000000b000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000117",
            INIT_2C => X"0000010500000000000000ad000000e800000000000000000000000d00000070",
            INIT_2D => X"0000000000000000000000000000000e000000000000007b0000002f00000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000007c000000bc0000000000000014000000a1",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"000000000000000000000000000000000000007b000000000000000000000014",
            INIT_33 => X"000000210000000000000016000000000000000c000000000000007600000081",
            INIT_34 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_35 => X"000000000000000000000000000000000000006a000000440000000000000062",
            INIT_36 => X"0000007d00000000000000000000003d0000005b000000000000008400000061",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"00000000000000a7000000d10000002d00000000000001240000001b00000012",
            INIT_39 => X"0000011200000025000000570000005d0000008f0000006b0000004b0000007d",
            INIT_3A => X"000001ad0000005700000084000000000000019c000001b100000000000000b9",
            INIT_3B => X"000001f500000091000000eb000001d2000000ae000000b6000000790000007f",
            INIT_3C => X"000001390000005800000095000000fd0000009300000000000000000000003f",
            INIT_3D => X"0000004b000000000000001000000000000000000000000000000016000000dd",
            INIT_3E => X"0000006a0000000000000000000000a900000000000000000000003e00000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY8;


    MEM_GOLD_LAYER0_ENTITY9 : if BRAM_NAME = "gold_layer0_entity9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000140000000a900000035000000a20000004700000045000000af00000049",
            INIT_01 => X"0000009200000000000000000000000000000000000000000000003300000000",
            INIT_02 => X"00000062000000000000000000000000000000aa00000000000000000000001d",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000002e00000050000000000000000000000000",
            INIT_06 => X"000000000000000000000025000000340000001c000000000000000000000033",
            INIT_07 => X"000000000000000000000000000000120000004900000016000000b900000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"00000000000000cf0000009d000000f5000000bc0000001b0000007800000000",
            INIT_0B => X"0000003c0000006400000177000000b10000010c00000101000000db000000ec",
            INIT_0C => X"000000aa000000b800000056000001370000007a00000131000000e8000000a0",
            INIT_0D => X"00000000000000fd0000000e0000007200000020000000a7000000000000000f",
            INIT_0E => X"0000005c00000000000000000000001500000088000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000014b0000001a",
            INIT_10 => X"0000004500000000000000000000000000000000000000000000004d00000018",
            INIT_11 => X"0000000000000000000000000000001200000086000000330000004100000009",
            INIT_12 => X"000000000000000000000005000000000000000000000000000000000000003e",
            INIT_13 => X"000000000000002200000018000000f1000000390000001c0000000000000000",
            INIT_14 => X"0000000000000032000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000450000003000000000000000000000006500000000",
            INIT_17 => X"0000000000000023000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000003200000046",
            INIT_19 => X"0000000000000000000000170000002400000000000000000000000000000060",
            INIT_1A => X"000000000000000000000000000000000000000000000023000000aa00000008",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"000000000000014e0000011a000001730000010d000000bb0000000100000069",
            INIT_1D => X"0000007b0000011e0000000000000000000000480000004b0000000b00000049",
            INIT_1E => X"0000012600000150000000a40000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000120000000b00000021",
            INIT_21 => X"000000dd000000a40000006d00000035000000ab000000a90000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000650000000000000000000000000000000000000000",
            INIT_25 => X"00000007000000100000002f00000064000000e9000000ca0000000000000108",
            INIT_26 => X"000000c00000008a000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000004e00000082000000ab000000cc00000081",
            INIT_28 => X"000000530000006d000000b80000008100000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000001d10000003a000000e6",
            INIT_2A => X"0000008a00000050000000710000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000041000000000000000000000016000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000008400000000000000000000004500000000",
            INIT_2D => X"000000000000000000000089000000920000006800000087000000ce00000033",
            INIT_2E => X"0000000000000021000000b30000000000000056000000460000003600000067",
            INIT_2F => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000004700000000000000000000000000000000",
            INIT_31 => X"00000002000000000000000000000000000000f60000010b000001130000010e",
            INIT_32 => X"0000004c000000000000009f0000000600000048000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000000000000000000000000000c600000000",
            INIT_34 => X"00000026000000a20000000000000027000000770000000000000000000000dc",
            INIT_35 => X"000000b50000019f000000000000001800000000000000490000000f00000069",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000054000000190000000000000000",
            INIT_3B => X"000000550000003c000000000000003800000003000000000000000000000000",
            INIT_3C => X"0000009500000062000000020000000000000010000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000003500000000000000000000004c00000098",
            INIT_3E => X"0000000b000000190000000000000000000000b5000000000000001b00000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY9;


    MEM_GOLD_LAYER0_ENTITY10 : if BRAM_NAME = "gold_layer0_entity10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_01 => X"000000000000001d0000009000000088000000f200000000000000800000006f",
            INIT_02 => X"000000aa000000ef000000f50000000000000000000000000000000000000000",
            INIT_03 => X"00000022000000000000000000000001000000000000000e00000000000000a9",
            INIT_04 => X"0000004b000000970000008a000000a2000000d600000000000000b800000000",
            INIT_05 => X"0000000000000043000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000005800000000000000000000005300000048000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000014100000000000000000000019b0000000e000000000000004e0000010a",
            INIT_09 => X"00000075000000320000004d000000000000013a000001560000012200000000",
            INIT_0A => X"00000172000001d4000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000006000000ce0000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"000000000000000000000000000000000000000000000000000000aa000000c8",
            INIT_0E => X"00000000000000bb000000000000000000000000000000000000016000000044",
            INIT_0F => X"000000000000011c0000000000000000000000000000002c0000006200000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"000000000000000000000000000000000000000000000000000000000000002c",
            INIT_12 => X"00000000000000b30000000000000000000000e5000000000000000000000060",
            INIT_13 => X"00000058000000ec00000000000000000000017400000000000000000000002e",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000057000000000000000000000000000000000000000000000000",
            INIT_16 => X"00000000000000000000002e0000000000000000000000000000000c00000000",
            INIT_17 => X"00000012000000000000006b0000000000000009000000000000000000000000",
            INIT_18 => X"000000000000006c00000021000000290000006e00000082000000000000005f",
            INIT_19 => X"0000008a00000092000001790000017400000191000000bb0000005300000000",
            INIT_1A => X"0000004b00000041000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"00000000000000000000000000000000000000000000003f0000005800000048",
            INIT_1D => X"00000000000000000000000000000000000001730000000000000000000001f8",
            INIT_1E => X"000001ce000000000000009a00000083000000000000003c0000006900000000",
            INIT_1F => X"0000006200000000000000000000000000000000000000000000002c00000000",
            INIT_20 => X"00000000000000150000008900000000000000b8000000ac000000540000006f",
            INIT_21 => X"00000000000000de0000015a000001d9000000c6000001220000008100000019",
            INIT_22 => X"000000000000000000000000000000220000009f000000000000000000000144",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"00000000000000000000000000000000000000920000000000000000000000fb",
            INIT_25 => X"00000000000000000000016900000056000000cb0000018c0000000700000000",
            INIT_26 => X"000000d9000000440000003c0000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"000000000000000000000000000000000000000000000110000000f900000077",
            INIT_29 => X"0000016a0000004300000000000000d700000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000009f0000000000000000000000420000013400000000000000fb000000a9",
            INIT_2C => X"000000000000005400000000000000000000004b000000190000004c00000000",
            INIT_2D => X"0000005800000000000000650000002900000000000000000000000000000063",
            INIT_2E => X"00000000000000000000000000000000000000000000003c0000000000000000",
            INIT_2F => X"0000002b00000004000000810000006400000077000000f20000003800000000",
            INIT_30 => X"00000000000000d7000000000000000000000000000000000000000000000000",
            INIT_31 => X"000000000000000000000000000000000000000000000000000000530000007c",
            INIT_32 => X"00000000000000000000007b0000001a00000054000000000000016100000040",
            INIT_33 => X"0000000000000174000000420000000000000000000000850000000000000017",
            INIT_34 => X"000000180000004a0000002e000000000000004d000000ea0000000000000000",
            INIT_35 => X"0000000f000000000000001a0000000000000098000000000000000000000000",
            INIT_36 => X"000000000000008e000000000000000b00000000000000350000015200000000",
            INIT_37 => X"0000000000000124000000b90000000000000000000000d20000000000000000",
            INIT_38 => X"000000980000000000000074000000520000000b0000005c000001d10000009e",
            INIT_39 => X"0000013100000040000001110000010b00000027000000000000000000000000",
            INIT_3A => X"0000000000000015000001570000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000055000000000000000000000000000000000000000000000000",
            INIT_3D => X"000000000000010d000000000000000000000000000000c70000005d0000004a",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"000000080000000000000000000000000000000000000021000000c200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY10;


    MEM_GOLD_LAYER0_ENTITY11 : if BRAM_NAME = "gold_layer0_entity11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004f0000004300000000000000000000000000000000000000b90000004e",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000006900000000",
            INIT_04 => X"00000000000000db0000010a000000000000000000000000000000000000004d",
            INIT_05 => X"00000000000000be000000220000004800000000000000690000014400000000",
            INIT_06 => X"00000000000000c40000000000000026000000ef000000000000011e00000055",
            INIT_07 => X"00000000000001270000000000000000000000870000004e000000580000007f",
            INIT_08 => X"0000001f00000000000000cf00000000000000aa000000d30000002200000000",
            INIT_09 => X"0000005600000000000000e4000001a8000000ca000001290000017c00000141",
            INIT_0A => X"000000c000000169000001840000000000000000000000000000000000000000",
            INIT_0B => X"000000000000000000000000000000000000000000000000000000000000006f",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000037",
            INIT_0D => X"000000000000000000000000000001020000005e000000000000000000000082",
            INIT_0E => X"0000006400000000000000dc0000000000000000000000000000000000000000",
            INIT_0F => X"000000f90000000000000000000001ba0000018400000000000000ac000000a4",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY11;



end a1;