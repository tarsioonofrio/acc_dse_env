library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package inmem_package is
  type mem is array(0 to 4000000) of integer;

  constant input_mem : mem := (
    -- bias
    -6075, -1035, 250, 3118, 4061, -3808, 5166, -6103, 1262, -3443,

    -- weights
    -- filter=0 channel=0
    0, -2, 3, 7, -1, 2, -2, 5, 7, 5, 2, 3, 1, 2, 4, -2, 3, 1, -7, -2, -3, 7, 0, -2, 0, -3, 0, -5, 7, 2, 0, -3, 7, 1, -8, -10, 0, -5, -2, -9, -3, -5, 1, -3, 0, 3, 6, 3, 1, -24, -25, -17, -13, -28, -9, -18, -9, -26, 14, 2, -8, -26, -12, -21, -11, 3, 7, 9, -8, 3, -1, 9, -4, 15, -12, 7, -2, -4, 2, 10, -3, 4, 7, 2, -3, 1, 4, -3, -6, 3, -3, -4, 5, 1, -2, -6, 15, -11, 0, 0, 4, -3, -10, 6, 7, -2, 0, -10, 7, -12, 20, 6, -2, 1, -10, -10, -6, 0, -4, 0, -2, 7, 1, -6, -6, -1, 4, 5, -7, -2, -10, 0, -3, -1, -3, -6, -9, -10, -13, -2, -2, -11, -12, 4, 6, 2, -10, 1, -10, -6, -11, -14, -7, -9, 2, -18, -5, -8, -9, -23, -13, 0, 11, 27, -20, -10, -16, 25, -21, -18, -14, 15, -8, 0, 4, 21, -7, -13, -8, -15, -15, 14, 9, -2, -23, 4, 1, -9, -17, -28, -15, 11, 6, 5, -3, 5, 3, 7, 0, -8, -6, 4, -3, 0, 3, 4, 0, 7, 2, 4, -3, 4, -5, 0, 7, -2, 2, 5, 6, 5, 6, 7, 0, -5, 1, 10, 3, 16, -2, -5, -12, -11, 3, -11, -19, 7, 0, -12, -4, 8, 14, 8, 7, 15, 16, -2, -5, 1, 19, 12, -8, 15, 4, 2, 7, 20, -5, -2, -5, 7, 6, 0, -1, 1, -5, 6, -6, -3, -6, 3, -4, -4, 0, 4, 0, 0, -4, -14, -4, -2, 1, -5, -7, 19, -13, -3, -8, 5, 12, -1, 9, 0, 6, 0, -16, -4, 13, 1, 0, -6, 12, 7, 14, 6, 10, -2, -21, -10, -5, -2, -2, -3, -6, -13, 15, 14, -10, -14, -10, 2, -7, -9, -3, 1, -8, -15, -2, -7, -20, -23, -5, -3, -11, -3, -9, 7, 0, 3, -5, -4, -4, 8, 15, 7, 0, 11, -2, 14, 3, 5, -1, -9, 20, 5, 13, 4, 13, 4, 5, 10, 8, 3, 0, 18, 11, 0, 3, 3, -7, -2, 10, 4, -4, 12, 3, 0, 0, 4, -1, -5, -7, 0, -1, 1, -4, -4, -6, 5, -4, -7, 0, -4, 6, -5, 0, -4, 3, -9, -4, 1, -2, -1, -2, 5, 6, 1, -3, -9, 3, -3, -3, 6, -6, 2, 6, -4, -4, 3, 6, 14, -7, -6, 6, -2, -10, 0, -8, -9, -8, -8, -4, 0, -15, -13, -11, 5, -6, -10, -13, 3, -15, -13, -3, -6, 2, -16, -10, 1, -5, 3, -2, -1, -10, -4, -7, 0, 0, -5, -6, 1, -7, -4, -2, -5, 1, 5, -14, -4, -7, -2, 7, 17, -4, -5, 3, 22, -3, -10, -11, -7, 22, -3, 3, 27, 25, 6, -10, 25, 21, 15, -11, 19, 14, -2, 9, 25, 2, 6, 0, -7, 4, 1, -6, -2, -5, 4, -4, -6, -6, 5, 7, 6, -9, -3, -13, 6, -21, -13, -5, 8, -22, -23, -9, 1, -3, -7, -7, 17, -6, 0, 0, -5, -10, -2, -4, -6, -9, 2, -3, -4, -12, 2, -5, 1, -2, -7, 1, 0, 6, 2, 5, -5, 4, 6, -4, -3, -1, -3, 5, -3, -14, 2, -3, 8, -15, -13, 2, 2, -14, -12, -11, 5, -7, -13, -7, 10, 0, 1, -5, -4, -6, 5, 1, -1, -6, -4, -7, 1, -3, -3, 1, 2, 9, 1, 3, 1, 15, 1, -2, 11, 5, 8, -1, 5, 8, 0, 7, 4, -10, 7, 4, -6, 3, 4, 3, -8, 0, -5, 0, -1, -4, 1, 1, 4, 0, 1, -18, -17, -3, 2, 1, -14, -8, 0, -17, -3, 5, 2, -5, 8, 21, 12, 23, 5, 10, 5, -1, 8, 4, 6, -4, 0, 9, 0, 2, -12, 1, 0, 5, 13, -12, -15, -4, -1, -6, -8, -8, -6, -1, 4, 5, 2, -13, -18, -13, 8, -37, 28, -3, 5, -41, 32, -9, 7, -18, -21, -24, 22, -10, 0, 13, 32, -12, -12, -6, 13, -6, -3, -15, 10, 0, -1, 6, 32, 6, -8, 0, -7, -7, 1, 3, -5, -1, 13, 7, 9, 2, 6, -12, 7, 14, -6, 0, 2, 0, -8, -11, 10, 15, 0, -10, 0, 10, -2, 4, 19, 12, 8, 5, 24, -3, -4, -13, 15, 8, -9, -18, 17, 0, -3, 2, 13, -2, -4, -9, -12, -2, -20, 8, -3, 0, -17, 4, 4, -8, -2, -8, -7, -3, -7, 2, 8, -19, -15, -11, 8, -14, -15, -6, 4, -12, -7, 6, 19, -8, -9, 0, 1, -7, -13, -8, 3, -15, -10, -6, -5, -7, -7, -16, -5, 9, 1, 11, 7, 4, -7, -6, -4, -2, -15, 4, -2, 2, -9, -3, -4, 11, -3, 6, 18, 15, 12, -17, 14, 5, 4, -9, -12, 2, 7, 14, 2, -4, -3, 3, 0, -7, -2, 5, -3, -4, -15, -9, 1, -14, -1, 9, 12, -7, 5, -4, -6, 4, -4, 2, -3, -3, -1, -7, -6, 0, 3, 5, 0, -4, 1, -2, 1, -3, 0, 2, 6, 3, 5, 5, -5, 4, 0, 3, 1, -12, -16, -5, 1, -12, -11, -12, 11, -22, -21, -8, -3, -9, -16, -3, 16, -1, -5, 0, -5, -20, 0, 8, -11, 0, 0, -26, -1, 11, -2, 4, 11, -6, -1, -3, 6, 0, 0, 4, 0, -2, 0, -4, 4, -7, 3, -7, 6, -6, 2, 8, 3, -7, -2, 6, 0, 0, -4, -3, -8, 0, 2, -7, -4, -14, -5, -2, 8, -22, 20, 6, 4, -22, 17, -5, 4, -12, 0, -17, 17, 20, 8, 11, 21, 19, 1, -8, 21, 4, 8, -17, 18, 5, 1, 6, 16, -6, -13, -9, -11, -11, -4, 12, -9, -12, -6, 9, -6, 1, -7, -11, -9, -3, -1, -7, 0, -5, 9, 2, -8, 0, 0, -10, -11, -5, 0, -16, -3, 2, -2, 5, 5, 11, 1, 8, -6, 10, 0, 1, -4, 3, 5, -2, -11,
    -- filter=0 channel=1
    7, -4, -8, -4, 0, 2, -2, -9, -3, -5, -1, -7, 3, 2, -2, 0, -1, -4, -1, 4, 1, -3, -7, -3, 6, 7, 5, -3, -6, 0, 6, -7, -4, 2, 2, -3, 1, 2, -2, -1, -9, -5, 8, 3, 3, 5, 1, 1, 11, 14, 10, 7, 9, 0, -4, 11, -5, -2, 7, 11, 7, 5, 17, 25, 12, 0, -3, 1, 10, -21, -7, -6, 1, -13, 1, -10, 6, 8, -12, -3, 5, 4, -6, 3, 4, 6, -5, -1, 4, 2, -6, 6, 1, 0, 2, -3, -13, -12, 2, -19, 10, 9, 7, -13, 1, 23, -5, -24, -12, 5, 5, 5, 6, 0, 0, 3, 7, -9, -1, -1, 0, -10, -6, 0, 1, 7, 2, 5, 11, 0, 5, 7, 8, -12, -20, -2, 12, -7, -2, -1, 6, 3, -9, 0, 8, 0, 3, 0, -12, -16, -26, -11, 4, -5, -17, -5, -2, 7, 0, 0, 23, 16, 9, 10, 10, -28, -30, -27, -4, -34, -32, -13, 22, -9, -3, -5, 3, 6, 16, 4, 11, -7, 19, 0, 14, 7, 14, -3, 2, 19, 26, -2, 4, 0, -2, -7, -2, 2, -9, -7, -7, 0, -8, 3, 9, 9, -4, -8, 7, 1, 0, -3, -6, 0, -7, 0, -5, 6, 0, 0, -2, 3, 8, 8, 15, 8, -1, 12, 8, -24, -20, -16, 5, -22, -25, -25, 15, -16, -33, -17, -14, -3, -3, -22, -7, 18, 22, -13, -7, 31, 27, -19, -11, 0, 10, 0, 0, 6, -8, 5, -7, -3, -7, -2, -7, -7, -2, 0, 7, 0, -4, 2, 0, 7, 9, 21, -3, -24, 0, 2, 5, -9, -15, -3, 8, -23, -19, -4, -9, 0, 1, -6, 2, 12, 23, -16, 1, 23, 2, -30, -7, 11, 16, -5, 9, 3, 23, 29, 5, 0, 19, 13, -12, 15, 7, 13, 5, -7, 0, 19, 7, 7, 13, 4, 1, -16, -8, 7, -1, -14, -16, -6, 8, 7, 1, 0, -7, 7, 1, 8, -8, 31, 8, -10, -6, 25, 5, 13, 0, 22, 3, 8, -21, 13, 7, 6, 2, 39, 16, -11, -20, 28, 12, 0, -23, 13, 12, 22, -2, 16, 20, 6, -1, 24, 19, 14, 0, 10, 16, 5, -5, -1, 8, 5, -2, -1, 0, 2, 0, -7, -9, -1, -5, -1, -1, -10, -8, -9, -6, -6, 4, 5, -3, -3, -5, -7, -10, 0, 1, -8, 3, -8, -6, 1, -3, 2, 2, -2, 4, 7, 0, -7, -2, 1, -3, -13, -15, 6, -5, 4, 3, 9, 11, 0, 2, 3, 4, -7, -10, -9, 12, 0, -22, -6, 4, 6, -18, -15, 7, -2, -1, -8, -5, 3, 2, 2, -2, 4, 2, 4, 10, 5, 1, 2, 12, 4, 11, 8, 6, -2, 1, 12, -10, 6, 0, 9, 0, -7, 9, 27, -21, -13, -1, -7, -6, 26, 29, -21, -7, 40, 23, -25, -13, 7, 13, -7, -3, 3, 9, -3, -5, 6, -5, -3, -3, 4, 2, 5, -4, 4, -3, -5, 27, 5, -5, 5, 0, -18, -22, -22, 9, -16, -24, -12, 15, 6, -15, 1, 9, 16, 8, 7, 0, -10, -13, -1, -3, -12, -10, -2, 16, -1, -7, -1, -2, -2, 0, -3, -6, -4, 1, 4, -4, 3, -1, -2, -7, 1, 1, -3, 10, 6, 15, 2, 5, -10, -1, 2, -2, 1, -8, 1, 8, 12, 0, 2, 2, -2, 5, 2, 1, -7, 0, 0, 6, 2, 3, -2, 1, -2, 6, 0, -8, -4, 1, -15, -5, 26, 13, -1, 1, 30, 9, -4, -13, 0, -6, 3, -3, 1, 8, 0, 0, 6, 3, -6, 1, 3, -4, 7, 0, -5, -6, 0, 8, -4, -16, 2, 0, -4, -24, -5, -3, -10, -15, 0, 4, 5, 1, 9, -6, 20, 18, -1, -7, 43, 16, -6, -13, 37, 7, -9, -19, -8, 1, -3, 5, 2, 0, -6, -8, -18, -17, -7, -5, -24, -26, -1, 10, -6, 2, 13, 1, 18, 41, 11, 21, 4, 43, -11, 17, 23, 49, -7, 1, 36, 42, 0, 27, 4, 5, 7, 18, -40, -27, -30, -5, -26, -21, -35, 26, -3, -21, -17, -6, 1, 2, 0, 7, -3, 1, 7, 10, -4, 4, 5, 5, 3, 8, -3, -18, -15, -9, -3, 3, 9, -4, -18, -3, 9, 22, -20, -11, -13, -11, -5, 7, 5, -3, 0, -8, 2, -9, -15, -6, -7, 0, -14, 3, -2, -5, -11, -2, 17, 21, 17, -3, 11, 8, 9, -6, 9, 6, 1, -2, 0, 7, 17, 19, 4, -6, -2, 11, -18, -26, -23, 10, -14, -26, -18, 21, 7, -7, -1, 10, 11, -2, -4, 9, -4, -27, -13, -2, -11, -27, -10, 15, -6, -6, -18, 0, -13, -16, -11, 6, -6, -9, -20, -5, -7, -18, -8, 3, 0, 5, 0, -6, -5, 0, -9, -5, 9, 8, -3, 0, -4, -8, -11, -10, -8, 8, 13, 9, 4, -3, 7, 16, -13, -19, -6, 3, -5, -4, -12, 5, 6, 3, 18, 1, 7, 5, 6, -2, 0, -1, 3, 0, -5, -1, -5, 5, 5, 3, 1, -5, 0, 0, -5, -3, -2, 5, -6, -2, -7, 5, -4, -4, 3, -5, 0, 24, 8, -5, -7, 4, -8, -28, -23, 0, -11, -25, -15, 22, 17, -4, -15, -11, -8, -5, 11, 12, -8, 6, -2, 0, 1, 23, -8, -1, -2, -8, -8, -2, 0, -1, -7, -4, -7, 5, 0, 2, -4, -5, 7, 3, -5, -4, -3, -10, 3, 4, 10, 11, 6, 8, -1, 1, 11, 13, 2, 2, 0, 5, 2, 3, 14, 20, 6, 17, -10, 9, -3, 13, 2, 21, -2, 6, 11, 21, 2, -23, -10, -6, -5, -11, 19, 20, -9, 0, 21, 33, -18, -11, -3, 7, -9, 4, 7, 10, 14, 7, 24, -1, 8, 1, 12, 9, 12, 0, 16, 6, 22, 3, 2, 3, 17, -9, 15, 8, 21, -10, 19, 5, 24, 2, 7, 20, 18, 0, 4, 2, -4, 3, -5, 4, 0, 5, -7, -3, -4, -6, -5, 0, 5,
    -- filter=0 channel=2
    12, 8, 1, -2, 6, 0, 5, -5, 9, 2, -1, 0, 4, 2, 1, 2, 4, 7, -1, -6, 2, -7, -5, 0, -6, 1, 1, -4, 1, 3, -5, 4, 3, -7, 3, -1, -6, 6, -5, 4, 6, 4, 0, 0, 2, 4, 4, -1, 9, -8, -1, 0, -9, -12, -9, -7, -4, -3, 0, -12, 3, -3, -7, -7, 11, 4, 3, 8, -3, 1, -3, 7, 9, 7, -1, -2, 0, 0, 0, 5, 9, -3, 9, 1, 3, -3, -7, 6, 7, -4, -4, 7, -2, -2, -7, -1, -2, -9, -4, -7, 6, 2, 4, 4, -2, 2, 7, -1, -3, 1, -6, 2, 3, -3, -9, 0, 4, 10, 2, -1, -3, -1, -8, 0, -1, 0, 2, 4, 7, 0, 3, 8, 0, 1, -2, 1, -1, -5, -4, -7, 1, 0, -2, 6, -5, -10, 0, 0, 6, 9, 0, -4, 6, 11, 7, 1, -4, 1, -9, 1, 18, 11, 10, 7, 7, -2, 7, 9, -1, -12, -11, -7, 10, 7, 4, 10, -6, -15, 0, -5, -5, 3, -3, 0, -7, -6, -9, 4, -7, -7, -3, 0, 3, 1, -5, -4, 2, -2, -2, 5, -1, -4, 0, 0, -2, 0, 2, 3, 6, 7, -6, -4, -4, 1, -7, -6, 4, 2, -5, -5, 4, -3, 0, 0, 6, 12, 12, 1, -1, 9, 5, -1, 0, 2, -5, 0, 11, 13, 4, 5, -1, 0, 2, 0, -4, -8, 2, 0, -5, 0, 7, -2, -9, -4, 8, -4, -6, 2, -6, 1, 7, 1, -6, 7, 5, -6, 5, -5, 3, -3, 2, -4, 7, 1, -4, -8, 2, 0, 6, -7, -4, 2, 3, 2, 2, -9, -10, 2, -11, -11, -6, -4, 3, -2, -5, -9, 2, 5, 5, 9, -6, 0, 5, -5, 10, -9, -15, -1, -4, -13, -6, -9, 3, -13, 4, -4, -2, -3, -8, 2, 9, 1, -2, -3, 6, 0, 6, -8, 6, -11, 4, 4, 0, 0, -8, -4, -7, 0, 0, -1, -4, -1, 0, -3, -3, 7, 4, 0, -4, -4, -4, -1, -8, -6, 2, -1, -5, 1, 0, -6, -3, -1, -4, 7, -11, 1, 5, -7, 0, 0, -8, -3, 1, 2, -1, 0, -7, 0, 5, -6, -4, -8, -8, 2, 5, 7, 4, 2, -4, 4, 5, 0, -5, -3, -3, 3, 0, -7, -5, -4, 4, -2, 3, -5, -5, -2, -1, -5, 0, -1, -4, -4, -6, 2, -2, -5, 1, 9, 2, 3, 6, 4, 6, 2, -2, 5, 8, 3, -5, -5, 5, 0, 7, 4, 10, 8, -1, 10, 11, -1, 2, 2, -3, 0, 6, 1, -3, -7, 0, -1, -6, 8, -7, 3, -3, 6, -3, -7, -4, 2, 3, 0, -5, 7, -3, -6, -8, -5, -2, 0, -6, -6, 0, -5, 3, 2, -4, -4, -7, -10, -3, -5, 1, -3, 0, 0, 5, -6, -3, 6, 2, 5, -4, 8, 3, -3, 6, -5, 5, 0, 3, 6, 1, 4, 0, 5, -4, 1, 4, 4, 2, -6, 17, 11, 6, 9, 4, -2, 5, 2, 0, 4, -3, -3, 18, 7, 5, 4, 5, -2, 8, -4, 11, 14, 1, 10, -1, -8, 3, -9, 6, 9, 3, 6, -1, -6, 3, 7, 2, -3, 2, 6, -7, 4, 5, 0, 0, 0, 3, 2, -2, 3, 7, 3, -7, -9, 7, 4, 3, -8, -2, -7, -1, -3, -6, -3, -6, 7, 2, -5, -5, -5, 5, -1, 2, 5, 7, 1, 7, -2, 5, -7, 0, -6, 6, 0, 4, 1, 0, 5, 1, 2, 3, 7, -8, 0, -5, -4, 4, 1, -7, -7, -7, 10, 0, -7, -6, 2, 4, -4, 5, -3, 6, -4, -3, -5, -7, -1, 3, 3, 12, -2, -1, 0, -2, -7, 4, 3, 8, -6, -7, 0, -4, 4, -3, 2, 9, 5, 5, -1, 1, -2, -12, 1, -9, 5, -3, 5, -1, 2, 2, 2, 8, 0, 7, 13, 5, 2, 3, -4, -9, 1, -10, -29, -15, 5, -14, -13, -7, 4, -11, -7, -5, 5, -15, -20, -15, 9, 26, 23, 19, 19, 17, 10, 9, 3, 15, -11, -10, 2, 16, 10, 9, 10, -5, -4, 0, -1, 5, -4, 5, 2, 5, -5, -4, 3, 7, 0, 5, -3, 3, -2, -6, -7, -4, 11, 15, 4, -2, 9, -1, -5, -4, -8, 1, 8, 11, 10, 6, -1, -4, -5, -6, 4, -2, 7, 0, 1, 2, -2, -2, -5, 1, -7, -1, -12, 0, -3, -5, 2, -9, -8, -8, 0, -7, -13, -11, -7, 5, 10, 18, 9, 10, 7, 7, -4, -2, -1, 0, 0, 15, 11, 13, -2, 12, 13, 1, -2, 3, 8, 1, -4, 2, -5, -2, 5, 1, 8, 1, 4, -2, -3, -5, -8, -8, 1, 7, 2, -3, 10, 21, 10, 2, 1, -5, -8, -3, 5, -8, -1, 3, 2, 2, -4, -1, 12, 7, 2, 2, -2, -3, -1, 12, 7, 3, -5, 4, 4, 6, 2, -2, 2, -9, 3, 8, 5, 0, 2, -3, -2, 5, 4, -2, 5, 4, -1, 0, 5, 3, -2, -7, 4, 3, -4, -2, 1, -4, -6, -1, 0, -3, 3, 4, 4, 5, -7, 0, 6, -2, -4, 9, 13, 11, 13, 7, -1, 14, -2, -5, 0, -1, 5, 9, 7, -3, 4, -10, -4, 0, -6, -3, 14, 8, 8, -9, -4, -4, -8, 6, -3, 3, -2, -1, -2, -5, -5, 3, 3, -4, 1, 6, -2, -4, 0, 4, -1, 5, -3, -3, -7, -2, -3, -8, 2, -6, 7, -4, -2, -3, 3, -1, -12, 0, 3, -10, -14, -10, 0, 5, -9, -4, -3, 2, -6, -2, 0, -5, -11, -2, 9, 0, -6, -7, 3, -8, -6, -2, 1, -2, -2, -7, 1, -3, 4, 2, 6, 3, -3, -3, -7, 0, -10, -3, 0, 0, -10, 5, -8, -6, -13, -15, 2, -9, -7, -9, -9, -5, -2, 5, -2, -3, 0, -7, -3, -9, -15, -2, -5, 4, -4, 0, -3, 4, 1, 7, 6, -7, 6, -4, 4, 6, 0, 2, -5,
    -- filter=0 channel=3
    -2, 7, 4, -9, 2, 4, 4, 7, 0, 2, -10, 3, -4, 5, -5, 0, -7, 2, -6, 0, -3, 3, -7, -5, 0, 3, 4, 7, 4, 7, -2, -6, -1, -3, -4, -5, -3, 5, 4, 0, 4, -6, -7, 5, 7, 6, 9, 4, 8, -25, 1, 5, 4, 4, 0, 12, 0, 12, -12, 5, -5, -14, -5, -3, 0, -2, 1, -5, 0, 0, 1, 8, 3, -10, -6, 9, 2, -2, -12, 0, 0, -2, 2, -11, 7, 3, 0, -2, -1, 0, -4, 4, 3, 0, 0, 0, 6, 17, 18, 12, -12, -6, 15, 30, -7, 3, 17, 24, 3, 9, 8, 9, 5, 7, 4, 10, 13, 8, 2, 4, 7, 1, 6, 3, -4, 0, -2, -14, 9, 5, 6, -7, 8, 3, 0, 5, -1, 0, 4, 4, 8, 6, 2, 6, 4, -8, 0, -1, 13, 31, 32, 21, 26, 21, 19, 19, 13, 4, 7, 4, 0, -23, -17, -29, -1, 14, 15, 12, 0, 3, 19, 8, 4, -11, -24, -26, 6, 15, -5, 9, 6, -12, -1, 0, 10, -1, 0, 6, -1, 4, 3, -9, 0, 1, 8, 0, -4, 7, 6, 8, -2, 0, -2, 9, -5, -4, 2, -4, 7, -5, -5, 1, -4, -4, 7, 0, -3, 6, 0, 0, 7, -2, 2, 0, -1, 2, 0, -10, 14, 17, 15, 11, -20, 7, 15, 10, 14, 12, 12, 1, -4, 6, 5, 9, -18, -4, 1, 16, -9, -7, -7, 9, -8, 0, 0, 17, 0, 2, 0, -3, -4, 6, -3, 0, 1, -7, 5, 5, 6, 4, -7, -5, -6, -5, -8, -20, 10, 13, 7, 1, -14, 14, 14, 8, 12, 0, 10, 4, 11, 9, 10, 19, -29, -6, 7, 20, -10, -9, 3, 17, -3, 5, -11, 2, 0, -10, -14, -1, 4, -4, -7, 9, -27, 6, -2, 8, 10, -4, 1, 16, 13, -8, -11, -10, 14, 8, -6, 7, -1, 13, 11, 0, 8, 0, -7, 8, 8, -9, 8, 8, -18, 4, 4, 13, -3, -4, 3, 10, 3, -9, 0, 0, -3, -6, 4, 9, -21, -15, 6, 12, -29, -17, 10, 15, -12, -12, -13, 4, -6, -6, -8, -3, -3, -4, -9, 9, -7, -15, -6, 15, 7, -1, 5, 4, -3, 0, 4, 0, 0, -4, -6, -1, 4, 1, 9, 3, -1, 0, 11, 6, 7, -5, -4, 4, 4, -6, 0, 1, 10, 2, -3, -3, -5, 0, -5, -7, 1, 1, -6, -5, 2, 4, 6, 0, 2, 8, 12, -4, 5, -4, 8, -9, -2, -4, 0, -13, 17, 11, 0, 8, 6, 16, 6, 0, 8, 9, 4, 12, 7, 6, 12, 8, 10, 5, 0, 3, 12, 2, 0, -1, -4, -5, 5, 3, 0, -18, -5, -1, -5, -2, -3, 4, -18, 9, -11, 9, 0, -14, -8, -6, 2, 2, 12, 6, -29, -5, 10, 23, -31, -28, 6, 28, -1, 2, 3, 5, -7, 5, 1, 5, 5, 7, 1, 0, -7, -7, -1, 7, 1, -1, -6, -3, -2, -16, -5, -2, 7, 11, 12, 14, 6, 14, 8, -5, 7, -16, -12, -9, 8, -5, -3, -10, 7, 10, 6, -5, -1, 16, 19, 20, 3, -3, -1, 0, 0, 4, 0, -7, -2, 2, -1, 6, 3, -7, 0, -2, -7, -2, 5, -3, 1, 0, -2, 0, 9, 11, -4, 13, 1, -1, -2, 2, -1, -8, -5, -4, -7, 0, -7, 6, -2, 4, 2, -7, 5, 1, -6, -1, 6, -6, -6, 0, -6, 7, 0, 3, -13, -11, -4, 9, -17, -14, -3, 0, 0, 5, 3, 1, -6, -1, -3, -3, 6, 0, 2, -6, 0, -5, -5, 8, 2, -4, 7, 3, 11, 11, 5, 10, 16, 10, 10, 8, -1, 22, 14, 28, -4, -1, -4, -4, -5, -8, -10, -5, -22, -20, 0, 12, -19, -23, 11, 28, -11, -6, 4, 0, 0, -6, 7, 8, -15, 17, 17, 9, 13, 18, 5, 7, 10, 3, -10, -14, -10, 2, 12, -27, 7, -23, -4, 25, 3, -23, -14, 26, -6, 22, 2, -20, -5, -5, -22, -35, 14, 8, 2, 8, -12, 0, 15, 6, -4, -10, -12, -14, 0, 4, -3, 5, 4, 1, 6, 0, -3, -6, 0, 0, -3, -2, 0, -4, 8, 7, 10, 19, 12, 6, 7, 26, -18, -8, 21, 29, -1, 6, -4, 9, 0, 2, -12, -4, 0, 0, 5, 11, -25, -12, 11, 7, -9, -3, -9, 2, 6, -13, -9, 9, -1, -9, -9, 6, -10, 7, 11, 15, 8, -9, -7, -1, 3, -14, -5, -16, 1, 1, 9, -1, 4, 9, 10, 2, -2, -4, -14, -21, 0, -12, -6, -8, 13, 12, 11, 0, 10, 8, 6, 1, 9, 3, 4, -1, 5, -4, -4, 12, -7, 7, 34, 32, 15, 21, 23, 15, 6, 6, 10, 8, -5, 9, 15, 3, -22, -8, -2, 0, 1, -4, -3, 18, 6, 4, -4, -10, 13, 0, 2, -10, 10, 16, 4, -4, -1, 6, 6, 15, 5, 0, 1, -2, -1, 6, 7, -3, 2, 3, 3, 2, -4, -7, -5, 2, 6, -7, 5, 2, 3, 4, -6, 1, 7, 6, -5, -5, -7, -2, 1, -3, -1, 2, -6, 5, 0, -3, 3, -5, 3, 13, 13, 6, 4, 6, 8, 2, 7, -6, 4, 3, 6, 20, 17, 12, 16, 9, 8, 11, -3, 6, 14, 21, 2, 0, -2, 1, -3, -2, 4, -7, -5, -3, 0, 0, -7, 4, 1, 0, -5, -3, 7, -1, 11, 9, 2, 9, -3, -5, 0, 12, -2, -11, 7, 17, -4, -8, -7, 9, -2, 8, 2, -11, 13, -13, -9, 14, -3, -18, -1, 7, 5, 1, 3, -8, -6, 5, 0, 4, -11, -8, 13, 12, -17, -22, 3, 25, -9, 6, -3, 7, 13, -16, 1, 1, 0, -6, -10, 10, -2, 2, -9, 7, 4, -21, -9, 10, -5, -9, -10, 1, -8, 1, -15, 0, 1, 0, -12, 8, -3, -17, -10, 0, -4, -1, 5, 6, -12, 7, 0, 2, 2, 1, -1, 3, 0, -2, 6, 4,
    -- filter=0 channel=4
    0, -11, 5, 11, -1, 3, -5, 5, -4, -1, -3, 2, -1, -9, -2, 1, 2, 1, -5, 2, 0, -3, 6, -6, 3, -1, 2, -6, -4, 1, 0, -2, -3, 4, -7, 1, 0, 2, -6, -3, 3, -2, 1, -1, -3, -4, -2, -4, -5, 14, 9, 3, -4, -6, -12, 12, -14, -15, 0, 32, 1, 13, 11, 14, -15, 2, 8, 7, -11, 1, -1, 7, -15, 7, 0, 5, -6, 9, -3, 7, -10, -1, -1, 0, 0, 4, 2, -5, 0, 0, 5, -6, 6, 0, -3, 5, 8, -7, 2, 2, -12, -22, -7, 0, -13, -23, -13, -4, -13, -5, -7, 3, -13, -16, -2, -3, -9, -4, 2, -3, 2, -2, 0, 7, -2, 7, -2, 4, -4, -2, 12, 12, -8, -12, 0, 11, 0, 6, -5, 5, -1, 3, -1, 12, -6, -3, -3, 0, -20, -14, -1, 0, -19, -6, -2, -7, -13, -13, -4, 2, -6, 8, 20, 26, -14, -3, 2, 36, -17, 7, -13, 30, -7, 22, 28, 29, 1, 0, 8, 9, -15, -3, 1, -7, -25, -14, 2, -9, -9, -14, 1, 6, 5, 5, 0, -3, 5, 6, 0, 0, 2, -1, -5, -7, 1, -10, -2, 6, 2, -6, -2, -7, 3, -3, 0, -1, 7, -5, 6, 5, -1, -6, 4, 7, -16, 0, 5, 8, -3, -1, -4, 1, 4, 3, -4, 2, -8, -6, 7, 13, -7, -2, 5, 4, 0, 0, -1, 0, 5, -7, -4, -2, -9, 0, 0, 0, -1, 7, -1, 0, -7, 0, 3, 1, -2, 6, 2, 7, 6, 4, -3, 2, -18, 7, 1, -3, -7, -8, -3, 15, -1, -12, 0, 8, -21, -2, 0, 5, -12, 0, 2, 0, -5, -20, -15, 0, -11, -21, -14, 1, -15, 1, -1, 2, -4, 20, 0, 4, -8, -5, 3, 0, -6, -8, 0, 10, -5, 19, 8, -5, 0, 10, -1, 13, -12, -5, 6, 11, -8, -10, -6, 30, -11, 13, 11, 18, -1, 8, -2, -7, -13, -8, -10, -1, -13, -7, -5, -15, -13, -1, 0, -9, -7, 11, 3, 0, -13, -18, -4, -10, -5, -15, -5, -13, 0, 12, -6, -10, -4, -4, 3, 0, 0, -2, 6, -16, -2, 0, -5, -5, 5, 0, 0, 9, -6, -12, 0, 3, -14, 1, 0, -4, 0, -4, 2, 8, -6, 0, -8, -5, 5, -6, -1, 6, 8, -4, -7, 1, -9, -7, 2, -4, 4, -7, -3, -8, -3, 0, -3, 8, 2, -6, -12, 5, -5, 2, 7, 2, 2, -3, 5, 4, -2, -2, 13, 12, 0, 0, -6, 13, -12, -3, -2, 7, -10, 1, 3, 5, 2, -3, 2, 7, 0, -7, -1, 11, -3, -3, 4, 7, 5, -2, 8, -2, -9, 8, 6, -7, -7, -2, -2, 2, -3, -14, 4, 17, -13, 5, 5, -10, -11, -2, -2, -9, -10, -16, -12, -9, -3, -17, -11, 3, -11, -5, 6, -4, -8, 7, -4, 1, 5, 1, 4, -1, -7, -4, 2, -2, 4, -7, 2, -1, -11, -2, 8, 26, 0, -2, -7, 22, -6, 0, -4, 25, -11, 4, 9, 31, -13, -18, 0, 10, -4, -3, 10, 6, 3, -1, -16, 6, -10, 4, 19, 10, 0, -3, 7, -5, -5, 7, -4, 2, -7, 1, 0, 4, -6, -4, 5, 5, -1, -4, 5, 17, -11, 2, -9, 11, -9, -5, 1, 14, -5, 3, 4, 8, 6, 0, 6, -4, 7, -3, 5, -1, 7, 0, -5, 0, -4, 0, 6, -6, 7, -4, -7, 5, 0, -1, 0, -7, 7, 3, -4, -8, 0, 0, -3, -5, -4, 2, 5, -1, -1, 0, -1, -2, -2, -2, 1, -6, 4, 0, -7, 6, -13, -5, -11, -11, -14, -7, 3, -5, -5, -21, -17, -4, -9, 0, 9, 3, -10, 4, 0, -6, -13, -10, 5, -13, -15, -17, 2, -12, -8, 7, 7, -7, -8, -5, 1, 4, -5, -5, -10, 8, -19, 0, 2, 11, -11, 11, 7, 9, -13, -21, 9, 5, -36, -29, -13, -6, -27, -31, -22, 1, -23, -28, -2, 2, -15, -1, 27, 24, -11, -3, 0, 26, -6, 12, -6, 30, -15, 0, 27, 37, 0, 4, -8, -6, -5, -5, -2, -3, -7, -6, 0, -6, -1, 2, 0, -2, -7, -12, -9, -3, 3, -15, -2, 6, -8, -13, -5, -2, -3, 4, 12, -5, 2, -3, 6, 5, -5, -4, -6, -4, 7, -7, -13, 0, 3, 12, 13, 9, 2, 11, 1, -5, -9, -2, 9, 0, -1, -13, 0, 16, -5, 10, 7, -10, 1, 12, 16, 18, 1, 1, -10, 19, -1, -1, -13, 27, -13, 15, 21, 32, -10, 3, 13, 16, 0, -14, -10, 17, 0, 2, 0, 16, 1, -7, 0, 10, -6, -1, 7, -4, -10, -17, -6, -10, -2, -21, -12, -1, -2, -6, -6, -13, -4, 2, 6, 4, -10, -4, 2, 6, 0, -14, 1, -12, -4, -7, -3, 2, -15, -5, -2, 3, -9, 0, 11, 6, -2, 3, -10, 6, -15, -2, 7, 18, -4, 5, -3, 8, -8, 2, 0, 7, -1, -5, 2, 1, 0, 6, 5, -4, 6, -7, 5, -1, 5, -5, 4, 0, 6, -1, 4, -7, -5, 0, 6, -4, -6, 2, 14, 32, -16, -6, -9, 38, -3, 7, -5, 23, -7, 7, 6, 20, -17, -23, -10, -16, -4, -15, 4, -1, -2, -29, -20, -7, -9, -4, 2, -3, 2, -1, 1, -3, -1, 3, 6, 0, -3, 0, 0, 0, 5, 7, -4, -6, 1, 0, 4, -3, 0, -9, -2, -3, -9, -11, 0, -10, -7, -1, 4, -5, -7, -8, 4, 5, -28, -7, -1, 3, -23, -10, -8, 10, 0, -17, 5, 4, 1, 2, 2, 1, 3, -15, -4, -3, -5, -13, -10, -8, -5, -6, 5, 0, 10, -3, -3, -2, -3, -3, -1, 11, -5, 1, 2, 9, -8, 6, -7, -7, -9, 10, 0, -6, -5, -2, 0, 8, -3, 1, -4, -3, 6, 20, 2, 2, 0, -1, 0, -5, -2, 0, 0, -7, 3, 4, -1, 6, 4, 1, 6, 2,
    -- filter=0 channel=5
    8, 13, 12, -6, -4, 0, -1, 6, 8, 5, -7, -4, 1, 4, -5, 2, -4, -6, -2, -4, -5, 2, 4, 4, 0, 0, -2, -6, -3, 7, 0, -7, 3, 4, -1, -8, 6, -6, 4, -9, 6, 1, 6, 0, 0, 7, -8, -5, -4, -4, -13, 3, 15, -6, -1, -10, 23, 0, 0, -9, 0, -3, 0, -26, -9, -12, -8, -7, 7, -2, 1, 18, 5, 5, 5, 13, -5, 7, 14, 12, 8, 2, 7, 0, 7, -1, 7, 2, 5, 7, 6, 0, 6, 0, -4, 4, -21, 2, 15, 13, 16, 10, 10, 11, 6, 27, 14, 15, -20, -14, -11, -6, 9, 2, -7, 6, 13, 11, 0, 9, 15, -4, -3, 3, -4, -9, 2, 1, 4, 2, -6, -13, 14, 5, -11, 2, 17, 0, -5, -1, 12, 2, -4, 3, 3, 11, 11, 6, 19, 7, 5, 12, 14, 15, 5, 19, 0, 0, 0, 6, 2, -13, -14, -5, 27, -18, 0, 16, 25, -11, 9, 22, 9, -14, 9, 4, -15, -3, -17, -6, 5, 22, -30, -1, 1, 13, -22, 6, -7, -6, -19, -12, 1, 2, 6, 6, 2, 0, -6, 0, 0, 8, 0, -5, 0, 1, 0, 2, -1, -2, 1, -2, -7, 0, -6, -4, -5, -5, -5, 0, 6, 6, 3, -7, -27, -11, -22, -18, -5, 19, 23, 33, 22, 11, 17, 25, 13, 10, 26, 14, -15, -9, 0, 2, -2, 4, 5, 16, 9, 2, 10, 16, -12, -5, 1, 1, -8, -1, 2, -2, -5, 4, -2, -3, 0, -7, 1, 4, 4, 4, 1, 6, -9, -22, -24, -14, 9, 1, 8, 19, 20, 4, 10, 20, 17, 18, 27, 16, -26, -19, -10, -2, 23, 7, 13, 23, 10, 13, 9, 33, -28, -14, -5, -7, -26, -12, -27, -23, 27, 0, 12, -5, 39, -1, 12, -6, 17, -2, 13, -3, -9, 4, -17, -13, 7, 7, 5, -3, 23, 0, -4, -8, 1, -10, -3, 3, -7, -8, -16, 0, 35, -2, 4, 11, 14, 1, 15, 2, -26, -5, -5, -5, -21, -12, -2, 2, 24, 1, 6, 5, 29, -3, 22, 4, -31, -20, 0, -1, -7, -17, -12, -16, 13, -14, -7, -7, 4, -7, -3, -8, 0, -4, -12, -13, 6, 8, -3, -3, 11, 1, 9, -4, -2, 0, -4, 2, 10, 0, 3, 7, 6, 0, -3, 0, 8, 7, 3, 0, 2, -6, -1, 11, -2, 4, 9, -8, 5, -5, 10, 10, 12, 6, 0, 6, -5, 10, -2, 9, -3, -7, 2, -12, 9, 0, -14, -12, 7, 12, 0, -1, 15, 3, 3, 0, 14, 2, 0, 12, 7, 0, 7, 0, 1, -6, -8, 1, -3, -8, -4, -12, -3, 0, -6, -5, -17, -6, -10, -4, 18, -4, 12, -6, 22, 0, 5, -6, -5, -14, 8, -14, -15, -12, 2, 9, 15, 0, 19, 27, 20, 8, 19, 25, -16, -2, 9, 0, 0, 1, -9, 4, 3, -4, 7, 0, -4, -4, 0, -7, 4, 4, -2, -1, 14, -2, -4, -8, 15, 5, 1, -1, 5, 4, 6, -1, 2, -8, -12, -5, -3, 0, -2, -17, 10, 14, 3, 4, 18, 4, -12, -2, -4, -6, 1, -5, 6, -7, 4, -7, 1, -7, 3, -7, 5, -3, -5, -5, 1, -8, 4, 0, -5, -5, -5, -12, 13, 0, -8, -3, 10, -11, 1, -8, 8, -7, -2, -2, -7, 6, -7, 0, 4, -7, 1, 2, 7, -7, 6, -3, 0, 3, 2, -7, -7, 0, -3, -1, -11, -6, -4, 9, -3, 0, -3, 12, 1, -1, -3, -1, -8, 0, -7, -4, -3, 3, 3, 6, 3, 2, -8, -6, 1, 3, 8, 11, 0, 3, 5, -4, 8, 22, 15, 7, 22, 13, 16, 19, 4, -11, -4, -6, -27, -32, -15, -13, 16, -2, 9, 9, 25, -8, 12, 11, -21, -2, 2, 2, 4, 0, 12, 6, 24, 10, 11, 9, 2, 7, 17, 6, -22, -10, -7, -19, -16, -18, -20, -27, 15, 0, -28, 3, 0, 2, -33, 3, -18, -22, -14, -9, -24, -17, -10, -4, 11, 13, 8, 33, 20, 6, 4, 22, -7, 1, 11, 18, 9, -1, 0, 4, 4, -5, 0, -5, 10, -9, 7, -1, 7, 0, 6, 3, -20, -9, -11, -10, 4, 17, 11, 28, 17, 15, 15, 22, -15, -6, 5, 0, -27, -13, -13, -12, 0, 12, 14, 24, 13, 12, 16, 33, -2, -1, 10, 10, -25, -7, -9, -14, 11, 10, 10, 6, 40, -5, 18, 1, -3, -11, 0, -16, 0, -4, -11, -11, 15, -5, -5, 4, 15, -5, -6, 4, 5, -4, -4, -2, 7, 4, -1, -6, 2, -5, 8, -6, 6, 7, 3, -7, 14, 6, 11, 4, -8, 4, 0, 4, 19, 16, 17, 15, 11, 19, 25, 13, -7, -8, 1, -1, -5, -7, 6, 1, 0, 9, 8, 20, 6, 19, 15, 25, -27, -8, -14, -10, -3, 3, -7, -11, 11, 3, 3, 9, 14, 2, 0, 0, -4, -3, -6, -13, 9, 5, 2, -6, 7, 2, -5, 2, 4, 5, 5, -6, -6, 3, 0, -2, 2, -3, 6, -3, -4, -1, 0, 0, -5, 0, 4, 3, -7, -5, 0, -1, 1, 0, -11, -8, 18, 4, 5, 0, 15, -3, 5, 4, 3, -3, 8, 0, -5, -10, -13, -11, -6, 7, 11, 12, 6, 15, -3, 13, -27, 0, -5, 2, 0, 4, 6, 1, -7, -5, 3, 6, -1, 3, 1, -5, -5, 0, -5, -2, 1, -3, -12, -14, 13, 0, -6, -3, 22, 2, 1, 6, 0, -3, -9, -9, -3, -12, -17, -15, 8, 14, -13, 2, 4, 9, -22, 16, -4, -5, -1, -4, -16, -12, -10, 5, 9, -6, 6, 10, 15, 9, 16, 13, -11, -6, 1, 0, 0, -4, -14, -6, 25, -5, -18, -5, 25, -2, -7, -11, 12, -5, -11, -8, 11, -5, -17, -14, 16, 2, -20, -10, 19, -6, -13, -9, -6, -4, -18, -11, -2, 2, 3, 7, 5, 1, 6, 1, -4, 7, 2, 5, 0, 1, -2, 2,
    -- filter=0 channel=6
    -6, -4, -6, -10, 0, -3, 4, -6, 4, -5, 16, -3, -5, 0, 3, 1, 4, -1, 0, 4, 7, -6, 3, 1, 1, 7, 4, -7, -6, 0, 6, 4, 0, -4, 2, -3, 0, 1, -5, 11, 5, 2, -8, 2, -6, -6, -2, 0, 0, 2, 3, -10, 10, 37, 16, 9, 0, 25, -15, 11, 3, 0, -6, 9, -2, 4, -8, -9, -8, 3, 10, -17, 6, 10, -6, -16, 6, -7, -3, 0, -1, -7, -2, -3, -4, -1, 0, 0, 7, 0, -6, -3, -6, 0, 0, -1, -2, -9, -9, 0, -18, -19, -19, -12, -6, -2, -4, -3, -7, 8, 14, 5, -2, 12, -3, 0, -9, -8, 1, 0, -7, 0, 4, 5, 0, -7, 5, 6, 9, 1, -11, 0, 9, 2, 15, 8, -3, 9, 30, 7, -8, -5, 10, 7, 0, 8, 0, 0, -18, -3, 1, 5, -18, -15, 1, 1, -8, 23, 8, 1, -2, -21, -29, -15, 12, 48, 9, -19, 16, 56, 21, -16, 4, -6, -24, 8, 0, 0, 2, 9, 3, 3, 7, 4, 20, 9, -12, 3, 3, 2, -19, 13, -1, 1, -6, 3, 0, 7, 4, -5, -4, 1, -1, 4, -5, -6, -2, -1, -8, 0, 6, 0, 4, -7, -4, 4, 4, -6, 2, -1, 0, 2, 0, -5, 11, 3, 1, 4, -5, -7, -11, -15, -14, 11, 3, -25, 2, -5, -12, 0, -5, -8, -3, 5, -8, -13, -6, -8, -10, -14, -8, 0, -11, -9, 1, 2, -3, -4, 0, 0, 3, 0, 2, -3, 2, -4, -1, 4, -2, -2, -3, -6, 6, -6, 0, 2, 1, -6, -9, -6, -5, 6, -5, -16, 7, -6, 0, 0, 0, 14, -7, 0, -10, -17, -13, 0, -8, -19, -23, -1, 5, 11, -5, 11, 10, -16, 1, 11, -7, 0, -19, 17, -11, 16, -35, -1, 0, -4, 1, 8, 16, 3, -3, 6, 14, 19, 9, 6, 18, 31, 3, 0, 9, 0, 0, 0, -8, 6, 4, 11, -12, -21, -19, 5, -11, -15, -26, -5, 4, -2, -12, 15, 11, -9, -16, 4, -6, -31, -15, -6, -11, -25, -25, 0, -2, -3, 2, 14, -1, 1, -8, 7, -3, -9, -7, 10, -5, -15, 0, 5, -9, 12, 3, 1, 7, 0, -5, 0, -10, -21, 1, 8, 0, 8, 3, 2, 3, -6, 0, 2, 6, -11, 0, 2, -11, -4, 5, 0, -6, -4, 0, -7, -1, 1, 0, 2, 3, -2, -1, 1, -8, 5, 11, 1, -8, -8, -2, 4, -5, 0, 0, -2, 3, 0, -1, 0, 8, 17, 4, -2, 5, 18, 21, 3, 1, -1, -1, 5, 0, 8, 3, -5, 6, 10, 10, -4, 13, -1, 10, 15, 3, -14, 9, 4, -7, -21, 0, -3, -1, 6, -22, 1, 1, 21, -18, -8, 3, -10, -2, 14, -6, 1, 0, 16, -4, -12, -22, -11, -7, -9, -19, -10, -6, -7, -7, 21, -2, -6, 3, 5, 5, 4, -4, 6, -5, 0, 4, 3, -3, 6, 0, 0, 8, -1, -5, -13, 13, 35, 24, -3, 16, 33, 27, 6, 2, -12, -6, 1, 10, -5, -1, -5, 3, -4, -16, 6, -3, 14, 19, -4, 3, -4, -6, 0, -2, 4, 1, 3, 0, 6, 0, -1, -2, -2, 2, 0, 5, 3, -6, 4, 6, 2, 8, -4, -4, 21, 6, 0, 4, 21, 3, 12, 4, -7, 9, 4, -7, 4, -7, 3, 1, 1, -2, 0, 7, -2, -7, -3, 0, -1, -7, -4, -14, -7, -9, -5, -11, -10, 3, -1, -1, 1, -1, -1, -4, 0, -4, 8, 0, -2, -3, 9, 6, -4, -2, 5, 4, 6, 3, 4, -4, -6, -7, -2, 1, 17, 16, 19, -9, -21, -6, -8, -10, -15, 9, -7, 3, 1, 5, 11, 7, -13, -3, 16, -11, -28, -24, 6, -8, -19, -23, -9, -5, 12, -3, 1, 0, -5, 2, -1, -12, 10, 3, -6, -1, 6, -1, -9, 0, 9, 14, 9, -20, 6, -30, 30, 39, 15, -24, 5, 29, 8, -4, -3, -20, -3, -22, 12, 15, -18, -23, 0, 4, 21, 22, -12, 0, 45, 26, -21, 2, -11, -28, -17, 5, 8, 0, 2, -6, 0, -2, 2, -1, 4, -3, 6, -6, -6, 7, 0, -2, 12, 11, 15, -11, -16, -17, -7, -16, -23, -19, -15, 8, 11, 2, 7, 3, 6, 4, 11, -9, -1, -7, -7, -2, 3, -8, -20, -5, -17, -18, 0, 0, 1, 8, 14, -13, 2, -7, 17, 0, 5, -23, -8, -1, 1, -3, 16, -2, -7, -16, -4, 6, 31, 22, -7, 12, 40, 22, -6, 2, -18, -13, 7, 3, 2, -3, -6, 10, 29, 0, -4, 0, 18, 12, 4, 2, 1, -5, 2, 5, 0, 5, 2, -7, -22, -8, -10, -11, -8, -6, 7, -2, 12, 24, 17, -13, -10, -20, -9, -4, -16, -10, -4, -7, 0, -15, 1, 14, 16, 16, 10, 3, 0, -10, 14, -11, 2, -8, 4, 2, 21, 24, 2, 10, 4, -12, 9, 0, -4, 2, 0, -7, -3, -4, -6, -7, 5, -1, 3, 4, -3, -7, -1, -3, -4, 0, -1, 2, 6, 2, 0, -3, 2, 0, 5, 1, 5, -3, 7, 3, -5, -22, 2, -1, 41, 5, 1, 13, 40, 31, 11, -1, -11, -9, 5, 8, 25, 14, 11, -13, -14, -25, 2, -14, -19, -1, -5, -1, 2, -4, 4, 0, 7, -5, 7, 4, 3, -2, 0, 0, -7, -1, 7, -3, 0, 0, 2, 7, 11, -2, 14, -10, -17, -8, 13, -8, 0, -3, 0, -1, 20, 2, 11, -7, 12, -15, 20, 19, 6, -12, -7, 9, -5, 7, -1, -11, -4, -9, 7, -5, -6, 3, 3, -6, -16, -3, 0, -4, -12, -16, -9, -8, -1, 6, 10, 5, 8, -4, 5, -7, 8, -12, 8, -4, 2, -2, 18, -3, 0, 10, 13, 7, -10, -2, -3, 5, -3, -23, 0, 9, 4, -14, 10, -4, -8, 8, 6, -4, -5, -5, 6, -3, 4, -6, -4, -4, -1, 8, -4, 0, 2, -3, 6,
    -- filter=0 channel=7
    -11, -5, 7, 2, -10, -2, 2, 4, -1, 4, -10, 4, -5, -2, -2, 5, 4, -5, 0, 4, -7, 3, 2, 2, -6, 2, 1, 6, -7, 4, 7, 6, 2, 1, 4, -2, -5, -8, -1, -10, -5, 5, -2, 4, -7, 3, 4, 0, -14, 20, -4, -3, -9, 9, 7, -14, 5, 3, 16, -19, -5, 24, 4, -9, 0, -6, -2, 14, 0, -9, 4, 2, -14, -5, 11, 11, -4, 14, 11, 6, 0, 2, 6, 10, -5, 4, 0, 6, 1, 5, -5, 5, 1, 5, 2, 6, -10, -1, 5, -15, 5, 3, -9, -14, -7, 6, -1, -25, 10, 1, -2, -11, 6, 6, 5, -9, 0, 10, 3, -11, 5, 10, -3, -2, -5, 13, 9, 0, 0, -1, 9, 12, -9, -15, -5, 3, -6, -18, -9, 4, -4, 5, -6, 3, 1, 4, -2, -7, 25, 16, -2, -14, 18, 21, -6, -19, 4, 22, -7, -11, -14, 13, 13, 26, -31, -38, 1, 29, -16, -43, 0, 29, -20, 3, 27, 30, -11, 8, -9, -12, 1, 22, -17, -11, 5, 24, -1, -19, 9, 6, -7, -6, -7, -7, -5, 2, 7, -2, 4, 0, -2, -3, -4, -3, -8, 3, -2, 2, 3, 1, 0, 2, 1, 4, 4, 2, -2, -1, -4, 1, -7, -2, 6, -6, -12, 16, 22, 2, -11, 8, 20, 23, 0, -10, 8, 12, -12, 7, 23, 5, -2, -15, -12, -13, 5, 0, -14, -6, 0, -9, -9, 0, -1, -15, -2, -3, 7, -4, -1, 3, 6, -6, -2, 4, 3, 7, 1, 0, -1, -2, -1, 5, 8, 12, 3, 0, 7, 15, 12, -8, 11, -8, 19, 2, -11, 16, 13, -5, -14, 0, -3, -20, -6, 29, -3, -16, -15, 15, -2, -26, -1, -6, -12, -23, -11, 18, -14, -20, 5, 36, 12, -30, 6, 0, 25, -36, 2, 22, -5, -20, 0, 13, 4, -7, 8, -10, 4, -8, 0, -12, 1, -4, -4, 4, 6, 11, -1, 8, -10, -19, 4, 15, 9, -9, 1, 24, -3, -20, -3, 5, -2, -14, -10, 5, -6, -12, 9, 15, -9, -18, 0, 20, -4, -17, 0, -1, -16, -20, 3, -3, -18, -10, -2, 11, -9, -11, 7, 12, -17, -22, 10, -1, -10, -5, -5, 5, -1, 0, -3, 0, -13, 0, 4, -8, -9, 1, 3, 5, 1, -7, -11, 7, 5, -3, -1, -2, 6, 5, 4, 3, 4, -4, -5, 1, 9, -4, -6, 11, 9, 5, -7, -4, 4, 8, -9, -1, -3, 1, 7, 8, 0, 9, -8, 15, 11, 2, -7, -12, 12, 2, -5, -14, 1, 5, -12, 6, 5, 5, -12, 0, 0, -7, -9, -5, 6, 3, 0, 3, 5, -9, -4, 3, -10, 2, 1, 20, -2, -2, 7, 13, 6, -16, 0, 9, 10, -11, 2, 14, 0, -18, -12, -17, -2, -19, -10, 4, -4, -8, 5, 6, -4, -14, 6, -18, 2, -14, -4, -4, -4, -3, -4, 0, 7, -6, 0, 1, 0, -2, 7, -6, 1, -6, -14, 6, 6, 12, -10, -29, 8, 11, 2, -17, 9, 8, -4, 17, 3, 22, 1, 11, 6, 2, -2, 7, 1, -6, -14, -7, -4, 7, -11, 6, 3, 8, -5, 2, 5, -6, 3, 3, -6, 4, 5, 3, -7, 3, -5, 0, -6, 7, 10, 7, -7, 0, 8, -14, 6, -9, -1, -8, 0, -1, 0, 3, 0, 3, -3, 1, 1, 1, 0, 0, -5, 0, 0, -3, 0, -4, 5, -5, 4, -5, 2, -11, -1, -4, 0, -14, -2, 4, -7, -8, -13, 0, -4, -9, 1, 0, 5, 6, -4, -4, 12, 0, 10, -12, 15, 6, 6, -7, 11, 7, -1, -3, 3, 9, 0, -15, 18, 9, 6, -1, 12, 17, -1, -4, -1, 8, 2, -6, -5, -5, 0, -19, -1, 8, -4, -9, 7, 16, -15, -15, 2, -7, -8, -14, 0, 9, 9, -8, 7, 1, 0, 2, 6, 6, 2, 8, 6, 6, 9, 7, 27, 5, -24, -23, 13, 49, -4, -33, 22, 51, -14, -47, 28, 9, -24, -11, -24, 19, 19, 35, -43, -17, 13, 39, -18, -36, -6, 26, -23, 0, 19, 32, 10, 8, 3, 2, 7, 1, 8, -7, 10, 10, 1, -8, 3, 8, 0, -9, 0, -10, -1, -14, 2, 2, 12, -12, 8, 19, -6, -7, -18, 1, -6, -4, -4, -4, 14, 3, -3, -6, 20, 0, 6, 4, 0, -5, -11, 0, 14, 11, 3, 22, -16, -27, 10, 29, 15, -20, 7, -1, 17, -13, 3, 29, -6, -13, -3, 3, 2, 15, -8, -19, 4, 17, -12, -35, 8, 11, 0, 5, 17, 16, -2, 3, 17, 11, 0, -8, 15, 7, 0, -16, 0, 6, -2, 3, 0, 4, -13, 7, -2, -1, -4, 13, 9, -12, 16, 9, 14, -19, 10, 8, 2, -14, 4, 12, 13, 6, 2, 3, -1, -9, -8, 6, 14, -7, -6, -11, -9, -11, -1, 18, 14, -9, -1, 3, 11, -6, -5, -11, 10, -3, 0, 18, -2, -3, 6, -1, 4, 3, 0, -5, 7, -7, -3, 7, 5, 5, 6, -3, 4, 5, 6, 2, -5, -2, -3, 2, 3, -5, 2, -1, 4, 7, 5, 6, -1, 0, 4, 7, 16, 15, -6, -31, 12, 13, -3, -16, 5, 9, 0, -8, -4, 16, 17, 9, -7, -11, 14, 17, 7, -13, 16, 37, -8, -20, -9, 5, 2, -22, -4, 4, 2, 0, -1, -1, 4, 3, -6, -3, -4, 5, 4, 0, 5, 6, 1, 8, -7, -2, 9, 10, -1, -11, 5, 12, -13, -12, 3, 0, -5, -14, 22, 7, 1, -13, 10, 22, 7, -16, 11, 33, -1, -19, 11, 9, -4, 4, 3, -11, -12, -13, 1, -2, -1, -13, 3, 3, -9, -14, 0, -7, -7, -8, 5, 13, -2, -4, 8, 15, 9, -17, 9, 5, 8, -28, 8, 20, -18, -12, 27, 24, -4, -5, 30, 13, 11, -15, 25, 25, 1, -25, 7, 13, -11, -14, -9, 6, 0, -7, 2, -2, 4, 0, -7, -6, 4, 0, 5, 0, 6, 1,
    -- filter=0 channel=8
    3, -4, -2, -6, 2, 0, 7, -3, 0, 0, -2, 1, 5, 0, 2, -2, 5, 7, 4, 4, 0, 0, 6, -6, -1, -7, 2, 0, 2, -7, 5, 7, 7, 8, 5, -5, -3, -1, 7, 7, -1, 0, 9, 10, 3, 2, -2, 6, 1, 24, 15, -30, -7, 15, 15, -16, -5, 5, -4, -22, 5, 16, -2, -36, 0, 15, 5, -2, -2, 5, -3, -13, -13, 14, 6, -17, -9, -12, 0, -27, 2, 0, 4, 0, -3, 7, -5, -5, -3, -7, -2, -3, -4, 0, -6, 0, 20, 9, 1, 30, -3, -13, -15, 20, -17, -37, -17, 20, 6, -3, -8, 19, -6, -12, -2, 4, -20, -7, 0, 0, -10, -8, 2, 0, 1, 0, -4, -2, -5, -9, -7, -20, -3, -2, 5, -3, -13, -2, 12, -14, -7, -13, 4, -21, 0, 13, 0, -2, -29, -21, 1, -5, -26, -36, -12, 17, -10, -19, 16, 18, 2, -3, -17, -48, 0, 41, 9, -25, -2, 46, 24, -33, 0, 3, -2, -59, 20, 0, 0, 1, -12, -10, 19, 9, -18, -11, 2, 12, 17, 5, 2, 5, -1, 4, -5, -3, -3, -4, 0, 5, -2, 2, -2, 0, -8, -11, -9, 2, -5, 3, -7, -3, -6, 7, -3, -2, -4, 4, -6, -7, -5, 3, 1, 4, 11, -11, 0, -6, -12, -12, -6, 0, 11, 8, -6, -7, -9, -4, 4, -15, 12, 22, 26, 26, 0, 0, -13, 4, 2, -3, -15, 16, 5, 4, 0, 20, 8, 1, 0, -5, -9, -4, -1, -8, 0, -4, -1, 2, 2, -6, -6, -3, 2, -10, 0, -20, -18, -4, -2, -14, 0, 3, -7, -25, -15, -3, 8, -17, 20, 0, 8, 21, -6, 8, -17, -2, -9, -16, -16, 19, 21, 3, 7, 7, 20, 14, 11, -11, -9, 6, 2, -22, -4, 10, 0, -33, 0, 7, 25, -30, -7, 6, 2, -32, -10, 4, 2, -15, -13, 15, 1, -17, -1, 0, 2, -35, 3, 9, 12, 0, 8, 4, -10, -5, 0, 0, 3, -17, 18, 0, -2, -5, 32, 10, 8, 20, -2, 4, -29, -5, 0, 2, -23, -3, 24, 22, 7, 0, 19, 0, 0, 8, -2, -15, 1, 5, 0, -2, 2, 0, 9, -3, 12, -2, 1, -4, 9, 3, 3, 0, 3, 7, 0, -4, 0, -5, -7, 1, -4, -2, -1, 2, -7, -13, -9, 1, -1, 4, -1, 2, -10, 0, -3, -7, 1, 7, -2, 0, 4, -12, 0, -12, -1, 3, -9, -9, -5, 3, 1, -9, 5, -2, 0, -6, 3, -17, -17, -6, 6, -1, -12, -8, 0, -13, -9, -17, -7, -22, -7, 4, -7, -5, -9, 6, 0, 3, -14, 0, 5, -2, -10, -1, -8, -13, 4, 7, 6, -18, -3, 8, -4, -28, 8, 2, 4, -20, 3, 6, 8, -21, 23, 22, 16, 19, -2, 7, -31, 0, 0, 4, -20, -3, 31, 23, -11, 0, -3, -2, -5, -5, 1, -5, 5, 5, -1, 7, 4, 7, 6, -1, -5, -4, -10, 3, 0, -37, -23, -2, 16, -13, -23, 0, 6, -23, -17, -1, -1, -51, -13, -10, -2, -7, -19, -13, -4, -6, -7, -4, -6, 3, 3, -3, 1, -19, -2, 0, -1, -7, 0, 4, -6, -7, -6, -7, 2, -2, 5, -7, -7, 1, -11, 0, 0, -29, -13, 0, 15, -11, -12, 8, 7, -22, -16, 4, -1, -21, 0, -2, 7, -5, 5, 3, -6, 0, -7, 6, -2, -2, 0, -7, 7, -4, 12, 11, -3, 18, 4, -10, -9, 4, -1, -3, -11, 8, 18, 19, -5, 9, 3, -1, 8, -6, -11, 0, 2, 1, -13, -5, 6, 4, -4, 0, -2, -3, -5, -18, 0, 18, -17, -28, -19, -11, -16, -18, -1, 0, 8, -1, -6, -2, 26, 17, -17, 11, 10, -6, -31, 1, 0, 7, -18, 0, 24, 22, 10, 17, -1, 5, -6, -20, -5, 8, -7, -10, -13, -11, -2, -6, -1, 4, 11, -6, 35, 36, 23, 16, -31, -2, 25, 16, -18, -17, 26, 15, 23, 23, 21, -2, 0, -14, -7, -49, 0, 7, 21, -20, 8, 13, 27, -13, 1, -5, -4, -39, -5, -7, 3, -1, 2, -4, 3, 0, -11, 0, -6, -8, -6, -1, 0, 0, 5, 1, 3, 14, -14, -21, -26, -4, -3, -3, -5, 2, 20, 4, 7, 22, 13, 12, 3, -14, -2, -1, 4, -18, 11, 18, 0, -26, 1, 4, 2, -22, 11, -1, 14, -4, -15, 0, -16, -6, 1, 7, -2, -18, -2, 5, 4, -23, -9, -3, -3, -39, -13, 10, 17, -11, -15, 19, 12, -18, -8, 1, -3, -43, -10, -10, -12, -11, -7, -15, -2, 1, -16, 2, -4, -4, -14, -5, 0, -16, 15, 7, 8, 16, -4, -14, -16, 10, -27, -35, -30, -4, 3, -17, -3, 17, 14, 12, -3, -5, -1, 0, -10, -12, -7, -13, 1, 3, 13, 3, 20, 11, 4, -10, -4, -28, -3, -4, 3, -19, -6, -1, 4, -12, 9, 3, 10, -39, -2, 3, 6, 6, -4, 5, 5, -5, -5, 0, -8, 2, 2, 1, 4, 1, 3, 5, -7, -7, 5, 3, 0, 3, -2, 0, 4, -3, -2, 0, 1, -5, -11, -8, 2, -32, -16, -1, 19, -10, -17, -2, 20, -13, -19, -8, -7, -33, -7, -6, 28, 31, -32, -33, -27, 0, -15, -21, -4, -10, 12, 8, 6, 8, 0, 0, 3, -4, 3, 3, -2, -2, -3, -3, -3, -1, -2, 0, 1, 5, 0, -6, 10, 0, -11, -5, -13, -2, -9, -3, 2, -4, 0, -2, 11, 10, 17, 15, 16, 0, -14, 0, 7, -2, -7, -3, 14, -7, 19, 12, 17, -9, 15, 21, 16, 12, -4, 1, -13, 0, 3, 7, -16, -10, 6, 3, 4, 13, -2, 14, 12, -6, -20, -6, 8, 4, -8, -3, 4, 1, -5, 0, 14, -13, -7, 6, 14, -22, -12, -17, 16, -9, -22, -5, 23, -20, 0, 2, 2, -24, 10, -3, 2, 5, 6, -7, -4, 7, 3, 0, 0, -2, 5, -6, -1, 8,
    -- filter=0 channel=9
    0, -5, 4, 0, -5, 10, 1, -8, -4, 2, 10, -10, -4, 0, 7, -4, 5, 3, -3, 3, 3, -5, 2, 2, 0, 2, -4, 0, 5, -5, 5, 0, -7, 4, 8, 6, 5, 0, 5, 9, 0, 4, 0, 4, 3, 3, -4, -2, -6, -9, 21, 28, 0, -5, -13, 17, 3, -7, -9, 14, -20, -5, 15, 30, -3, 7, -7, -6, 10, 1, -12, -6, 8, -5, -6, 0, 9, 7, -7, -8, -6, 0, 0, 6, 3, 1, -6, 2, -2, -4, 5, 7, 2, 0, 7, -5, 25, 17, -13, -36, 18, 7, 20, -1, 33, 3, 1, -12, 19, -11, -27, -24, 2, 9, 8, 11, 8, -3, -1, 8, 6, 5, -8, 5, -4, -2, -5, -4, -6, -1, -10, 2, 6, 9, 5, -18, 5, 9, 12, -6, -2, 21, 14, 1, 3, -11, 0, -5, 25, 7, 0, 2, 15, 13, -1, 2, 19, -9, 1, 0, -4, -14, -13, 3, 5, 0, -13, -33, 6, 8, -11, -44, 1, -7, -8, -7, -3, 10, 15, 6, 7, -17, -6, 5, 13, -14, 4, 9, 14, 16, 18, 11, -4, 2, 2, 1, -5, -3, -6, -4, -1, 6, 1, 1, -5, 4, 9, -3, 0, 1, 0, -4, -3, 2, -2, -1, -5, 2, -6, 0, -7, 5, -3, 0, 4, 7, -3, 0, 10, 13, -4, -28, 4, 6, 5, -28, 9, 12, -17, -28, 7, 3, -13, -26, 10, 1, 12, -7, 6, 1, 22, -8, 21, -2, -6, -20, 8, 0, -1, -8, -6, 1, -6, 7, 10, 1, 5, -2, -2, 0, 3, -3, 6, -8, -7, 19, 15, 3, -14, -3, 10, 2, -9, -3, 10, 7, 1, -2, 14, 19, -13, -27, 11, 0, 9, -7, 28, -3, 0, -18, 11, -1, -11, -14, -5, -4, 23, 39, 12, -23, 2, 14, 11, -17, -15, 24, -3, -3, 4, 27, -1, -13, 10, 21, 12, 2, -12, -5, 0, 7, 0, -9, -6, 3, 5, 0, 16, -14, -1, 2, 4, -6, 19, -3, 11, -1, 12, 4, 7, 4, 7, 11, 14, -5, 1, -18, 6, 1, 28, -11, 18, -9, 12, -11, 12, -18, 2, -9, 6, 3, 5, 8, 8, -5, 9, 6, 8, 0, 12, -1, 2, -8, -1, 7, -5, -1, 11, 11, 0, 3, 16, -6, -2, 3, 13, 0, 0, 2, -4, -9, 0, 3, 5, 4, -4, 6, 2, 3, -1, -1, -3, -1, 6, -7, 0, 5, -6, -3, -1, -1, 8, 8, -6, -13, 6, 11, 1, 0, -1, 8, -7, 9, -3, -5, -4, 9, 2, 9, -9, -1, 9, 17, 5, -4, 1, 10, 1, -5, -8, 6, -5, -2, 7, 2, -1, -3, -2, 4, 4, -3, 0, 6, 5, -3, 5, -13, 4, 20, -1, -15, 4, 13, 14, -4, -4, 22, -5, -6, -2, 19, 25, 9, -24, -44, 9, -1, 18, -28, 10, -1, 24, -22, 19, 0, -15, -35, 6, -7, 2, -6, 0, 0, 5, -5, -6, -5, -2, -3, 0, -3, -6, -2, -6, -2, -2, -8, 3, 12, -11, -17, 10, 5, -10, -20, -9, 3, 10, 8, 12, -2, 6, 11, 1, 3, 3, -2, 3, 8, 0, -11, -7, -1, -6, 1, 7, -2, 7, 2, 0, -6, 4, -1, 1, 0, 5, -7, 0, -2, -3, -7, 1, -9, 5, 13, 2, 3, -10, 6, 3, 10, -5, 4, -3, 0, 0, 7, 6, -7, 0, 4, -3, 7, 5, 7, -6, 3, -4, 7, 2, -1, -3, -7, 1, 0, -7, -13, 12, 4, 14, -5, 14, 4, 12, -4, 3, -8, -4, -13, 0, -7, 0, 10, 9, -5, 7, -6, 2, 7, 10, 7, 2, 6, 1, -8, 22, 9, 0, 4, 10, 2, -4, -4, 15, 17, -5, -1, 4, -6, -10, 4, 8, -8, 4, -20, 21, -4, 30, -7, 16, -5, 18, -5, 8, -11, 0, -14, 5, -6, 0, -9, 13, 6, 6, -5, 19, 1, -12, -10, 16, -2, -7, 6, 21, 6, 32, -3, 23, -27, 8, -2, 20, -33, 11, 1, 27, 6, 42, 3, 4, 1, -20, -17, 8, 11, -19, -50, 8, 19, -4, -47, 0, 8, -19, -38, -1, 1, 4, -1, 0, 1, 0, 0, 0, -7, -3, 0, 6, 5, 7, 6, 22, 7, -16, -34, 25, 3, 10, -18, 8, -4, 7, -10, 17, 5, -13, -37, 14, -8, -15, -7, 18, 12, -15, -20, 1, 1, -9, -7, 11, -1, -23, -21, 0, 1, 1, 23, 1, -5, -5, 10, 4, -5, -6, 22, 9, -16, 11, 18, -9, -9, -9, 9, 11, 0, -15, -17, 5, 4, -1, -30, -4, 4, -12, -8, -7, -11, 3, 0, -3, 1, -7, -10, 7, 17, -8, -3, 0, 8, 6, -1, 14, 8, -17, -13, 10, 6, 12, 2, 10, 12, -4, -10, 23, 4, -10, -4, -3, 0, -7, -22, 1, 6, 13, -5, 14, 16, 0, -16, 0, -7, -13, -18, 2, 5, 0, 14, 2, 9, 5, 5, 3, 15, 3, 1, 0, -7, 5, 1, 8, -4, 4, 7, 3, -6, 0, -3, -7, -3, -2, -5, -4, 6, -5, -2, -4, 3, -1, 0, 6, 5, 4, 2, 5, -4, 4, 1, 8, -4, 4, 1, 6, -6, -2, 2, 2, 11, -11, -26, 0, 6, 0, -17, -5, 5, 9, -6, 30, 15, -10, -1, 16, 13, 7, -2, 9, 1, 2, 15, 11, 6, -18, -16, -5, -6, 4, 1, -2, -2, 6, -7, -4, 0, 0, 3, -1, 3, 5, -4, 11, 5, 0, -6, -7, -4, 9, 11, 9, -5, -1, 6, 10, 3, 0, -11, 11, -3, 13, 3, 9, -7, 8, -6, 22, -7, 8, -5, 5, 9, 21, -12, 28, 6, -13, -36, 8, 5, 8, -12, 6, -11, 11, -11, 20, 6, -8, -25, -8, 7, 16, 17, -3, -15, -6, 11, -7, -19, -2, 22, -1, -4, 27, 15, -7, -12, 21, 11, 2, -17, 3, 30, -2, -23, 7, 24, -5, -7, 31, 31, 4, 0, -5, 4, 0, 7, 5, 8, 3, 8, -2, -1, 11, 8, -7, -5,

    -- ifmap
    -- channel=0
    174, 174, 112, 165, 0, 32, 0, 109, 0, 0, 0, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 78, 0, 0, 6, 89, 5, 88, 50, 50, 0, 161, 63, 68, 812, 370, 192, 154, 921, 191, 41, 0, 1072, 0, 0, 0, 1094, 0, 0, 0, 316, 124, 26, 21, 265, 117, 47, 99, 166, 31, 40, 97, 0, 23, 0, 158, 27, 35, 3, 77, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 277, 252, 344, 4, 462, 292, 386, 57, 866, 784, 959, 1204, 443, 558, 1184, 1304, 0, 0, 0, 19, 0, 92, 95, 0, 0, 76, 12, 1, 612, 445, 463, 482, 349, 369, 248, 370, 67, 126, 101, 281, 0, 0, 0, 106, 0, 0, 0, 0, 770, 711, 625, 346, 570, 516, 433, 136, 564, 388, 675, 859, 0, 0, 406, 349, 912, 812, 445, 374, 779, 667, 341, 285, 506, 336, 152, 198, 93, 0, 0, 0, 225, 347, 259, 540, 287, 247, 217, 599, 121, 319, 145, 600, 0, 134, 0, 738, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 0, 0, 0, 90, 206, 59, 535, 564, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 465, 359, 361, 391, 804, 742, 997, 1147, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 122, 0, 0, 10, 133, 196, 23, 0, 57, 153, 101, 0, 0, 0, 179, 128, 91, 208, 0, 0, 0, 126, 157, 199, 78, 529, 370, 360, 178, 953, 856, 683, 807, 828, 719, 1036, 1228, 503, 0, 0, 0, 756, 0, 0, 0, 1078, 0, 0, 0, 1340, 0, 19, 4, 522, 381, 224, 279, 323, 195, 68, 93, 0, 0, 0, 0, 147, 0, 0, 0, 241, 160, 115, 0, 616, 80, 27, 0, 898, 0, 157, 278, 790, 302, 535, 574, 0, 0, 0, 0, 722, 166, 145, 0, 1188, 474, 652, 713, 1334, 655, 1163, 1215, 267, 169, 336, 166, 628, 297, 375, 155, 618, 463, 413, 663, 605, 654, 424, 774, 34, 118, 62, 136, 0, 22, 12, 86, 0, 104, 180, 84, 23, 0, 0, 0, 140, 151, 131, 128, 74, 62, 80, 45, 0, 111, 7, 88, 0, 0, 0, 0, 273, 330, 267, 238, 160, 150, 88, 109, 4, 159, 47, 275, 0, 0, 0, 11, 350, 327, 187, 343, 31, 74, 61, 269, 0, 0, 0, 155, 0, 0, 0, 0, 351, 245, 149, 122, 189, 59, 8, 82, 40, 0, 0, 36, 0, 0, 0, 0, 304, 106, 41, 0, 598, 154, 0, 0, 882, 53, 42, 197, 958, 0, 129, 156, 0, 0, 0, 0, 125, 0, 0, 0, 581, 289, 229, 334, 829, 710, 1194, 1327, 87, 51, 62, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 904, 878, 598, 564, 483, 512, 269, 386, 0, 0, 0, 101, 0, 0, 0, 0, 0, 0, 0, 100, 0, 16, 0, 66, 0, 22, 149, 112, 315, 350, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 607, 460, 381, 388, 430, 384, 255, 298, 35, 92, 58, 102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 239, 81, 74, 0, 611, 530, 618, 573, 750, 845, 1018, 1057, 166, 92, 124, 11, 139, 85, 84, 1, 129, 50, 137, 139, 203, 106, 71, 0, 0, 0, 0, 0, 0, 0, 10, 26, 6, 0, 0, 0, 1257, 1314, 1106, 1189, 107, 0, 105, 0, 934, 211, 150, 0, 1217, 559, 870, 904, 1403, 903, 1146, 1220, 628, 538, 378, 203, 430, 343, 198, 132, 275, 198, 230, 395, 0, 0, 0, 0, 0, 287, 296, 781, 312, 339, 615, 999, 228, 723, 334, 1632, 83, 941, 0, 2184, 525, 597, 393, 461, 294, 417, 411, 429, 0, 263, 244, 124, 0, 0, 0, 0, 144, 9, 14, 54, 90, 47, 59, 92, 84, 62, 0, 37, 98, 59, 0, 340, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1473, 1368, 1304, 1434, 43, 0, 0, 0, 80, 80, 32, 0, 118, 129, 134, 63, 232, 245, 98, 66, 38, 0, 0, 0, 346, 0, 0, 0, 788, 0, 0, 0, 994, 0, 204, 226, 761, 726, 500, 551, 387, 449, 235, 326, 0, 12, 0, 61, 0, 0, 0, 0, 278, 280, 164, 143, 0, 40, 0, 66, 0, 0, 0, 16, 0, 0, 0, 0, 570, 470, 403, 280, 614, 412, 365, 82, 374, 482, 349, 687, 0, 0, 242, 350, 272, 191, 230, 0, 421, 236, 176, 77, 660, 563, 760, 807, 389, 591, 785, 713, 74, 119, 51, 353, 0, 62, 64, 196, 0, 0, 0, 27, 26, 0, 0, 0, 93, 0, 36, 0, 93, 0, 0, 0, 143, 0, 4, 52, 0, 11, 16, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 706, 688, 418, 349, 424, 425, 136, 306, 0, 0, 0, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 116, 0, 0, 0, 0, 1452, 1332, 1077, 1205, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 141, 111, 160, 131, 189, 131, 174, 201, 53, 221, 514, 416, 427, 517, 0, 161, 120, 438, 205, 205, 309, 497, 110, 409, 278, 829, 52, 506, 0, 1064, 0, 0, 0, 0, 130, 0, 0, 0, 453, 40, 126, 167, 741, 615, 941, 1077, 444, 222, 316, 27, 474, 267, 326, 0, 632, 70, 96, 217, 660, 45, 179, 125, 418, 141, 276, 26, 374, 165, 316, 113, 458, 0, 272, 239, 285, 189, 348, 129, 0, 0, 18, 0, 80, 0, 0, 0, 99, 0, 61, 178, 84, 0, 119, 105, 
    
    
    others => 0);
end inmem_package;
