LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE inmem_package is
		type padroes is array(0 to 4000000) of integer;

		constant input_mem: padroes := ( 
					-- bias
					-- layer=0
					-4005, 1278, -1449, 2196, 29, 2212, 4394, 6249, -784, -8468, -326, 5074, 6285, 2635, -12384, 7587,

					-- weights
					-- layer=0 filter=0 channel=0
					31, 34, 10, -9, -54, -27, 0, 4, 3,
					-- layer=0 filter=0 channel=1
					44, 46, -45, 56, -1, -35, 24, 53, 33,
					-- layer=0 filter=0 channel=2
					32, 24, -55, -52, -61, -19, -58, -38, 11,
					-- layer=0 filter=1 channel=0
					-26, 27, 31, -45, -64, -58, -30, 16, -11,
					-- layer=0 filter=1 channel=1
					23, 24, 37, 15, -40, -40, -10, -45, 7,
					-- layer=0 filter=1 channel=2
					7, 50, -13, 38, 29, 51, -40, 6, 12,
					-- layer=0 filter=2 channel=0
					-49, 19, -13, 32, 5, 36, -1, -5, 11,
					-- layer=0 filter=2 channel=1
					-21, -33, -6, -63, -36, -12, -20, 14, -37,
					-- layer=0 filter=2 channel=2
					50, 9, 39, -31, 6, 55, 45, 24, 36,
					-- layer=0 filter=3 channel=0
					18, 2, -26, 33, 45, -18, 22, -25, -58,
					-- layer=0 filter=3 channel=1
					-8, -5, -62, 55, -4, -46, -26, 30, -62,
					-- layer=0 filter=3 channel=2
					64, 31, 0, 52, 16, -11, 82, 30, -52,
					-- layer=0 filter=4 channel=0
					-27, -58, -26, -10, 43, -21, 77, 43, -6,
					-- layer=0 filter=4 channel=1
					-66, -81, -4, -51, -3, 43, 34, 68, 57,
					-- layer=0 filter=4 channel=2
					-31, -62, -31, 1, 57, 11, 51, -6, -7,
					-- layer=0 filter=5 channel=0
					44, 40, 38, 31, 47, 59, 69, 47, -6,
					-- layer=0 filter=5 channel=1
					27, -17, -16, -26, 24, -28, 33, -8, -43,
					-- layer=0 filter=5 channel=2
					-42, -46, 4, -27, -54, -58, -12, -23, -42,
					-- layer=0 filter=6 channel=0
					25, 0, 28, 4, 48, 51, -42, 13, 68,
					-- layer=0 filter=6 channel=1
					-66, -4, 5, -77, -63, 34, -16, -48, -11,
					-- layer=0 filter=6 channel=2
					9, -28, 28, -68, 16, 37, 15, 0, 14,
					-- layer=0 filter=7 channel=0
					38, 64, 17, 51, 45, -22, 31, 52, 0,
					-- layer=0 filter=7 channel=1
					-16, -51, -10, -11, 9, -55, -60, -69, -45,
					-- layer=0 filter=7 channel=2
					33, 28, 10, -57, -70, 0, -14, -58, 40,
					-- layer=0 filter=8 channel=0
					21, 45, -1, 52, 60, 51, -9, -53, -57,
					-- layer=0 filter=8 channel=1
					47, 3, -34, -8, -9, 23, -47, -55, -59,
					-- layer=0 filter=8 channel=2
					-8, 10, -4, 11, 57, 28, -9, -43, -7,
					-- layer=0 filter=9 channel=0
					3, 2, -5, -6, -8, 22, -63, -59, -16,
					-- layer=0 filter=9 channel=1
					43, 30, -33, 29, 27, 23, 49, 45, -13,
					-- layer=0 filter=9 channel=2
					32, 59, 40, -23, 41, 6, -9, 44, 39,
					-- layer=0 filter=10 channel=0
					20, 61, 37, 37, -11, -46, -15, -40, -56,
					-- layer=0 filter=10 channel=1
					29, 16, 49, 30, -28, 18, 33, -65, -82,
					-- layer=0 filter=10 channel=2
					-26, 29, 69, -13, -36, -38, 53, 16, -53,
					-- layer=0 filter=11 channel=0
					-19, -35, 28, -48, -9, -26, -43, -20, -32,
					-- layer=0 filter=11 channel=1
					-39, -3, 38, -29, -30, -7, 21, 1, 31,
					-- layer=0 filter=11 channel=2
					47, 22, 51, -22, 44, 51, -27, -5, 51,
					-- layer=0 filter=12 channel=0
					-59, -37, 62, -32, -7, 27, -41, 40, -8,
					-- layer=0 filter=12 channel=1
					-41, 5, 38, 3, 10, 75, -13, 58, 48,
					-- layer=0 filter=12 channel=2
					-40, -2, -7, -57, 41, -1, -41, -21, -6,
					-- layer=0 filter=13 channel=0
					-35, -55, -39, -33, -28, 52, -7, 77, -2,
					-- layer=0 filter=13 channel=1
					-42, -1, -65, -20, 25, 19, 61, 3, 27,
					-- layer=0 filter=13 channel=2
					-37, -14, -68, -23, 7, -1, 54, -24, 62,
					-- layer=0 filter=14 channel=0
					-5, 56, 15, 36, 18, 10, 35, 45, 10,
					-- layer=0 filter=14 channel=1
					-28, 16, -6, 21, 41, -47, -9, -3, -47,
					-- layer=0 filter=14 channel=2
					-33, -32, 9, 25, -38, 16, -9, 26, -21,
					-- layer=0 filter=15 channel=0
					-11, 13, -35, 24, -31, -17, 19, -28, -46,
					-- layer=0 filter=15 channel=1
					2, 49, 20, 70, 38, -16, 66, 43, -11,
					-- layer=0 filter=15 channel=2
					-37, -49, -8, -9, -28, -38, 35, -14, -52,

					-- test image
					-- image=0 channel=0 column=0
					40448,40704,42240,42496,40960,39936,41472,40704,40448,40704,41216,40960,41216,42496,43264,43520,42752,41472,40960,40960,39936,38144,38400,37888,38144,36608,35840,36096,36608,35072,32256,29696,
					-- image=0 channel=0 column=1
					38912,38656,40704,42496,41472,40960,41984,41472,41728,39936,39680,40704,41728,43520,43776,43776,43264,40960,39424,38656,37120,35584,35840,36096,38144,37632,37120,36352,36608,34816,32000,30464,
					-- image=0 channel=0 column=2
					38656,38656,40448,42752,40960,41728,42240,42240,41728,41472,40448,40192,41216,42496,42752,43264,43520,40704,37120,30976,28160,25088,25856,29184,30720,34304,36608,35840,36352,35584,33280,30720,
					-- image=0 channel=0 column=3
					39680,39680,40960,44544,42752,42752,43264,43264,42240,42240,42752,48896,45312,40192,41472,41984,40448,38144,26624,26368,25088,23552,20480,18944,22016,21248,28928,33792,35840,35840,34816,32512,
					-- image=0 channel=0 column=4
					39680,39936,41216,43520,43264,41728,43264,42496,41984,41984,44288,62976,49920,38656,37376,36352,28416,19968,21760,28928,28672,27136,24832,23808,18944,21504,21760,26880,32768,35328,34048,33024,
					-- image=0 channel=0 column=5
					37888,34048,33280,37632,41216,42240,42752,42752,41728,42240,41728,46080,40192,32768,24832,16896,17664,16896,22784,30208,31232,30464,29184,24064,25344,23296,14848,17152,27648,35840,35328,34304,
					-- image=0 channel=0 column=6
					32512,27904,12032,22528,39168,43520,43008,43520,43264,42496,41984,37632,33024,32512,25600,17408,19968,18432,21248,33792,37376,31744,26880,27392,29440,21760,16128,11776,20224,33792,36096,34304,
					-- image=0 channel=0 column=7
					33536,25344,10752,17920,36608,42752,42240,43008,43776,41216,35840,30720,33280,36864,29696,22528,23296,21760,19712,31744,41728,34816,26112,27136,25600,21760,13824,12544,14592,27392,35328,34816,
					-- image=0 channel=0 column=8
					43520,26368,13824,31744,39168,41216,41728,42496,42240,44544,28928,32000,40192,39936,30976,22016,20992,21504,20480,20736,35328,37376,28928,22272,21248,22016,18176,14336,10240,18944,34048,35072,
					-- image=0 channel=0 column=9
					46080,34304,24064,39424,44544,40448,39936,39168,52992,60672,52992,39936,44544,37888,32000,23808,22016,18944,15104,19456,35072,36608,34048,27136,22016,22272,21504,19200,12800,10240,24320,33792,
					-- image=0 channel=0 column=10
					46848,27648,36352,42240,45312,39680,40704,31232,54528,60672,56320,41984,46848,39936,32000,30720,19968,20480,11520,23296,44800,40192,39680,27392,22272,26368,22528,19968,15104,10496,15104,26624,
					-- image=0 channel=0 column=11
					48128,25600,34560,43520,47872,42496,44288,34304,29952,49664,50944,43520,47360,48384,34304,29952,26112,21504,9728,32000,53760,40960,37376,23808,21248,24064,26624,21760,18688,14080,15872,19456,
					-- image=0 channel=0 column=12
					48384,23040,32512,44800,44544,42496,45568,40704,24832,43008,43008,35072,47616,55296,40960,31488,30720,29440,12800,38400,49664,39680,31488,23296,21504,21504,24320,22016,21504,18688,20224,18688,
					-- image=0 channel=0 column=13
					48384,23808,38912,47360,30464,34816,44288,42752,26368,37632,37120,42752,48384,57856,46080,36096,32256,29952,18176,39424,47616,38144,29184,22272,20480,18432,20480,25344,25600,23040,24832,24064,
					-- image=0 channel=0 column=14
					49664,27648,43008,47616,26880,25344,39936,42752,25600,29440,35328,50688,48640,44032,37120,39424,37376,26368,18176,38912,45824,35072,33280,28160,21760,23296,24320,27904,29440,25600,24832,29952,
					-- image=0 channel=0 column=15
					50432,33792,44032,47104,33280,19968,35840,39680,29440,33280,36608,58880,61952,37120,34560,33536,30976,27648,24320,36864,43008,38912,28672,22272,18176,22272,26880,28672,30720,26368,30976,34816,
					-- image=0 channel=0 column=16
					51968,37376,43008,48896,43008,19968,32256,35328,35328,24576,39424,44288,41472,35840,28928,28928,25856,26880,28672,43776,39936,37888,34560,27904,19968,20224,24064,25856,27392,32000,38656,36864,
					-- image=0 channel=0 column=17
					54784,41728,41984,46848,45056,24064,24576,39936,37888,27136,33024,30208,29184,29696,26112,29440,22016,25856,36864,30208,17408,32768,34048,19200,15360,14848,18176,26112,29696,36608,38400,35840,
					-- image=0 channel=0 column=18
					54272,45568,42752,44288,45056,31744,22016,36096,39168,34560,26624,19712,34304,31744,33024,37632,21760,23552,38400,33792,29952,27392,19200,16384,11264,16640,22016,34048,39680,40960,39424,38656,
					-- image=0 channel=0 column=19
					50944,47872,43776,44544,45312,36864,22016,30464,31232,35072,36864,17920,33024,27648,37120,47104,29696,18688,33536,35072,34304,22784,13056,13312,12032,23040,30976,41728,43776,41984,40448,38144,
					-- image=0 channel=0 column=20
					42240,49920,45824,45312,46336,38912,25344,33536,43776,26368,23808,20480,23808,31232,45568,48896,38400,25600,22784,22272,15360,11776,9728,6144,11776,15360,27648,36864,36864,32768,32512,30720,
					-- image=0 channel=0 column=21
					29952,49920,45312,45568,46336,35328,21248,38400,62720,56064,34048,34304,38144,45056,48640,49664,43008,32000,28160,15616,8960,8704,12544,14848,15616,14848,17664,18432,19968,17664,15104,14080,
					-- image=0 channel=0 column=22
					20224,44800,44544,45056,45312,35840,27904,54016,64768,64512,53248,31744,29184,31744,29696,31232,26624,17408,17408,15360,13312,12800,13056,14336,14336,13056,11008,13056,15104,12288,11008,10752,
					-- image=0 channel=0 column=23
					10496,24576,36864,43008,45568,42240,42240,62976,64768,58112,28160,15360,13568,12544,12544,12288,11520,10752,11776,10752,9728,11776,11776,11008,10752,11776,11776,12800,14080,13568,13056,11520,
					-- image=0 channel=0 column=24
					7424,7424,15104,33536,42496,33792,49664,65024,61696,36096,15616,12800,12800,13056,12544,12800,12032,10752,9984,8704,8960,9984,9728,10752,11520,14336,15872,15104,14336,12800,11776,13056,
					-- image=0 channel=0 column=25
					12288,7680,8704,18688,32768,32768,55040,65280,47872,16896,13824,12800,13312,13312,11776,11520,11008,10496,9216,9984,10240,10240,11008,11776,15104,15872,16384,15104,13824,12800,17920,21248,
					-- image=0 channel=0 column=26
					13312,8960,7936,10496,16896,32768,57344,61440,31744,14848,12544,14336,13824,11264,11264,12032,11776,11008,11008,11264,11264,11520,13824,14848,13824,11776,11008,9216,13056,18688,21760,19456,
					-- image=0 channel=0 column=27
					12800,8960,7424,8960,11264,19968,51712,54016,24832,16640,13824,12288,14848,12288,10240,11520,12032,12288,12032,11776,13056,9984,9984,12288,12032,9984,7168,10240,17152,17152,11776,13056,
					-- image=0 channel=0 column=28
					12800,8960,8192,8448,10496,11776,26624,43520,16384,13824,13312,13568,15616,14848,13824,11520,10752,10496,11776,12544,11776,10752,10240,9984,9472,10240,11264,16128,12032,7936,3840,13056,
					-- image=0 channel=0 column=29
					17408,10752,7936,9728,9472,11008,10752,18176,12544,7936,6912,9728,12544,14336,14848,13568,14336,15360,14592,13568,12800,11520,9984,8448,10752,15872,20224,18688,14336,9728,3328,10240,
					-- image=0 channel=0 column=30
					15616,12544,8960,11008,9984,10752,11264,10240,10752,6912,5888,7680,6912,7424,9216,12032,14336,15872,16896,19200,17664,12544,11008,11008,15360,21760,27904,23808,15360,6656,7424,5120,
					-- image=0 channel=0 column=31
					13824,14336,11520,11008,10240,10240,10240,9728,9216,6656,5632,7424,6400,7424,4864,4608,8192,12032,15616,18944,16896,13568,13312,11520,17152,22784,26880,22784,12288,6144,8704,5376,
					-- image=0 channel=1 column=0
					28672,28416,29696,30208,28672,27904,29440,28928,28416,28928,29696,28416,28416,29952,29952,30464,29952,28928,28416,28672,27904,27392,27392,27136,27392,25856,25088,24832,24832,24320,23296,21760,
					-- image=0 channel=1 column=1
					28672,28160,29184,29696,28672,28928,29952,29184,29696,28160,28416,28160,28928,30464,29952,29440,29440,28416,28672,29440,28160,26624,26112,25600,26880,26112,26112,24832,25088,24320,23296,22528,
					-- image=0 channel=1 column=2
					28160,27904,28416,28416,27136,29440,29952,29952,29440,29440,29184,27904,28416,29440,29184,28928,29696,29184,28416,24576,23040,19968,19712,21760,22016,24576,26368,25344,25344,25088,24320,22784,
					-- image=0 channel=1 column=3
					27392,28160,27904,28672,28160,29952,30720,30464,29440,29952,31488,37376,33280,28416,29440,29184,28672,28416,20480,22272,23040,23040,19200,16128,17920,15872,21760,25088,26112,25856,25344,24064,
					-- image=0 channel=1 column=4
					27392,29184,29440,29184,29184,28928,30720,29696,28928,29696,32768,54784,39936,29184,28416,27648,20480,13568,17664,26368,28160,29184,26112,24064,18432,19968,18688,21248,24576,25856,24064,23808,
					-- image=0 channel=1 column=5
					27904,26624,25600,28672,29440,28928,29696,29440,28416,29696,30208,35328,31232,26112,19200,12800,14848,14336,21248,28928,30976,31232,29696,24576,25600,23296,14848,14848,21504,26880,25088,24320,
					-- image=0 channel=1 column=6
					25600,24320,9472,18944,29952,30208,29440,30208,29952,29696,30720,27392,25088,27648,22272,17152,21248,19200,21504,33280,36352,30208,25344,26112,28416,21248,18176,12032,15616,25088,25344,23808,
					-- image=0 channel=1 column=7
					29440,24576,11008,16384,28416,29952,29184,29696,30464,28928,27904,24064,28160,33536,27136,22272,24320,22528,19712,30208,39168,31744,23808,25088,23808,20736,15360,13568,12032,21248,26368,24832,
					-- image=0 channel=1 column=8
					41216,26880,14848,30976,31744,28928,29952,31232,30976,34560,22784,26880,36096,36608,28416,20480,20736,21760,19968,18176,32000,34560,26368,20224,19712,20992,18688,14592,8960,15104,27136,26368,
					-- image=0 channel=1 column=9
					45056,35584,25600,39424,38144,29696,29696,30208,46080,54784,46080,33536,39168,33536,28160,21760,21504,18944,14592,17408,32000,34048,31744,25088,20736,21760,21760,19456,12544,7680,19200,26368,
					-- image=0 channel=1 column=10
					46848,29696,38656,43264,39936,28672,30208,22784,50432,57344,48896,34560,40704,35072,27648,28416,19456,20480,11264,21760,42240,37632,37632,25600,21248,26112,22528,20224,15104,9216,11776,20736,
					-- image=0 channel=1 column=11
					48896,27648,36864,44800,42752,30720,31488,23808,24320,46592,43776,36352,41216,43776,30464,27392,25088,21504,9728,30976,51456,38912,35584,22784,20480,23808,26624,22272,19200,13568,14080,14336,
					-- image=0 channel=1 column=12
					49664,24576,34304,46080,39936,31488,31488,27904,17408,39424,36864,29184,42496,51712,38144,28928,29184,29184,12800,37632,47872,38144,30208,22528,21248,21504,24320,22272,22272,18688,18944,14080,
					-- image=0 channel=1 column=13
					49152,24320,39424,48128,28160,27136,31744,29696,18432,33792,32000,38144,44544,55296,44032,33536,29952,29184,18176,38912,46336,36864,28160,21760,20480,18688,20480,25600,25856,22528,22784,18688,
					-- image=0 channel=1 column=14
					50176,27392,42752,47616,27904,22784,30464,31232,18944,27136,31488,47360,46080,42240,35840,36608,34816,25600,18176,38912,44800,34048,32768,27904,22016,23808,24576,28160,29696,24576,21760,24320,
					-- image=0 channel=1 column=15
					50432,33024,42752,45568,35072,21248,30720,32000,24064,30720,33536,56576,60416,35328,33280,30976,28672,26624,22528,34304,40704,37632,27648,21760,18432,22528,26624,27904,28160,22016,24576,26624,
					-- image=0 channel=1 column=16
					51968,37376,41984,46592,43520,22016,32000,32256,30976,20480,36608,41728,38912,33792,27136,27136,25856,25856,23040,36608,35328,36096,33280,26880,19456,20224,23808,23296,21248,22528,27648,26624,
					-- image=0 channel=1 column=17
					55040,42496,42752,47104,46592,26112,24576,38144,35072,23808,29696,26880,26112,26880,23296,28160,23296,26368,32768,24576,14336,30720,32256,17664,14336,14336,17920,23808,24064,28672,29696,28160,
					-- image=0 channel=1 column=18
					54016,47104,44800,46336,47104,33536,22528,35584,37888,32768,23040,16384,30976,28416,29952,36608,23552,24576,35584,29952,27904,25344,17408,15104,10496,15872,17664,26880,30464,30720,29440,28416,
					-- image=0 channel=1 column=19
					49152,48384,45056,45824,46592,38144,23040,30976,31744,34816,34304,15104,30208,24832,34304,45056,30208,19200,30464,31744,33024,22016,12544,13056,12544,23040,23296,30208,30976,28928,28416,27392,
					-- image=0 channel=1 column=20
					39936,49408,45568,44288,46336,40192,26368,34560,44800,26880,23040,19712,23040,30208,44288,46592,37888,25600,19968,19712,15616,13312,11776,8448,14592,18176,25600,32000,31488,27904,28928,26880,
					-- image=0 channel=1 column=21
					30720,51200,45568,43264,45824,36864,22272,39168,63232,56832,35840,36096,39936,46592,50176,49152,44032,34048,27904,15872,12544,13824,17920,20736,21760,21504,25344,25856,26624,24576,23552,23040,
					-- image=0 channel=1 column=22
					26880,50432,46848,44032,45312,37376,28672,54016,64512,64768,57344,36608,33792,36096,34048,34048,31744,23808,22272,20992,21504,21504,21760,23808,24064,23296,24576,26624,27648,24832,24832,24320,
					-- image=0 channel=1 column=23
					22784,35072,43008,44544,46592,43520,42496,62720,64256,59136,34816,22528,20480,19456,19200,18432,20224,20736,20736,20992,22016,23040,22784,22272,22784,23808,24064,24576,24576,24064,24320,23040,
					-- image=0 channel=1 column=24
					23296,22272,26112,39168,45824,34816,48384,64000,62720,40704,24064,21504,21504,21760,21248,21504,22016,21504,20992,20224,21248,22016,21760,22784,23552,26368,26368,25856,26112,25344,24064,26368,
					-- image=0 channel=1 column=25
					28416,24064,21760,27136,37888,34816,54528,64768,50688,23808,23296,22528,23040,23040,21248,20992,20992,20736,20480,21248,22016,22784,23552,24320,27648,28160,27904,27648,27648,26880,31488,35072,
					-- image=0 channel=1 column=26
					29184,25344,22016,21248,24320,37120,58624,62720,36608,23552,22272,24064,23552,20992,20992,21248,21504,21248,22016,22528,23040,24832,27136,28160,26880,24832,24320,23296,27648,33280,35328,32000,
					-- image=0 channel=1 column=27
					28160,25088,22784,22016,21248,27136,56064,58368,32256,26624,24064,22272,24832,22272,20480,20992,21504,22272,22784,22784,24832,23552,23808,26112,25856,23808,21760,25856,33024,32256,25088,24576,
					-- image=0 channel=1 column=28
					27648,24832,23552,22528,22528,21504,34048,50432,25600,24832,24064,24320,26368,25600,24576,21248,20224,20480,22528,23552,23552,24320,23808,23552,23040,23808,26112,32000,28160,23040,15360,23808,
					-- image=0 channel=1 column=29
					31744,25600,22528,23296,22272,22784,20224,27392,22784,19712,18176,20992,23808,25600,26112,23552,24064,25344,25344,24832,24320,24064,22528,21248,23296,28672,33792,33536,29696,24832,16384,21760,
					-- image=0 channel=1 column=30
					29696,26112,21760,23296,23040,23552,22528,20736,21760,18432,17152,18944,18176,18688,20480,22016,24320,25856,27904,30464,28928,24320,22528,22528,26880,33280,39936,37120,29440,20992,20992,16384,
					-- image=0 channel=1 column=31
					27392,26880,22784,22016,22784,23552,22272,20736,20224,17664,16896,18688,17664,18688,16128,14848,17920,22272,26624,30464,28416,24576,24320,22272,27904,33536,37376,34560,25344,19712,21504,17152,
					-- image=0 channel=2 column=0
					12544,12032,13056,13568,11776,10496,12032,11520,11264,10496,10496,13312,12544,10496,11520,11264,10240,9728,9984,11008,11264,11520,11520,11008,11264,9984,11008,10496,9728,9216,9216,8448,
					-- image=0 channel=2 column=1
					13056,10240,11520,14336,12544,11008,12032,11520,11776,9728,10496,13824,13312,10496,10240,8448,7680,8448,10496,12800,13568,14080,13312,12288,12800,11776,11520,9728,8704,7936,8192,8704,
					-- image=0 channel=2 column=2
					12032,8448,9216,12288,10752,11264,11520,11520,11008,11008,12288,14592,13056,9728,9472,8960,9984,12032,13824,12544,13312,12800,12032,12800,12288,14080,13056,9984,8960,8704,8704,8448,
					-- image=0 channel=2 column=3
					10240,8192,7936,11264,11008,11776,12288,12288,11264,11520,14592,24320,19200,10496,12032,13824,14848,17152,12032,16640,19456,21504,16896,12800,13312,9984,11520,11776,11008,9984,9984,9216,
					-- image=0 channel=2 column=4
					10496,12288,12544,12032,11008,10240,12032,11264,10496,10752,15104,41984,27392,14336,15360,18176,12800,7936,14336,25088,28416,30208,26880,23808,17152,17920,12032,11520,12288,11776,9216,9216,
					-- image=0 channel=2 column=5
					13824,16384,14592,13568,11264,9984,10496,10496,9472,9984,10752,21760,19968,14848,11008,7936,11008,11520,19456,28160,30720,31232,29696,24576,24832,22016,12032,9472,12544,14848,11264,10240,
					-- image=0 channel=2 column=6
					14592,20480,4352,7168,12288,11008,10240,11008,10752,9472,9984,13312,15104,19200,17920,14592,18432,16384,18944,30976,33792,27648,23040,24064,26368,19712,17664,9984,9216,14848,12288,9984,
					-- image=0 channel=2 column=7
					23040,23552,9728,10496,14336,10752,9216,9984,12544,13056,13056,12544,19712,27392,23808,20224,22528,20992,17664,27392,35840,28672,20736,22528,21504,18944,14848,12544,8192,12800,13056,9984,
					-- image=0 channel=2 column=8
					36864,26880,15104,28928,20992,11008,10496,12800,16896,24320,15104,19968,30976,32768,25856,18944,19712,20992,18688,15616,28672,31488,23808,17920,17664,19456,17152,13568,6912,8960,15104,11520,
					-- image=0 channel=2 column=9
					41728,36608,26880,38144,28672,13056,12032,15360,37376,50688,42496,30464,37120,32000,27392,20224,20224,18176,13568,14848,28672,31232,29184,22784,18944,19968,19968,18176,11008,3840,11264,14592,
					-- image=0 channel=2 column=10
					44800,31232,40448,43008,31232,12800,13056,12032,45824,57856,48128,33536,39680,33792,26624,26624,17664,19712,10240,19712,39424,35072,35328,23552,19712,24576,20224,18688,15104,8448,7936,11776,
					-- image=0 channel=2 column=11
					48384,29696,39168,45568,34816,15104,14080,11264,20480,48128,41984,34048,38656,40704,27136,24320,22784,20224,8704,28928,49152,36352,33280,20992,19200,22528,24064,20736,19968,14080,12288,6656,
					-- image=0 channel=2 column=12
					49664,26880,36864,47360,34048,17408,13568,12032,11264,38912,32256,24064,37888,46848,33024,25088,26880,27904,12032,35840,45568,35840,28416,21248,20224,20480,21760,20736,22784,18688,16384,6144,
					-- image=0 channel=2 column=13
					49408,26368,41728,49152,25088,16896,14848,12800,9984,30720,26368,32512,39680,51200,40192,29952,27392,27904,17408,37632,44544,34816,26624,20480,19456,17920,18432,24064,25344,20736,17664,8704,
					-- image=0 channel=2 column=14
					50176,28672,44032,48128,27904,17152,15872,14080,8704,22528,26368,43264,43264,40704,35840,34304,32000,24320,17920,38144,43520,32512,31232,26880,21248,23296,23040,26624,28416,20480,13568,12032,
					-- image=0 channel=2 column=15
					50432,34816,44544,46336,36352,19712,22528,19712,13312,23808,29696,54016,58880,35072,33280,28672,25856,24320,19200,30208,37376,35328,25856,20480,17408,22272,25344,25344,23808,13824,12288,12288,
					-- image=0 channel=2 column=16
					52224,40960,45568,48128,44032,23040,32256,28928,20992,9472,34048,39680,36096,29952,22528,23040,23552,22272,14848,26624,27904,32256,30208,24832,18432,19712,24064,20992,14080,11520,14080,11776,
					-- image=0 channel=2 column=17
					55040,46080,47104,49664,47616,26880,26112,37120,28416,15616,26880,24320,22784,22784,18688,25088,22528,24320,26112,16384,8192,26880,29440,15616,13056,13568,16640,19968,16384,17408,16384,13824,
					-- image=0 channel=2 column=18
					52480,49152,48384,49408,48128,34048,24576,36608,36096,28416,20480,14080,27648,24576,25600,34048,23808,23808,30720,23808,23552,22016,14848,13312,9984,15360,10240,15104,15872,13824,11520,11776,
					-- image=0 channel=2 column=19
					46080,47872,46336,47360,47104,38912,25344,33792,33280,34560,32256,13056,27648,22016,31488,43008,30208,18688,26368,26880,30208,19968,11264,12800,13312,23808,15360,17408,16384,13312,12800,11776,
					-- image=0 channel=2 column=20
					37376,47872,44800,44032,46080,40960,28416,37376,47360,28416,22272,18688,22016,29696,44288,45312,37888,25856,16896,16128,14592,13824,13056,10496,17664,21248,19200,20992,19456,15616,17664,16128,
					-- image=0 channel=2 column=21
					31744,51200,45056,43008,45824,37632,23296,40704,64000,57600,36864,37632,41984,49152,53248,50432,46336,36608,27904,15872,14848,17408,22272,26112,28160,28416,31232,30464,30720,28672,28672,29440,
					-- image=0 channel=2 column=22
					34048,54528,49152,45312,46592,38400,28928,53504,63232,64512,59392,40192,38144,41472,39936,38912,37888,30464,26624,25856,28416,28160,29440,32000,33536,33280,34560,36096,36352,33792,35072,33792,
					-- image=0 channel=2 column=23
					34560,43008,48128,48128,49152,44544,41984,60672,61696,58368,39168,28416,26880,26880,27392,25856,29440,30720,28928,29696,32000,32000,32256,32768,33792,35584,35072,35072,34560,34304,35584,34048,
					-- image=0 channel=2 column=24
					36096,33280,34304,45056,48896,35072,46336,61952,62720,44800,32512,30208,30464,30976,30720,29696,29952,29952,29440,28928,30720,32000,32000,33280,34304,37120,36352,36352,37376,36864,35840,38144,
					-- image=0 channel=2 column=25
					41472,35840,31744,34816,42752,36608,53504,63744,52480,30208,32768,32000,32512,32512,30976,29440,28928,28672,28928,29952,31488,33536,34304,35328,38400,38912,37632,38144,39424,38912,42752,46592,
					-- image=0 channel=2 column=26
					42240,37632,33280,31232,32256,41984,59904,63232,39168,29184,31488,33536,33024,30464,30464,30464,30464,30464,31488,32512,33536,36096,38400,39424,38400,36096,35840,35328,40448,45568,46592,43264,
					-- image=0 channel=2 column=27
					41472,38144,35328,34048,32256,35328,59648,59904,35840,32256,33024,31744,34048,31488,29696,30464,31232,32256,33280,33792,35840,35328,35584,37888,37632,35584,34048,39168,46592,45056,36352,35584,
					-- image=0 channel=2 column=28
					41216,37632,36608,36096,35328,32000,40704,54016,30464,30976,32768,33280,35584,34560,33536,30720,30208,30720,33280,34560,34816,35584,35328,34816,34560,35328,38656,45568,41984,35840,26368,34816,
					-- image=0 channel=2 column=29
					45312,37888,35072,37376,35584,33792,28928,34048,29184,26880,26880,29952,32768,34560,35072,32768,33536,35072,35584,35328,35072,34816,33536,32000,34048,39424,45824,46336,43008,37376,27648,32512,
					-- image=0 channel=2 column=30
					43008,37888,33792,36608,35584,34304,32000,28672,29440,26624,26112,27904,27136,27648,29440,30720,32768,34560,36864,39936,38912,34304,32512,32512,36864,43520,50432,48640,41984,33280,32256,27392,
					-- image=0 channel=2 column=31
					40960,38144,33792,34304,34304,33792,31488,29440,29184,26880,25856,27648,26624,27648,25088,22784,25600,30208,35072,38912,37120,33536,33280,31488,37120,42752,46592,44800,37120,31744,33024,28160,

					others=>0 );
END inmem_package;
