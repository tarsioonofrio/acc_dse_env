LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE gold_package is
		type padroes is array(0 to 4000000) of integer;
		constant gold: padroes := ( 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 26, 26, 5, 3, 12, 0, 8, 23, 17, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 11, 18, 27, 23, 27, 26, 30, 
		39, 0, 0, 0, 2, 25, 24, 20, 20, 27, 32, 40, 35, 32, 45, 
		46, 34, 0, 0, 14, 25, 25, 25, 26, 32, 28, 31, 32, 49, 28, 
		45, 39, 10, 0, 9, 16, 24, 30, 29, 31, 30, 29, 38, 48, 46, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 2, 1, 0, 0, 48, 9, 0, 0, 0, 23, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 7, 11, 16, 0, 0, 
		13, 44, 6, 0, 0, 0, 32, 10, 4, 0, 0, 0, 0, 0, 1, 
		27, 92, 15, 16, 112, 66, 0, 0, 0, 10, 23, 15, 11, 17, 0, 
		0, 10, 5, 0, 0, 0, 21, 13, 14, 61, 0, 0, 0, 9, 30, 
		0, 3, 0, 0, 0, 15, 0, 6, 0, 39, 0, 0, 0, 14, 20, 
		0, 15, 20, 23, 23, 26, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
		0, 9, 0, 17, 0, 0, 0, 0, 21, 0, 0, 0, 0, 9, 30, 
		0, 0, 0, 19, 0, 0, 4, 57, 0, 0, 0, 0, 42, 37, 0, 
		0, 0, 0, 67, 119, 92, 46, 0, 0, 2, 25, 57, 32, 0, 0, 
		0, 0, 25, 70, 0, 0, 0, 0, 0, 0, 2, 0, 4, 0, 0, 
		9, 0, 0, 0, 0, 0, 2, 0, 0, 6, 14, 20, 6, 0, 26, 
		0, 5, 0, 0, 0, 4, 9, 1, 0, 4, 0, 0, 0, 14, 0, 
		0, 0, 0, 0, 0, 0, 0, 2, 23, 19, 2, 0, 42, 27, 3, 
		
		28, 24, 23, 25, 24, 25, 29, 29, 21, 19, 21, 20, 21, 29, 21, 
		24, 27, 22, 27, 18, 0, 44, 22, 24, 4, 18, 29, 27, 22, 20, 
		17, 20, 26, 29, 20, 14, 37, 41, 10, 0, 5, 9, 21, 23, 14, 
		48, 0, 37, 22, 18, 12, 3, 5, 0, 0, 22, 6, 13, 22, 4, 
		39, 0, 51, 0, 0, 10, 31, 17, 11, 0, 16, 28, 0, 17, 12, 
		33, 0, 59, 0, 0, 26, 19, 23, 24, 0, 27, 38, 0, 8, 21, 
		37, 12, 53, 31, 0, 0, 1, 19, 31, 0, 43, 24, 3, 0, 18, 
		21, 14, 47, 31, 0, 0, 37, 13, 24, 0, 17, 31, 0, 0, 27, 
		16, 0, 44, 0, 9, 22, 31, 0, 6, 33, 0, 34, 0, 12, 14, 
		0, 0, 41, 0, 33, 6, 0, 0, 17, 0, 27, 9, 0, 0, 25, 
		0, 0, 46, 0, 17, 1, 0, 0, 28, 17, 0, 0, 0, 4, 14, 
		0, 0, 20, 0, 33, 35, 6, 5, 3, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
		
		22, 20, 25, 18, 19, 21, 22, 23, 18, 10, 12, 23, 20, 14, 13, 
		19, 24, 27, 16, 30, 8, 0, 9, 11, 18, 0, 0, 13, 23, 11, 
		0, 50, 22, 19, 25, 34, 0, 0, 10, 39, 0, 0, 0, 15, 27, 
		0, 47, 11, 29, 0, 34, 0, 0, 0, 65, 0, 0, 0, 0, 61, 
		0, 0, 0, 89, 0, 2, 0, 0, 0, 87, 0, 0, 0, 0, 31, 
		0, 0, 0, 31, 52, 15, 0, 0, 0, 124, 0, 0, 9, 0, 0, 
		0, 0, 0, 0, 64, 35, 0, 0, 0, 99, 0, 0, 2, 4, 0, 
		0, 0, 0, 0, 53, 40, 0, 0, 0, 71, 0, 0, 18, 0, 4, 
		0, 0, 0, 11, 0, 28, 0, 0, 19, 0, 0, 0, 22, 22, 17, 
		0, 0, 0, 43, 0, 21, 41, 0, 0, 0, 0, 4, 19, 33, 5, 
		22, 0, 0, 99, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 
		29, 21, 0, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 29, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 4, 1, 0, 0, 0, 
		0, 0, 0, 0, 0, 26, 0, 0, 1, 20, 19, 0, 0, 2, 0, 
		0, 9, 0, 0, 0, 20, 0, 0, 14, 64, 46, 34, 11, 6, 4, 
		0, 26, 0, 0, 0, 16, 30, 24, 25, 79, 27, 33, 11, 0, 23, 
		47, 76, 0, 59, 83, 58, 32, 12, 8, 68, 49, 16, 24, 3, 3, 
		63, 90, 0, 9, 110, 76, 51, 26, 0, 125, 50, 13, 38, 22, 6, 
		66, 66, 17, 0, 70, 89, 87, 41, 12, 121, 41, 17, 27, 46, 17, 
		86, 72, 36, 0, 60, 131, 34, 44, 19, 78, 51, 10, 46, 38, 5, 
		96, 109, 30, 76, 22, 47, 26, 29, 54, 0, 47, 0, 19, 22, 10, 
		101, 108, 36, 89, 46, 30, 62, 60, 32, 39, 2, 11, 45, 26, 1, 
		124, 99, 33, 154, 88, 74, 125, 96, 50, 9, 32, 57, 66, 54, 41, 
		119, 123, 89, 170, 83, 48, 57, 54, 58, 60, 70, 74, 79, 81, 77, 
		76, 105, 135, 117, 30, 69, 67, 62, 62, 70, 80, 86, 90, 94, 100, 
		80, 80, 143, 72, 63, 74, 64, 66, 73, 78, 81, 87, 81, 106, 90, 
		75, 86, 80, 55, 51, 72, 78, 72, 82, 79, 74, 77, 112, 97, 64, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 66, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
		0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		
		9, 0, 2, 6, 6, 0, 7, 8, 6, 13, 20, 5, 5, 13, 12, 
		1, 0, 0, 8, 0, 0, 45, 8, 37, 0, 3, 8, 0, 0, 7, 
		25, 0, 4, 5, 1, 0, 47, 22, 0, 0, 26, 16, 40, 0, 0, 
		79, 0, 10, 0, 7, 0, 0, 40, 14, 0, 54, 18, 36, 30, 0, 
		97, 0, 65, 0, 0, 42, 52, 47, 26, 0, 4, 70, 0, 34, 0, 
		121, 0, 84, 35, 0, 55, 27, 37, 45, 0, 91, 88, 0, 25, 28, 
		116, 13, 31, 48, 0, 0, 8, 57, 59, 0, 95, 50, 0, 0, 38, 
		88, 10, 67, 21, 0, 0, 124, 26, 44, 0, 49, 54, 0, 7, 27, 
		72, 0, 137, 0, 54, 17, 23, 0, 0, 34, 0, 83, 0, 0, 0, 
		12, 3, 104, 0, 57, 51, 0, 0, 45, 29, 76, 8, 0, 0, 28, 
		0, 14, 101, 0, 82, 39, 0, 40, 101, 47, 0, 0, 0, 0, 14, 
		0, 0, 51, 0, 148, 90, 3, 5, 18, 3, 0, 0, 0, 0, 12, 
		34, 0, 0, 5, 163, 5, 13, 6, 6, 0, 0, 0, 9, 7, 0, 
		34, 1, 0, 62, 51, 0, 19, 6, 0, 0, 6, 1, 13, 0, 41, 
		50, 0, 8, 0, 27, 0, 5, 10, 0, 0, 20, 0, 0, 15, 63, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 6, 8, 12, 0, 0, 
		0, 5, 0, 0, 0, 2, 0, 0, 9, 64, 7, 9, 0, 19, 0, 
		0, 55, 0, 0, 0, 0, 0, 0, 17, 78, 0, 14, 0, 0, 43, 
		0, 56, 0, 20, 5, 0, 0, 0, 9, 76, 2, 0, 19, 0, 32, 
		0, 49, 0, 0, 83, 0, 0, 0, 0, 146, 0, 0, 33, 6, 0, 
		0, 29, 0, 0, 73, 45, 22, 0, 0, 147, 0, 0, 25, 30, 0, 
		0, 13, 0, 0, 31, 93, 0, 21, 0, 85, 0, 0, 42, 23, 0, 
		7, 57, 0, 51, 0, 27, 0, 13, 35, 0, 26, 0, 30, 3, 0, 
		30, 45, 0, 88, 0, 20, 42, 8, 13, 15, 0, 22, 49, 19, 0, 
		110, 40, 0, 139, 0, 13, 105, 56, 0, 19, 47, 67, 84, 87, 56, 
		162, 98, 5, 137, 0, 20, 75, 70, 56, 75, 85, 90, 85, 87, 78, 
		84, 141, 103, 64, 0, 72, 71, 72, 71, 80, 91, 94, 95, 97, 101, 
		79, 98, 177, 34, 40, 83, 64, 73, 82, 87, 93, 97, 88, 119, 98, 
		70, 97, 96, 80, 65, 92, 87, 75, 83, 81, 72, 85, 111, 86, 53, 
		
		109, 113, 116, 114, 115, 108, 117, 127, 115, 82, 65, 76, 86, 97, 98, 
		113, 119, 123, 115, 120, 103, 94, 84, 53, 47, 14, 22, 46, 72, 88, 
		49, 78, 118, 121, 123, 105, 51, 40, 33, 41, 14, 18, 1, 37, 75, 
		0, 70, 100, 121, 88, 78, 36, 19, 8, 54, 12, 24, 6, 6, 69, 
		0, 35, 78, 128, 41, 51, 22, 14, 3, 68, 35, 8, 20, 0, 41, 
		2, 20, 71, 93, 63, 53, 22, 29, 0, 85, 6, 3, 24, 7, 9, 
		18, 0, 54, 68, 74, 65, 17, 16, 0, 63, 0, 8, 21, 23, 16, 
		13, 2, 23, 32, 76, 48, 0, 22, 15, 80, 17, 9, 26, 24, 66, 
		0, 8, 0, 26, 31, 42, 36, 21, 37, 37, 40, 0, 28, 66, 92, 
		19, 21, 0, 33, 0, 30, 51, 9, 24, 18, 0, 2, 21, 74, 78, 
		8, 19, 0, 82, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 5, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
		3, 3, 0, 0, 0, 39, 19, 0, 0, 9, 34, 23, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 5, 13, 10, 0, 0, 11, 0, 0, 
		33, 32, 4, 2, 9, 13, 29, 4, 0, 0, 0, 0, 0, 0, 0, 
		29, 38, 10, 11, 55, 46, 7, 5, 0, 10, 30, 20, 6, 10, 0, 
		0, 0, 4, 0, 0, 0, 20, 20, 23, 11, 0, 0, 0, 5, 25, 
		20, 0, 0, 0, 0, 14, 0, 9, 3, 0, 0, 15, 9, 12, 7, 
		21, 9, 34, 25, 2, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
		12, 0, 13, 0, 21, 0, 1, 17, 2, 26, 0, 0, 0, 0, 5, 
		0, 0, 8, 20, 0, 0, 12, 38, 9, 0, 0, 0, 5, 9, 0, 
		0, 3, 3, 29, 80, 60, 0, 0, 0, 21, 35, 33, 13, 2, 5, 
		0, 0, 2, 16, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 
		3, 0, 0, 0, 0, 0, 0, 0, 0, 4, 8, 10, 0, 0, 14, 
		0, 3, 0, 0, 0, 1, 10, 1, 0, 0, 0, 0, 0, 5, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 5, 15, 1, 0, 21, 15, 0, 
		
		68, 72, 68, 71, 68, 65, 76, 71, 68, 70, 59, 53, 51, 59, 51, 
		63, 68, 74, 76, 68, 74, 90, 77, 59, 20, 36, 35, 31, 41, 53, 
		79, 39, 68, 71, 72, 100, 59, 21, 9, 34, 78, 46, 50, 25, 40, 
		64, 8, 73, 69, 76, 29, 70, 45, 34, 51, 78, 56, 28, 19, 19, 
		79, 86, 93, 51, 123, 108, 101, 52, 36, 0, 82, 66, 30, 26, 15, 
		94, 106, 96, 75, 95, 100, 107, 67, 46, 20, 127, 58, 38, 35, 14, 
		80, 134, 68, 71, 60, 72, 147, 80, 72, 57, 104, 50, 25, 31, 50, 
		103, 108, 75, 61, 53, 137, 127, 79, 48, 73, 88, 56, 31, 60, 41, 
		127, 120, 91, 60, 70, 60, 56, 56, 38, 68, 65, 43, 7, 31, 69, 
		116, 121, 107, 47, 103, 43, 33, 96, 75, 75, 43, 0, 17, 63, 75, 
		86, 116, 105, 52, 137, 102, 110, 129, 85, 19, 0, 9, 32, 44, 38, 
		78, 85, 101, 149, 201, 44, 31, 28, 23, 18, 21, 22, 22, 33, 31, 
		38, 57, 52, 199, 75, 24, 30, 20, 16, 14, 17, 28, 45, 34, 28, 
		34, 24, 64, 147, 34, 26, 26, 25, 21, 25, 29, 34, 22, 27, 69, 
		43, 23, 31, 48, 20, 18, 30, 24, 27, 30, 35, 16, 22, 69, 37, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		
		50, 42, 46, 51, 52, 41, 54, 54, 54, 57, 45, 35, 36, 47, 48, 
		48, 47, 51, 55, 48, 11, 76, 53, 49, 0, 20, 28, 20, 29, 47, 
		56, 22, 49, 50, 53, 42, 24, 23, 11, 0, 25, 10, 39, 28, 18, 
		66, 0, 60, 46, 51, 17, 33, 33, 15, 0, 19, 20, 7, 20, 5, 
		40, 19, 76, 27, 36, 56, 34, 19, 17, 0, 21, 45, 8, 26, 24, 
		34, 0, 62, 31, 0, 0, 8, 33, 35, 0, 46, 25, 9, 20, 19, 
		19, 19, 26, 59, 0, 0, 35, 19, 44, 0, 32, 21, 1, 0, 31, 
		9, 4, 48, 51, 25, 12, 44, 8, 12, 0, 5, 22, 0, 17, 14, 
		8, 0, 34, 0, 39, 0, 3, 9, 0, 43, 4, 21, 0, 0, 40, 
		0, 0, 31, 0, 49, 19, 0, 24, 37, 23, 30, 6, 0, 30, 53, 
		0, 1, 31, 0, 32, 62, 14, 18, 34, 21, 0, 0, 4, 12, 21, 
		0, 0, 17, 0, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 29, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 10, 8, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 30, 11, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 2, 
		0, 0, 0, 13, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 10, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 1, 0, 0, 
		0, 0, 1, 0, 1, 14, 9, 10, 0, 11, 27, 11, 22, 0, 0, 
		0, 0, 0, 7, 0, 0, 0, 0, 1, 0, 0, 10, 0, 0, 0, 
		10, 0, 2, 0, 0, 0, 0, 0, 0, 15, 25, 0, 7, 23, 30, 
		41, 0, 0, 0, 19, 65, 70, 70, 40, 34, 27, 35, 35, 30, 34, 
		26, 39, 0, 5, 52, 26, 23, 28, 31, 30, 29, 29, 20, 28, 29, 
		33, 28, 32, 15, 27, 27, 26, 28, 25, 29, 38, 39, 38, 42, 33, 
		30, 32, 35, 60, 44, 42, 25, 17, 17, 28, 32, 33, 21, 26, 18, 
		
		others=>0 );
END gold_package;
