-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use IEEE.std_logic_arith.all;

-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity bram_single is
    generic (
        DEVICE     : string := "7SERIES";
        BRAM_NAME  : string := "default"
        );

    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic;
        DI   : in std_logic_vector(36-1 downto 0);
        ADDR : in std_logic_vector(9-1 downto 0);
        DO   : out std_logic_vector(36-1 downto 0)
    );
    attribute dont_touch : string;
    attribute dont_touch of bram_single : entity is "true";
   end bram_single;

  architecture a1 of bram_single is
    signal bram_wr_en    : std_logic_vector(8-1 downto 0);
    signal bram_addr     : std_logic_vector(9-1 downto 0);
    signal bram_di     : std_logic_vector(44-1 downto 0);
    signal bram_do     : std_logic_vector(44-1 downto 0);
    constant bram_par     : std_logic_vector(8-1 downto 0) := "00000000";

    begin
    bram_wr_en <= (others => '1') when WE = '1' else (others => '0');
    bram_addr <= ADDR(9-1 downto 0);
    bram_di <= bram_par & DI;
    DO <= bram_do(36-1 downto 0);


    MEM_IWGHT_LAYER0_INSTANCE0 : if BRAM_NAME = "iwght_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffff4d1ffffffffffffff0efffffffffffff684ffffffff00002b1d00000000",
            INIT_01 => X"0000047200000000fffff4ccffffffff000014280000000000000a8c00000000",
            INIT_02 => X"ffffac9cffffffff000023f300000000ffffde83ffffffff00000d3400000000",
            INIT_03 => X"fffff23cfffffffffffff67efffffffffffffe5affffffff000025ea00000000",
            INIT_04 => X"0000004700000000ffffffcfffffffff00000036000000000000003800000000",
            INIT_05 => X"0000009200000000000000150000000000000064000000000000007c00000000",
            INIT_06 => X"ffffff61ffffffffffffffb3ffffffff00000000000000000000007200000000",
            INIT_07 => X"ffffffb3ffffffffffffff28ffffffffffffff50ffffffffffffffa6ffffffff",
            INIT_08 => X"0000006e000000000000006700000000ffffff57ffffffffffffff9fffffffff",
            INIT_09 => X"ffffffe0ffffffffffffffecffffffffffffffecffffffff0000005800000000",
            INIT_0A => X"ffffffc4ffffffff0000003a00000000ffffffffffffffff0000003500000000",
            INIT_0B => X"ffffffd2ffffffff00000012000000000000005d000000000000002b00000000",
            INIT_0C => X"ffffffc7fffffffffffffff7ffffffff00000035000000000000000f00000000",
            INIT_0D => X"0000001d000000000000002e000000000000007c000000000000001b00000000",
            INIT_0E => X"ffffffc5ffffffffffffffcfffffffffffffffb8ffffffffffffffd4ffffffff",
            INIT_0F => X"000000ba00000000000000a7000000000000005b00000000ffffffaaffffffff",
            INIT_10 => X"ffffff5effffffffffffffd3ffffffff00000000000000000000002300000000",
            INIT_11 => X"ffffffe8fffffffffffffff8ffffffffffffff84ffffffffffffff63ffffffff",
            INIT_12 => X"0000008f00000000ffffffdcffffffff0000003c000000000000002000000000",
            INIT_13 => X"ffffffcaffffffff0000002c0000000000000017000000000000000500000000",
            INIT_14 => X"ffffff81ffffffffffffffddffffffff0000006500000000ffffffabffffffff",
            INIT_15 => X"0000007d00000000ffffff75ffffffffffffff87ffffffff0000006700000000",
            INIT_16 => X"ffffffc2ffffffff0000007f00000000ffffffd8fffffffffffffffcffffffff",
            INIT_17 => X"ffffff99ffffffffffffff8dffffffff0000007500000000ffffffcaffffffff",
            INIT_18 => X"0000001c000000000000008e0000000000000077000000000000005900000000",
            INIT_19 => X"0000000800000000ffffffafffffffffffffff28ffffffffffffffa4ffffffff",
            INIT_1A => X"0000006b00000000000000410000000000000051000000000000001d00000000",
            INIT_1B => X"ffffffbbffffffffffffff1affffffffffffff63ffffffff0000004900000000",
            INIT_1C => X"00000019000000000000004e000000000000003b000000000000003f00000000",
            INIT_1D => X"ffffff44ffffffffffffffa7ffffffff0000000d000000000000008f00000000",
            INIT_1E => X"0000003d0000000000000050000000000000004a00000000ffffff86ffffffff",
            INIT_1F => X"000000e80000000000000015000000000000005a00000000ffffffc7ffffffff",
            INIT_20 => X"ffffff28ffffffff0000001c00000000ffffff65ffffffff0000005b00000000",
            INIT_21 => X"ffffffe9ffffffff0000004500000000ffffffc0ffffffffffffffa4ffffffff",
            INIT_22 => X"0000002100000000ffffffa7ffffffff00000084000000000000009b00000000",
            INIT_23 => X"0000005a00000000ffffff9cffffffffffffffa9ffffffffffffff7cffffffff",
            INIT_24 => X"ffffffd2ffffffff000000830000000000000034000000000000001800000000",
            INIT_25 => X"0000002f00000000ffffffc7ffffffffffffff4bffffffff0000004000000000",
            INIT_26 => X"0000002b0000000000000075000000000000000800000000ffffffb9ffffffff",
            INIT_27 => X"ffffffabffffffff00000078000000000000000d00000000ffffffbcffffffff",
            INIT_28 => X"0000004f00000000ffffffe5fffffffffffffff4ffffffff0000003f00000000",
            INIT_29 => X"0000006a000000000000000e00000000ffffff99ffffffff0000000300000000",
            INIT_2A => X"ffffff8cffffffffffffffabffffffff0000002200000000ffffffbfffffffff",
            INIT_2B => X"ffffffebffffffffffffff87ffffffff0000001a000000000000003500000000",
            INIT_2C => X"fffffff9ffffffff0000006d00000000ffffff8bffffffff0000006c00000000",
            INIT_2D => X"000000a40000000000000089000000000000003800000000ffffffe5ffffffff",
            INIT_2E => X"0000000900000000ffffffcdffffffffffffff34ffffffffffffff59ffffffff",
            INIT_2F => X"0000006600000000ffffffecffffffffffffffe5fffffffffffffffeffffffff",
            INIT_30 => X"0000000100000000ffffff59ffffffffffffff94ffffffff0000008000000000",
            INIT_31 => X"0000008d00000000ffffff7effffffffffffffd8ffffffff0000001400000000",
            INIT_32 => X"ffffff7bffffffffffffffbbffffffff0000006a00000000000000a200000000",
            INIT_33 => X"ffffffe2ffffffffffffffaeffffffffffffffcaffffffffffffffdfffffffff",
            INIT_34 => X"ffffffe0ffffffffffffff8fffffffffffffffceffffffffffffffc0ffffffff",
            INIT_35 => X"fffffff5ffffffff0000000400000000ffffffb0ffffffff0000000f00000000",
            INIT_36 => X"ffffffc2ffffffff0000000a000000000000002a000000000000000400000000",
            INIT_37 => X"0000003300000000ffffffdfffffffff0000000b000000000000001e00000000",
            INIT_38 => X"0000008b00000000000000300000000000000012000000000000004c00000000",
            INIT_39 => X"00000033000000000000009e000000000000001200000000fffffff9ffffffff",
            INIT_3A => X"00000069000000000000006500000000ffffffeafffffffffffffff1ffffffff",
            INIT_3B => X"0000007100000000000000460000000000000015000000000000005b00000000",
            INIT_3C => X"fffffffffffffffffffffff7ffffffffffffffb4ffffffff0000006300000000",
            INIT_3D => X"0000000a00000000ffffffbcfffffffffffffffeffffffffffffffebffffffff",
            INIT_3E => X"0000002e00000000ffffffc2ffffffffffffffdbffffffff0000002200000000",
            INIT_3F => X"ffffffabfffffffffffffff5ffffffffffffffc3ffffffff0000000300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008900000000ffffffc8ffffffffffffffbeffffffffffffffa3ffffffff",
            INIT_41 => X"000000a300000000000000400000000000000074000000000000007600000000",
            INIT_42 => X"ffffff9cffffffff00000008000000000000001f000000000000004400000000",
            INIT_43 => X"ffffffa3fffffffffffffff7ffffffff0000001b000000000000001a00000000",
            INIT_44 => X"ffffff75ffffffffffffffb2ffffffff0000002000000000fffffff2ffffffff",
            INIT_45 => X"0000002a00000000fffffff8ffffffffffffffd0ffffffffffffffbbffffffff",
            INIT_46 => X"ffffff3fffffffffffffffa1ffffffffffffffedffffffffffffff8dffffffff",
            INIT_47 => X"0000001000000000ffffffbdffffffffffffffedffffffffffffff87ffffffff",
            INIT_48 => X"ffffff9afffffffffffffff6ffffffffffffff71ffffffffffffffbfffffffff",
            INIT_49 => X"0000006300000000ffffffd5ffffffffffffffccffffffffffffff99ffffffff",
            INIT_4A => X"000000ea0000000000000028000000000000002500000000000000a300000000",
            INIT_4B => X"0000004a00000000000000e80000000000000080000000000000000000000000",
            INIT_4C => X"ffffff83ffffffffffffffe4ffffffffffffffe4ffffffffffffff93ffffffff",
            INIT_4D => X"ffffffd7ffffffffffffffdaffffffffffffffb2ffffffff0000003d00000000",
            INIT_4E => X"000000260000000000000020000000000000001700000000ffffff89ffffffff",
            INIT_4F => X"0000000c000000000000003a000000000000004800000000ffffffc2ffffffff",
            INIT_50 => X"0000000d00000000ffffffe2ffffffffffffffe7ffffffff0000000e00000000",
            INIT_51 => X"fffffff9ffffffff0000004c000000000000000b000000000000001e00000000",
            INIT_52 => X"ffffffecffffffffffffffd8ffffffff00000019000000000000002500000000",
            INIT_53 => X"000000160000000000000025000000000000000c000000000000003100000000",
            INIT_54 => X"ffffffcdffffffff0000004200000000fffffffdffffffffffffffd9ffffffff",
            INIT_55 => X"ffffff91ffffffff0000003600000000ffffffdbffffffffffffffc7ffffffff",
            INIT_56 => X"0000009d0000000000000000000000000000000b000000000000004d00000000",
            INIT_57 => X"fffffff8ffffffffffffff94ffffffffffffffb2ffffffffffffffd3ffffffff",
            INIT_58 => X"fffffff3ffffffff00000078000000000000003900000000ffffffa1ffffffff",
            INIT_59 => X"ffffff7bffffffffffffff98ffffffffffffffbaffffffff0000005e00000000",
            INIT_5A => X"00000040000000000000005000000000ffffff42ffffffff0000002900000000",
            INIT_5B => X"00000005000000000000000a000000000000008f00000000ffffffecffffffff",
            INIT_5C => X"0000006e00000000ffffff4fffffffffffffff97ffffffff0000009400000000",
            INIT_5D => X"0000004d00000000ffffffb7ffffffffffffffe2ffffffff0000000f00000000",
            INIT_5E => X"ffffff0afffffffffffffff0ffffffff000000ca00000000fffffffbffffffff",
            INIT_5F => X"ffffffc4ffffffffffffff9cffffffff00000065000000000000007a00000000",
            INIT_60 => X"ffffffb4ffffffff000000c6000000000000001700000000ffffffefffffffff",
            INIT_61 => X"ffffffc7ffffffff00000040000000000000007f00000000ffffff5bffffffff",
            INIT_62 => X"0000001f00000000ffffffdaffffffff0000000000000000ffffff8effffffff",
            INIT_63 => X"fffffff6ffffffffffffffe5ffffffffffffffceffffffff0000000900000000",
            INIT_64 => X"000000180000000000000000000000000000002800000000fffffff5ffffffff",
            INIT_65 => X"ffffffe6ffffffffffffffe6ffffffffffffffd5ffffffffffffffefffffffff",
            INIT_66 => X"ffffffe1fffffffffffffff9ffffffffffffffdcfffffffffffffff1ffffffff",
            INIT_67 => X"00000018000000000000001b00000000ffffffdcffffffffffffffc5ffffffff",
            INIT_68 => X"ffffffceffffffff0000000900000000ffffffccffffffff0000002300000000",
            INIT_69 => X"ffffffc3ffffffffffffffbdffffffff0000003d00000000ffffffe4ffffffff",
            INIT_6A => X"ffffffdfffffffff00000051000000000000000000000000fffffff3ffffffff",
            INIT_6B => X"0000004e000000000000003b0000000000000051000000000000001000000000",
            INIT_6C => X"0000006900000000000000730000000000000024000000000000001900000000",
            INIT_6D => X"000000140000000000000006000000000000002b000000000000003200000000",
            INIT_6E => X"ffffff6affffffffffffff5affffffffffffffb4ffffffffffffffaeffffffff",
            INIT_6F => X"ffffffc5ffffffffffffff98ffffffffffffffedffffffff0000000a00000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER0_INSTANCE0;


    MEM_IWGHT_LAYER1_INSTANCE0 : if BRAM_NAME = "iwght_layer1_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000654b0000000000008bcd000000000000272900000000000003c600000000",
            INIT_01 => X"000000d900000000ffffe86afffffffffffff5cbffffffff0000046500000000",
            INIT_02 => X"0000333400000000000039d5000000000000283200000000ffff825dffffffff",
            INIT_03 => X"000081c200000000ffffd791fffffffffffff1ceffffffff0000132300000000",
            INIT_04 => X"ffffe18cffffffffffff340effffffff00006c670000000000001b2600000000",
            INIT_05 => X"000035a1000000000000525d00000000ffffe671ffffffff0000416b00000000",
            INIT_06 => X"fffff3e5ffffffffffffb86bffffffffffff795cffffffff0000aa3200000000",
            INIT_07 => X"00002c5500000000ffff5d14ffffffffffffc93dffffffff0000383600000000",
            INIT_08 => X"ffffffc4fffffffffffffff0ffffffff0000001700000000fffffffdffffffff",
            INIT_09 => X"00000004000000000000000200000000ffffffd6ffffffff0000005b00000000",
            INIT_0A => X"ffffffbeffffffff0000007700000000ffffffb8ffffffff0000001e00000000",
            INIT_0B => X"0000002500000000ffffff26ffffffff00000061000000000000003000000000",
            INIT_0C => X"ffffff79ffffffff00000071000000000000000600000000ffffff2dffffffff",
            INIT_0D => X"0000002a000000000000004b00000000ffffff9affffffff0000003000000000",
            INIT_0E => X"fffffff9ffffffffffffffb5ffffffff0000004800000000ffffffedffffffff",
            INIT_0F => X"00000056000000000000006000000000ffffffddffffffffffffffe0ffffffff",
            INIT_10 => X"fffffff5fffffffffffffff7ffffffff0000001b00000000ffffff54ffffffff",
            INIT_11 => X"000000a200000000ffffff22ffffffff0000003b00000000fffffff1ffffffff",
            INIT_12 => X"ffffffddffffffff0000005200000000ffffff94ffffffff0000009700000000",
            INIT_13 => X"ffffff94ffffffff0000003200000000ffffffbaffffffff0000007a00000000",
            INIT_14 => X"0000001a000000000000000d00000000ffffffa8ffffffff0000002000000000",
            INIT_15 => X"0000006700000000ffffffe7ffffffff0000001c00000000ffffffc3ffffffff",
            INIT_16 => X"ffffff9effffffffffffffebffffffff0000002300000000ffffffdfffffffff",
            INIT_17 => X"0000006b000000000000004e00000000ffffff40ffffffff0000000f00000000",
            INIT_18 => X"ffffff74ffffffff0000002c00000000ffffffacffffffffffffffccffffffff",
            INIT_19 => X"0000007700000000ffffffb5ffffffff00000000000000000000002500000000",
            INIT_1A => X"00000058000000000000001200000000ffffff7fffffffff0000005f00000000",
            INIT_1B => X"0000002b00000000ffffff43ffffffff0000006600000000ffffff46ffffffff",
            INIT_1C => X"ffffffdaffffffff0000004c00000000fffffffaffffffff0000007600000000",
            INIT_1D => X"0000002900000000ffffffd8ffffffffffffffc0ffffffff0000005e00000000",
            INIT_1E => X"ffffffa9ffffffff0000000e000000000000006800000000ffffff63ffffffff",
            INIT_1F => X"000000ac00000000fffffeb3fffffffffffffff9ffffffff0000003800000000",
            INIT_20 => X"000000690000000000000079000000000000008500000000ffffff74ffffffff",
            INIT_21 => X"fffffef8ffffffff0000008100000000ffffffb9ffffffffffffffb9ffffffff",
            INIT_22 => X"00000015000000000000004200000000ffffff97ffffffff000000a100000000",
            INIT_23 => X"ffffffc6ffffffff0000005500000000fffffec3ffffffff0000007f00000000",
            INIT_24 => X"ffffffe9ffffffff000000200000000000000063000000000000001d00000000",
            INIT_25 => X"0000001800000000ffffffd0fffffffffffffffaffffffff0000000d00000000",
            INIT_26 => X"fffffff9ffffffff0000002700000000ffffff94ffffffffffffffeeffffffff",
            INIT_27 => X"0000000800000000fffffffdffffffffffffffc6ffffffff0000001f00000000",
            INIT_28 => X"ffffffe9fffffffffffffff6ffffffff00000008000000000000001900000000",
            INIT_29 => X"0000006500000000ffffffeaffffffff0000000800000000ffffffe6ffffffff",
            INIT_2A => X"ffffffd0ffffffffffffff95ffffffffffffffb8ffffffff0000000800000000",
            INIT_2B => X"0000001f000000000000009400000000ffffff96ffffffff0000005400000000",
            INIT_2C => X"00000014000000000000008200000000000000d6000000000000007b00000000",
            INIT_2D => X"ffffff5cffffffffffffff84ffffffffffffff8affffffff0000002e00000000",
            INIT_2E => X"ffffffc8ffffffffffffffa2ffffffff0000000400000000ffffff55ffffffff",
            INIT_2F => X"ffffffcdffffffffffffffdfffffffff0000005300000000ffffffd6ffffffff",
            INIT_30 => X"000000d600000000000000e20000000000000042000000000000011400000000",
            INIT_31 => X"0000007500000000ffffffdfffffffff0000001400000000ffffffa2ffffffff",
            INIT_32 => X"ffffffceffffffffffffff67ffffffffffffff1dffffffffffffff44ffffffff",
            INIT_33 => X"000000890000000000000138000000000000001800000000ffffffccffffffff",
            INIT_34 => X"0000001800000000000000910000000000000034000000000000000e00000000",
            INIT_35 => X"0000002600000000000000b30000000000000076000000000000002600000000",
            INIT_36 => X"ffffff5fffffffffffffffa7ffffffff00000065000000000000004500000000",
            INIT_37 => X"0000002200000000fffffff2ffffffff00000024000000000000006400000000",
            INIT_38 => X"ffffff8dffffffff000000070000000000000067000000000000006000000000",
            INIT_39 => X"ffffffcafffffffffffffffaffffffffffffffb3ffffffff000000a900000000",
            INIT_3A => X"ffffff63ffffffff00000087000000000000007200000000fffffff6ffffffff",
            INIT_3B => X"ffffffe5ffffffff0000000e000000000000003600000000ffffffabffffffff",
            INIT_3C => X"ffffffefffffffff000000d6000000000000000300000000ffffffb7ffffffff",
            INIT_3D => X"00000005000000000000003f000000000000004200000000ffffff64ffffffff",
            INIT_3E => X"ffffffb2ffffffffffffffd3ffffffffffffffe7ffffffff0000004000000000",
            INIT_3F => X"fffffff8ffffffffffffffceffffffffffffffc3ffffffffffffff8affffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009800000000000000530000000000000051000000000000005200000000",
            INIT_41 => X"fffffea0ffffffffffffff7bfffffffffffffff0ffffffffffffffc8ffffffff",
            INIT_42 => X"000000ad000000000000002e00000000fffffe88fffffffffffffeedffffffff",
            INIT_43 => X"00000000000000000000000900000000ffffff92ffffffff0000002600000000",
            INIT_44 => X"0000000600000000fffffffdffffffffffffff5bffffffff0000003200000000",
            INIT_45 => X"ffffff94ffffffffffffffaeffffffffffffff68ffffffffffffff80ffffffff",
            INIT_46 => X"ffffffb1fffffffffffffff3ffffffffffffffd8fffffffffffffec5ffffffff",
            INIT_47 => X"fffffffcffffffff0000005300000000ffffffc8ffffffffffffffbdffffffff",
            INIT_48 => X"00000093000000000000001d0000000000000001000000000000007000000000",
            INIT_49 => X"ffffffafffffffff0000001100000000ffffffe3ffffffffffffffc7ffffffff",
            INIT_4A => X"0000002100000000ffffffeaffffffff0000002800000000000000ae00000000",
            INIT_4B => X"fffffffaffffffffffffffe3ffffffffffffff30fffffffffffffff4ffffffff",
            INIT_4C => X"000000070000000000000003000000000000001d00000000ffffffe9ffffffff",
            INIT_4D => X"ffffffe4ffffffff00000007000000000000000000000000fffffffaffffffff",
            INIT_4E => X"0000002a00000000ffffff69ffffffffffffffb1ffffffff000000b100000000",
            INIT_4F => X"fffffff0ffffffffffffff96ffffffff0000006000000000ffffff39ffffffff",
            INIT_50 => X"ffffffc0ffffffffffffff62ffffffff00000000000000000000005f00000000",
            INIT_51 => X"fffffee3ffffffff0000003f00000000ffffffc1ffffffffffffffd4ffffffff",
            INIT_52 => X"000000330000000000000043000000000000005300000000ffffff66ffffffff",
            INIT_53 => X"0000008f000000000000006600000000fffffff7ffffffff0000008d00000000",
            INIT_54 => X"fffffee5ffffffff0000003f000000000000004e00000000ffffffb4ffffffff",
            INIT_55 => X"ffffffbbffffffffffffffaeffffffff0000001900000000ffffff22ffffffff",
            INIT_56 => X"0000002900000000ffffffbeffffffffffffff8ffffffffffffffffdffffffff",
            INIT_57 => X"0000002e00000000ffffffccffffffff0000000300000000fffffff2ffffffff",
            INIT_58 => X"0000004a000000000000001200000000ffffffa1ffffffff000000bd00000000",
            INIT_59 => X"0000003500000000ffffff9fffffffffffffffb3ffffffff0000001b00000000",
            INIT_5A => X"ffffffd4ffffffff0000008900000000ffffff6dffffffff0000006000000000",
            INIT_5B => X"ffffff71ffffffffffffff9bffffffffffffff9cffffffff0000001d00000000",
            INIT_5C => X"0000002000000000ffffffe5ffffffffffffffacfffffffffffffeffffffffff",
            INIT_5D => X"000000f8000000000000004b00000000ffffffc1ffffffffffffff85ffffffff",
            INIT_5E => X"0000006f0000000000000021000000000000002500000000ffffffa3ffffffff",
            INIT_5F => X"ffffffb9ffffffff0000005d00000000ffffff81ffffffff0000004e00000000",
            INIT_60 => X"ffffffc1ffffffff000000850000000000000033000000000000001800000000",
            INIT_61 => X"ffffffb4ffffffffffffffa8ffffffff0000000d000000000000007b00000000",
            INIT_62 => X"0000000000000000ffffff12ffffffff0000008e00000000ffffff6effffffff",
            INIT_63 => X"fffffec8ffffffff000000290000000000000007000000000000004300000000",
            INIT_64 => X"fffffedfffffffffffffffe3ffffffff0000000a00000000fffffe4cffffffff",
            INIT_65 => X"ffffffc2ffffffff000000bb00000000ffffff57ffffffffffffff7affffffff",
            INIT_66 => X"00000047000000000000006b000000000000004500000000ffffff37ffffffff",
            INIT_67 => X"0000004e00000000ffffff5effffffffffffffcdffffffff0000000900000000",
            INIT_68 => X"ffffffc6ffffffff000000570000000000000095000000000000007400000000",
            INIT_69 => X"00000046000000000000005100000000ffffffc6ffffffff0000000300000000",
            INIT_6A => X"ffffffd6ffffffffffffffb2ffffffffffffffafffffffff0000001000000000",
            INIT_6B => X"ffffff72ffffffffffffffefffffffff0000004600000000ffffffe1ffffffff",
            INIT_6C => X"0000003d00000000ffffffe9ffffffff0000002e00000000ffffffe4ffffffff",
            INIT_6D => X"fffffff5fffffffffffffffbffffffffffffffc6ffffffffffffffa1ffffffff",
            INIT_6E => X"0000002300000000fffffff1ffffffffffffffe3ffffffff0000001900000000",
            INIT_6F => X"ffffffedfffffffffffffff8ffffffff0000001f000000000000008100000000",
            INIT_70 => X"ffffffefffffffffffffffe7ffffffff00000019000000000000000000000000",
            INIT_71 => X"ffffff79fffffffffffffff1ffffffff0000001800000000fffffff2ffffffff",
            INIT_72 => X"fffffff8ffffffffffffffcdffffffffffffffa5ffffffff0000008400000000",
            INIT_73 => X"fffffec5ffffffffffffffd8fffffffffffffff5ffffffff0000005900000000",
            INIT_74 => X"0000003100000000ffffffd6ffffffff0000005e00000000ffffff97ffffffff",
            INIT_75 => X"ffffff9affffffffffffffa4ffffffff00000055000000000000008d00000000",
            INIT_76 => X"ffffffa1ffffffffffffff55ffffffffffffffb4ffffffff0000004d00000000",
            INIT_77 => X"00000011000000000000004900000000fffffe6cfffffffffffffec0ffffffff",
            INIT_78 => X"0000003700000000ffffffacffffffffffffffe6ffffffffffffffe4ffffffff",
            INIT_79 => X"ffffffbbffffffff0000000e00000000fffffff9ffffffff0000001200000000",
            INIT_7A => X"ffffff9bffffffff000000d800000000ffffffc2ffffffff0000006d00000000",
            INIT_7B => X"fffffe79ffffffffffffff7afffffffffffffea2ffffffffffffff1affffffff",
            INIT_7C => X"ffffff9bffffffffffffff4efffffffffffffef8ffffffffffffff9effffffff",
            INIT_7D => X"fffffe1dffffffffffffffd9fffffffffffffc8afffffffffffffda4ffffffff",
            INIT_7E => X"ffffff55fffffffffffffe3affffffffffffffb0fffffffffffffee6ffffffff",
            INIT_7F => X"ffffffe6ffffffff0000000b0000000000000057000000000000009200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE0;


    MEM_IWGHT_LAYER1_INSTANCE1 : if BRAM_NAME = "iwght_layer1_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffff91ffffffffffffffefffffffffffffffd8ffffffffffffff72ffffffff",
            INIT_01 => X"fffffdf6fffffffffffffefeffffffff0000002800000000ffffffddffffffff",
            INIT_02 => X"fffffed4ffffffffffffff9bffffffffffffffd5ffffffff0000003f00000000",
            INIT_03 => X"ffffffb2ffffffff000000370000000000000000000000000000006900000000",
            INIT_04 => X"ffffffd5ffffffffffffffe8ffffffff0000005100000000ffffffd1ffffffff",
            INIT_05 => X"fffffffeffffffff0000002700000000000000a700000000ffffffb9ffffffff",
            INIT_06 => X"0000000300000000000000630000000000000012000000000000006200000000",
            INIT_07 => X"0000004f00000000ffffffc4ffffffff0000005200000000fffffff9ffffffff",
            INIT_08 => X"ffffff09ffffffff000000bb0000000000000038000000000000001e00000000",
            INIT_09 => X"ffffffa2ffffffff0000000500000000ffffffacffffffff0000003c00000000",
            INIT_0A => X"ffffffcaffffffff0000003200000000000000f600000000ffffff5effffffff",
            INIT_0B => X"fffffff0ffffffff0000001f000000000000001c00000000ffffffb3ffffffff",
            INIT_0C => X"0000003900000000ffffffc3ffffffff0000002500000000fffffff9ffffffff",
            INIT_0D => X"fffffffdffffffffffffffe5ffffffff00000080000000000000003000000000",
            INIT_0E => X"ffffffffffffffffffffffbfffffffffffffffedffffffff0000001400000000",
            INIT_0F => X"0000009600000000ffffff8bffffffff00000001000000000000011c00000000",
            INIT_10 => X"ffffffaeffffffffffffffd7ffffffff0000000500000000ffffffd0ffffffff",
            INIT_11 => X"ffffffd2ffffffffffffff70ffffffffffffffaeffffffffffffff12ffffffff",
            INIT_12 => X"ffffffc9fffffffffffffe57ffffffffffffffc0ffffffffffffffb3ffffffff",
            INIT_13 => X"fffffffdfffffffffffffff2ffffffffffffff56ffffffff0000003200000000",
            INIT_14 => X"ffffffe8ffffffffffffffe7ffffffff0000001600000000fffffff0ffffffff",
            INIT_15 => X"fffffffbffffffff0000000700000000fffffff0ffffffff0000001300000000",
            INIT_16 => X"ffffffe4ffffffffffffffcbfffffffffffffff0ffffffff0000003700000000",
            INIT_17 => X"ffffffeaffffffff0000002600000000ffffffb0ffffffff0000002500000000",
            INIT_18 => X"0000003700000000ffffffbbffffffffffffffa2ffffffff0000004900000000",
            INIT_19 => X"ffffffe5ffffffffffffffadffffffffffffffc9ffffffff0000006200000000",
            INIT_1A => X"0000007300000000ffffffeaffffffffffffffbdffffffff000000ab00000000",
            INIT_1B => X"ffffffa9ffffffff0000006800000000ffffffaaffffffffffffff87ffffffff",
            INIT_1C => X"0000009500000000fffffed2ffffffff0000000400000000ffffff84ffffffff",
            INIT_1D => X"0000003500000000fffffd89ffffffff0000002d000000000000004600000000",
            INIT_1E => X"ffffffa5fffffffffffffff8ffffffffffffff62ffffffff0000005400000000",
            INIT_1F => X"ffffff52ffffffffffffff4dffffffffffffffd4ffffffff0000004c00000000",
            INIT_20 => X"0000000300000000ffffff3cffffffffffffff9fffffffff0000005b00000000",
            INIT_21 => X"ffffff9cffffffffffffffe6ffffffff0000004b00000000ffffffdcffffffff",
            INIT_22 => X"0000001000000000ffffffe4ffffffffffffff8dffffffff0000007400000000",
            INIT_23 => X"ffffff58ffffffff00000065000000000000008b000000000000008f00000000",
            INIT_24 => X"0000000b00000000ffffff86ffffffff0000008c000000000000003d00000000",
            INIT_25 => X"0000001900000000ffffff63ffffffffffffffbdffffffff0000005100000000",
            INIT_26 => X"ffffffb1ffffffffffffff79ffffffff00000003000000000000001300000000",
            INIT_27 => X"0000006300000000ffffffddffffffffffffffd7ffffffffffffff87ffffffff",
            INIT_28 => X"0000004c00000000fffffffdfffffffffffffff8ffffffffffffff74ffffffff",
            INIT_29 => X"ffffffa5ffffffff0000001d000000000000005c00000000ffffff37ffffffff",
            INIT_2A => X"0000005d000000000000005e000000000000002b000000000000002b00000000",
            INIT_2B => X"ffffff53ffffffff00000047000000000000000000000000ffffff27ffffffff",
            INIT_2C => X"0000001c00000000ffffffb3ffffffffffffffc4ffffffffffffffecffffffff",
            INIT_2D => X"00000029000000000000005e000000000000005100000000ffffffc3ffffffff",
            INIT_2E => X"ffffffebffffffffffffffc5ffffffff00000018000000000000002f00000000",
            INIT_2F => X"ffffff8fffffffffffffff44ffffffffffffffa6ffffffff0000000b00000000",
            INIT_30 => X"0000002800000000ffffffa1ffffffff0000004a000000000000007900000000",
            INIT_31 => X"ffffffe4ffffffff000000b500000000ffffffbeffffffffffffffb1ffffffff",
            INIT_32 => X"fffffffcffffffff00000010000000000000001900000000ffffffb7ffffffff",
            INIT_33 => X"ffffffe1ffffffffffffff7effffffffffffffbeffffffff0000000600000000",
            INIT_34 => X"ffffffdeffffffffffffff78ffffffff0000004e00000000ffffff78ffffffff",
            INIT_35 => X"0000002300000000fffffff2ffffffff0000006100000000000000cb00000000",
            INIT_36 => X"fffffff4ffffffff00000094000000000000002900000000ffffffacffffffff",
            INIT_37 => X"0000000f00000000fffffff3ffffffff0000002400000000ffffffebffffffff",
            INIT_38 => X"0000000900000000fffffffffffffffffffffff0ffffffff0000000a00000000",
            INIT_39 => X"00000060000000000000001c0000000000000002000000000000001e00000000",
            INIT_3A => X"0000002400000000ffffffa6ffffffff0000004c00000000ffffffc7ffffffff",
            INIT_3B => X"0000002400000000fffffffdffffffffffffffcaffffffffffffffb0ffffffff",
            INIT_3C => X"0000003b000000000000001600000000ffffff74ffffffffffffffe6ffffffff",
            INIT_3D => X"ffffffb1ffffffff00000036000000000000000f00000000fffffff2ffffffff",
            INIT_3E => X"00000106000000000000001000000000ffffff69ffffffffffffffd1ffffffff",
            INIT_3F => X"000000a900000000fffffffeffffffffffffffceffffffff0000005a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000007000000000000000800000000ffffff95ffffffff0000006600000000",
            INIT_41 => X"ffffffe9ffffffffffffff62ffffffffffffffc4ffffffffffffffdbffffffff",
            INIT_42 => X"0000007d000000000000007a000000000000001b00000000ffffff7effffffff",
            INIT_43 => X"00000070000000000000003e00000000ffffffdfffffffff0000007f00000000",
            INIT_44 => X"fffffff9ffffffff000000730000000000000002000000000000006000000000",
            INIT_45 => X"0000000000000000ffffffd5ffffffff00000022000000000000008700000000",
            INIT_46 => X"0000001f000000000000001f000000000000009700000000000000ca00000000",
            INIT_47 => X"0000003e00000000ffffffa8ffffffffffffff88ffffffff0000001a00000000",
            INIT_48 => X"0000004500000000ffffffd0ffffffff0000007c00000000ffffffc0ffffffff",
            INIT_49 => X"00000074000000000000001c00000000ffffffecfffffffffffffff7ffffffff",
            INIT_4A => X"0000002400000000ffffffb8ffffffff0000003900000000ffffffe4ffffffff",
            INIT_4B => X"0000000600000000ffffffaaffffffffffffffa8ffffffff0000008e00000000",
            INIT_4C => X"ffffffebffffffff0000003900000000ffffffc4ffffffff0000009a00000000",
            INIT_4D => X"ffffffadffffffffffffffb8ffffffffffffffffffffffffffffffedffffffff",
            INIT_4E => X"ffffffc1ffffffffffffffe3ffffffffffffffcaffffffffffffffccffffffff",
            INIT_4F => X"ffffff97ffffffff000000740000000000000014000000000000009b00000000",
            INIT_50 => X"0000005a00000000ffffffe5ffffffff00000019000000000000002a00000000",
            INIT_51 => X"000000af0000000000000014000000000000008100000000ffffffd8ffffffff",
            INIT_52 => X"000000f2000000000000004c00000000ffffff41fffffffffffffff0ffffffff",
            INIT_53 => X"ffffff63ffffffffffffff50ffffffff00000001000000000000002800000000",
            INIT_54 => X"ffffffe5fffffffffffffffeffffffff0000000000000000ffffffc4ffffffff",
            INIT_55 => X"fffffffbffffffff00000032000000000000003e000000000000005700000000",
            INIT_56 => X"ffffffe4ffffffffffffff34ffffffffffffffe6ffffffffffffffb6ffffffff",
            INIT_57 => X"00000015000000000000007700000000ffffffd2ffffffffffffffc2ffffffff",
            INIT_58 => X"0000008500000000ffffffc9ffffffffffffffcaffffffff0000008600000000",
            INIT_59 => X"ffffffcfffffffff00000000000000000000001300000000fffffff1ffffffff",
            INIT_5A => X"fffffff8ffffffffffffff86ffffffff0000002000000000ffffffdbffffffff",
            INIT_5B => X"00000018000000000000000c000000000000000700000000ffffffa5ffffffff",
            INIT_5C => X"0000000b000000000000001800000000fffffffefffffffffffffffeffffffff",
            INIT_5D => X"fffffffbffffffffffffffe9fffffffffffffffbfffffffffffffffbffffffff",
            INIT_5E => X"0000004200000000ffffff7dffffffff00000002000000000000000000000000",
            INIT_5F => X"00000007000000000000003d000000000000002400000000ffffffc5ffffffff",
            INIT_60 => X"ffffff94ffffffff00000044000000000000006d000000000000004700000000",
            INIT_61 => X"ffffffc6ffffffffffffffceffffffff00000037000000000000007200000000",
            INIT_62 => X"00000003000000000000001500000000ffffffa5ffffffffffffff78ffffffff",
            INIT_63 => X"ffffffb5ffffffffffffffcfffffffff0000004d000000000000002e00000000",
            INIT_64 => X"0000003d00000000fffffff8ffffffff00000034000000000000009800000000",
            INIT_65 => X"fffffff7ffffffff0000002200000000fffffff9ffffffff0000006900000000",
            INIT_66 => X"fffffff8ffffffffffffff60fffffffffffffef2fffffffffffffff7ffffffff",
            INIT_67 => X"0000002a000000000000005500000000ffffffc1fffffffffffffff7ffffffff",
            INIT_68 => X"00000087000000000000000d0000000000000064000000000000007300000000",
            INIT_69 => X"0000002b00000000ffffff8effffffffffffffe1fffffffffffffffbffffffff",
            INIT_6A => X"0000002f00000000fffffffbffffffff00000021000000000000000900000000",
            INIT_6B => X"000000400000000000000035000000000000006800000000ffffffefffffffff",
            INIT_6C => X"0000002800000000ffffff87ffffffffffffffc0ffffffff0000002e00000000",
            INIT_6D => X"ffffffeeffffffffffffffe3ffffffffffffffdcffffffffffffff87ffffffff",
            INIT_6E => X"0000007c000000000000004f000000000000004a00000000ffffffb7ffffffff",
            INIT_6F => X"0000002c0000000000000023000000000000003c000000000000004600000000",
            INIT_70 => X"ffffffecffffffffffffffa9ffffffff0000000900000000ffffff85ffffffff",
            INIT_71 => X"fffffff9ffffffff0000000a000000000000001a000000000000004e00000000",
            INIT_72 => X"ffffffd7ffffffff000000ac0000000000000022000000000000009c00000000",
            INIT_73 => X"ffffffa5ffffffffffffffb6ffffffffffffffc1ffffffffffffffc0ffffffff",
            INIT_74 => X"0000006500000000ffffffa6ffffffff0000009400000000ffffffb7ffffffff",
            INIT_75 => X"00000001000000000000003b00000000ffffffb7ffffffff0000007100000000",
            INIT_76 => X"ffffff55ffffffffffffffb6ffffffff0000002300000000ffffff6cffffffff",
            INIT_77 => X"ffffff9affffffff0000003200000000ffffffbfffffffff0000004d00000000",
            INIT_78 => X"00000047000000000000009b00000000ffffff6dffffffff0000002c00000000",
            INIT_79 => X"0000001b0000000000000028000000000000007700000000000000c900000000",
            INIT_7A => X"ffffff5fffffffffffffff54ffffffffffffff98ffffffffffffffdbffffffff",
            INIT_7B => X"fffffff2ffffffffffffffe0fffffffffffffffdffffffff0000002e00000000",
            INIT_7C => X"00000084000000000000002d000000000000001400000000ffffffcdffffffff",
            INIT_7D => X"ffffffd3ffffffffffffffc0ffffffffffffffedffffffffffffffb7ffffffff",
            INIT_7E => X"00000022000000000000002300000000ffffffc7ffffffffffffff76ffffffff",
            INIT_7F => X"0000000200000000000000030000000000000008000000000000005700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE1;


    MEM_IWGHT_LAYER1_INSTANCE2 : if BRAM_NAME = "iwght_layer1_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff4ffffffffffffffffffffffffffffffeeffffffff0000000100000000",
            INIT_01 => X"000000dd000000000000000500000000ffffffebffffffff0000001500000000",
            INIT_02 => X"ffffff90ffffffff000000190000000000000093000000000000005400000000",
            INIT_03 => X"ffffffa9ffffffffffffff07ffffffffffffff45ffffffffffffff85ffffffff",
            INIT_04 => X"ffffffe9ffffffffffffff8bffffffff0000004b00000000ffffffc4ffffffff",
            INIT_05 => X"00000035000000000000002100000000ffffff80ffffffffffffffb7ffffffff",
            INIT_06 => X"ffffffa4ffffffff0000002100000000ffffff96fffffffffffffff4ffffffff",
            INIT_07 => X"0000002f000000000000008700000000ffffffa4ffffffff000000b300000000",
            INIT_08 => X"0000002000000000ffffff8fffffffff0000006d000000000000006000000000",
            INIT_09 => X"0000002f00000000ffffffe5ffffffff00000016000000000000001200000000",
            INIT_0A => X"0000002a00000000ffffffa6ffffffffffffffc7ffffffffffffffe7ffffffff",
            INIT_0B => X"00000094000000000000002e0000000000000089000000000000002000000000",
            INIT_0C => X"0000000700000000ffffffc3ffffffff0000001e00000000ffffff97ffffffff",
            INIT_0D => X"ffffffc5ffffffff000000190000000000000090000000000000007c00000000",
            INIT_0E => X"000000310000000000000021000000000000001c000000000000003b00000000",
            INIT_0F => X"ffffff9effffffffffffffcfffffffffffffffbdffffffffffffffd1ffffffff",
            INIT_10 => X"ffffff72ffffffff0000000200000000ffffffe6ffffffffffffff9affffffff",
            INIT_11 => X"fffffff8ffffffff00000026000000000000004e00000000ffffffe3ffffffff",
            INIT_12 => X"ffffff77fffffffffffffffcfffffffffffffffaffffffff0000004d00000000",
            INIT_13 => X"00000012000000000000001300000000ffffffffffffffffffffffdeffffffff",
            INIT_14 => X"ffffff9bffffffffffffffdbffffffff0000002b00000000ffffffddffffffff",
            INIT_15 => X"0000003c000000000000002000000000fffffff6fffffffffffffff1ffffffff",
            INIT_16 => X"ffffffe4ffffffffffffffd2ffffffffffffff60ffffffffffffffefffffffff",
            INIT_17 => X"fffffff9fffffffffffffffcfffffffffffffffaffffffff0000007500000000",
            INIT_18 => X"ffffffdbfffffffffffffff8ffffffff000000a5000000000000006f00000000",
            INIT_19 => X"ffffff93ffffffffffffffedffffffffffffff81ffffffff0000006500000000",
            INIT_1A => X"ffffffe1fffffffffffffffcffffffffffffffccffffffff0000003f00000000",
            INIT_1B => X"0000006a000000000000000400000000ffffffc9ffffffffffffff7affffffff",
            INIT_1C => X"fffffedfffffffffffffffabffffffff0000002700000000ffffffb6ffffffff",
            INIT_1D => X"0000003600000000ffffff86ffffffffffffffaeffffffffffffff59ffffffff",
            INIT_1E => X"000000cf00000000000000eb0000000000000066000000000000001400000000",
            INIT_1F => X"00000062000000000000006b000000000000001f00000000ffffff4affffffff",
            INIT_20 => X"0000011100000000000000aa0000000000000033000000000000004200000000",
            INIT_21 => X"0000000700000000000000220000000000000002000000000000004300000000",
            INIT_22 => X"ffffff87ffffffffffffff8ffffffffffffffffdffffffffffffffd1ffffffff",
            INIT_23 => X"ffffffd9fffffffffffffffbffffffffffffff6fffffffffffffff33ffffffff",
            INIT_24 => X"0000000500000000fffffff7ffffffffffffffe2fffffffffffffffbffffffff",
            INIT_25 => X"ffffffc4ffffffff000000140000000000000005000000000000000a00000000",
            INIT_26 => X"0000001000000000ffffff9effffffffffffffdfffffffffffffffecffffffff",
            INIT_27 => X"0000005d00000000000000760000000000000006000000000000005700000000",
            INIT_28 => X"ffffffd6ffffffff0000011c00000000fffffff8ffffffffffffff7dffffffff",
            INIT_29 => X"0000001600000000fffffffaffffffff00000099000000000000002d00000000",
            INIT_2A => X"ffffff9bffffffff0000001500000000ffffffe4ffffffffffffffb2ffffffff",
            INIT_2B => X"ffffffc4ffffffffffffffeaffffffff00000014000000000000005200000000",
            INIT_2C => X"ffffffe6ffffffffffffff0fffffffff0000004d00000000ffffffaaffffffff",
            INIT_2D => X"0000005e00000000ffffffccffffffff0000003700000000ffffffb1ffffffff",
            INIT_2E => X"0000001200000000ffffffd4ffffffff0000008700000000ffffffd3ffffffff",
            INIT_2F => X"0000011c00000000fffffff1ffffffffffffffaaffffffff0000019800000000",
            INIT_30 => X"0000004300000000000000710000000000000013000000000000009c00000000",
            INIT_31 => X"ffffffc0ffffffffffffff64ffffffff0000004c000000000000002000000000",
            INIT_32 => X"ffffffa8ffffffff00000018000000000000004f000000000000001300000000",
            INIT_33 => X"000000000000000000000047000000000000007700000000000000ad00000000",
            INIT_34 => X"ffffffeeffffffffffffffb1ffffffffffffff3afffffffffffffff2ffffffff",
            INIT_35 => X"ffffff35ffffffffffffffafffffffff0000000a000000000000000900000000",
            INIT_36 => X"ffffff69ffffffff000000430000000000000000000000000000004200000000",
            INIT_37 => X"ffffffeeffffffff000000e6000000000000001f000000000000008800000000",
            INIT_38 => X"ffffffccffffffff000000ba00000000ffffffa1ffffffffffffff37ffffffff",
            INIT_39 => X"0000002300000000ffffffbcffffffffffffffb4ffffffff0000006900000000",
            INIT_3A => X"0000001000000000ffffffc2ffffffff0000002a00000000ffffff4effffffff",
            INIT_3B => X"0000003300000000000000660000000000000039000000000000006e00000000",
            INIT_3C => X"000000620000000000000002000000000000007800000000ffffffdaffffffff",
            INIT_3D => X"fffffff5ffffffffffffffc6ffffffffffffffafffffffffffffffebffffffff",
            INIT_3E => X"0000008a00000000000000b100000000000000a4000000000000000300000000",
            INIT_3F => X"ffffffa0ffffffff000000d1000000000000004e000000000000004400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffffffffffffffffffbdffffffffffffffeaffffffffffffff82ffffffff",
            INIT_41 => X"00000022000000000000000300000000ffffff9affffffff0000005500000000",
            INIT_42 => X"ffffff6dffffffff00000014000000000000004500000000fffffff3ffffffff",
            INIT_43 => X"ffffff84ffffffff0000006e0000000000000062000000000000002500000000",
            INIT_44 => X"0000001400000000ffffff92ffffffff0000003b000000000000002300000000",
            INIT_45 => X"ffffff31ffffffff00000043000000000000006500000000ffffffacffffffff",
            INIT_46 => X"ffffffa3ffffffff0000002600000000ffffffeaffffffffffffffeaffffffff",
            INIT_47 => X"0000000900000000ffffffeaffffffffffffffb0ffffffffffffffe7ffffffff",
            INIT_48 => X"0000002100000000fffffff3ffffffff00000006000000000000001500000000",
            INIT_49 => X"fffffffeffffffff0000000f00000000fffffffcfffffffffffffff6ffffffff",
            INIT_4A => X"fffffff4ffffffff00000079000000000000007d000000000000003c00000000",
            INIT_4B => X"ffffff9dffffffffffffff1fffffffffffffff95ffffffffffffffedffffffff",
            INIT_4C => X"000000b8000000000000003400000000ffffff43ffffffff000000aa00000000",
            INIT_4D => X"ffffffa6ffffffff000000bd000000000000000800000000fffffe95ffffffff",
            INIT_4E => X"fffffff7ffffffffffffffe1ffffffff0000005f00000000ffffff47ffffffff",
            INIT_4F => X"fffffeeaffffffffffffffeffffffffffffffe74ffffffffffffff8bffffffff",
            INIT_50 => X"0000008f0000000000000036000000000000005500000000ffffff8bffffffff",
            INIT_51 => X"00000009000000000000003700000000ffffffc1ffffffff0000004000000000",
            INIT_52 => X"fffffffcffffffff0000005c0000000000000020000000000000001000000000",
            INIT_53 => X"0000000400000000fffffff1ffffffffffffff92ffffffffffffffe5ffffffff",
            INIT_54 => X"ffffffd3ffffffffffffffb4ffffffffffffffcaffffffffffffff26ffffffff",
            INIT_55 => X"0000003e00000000ffffffd6ffffffff00000058000000000000004e00000000",
            INIT_56 => X"ffffffe3ffffffff0000005100000000ffffffc4ffffffff0000001e00000000",
            INIT_57 => X"ffffffe5fffffffffffffee6ffffffff0000005a00000000ffffffabffffffff",
            INIT_58 => X"0000001300000000ffffffb0fffffffffffffe98ffffffff0000004400000000",
            INIT_59 => X"ffffff20ffffffff00000018000000000000002400000000ffffff50ffffffff",
            INIT_5A => X"0000004a00000000ffffffceffffffffffffff89ffffffffffffff68ffffffff",
            INIT_5B => X"ffffffa1ffffffff0000005700000000ffffffebffffffffffffffcbffffffff",
            INIT_5C => X"ffffffd5ffffffffffffff3affffffff0000001b00000000ffffffb2ffffffff",
            INIT_5D => X"0000009b00000000ffffffd2ffffffff0000002e000000000000007000000000",
            INIT_5E => X"ffffff94ffffffffffffffb5ffffffff0000004800000000ffffffebffffffff",
            INIT_5F => X"0000003400000000fffffffdffffffff0000000c00000000000000a100000000",
            INIT_60 => X"00000024000000000000002200000000fffffff5ffffffffffffffdeffffffff",
            INIT_61 => X"ffffff9dffffffffffffffa8ffffffff00000077000000000000001d00000000",
            INIT_62 => X"ffffffb3ffffffff000000480000000000000088000000000000003f00000000",
            INIT_63 => X"000000160000000000000025000000000000002d00000000ffffffe2ffffffff",
            INIT_64 => X"ffffff9bffffffffffffffd6ffffffffffffff70ffffffff0000003100000000",
            INIT_65 => X"0000001c00000000ffffffc8ffffffff0000008d00000000fffffff7ffffffff",
            INIT_66 => X"0000000e00000000ffffffd8ffffffffffffff78ffffffff0000005500000000",
            INIT_67 => X"00000005000000000000005e000000000000001e000000000000001b00000000",
            INIT_68 => X"00000014000000000000005f000000000000003000000000fffffffdffffffff",
            INIT_69 => X"fffffff9ffffffffffffffcfffffffffffffff7affffffff0000000e00000000",
            INIT_6A => X"0000009d00000000ffffffcbffffffff00000032000000000000001f00000000",
            INIT_6B => X"0000000800000000fffffff4fffffffffffffffbffffffff000000c500000000",
            INIT_6C => X"0000000a00000000fffffff5ffffffff0000001b000000000000000500000000",
            INIT_6D => X"ffffffdcffffffff0000000700000000fffffff8fffffffffffffff2ffffffff",
            INIT_6E => X"0000002f000000000000000b00000000ffffffe7ffffffff0000000400000000",
            INIT_6F => X"ffffffd3ffffffffffffffd6ffffffff0000001d00000000ffffffeeffffffff",
            INIT_70 => X"000000a600000000ffffffd1ffffffff00000033000000000000002e00000000",
            INIT_71 => X"ffffffefffffffffffffffb0ffffffffffffffe5ffffffffffffffb6ffffffff",
            INIT_72 => X"ffffff93ffffffffffffff7afffffffffffffff7ffffffff0000002300000000",
            INIT_73 => X"ffffffaaffffffff00000009000000000000003e00000000ffffffd6ffffffff",
            INIT_74 => X"ffffffd8ffffffff000000800000000000000072000000000000000200000000",
            INIT_75 => X"00000033000000000000000100000000ffffffa7ffffffffffffff75ffffffff",
            INIT_76 => X"0000000d000000000000003300000000ffffff87ffffffffffffff95ffffffff",
            INIT_77 => X"0000001300000000000000a000000000ffffff8dffffffff000000cd00000000",
            INIT_78 => X"0000003c00000000ffffffbfffffffffffffffbdfffffffffffffff2ffffffff",
            INIT_79 => X"00000091000000000000005d00000000000000cd000000000000004a00000000",
            INIT_7A => X"0000009d000000000000004c00000000000000b1000000000000011800000000",
            INIT_7B => X"0000000d00000000000000180000000000000018000000000000005800000000",
            INIT_7C => X"ffffffd9ffffffffffffffb1ffffffff0000001f000000000000002600000000",
            INIT_7D => X"ffffff85ffffffffffffffabffffffff0000000000000000ffffff8fffffffff",
            INIT_7E => X"ffffffcdffffffffffffff70ffffffffffffffaaffffffffffffffcaffffffff",
            INIT_7F => X"ffffff5fffffffff0000006700000000ffffffa8ffffffffffffff72ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE2;


    MEM_IWGHT_LAYER1_INSTANCE3 : if BRAM_NAME = "iwght_layer1_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002e00000000ffffffb0ffffffffffffffb1ffffffffffffffddffffffff",
            INIT_01 => X"0000004b000000000000004b00000000ffffffceffffffff0000008900000000",
            INIT_02 => X"000000c50000000000000018000000000000003a000000000000001900000000",
            INIT_03 => X"ffffffa5ffffffff0000001700000000ffffff42ffffffff0000008200000000",
            INIT_04 => X"fffffff9ffffffff00000007000000000000003500000000ffffffc5ffffffff",
            INIT_05 => X"00000006000000000000000d00000000ffffffd0ffffffffffffff65ffffffff",
            INIT_06 => X"ffffffebfffffffffffffffbffffffffffffff7affffffff0000001900000000",
            INIT_07 => X"ffffff97ffffffff000000180000000000000020000000000000001600000000",
            INIT_08 => X"0000001c00000000ffffffdaffffffff00000024000000000000003100000000",
            INIT_09 => X"0000001f00000000ffffff7bffffffff0000004d000000000000000e00000000",
            INIT_0A => X"fffffff8ffffffff0000001600000000ffffff9affffffff0000004800000000",
            INIT_0B => X"00000038000000000000002b000000000000006b000000000000008300000000",
            INIT_0C => X"00000013000000000000000f0000000000000041000000000000009100000000",
            INIT_0D => X"ffffff56ffffffffffffff0cffffffffffffffaaffffffff000000ba00000000",
            INIT_0E => X"ffffff57fffffffffffffeebfffffffffffffed0ffffffffffffffa1ffffffff",
            INIT_0F => X"ffffffedffffffff0000002000000000ffffff88ffffffffffffff32ffffffff",
            INIT_10 => X"0000001800000000000000220000000000000011000000000000000700000000",
            INIT_11 => X"0000002d000000000000001600000000ffffffe7fffffffffffffffeffffffff",
            INIT_12 => X"ffffffddfffffffffffffff1ffffffff000000ab000000000000000000000000",
            INIT_13 => X"fffffff9ffffffffffffffccffffffff0000004b00000000ffffff96ffffffff",
            INIT_14 => X"ffffffe3ffffffff0000004600000000fffffffeffffffffffffff82ffffffff",
            INIT_15 => X"ffffffb9fffffffffffffff5fffffffffffffff7fffffffffffffff4ffffffff",
            INIT_16 => X"00000061000000000000005f00000000ffffffb3fffffffffffffffbffffffff",
            INIT_17 => X"0000000e000000000000002e0000000000000024000000000000006800000000",
            INIT_18 => X"00000044000000000000002e0000000000000003000000000000001500000000",
            INIT_19 => X"fffffff6ffffffffffffff9dffffffffffffffa0ffffffffffffffb2ffffffff",
            INIT_1A => X"0000001700000000ffffff93ffffffffffffff9cffffffffffffff6affffffff",
            INIT_1B => X"0000004d0000000000000091000000000000002b000000000000000f00000000",
            INIT_1C => X"0000005800000000000000a8000000000000003b000000000000006a00000000",
            INIT_1D => X"ffffff9affffffffffffffe3ffffffffffffffc3ffffffff0000000600000000",
            INIT_1E => X"ffffff8affffffffffffffdafffffffffffffff6ffffffffffffffa0ffffffff",
            INIT_1F => X"00000008000000000000003a00000000ffffffffffffffffffffffb3ffffffff",
            INIT_20 => X"ffffffedffffffff00000003000000000000000f00000000ffffffc2ffffffff",
            INIT_21 => X"0000008e000000000000006a00000000ffffffe9ffffffffffffffbfffffffff",
            INIT_22 => X"0000001c00000000000000640000000000000070000000000000000900000000",
            INIT_23 => X"ffffff99ffffffff000000910000000000000072000000000000007b00000000",
            INIT_24 => X"0000001800000000fffffff4ffffffffffffffcdffffffffffffffb8ffffffff",
            INIT_25 => X"ffffffedffffffff00000032000000000000006200000000ffffffe5ffffffff",
            INIT_26 => X"fffffff0ffffffff0000004800000000fffffff3ffffffff0000002300000000",
            INIT_27 => X"00000023000000000000004400000000ffffffbdffffffff0000000b00000000",
            INIT_28 => X"ffffffd9ffffffffffffffd3ffffffff00000032000000000000004f00000000",
            INIT_29 => X"ffffffd4ffffffff00000016000000000000005b00000000ffffff2fffffffff",
            INIT_2A => X"0000002f000000000000003000000000ffffffb4ffffffffffffffe1ffffffff",
            INIT_2B => X"ffffffa7ffffffff0000003900000000ffffff9cfffffffffffffff7ffffffff",
            INIT_2C => X"ffffff6affffffff00000040000000000000000600000000ffffff8fffffffff",
            INIT_2D => X"00000003000000000000003800000000ffffff5fffffffffffffff41ffffffff",
            INIT_2E => X"0000009d00000000000000950000000000000078000000000000002300000000",
            INIT_2F => X"ffffffaaffffffffffffffe3ffffffff00000035000000000000004300000000",
            INIT_30 => X"ffffffb2ffffffffffffffd8ffffffffffffffc3ffffffffffffffeaffffffff",
            INIT_31 => X"0000004700000000000000400000000000000018000000000000000600000000",
            INIT_32 => X"ffffffd3ffffffffffffffdbffffffff00000033000000000000003300000000",
            INIT_33 => X"fffffffdffffffff0000000d000000000000005100000000ffffffddffffffff",
            INIT_34 => X"ffffffe5ffffffff0000000b0000000000000013000000000000000800000000",
            INIT_35 => X"0000000700000000000000170000000000000007000000000000000000000000",
            INIT_36 => X"ffffffc0ffffffffffffffa5ffffffffffffffbfffffffff0000001500000000",
            INIT_37 => X"000000640000000000000036000000000000008e000000000000005f00000000",
            INIT_38 => X"fffffffbffffffff0000003b000000000000002a000000000000001c00000000",
            INIT_39 => X"ffffffb2ffffffff0000001c0000000000000004000000000000001b00000000",
            INIT_3A => X"00000000000000000000005e00000000ffffffe1ffffffffffffffd5ffffffff",
            INIT_3B => X"0000004900000000ffffffffffffffff00000012000000000000005e00000000",
            INIT_3C => X"ffffff5bffffffffffffffd3ffffffffffffffdcffffffff0000002400000000",
            INIT_3D => X"ffffffd0fffffffffffffe31ffffffff0000006d00000000ffffff63ffffffff",
            INIT_3E => X"ffffffc3ffffffffffffff65ffffffffffffffdbffffffff0000009700000000",
            INIT_3F => X"00000032000000000000001200000000ffffffadffffffff0000000100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffe0ffffffff0000003300000000fffffff8ffffffffffffffc9ffffffff",
            INIT_41 => X"00000091000000000000000000000000ffffff4fffffffff0000000c00000000",
            INIT_42 => X"0000001a000000000000002c000000000000000100000000ffffff92ffffffff",
            INIT_43 => X"ffffffd2ffffffff0000004c000000000000007f00000000fffffffeffffffff",
            INIT_44 => X"ffffffddffffffff0000009d000000000000005e000000000000001400000000",
            INIT_45 => X"fffffff9ffffffff000000b1000000000000007900000000ffffffe3ffffffff",
            INIT_46 => X"ffffff28ffffffff00000021000000000000007900000000fffffff7ffffffff",
            INIT_47 => X"0000004000000000ffffffebffffffffffffff9affffffffffffffe8ffffffff",
            INIT_48 => X"00000004000000000000005400000000ffffffb9ffffffffffffffd8ffffffff",
            INIT_49 => X"000000550000000000000025000000000000004d00000000ffffff45ffffffff",
            INIT_4A => X"ffffff94ffffffff0000002200000000000000cf00000000ffffffeeffffffff",
            INIT_4B => X"ffffff5cfffffffffffffff7ffffffff0000003b00000000ffffffe3ffffffff",
            INIT_4C => X"0000003d00000000ffffffb5ffffffffffffffe8ffffffffffffffc5ffffffff",
            INIT_4D => X"0000001400000000ffffff72ffffffff0000004e00000000ffffff76ffffffff",
            INIT_4E => X"0000000a00000000ffffffe9fffffffffffffffdffffffffffffffe8ffffffff",
            INIT_4F => X"0000006e000000000000009700000000ffffff8dffffffffffffffc4ffffffff",
            INIT_50 => X"00000035000000000000006500000000ffffffa1ffffffffffffff96ffffffff",
            INIT_51 => X"ffffffcbffffffff000000a000000000ffffff32ffffffffffffffb3ffffffff",
            INIT_52 => X"ffffff8affffffff0000006b000000000000010800000000ffffff0fffffffff",
            INIT_53 => X"00000001000000000000002900000000ffffff92ffffffffffffff91ffffffff",
            INIT_54 => X"0000002e00000000ffffff72ffffffffffffffd4ffffffffffffffb4ffffffff",
            INIT_55 => X"ffffffd4ffffffffffffff58ffffffffffffffecffffffff0000002000000000",
            INIT_56 => X"0000000500000000ffffff64ffffffffffffff77ffffffffffffffdeffffffff",
            INIT_57 => X"0000001900000000ffffffe8fffffffffffffff6ffffffffffffffd2ffffffff",
            INIT_58 => X"0000001800000000ffffffe2ffffffff0000000f000000000000001a00000000",
            INIT_59 => X"00000001000000000000000000000000fffffff8ffffffff0000001400000000",
            INIT_5A => X"ffffffa7ffffffff0000000b000000000000005700000000ffffffdfffffffff",
            INIT_5B => X"0000003200000000ffffff82fffffffffffffff0ffffffff0000003400000000",
            INIT_5C => X"ffffffd4ffffffffffffffeaffffffff0000000800000000ffffffe2ffffffff",
            INIT_5D => X"ffffffe5ffffffff0000000000000000fffffff8ffffffffffffffecffffffff",
            INIT_5E => X"ffffffe4fffffffffffffff9ffffffff0000001200000000fffffffdffffffff",
            INIT_5F => X"0000001700000000ffffffe6ffffffffffffffe9ffffffff0000000c00000000",
            INIT_60 => X"0000001000000000ffffffdcffffffff0000000000000000fffffff2ffffffff",
            INIT_61 => X"fffffff1fffffffffffffff6ffffffffffffffe7fffffffffffffffdffffffff",
            INIT_62 => X"fffffff8ffffffffffffffe2ffffffff0000000a000000000000001500000000",
            INIT_63 => X"0000000100000000000000000000000000000007000000000000000d00000000",
            INIT_64 => X"fffffff9ffffffffffffffddffffffffffffffe7ffffffffffffffe5ffffffff",
            INIT_65 => X"fffffffcffffffffffffffdeffffffffffffffe2fffffffffffffff2ffffffff",
            INIT_66 => X"fffffff4ffffffffffffffebffffffff00000005000000000000001600000000",
            INIT_67 => X"0000000800000000ffffffecffffffffffffffeaffffffffffffffecffffffff",
            INIT_68 => X"ffffffd9ffffffff0000000e00000000fffffff5ffffffffffffffedffffffff",
            INIT_69 => X"fffffff9ffffffffffffffffffffffff0000000000000000ffffffe1ffffffff",
            INIT_6A => X"0000000b00000000ffffffe1ffffffffffffffe3ffffffff0000000600000000",
            INIT_6B => X"ffffffdbffffffffffffffe9ffffffff0000000b00000000fffffff0ffffffff",
            INIT_6C => X"fffffffeffffffffffffffdfffffffffffffffe5ffffffff0000000b00000000",
            INIT_6D => X"fffffff6ffffffffffffffe9ffffffffffffffeaffffffffffffffdfffffffff",
            INIT_6E => X"ffffffe9ffffffffffffffd8ffffffffffffffedffffffff0000000a00000000",
            INIT_6F => X"fffffff4fffffffffffffffffffffffffffffff3ffffffffffffffe7ffffffff",
            INIT_70 => X"ffffffeeffffffff00000000000000000000001100000000ffffffd0ffffffff",
            INIT_71 => X"fffffffffffffffffffffffdffffffffffffffe9ffffffffffffffeaffffffff",
            INIT_72 => X"fffffffeffffffffffffffe0ffffffffffffffeaffffffff0000000e00000000",
            INIT_73 => X"000000040000000000000002000000000000000400000000fffffffcffffffff",
            INIT_74 => X"ffffffeeffffffffffffffdcffffffff00000004000000000000000600000000",
            INIT_75 => X"ffffffecfffffffffffffff2ffffffffffffffe3ffffffffffffffdeffffffff",
            INIT_76 => X"ffffffeaffffffff000000120000000000000007000000000000001000000000",
            INIT_77 => X"0000000200000000ffffffe8ffffffffffffffdaffffffffffffffdbffffffff",
            INIT_78 => X"fffffffcfffffffffffffff7ffffffffffffffdeffffffff0000000400000000",
            INIT_79 => X"0000000900000000fffffffefffffffffffffffaffffffffffffffe3ffffffff",
            INIT_7A => X"0000001000000000fffffffeffffffff00000000000000000000001400000000",
            INIT_7B => X"00000019000000000000001400000000ffffffedffffffffffffffdeffffffff",
            INIT_7C => X"ffffffe7fffffffffffffff9ffffffff00000019000000000000000e00000000",
            INIT_7D => X"ffffffe3fffffffffffffff7ffffffffffffffeafffffffffffffff8ffffffff",
            INIT_7E => X"0000000b00000000ffffffe8ffffffff0000001200000000ffffffefffffffff",
            INIT_7F => X"fffffff3ffffffffffffffe6fffffffffffffff6ffffffff0000000c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE3;


    MEM_IWGHT_LAYER1_INSTANCE4 : if BRAM_NAME = "iwght_layer1_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffbaffffffff00000031000000000000003800000000ffffff92ffffffff",
            INIT_01 => X"ffffffdafffffffffffffff5ffffffff00000012000000000000004700000000",
            INIT_02 => X"ffffffbafffffffffffffff2ffffffffffffffbdffffffff0000005b00000000",
            INIT_03 => X"ffffffdeffffffffffffff53ffffffffffffff97ffffffffffffffe8ffffffff",
            INIT_04 => X"ffffffe0ffffffff0000003700000000ffffffb7ffffffffffffffd8ffffffff",
            INIT_05 => X"0000002100000000ffffffd7ffffffff00000065000000000000002800000000",
            INIT_06 => X"0000005700000000ffffffe6ffffffff0000001d000000000000000100000000",
            INIT_07 => X"ffffff1effffffff00000061000000000000001b00000000ffffffe8ffffffff",
            INIT_08 => X"fffffffeffffffffffffffafffffffff00000043000000000000006900000000",
            INIT_09 => X"0000002000000000000000b000000000ffffff78ffffffff0000004600000000",
            INIT_0A => X"00000016000000000000004b0000000000000085000000000000003e00000000",
            INIT_0B => X"fffffff0ffffffff0000006e00000000ffffffdbffffffff0000001100000000",
            INIT_0C => X"ffffffd3ffffffff000000a4000000000000007300000000ffffff69ffffffff",
            INIT_0D => X"ffffff99ffffffff0000006a000000000000007100000000ffffffeaffffffff",
            INIT_0E => X"ffffff74ffffffffffffffceffffffff0000004f00000000ffffffabffffffff",
            INIT_0F => X"0000001300000000ffffff7effffffffffffffccffffffff0000003600000000",
            INIT_10 => X"0000003100000000ffffffe7ffffffff00000005000000000000005300000000",
            INIT_11 => X"ffffffd8ffffffff0000004400000000ffffffbbfffffffffffffff4ffffffff",
            INIT_12 => X"ffffff93ffffffff0000001700000000ffffffe7fffffffffffffff5ffffffff",
            INIT_13 => X"ffffffbbffffffffffffffcfffffffff00000058000000000000004100000000",
            INIT_14 => X"0000002300000000ffffffe8ffffffff00000026000000000000002800000000",
            INIT_15 => X"ffffffc6ffffffffffffffebffffffffffffff85ffffffff0000005c00000000",
            INIT_16 => X"0000007c00000000ffffffcaffffffffffffff78ffffffff0000003800000000",
            INIT_17 => X"ffffffd8ffffffff000000c600000000ffffffbcffffffffffffffccffffffff",
            INIT_18 => X"fffffff5ffffffff0000001e000000000000006a00000000ffffff42ffffffff",
            INIT_19 => X"0000005f00000000ffffff97ffffffffffffffe4ffffffff0000008c00000000",
            INIT_1A => X"fffffff3ffffffff0000005600000000ffffff8affffffffffffffc3ffffffff",
            INIT_1B => X"ffffffc6ffffffffffffffd2ffffffff00000064000000000000003200000000",
            INIT_1C => X"0000001f000000000000000400000000ffffffa7ffffffff0000009d00000000",
            INIT_1D => X"0000002c000000000000003d000000000000002e000000000000000d00000000",
            INIT_1E => X"ffffffd6ffffffff000000760000000000000044000000000000003500000000",
            INIT_1F => X"0000001300000000000000070000000000000009000000000000003800000000",
            INIT_20 => X"000000050000000000000005000000000000000c000000000000001b00000000",
            INIT_21 => X"0000001a00000000fffffff4ffffffffffffffe9ffffffff0000000800000000",
            INIT_22 => X"ffffffc9ffffffff0000002d000000000000000f00000000ffffffddffffffff",
            INIT_23 => X"00000011000000000000004300000000ffffffe9ffffffffffffffa0ffffffff",
            INIT_24 => X"0000000100000000000000d3000000000000001200000000ffffff5bffffffff",
            INIT_25 => X"ffffff6cffffffffffffff66fffffffffffffffcffffffff0000003a00000000",
            INIT_26 => X"ffffffdaffffffffffffff3effffffffffffff64ffffffff0000006500000000",
            INIT_27 => X"ffffffb1ffffffffffffff36ffffffffffffffcdffffffffffffffd1ffffffff",
            INIT_28 => X"00000000000000000000001f00000000ffffffbafffffffffffffeacffffffff",
            INIT_29 => X"0000005400000000fffffff4fffffffffffffffdffffffff0000004100000000",
            INIT_2A => X"ffffffd7ffffffffffffff7cffffffff00000025000000000000002700000000",
            INIT_2B => X"ffffff50ffffffffffffff6effffffff0000002c00000000ffffffaaffffffff",
            INIT_2C => X"ffffff18ffffffffffffff72ffffffffffffffc0ffffffffffffff13ffffffff",
            INIT_2D => X"0000000500000000ffffffbcffffffffffffffa8ffffffffffffffe4ffffffff",
            INIT_2E => X"0000003800000000ffffffd2ffffffffffffff7effffffff0000002a00000000",
            INIT_2F => X"000000300000000000000034000000000000002000000000ffffffd5ffffffff",
            INIT_30 => X"0000004000000000ffffffdeffffffff00000031000000000000005e00000000",
            INIT_31 => X"ffffffe1ffffffffffffff7effffffffffffffbbfffffffffffffffcffffffff",
            INIT_32 => X"ffffff72ffffffffffffff93fffffffffffffea6ffffffffffffffe6ffffffff",
            INIT_33 => X"ffffffd6fffffffffffffff1ffffffffffffffddfffffffffffffed6ffffffff",
            INIT_34 => X"fffffff8ffffffffffffff6affffffffffffffffffffffff0000005700000000",
            INIT_35 => X"0000008e00000000ffffffe6ffffffff0000000600000000000000a400000000",
            INIT_36 => X"0000003f00000000ffffff97ffffffffffffffc1ffffffffffffff93ffffffff",
            INIT_37 => X"0000004b0000000000000014000000000000000900000000ffffff98ffffffff",
            INIT_38 => X"ffffffcaffffffff0000000000000000fffffff5ffffffff0000005300000000",
            INIT_39 => X"fffffff4ffffffff0000004100000000ffffff83ffffffffffffffa7ffffffff",
            INIT_3A => X"0000002600000000ffffffccffffffffffffffc7ffffffffffffffc7ffffffff",
            INIT_3B => X"fffffff9ffffffff000000820000000000000092000000000000000000000000",
            INIT_3C => X"0000009200000000ffffffbeffffffffffffffecffffffff0000001a00000000",
            INIT_3D => X"0000004a00000000ffffffe0fffffffffffffff9fffffffffffffffeffffffff",
            INIT_3E => X"ffffffefffffffffffffffa9ffffffffffffff9bffffffff0000008000000000",
            INIT_3F => X"0000000b00000000ffffffdeffffffffffffffefffffffffffffffc0ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffbefffffffffffffff1ffffffffffffff89ffffffff0000005200000000",
            INIT_41 => X"0000003f00000000ffffffe8ffffffff0000005100000000ffffff14ffffffff",
            INIT_42 => X"ffffffddffffffff000000150000000000000004000000000000000400000000",
            INIT_43 => X"0000001500000000ffffffe8ffffffff00000045000000000000006b00000000",
            INIT_44 => X"0000001300000000fffffffaffffffff0000000200000000fffffffeffffffff",
            INIT_45 => X"0000001e00000000000000140000000000000005000000000000000200000000",
            INIT_46 => X"fffffffbffffffff0000001100000000ffffffd9ffffffff0000009000000000",
            INIT_47 => X"ffffffa3ffffffff0000009700000000ffffffc7ffffffffffffff9bffffffff",
            INIT_48 => X"ffffff77ffffffffffffff90ffffffffffffffcfffffffffffffffc8ffffffff",
            INIT_49 => X"000000e200000000ffffffc4ffffffff0000002f000000000000002c00000000",
            INIT_4A => X"0000004a00000000fffffff3ffffffff0000000400000000ffffffe4ffffffff",
            INIT_4B => X"ffffffeaffffffff0000003f00000000ffffffc9fffffffffffffff7ffffffff",
            INIT_4C => X"ffffff3affffffffffffff5affffffffffffff8effffffffffffff92ffffffff",
            INIT_4D => X"ffffffb5ffffffff0000003000000000ffffffcbffffffff0000002300000000",
            INIT_4E => X"000000020000000000000014000000000000002300000000ffffff8fffffffff",
            INIT_4F => X"0000001c00000000000000560000000000000006000000000000006700000000",
            INIT_50 => X"ffffffa1ffffffffffffff6affffffff0000008f000000000000002600000000",
            INIT_51 => X"0000009000000000ffffffccffffffff00000010000000000000006100000000",
            INIT_52 => X"0000005800000000fffffffbfffffffffffffffcffffffff0000004700000000",
            INIT_53 => X"0000007a000000000000002e00000000ffffffceffffffff0000004900000000",
            INIT_54 => X"ffffffd7ffffffff0000004400000000ffffffebfffffffffffffff7ffffffff",
            INIT_55 => X"0000002100000000fffffffeffffffff0000003300000000fffffffeffffffff",
            INIT_56 => X"fffffffbffffffff0000005600000000ffffff78ffffffffffffffe5ffffffff",
            INIT_57 => X"0000001400000000ffffff7cffffffff0000001d00000000ffffff72ffffffff",
            INIT_58 => X"0000004800000000000000f700000000ffffffd3ffffffff0000003700000000",
            INIT_59 => X"ffffff0effffffffffffffd0ffffffff0000008500000000ffffffc0ffffffff",
            INIT_5A => X"fffffefdffffffff0000002a00000000ffffff88ffffffffffffff42ffffffff",
            INIT_5B => X"0000004500000000ffffffe1ffffffff00000085000000000000002d00000000",
            INIT_5C => X"ffffffbdffffffffffffff6affffffffffffffadffffffff0000015400000000",
            INIT_5D => X"fffffd68ffffffff0000005500000000ffffff35fffffffffffffe94ffffffff",
            INIT_5E => X"ffffffc8ffffffffffffff89ffffffff0000011e000000000000010400000000",
            INIT_5F => X"ffffffadffffffff0000009300000000ffffff9cffffffff0000002200000000",
            INIT_60 => X"00000006000000000000002700000000fffffff0ffffffff0000004700000000",
            INIT_61 => X"0000001c00000000000000190000000000000031000000000000005a00000000",
            INIT_62 => X"ffffff3dffffffffffffff71ffffffffffffff9affffffff000000ac00000000",
            INIT_63 => X"ffffff62ffffffffffffff5fffffffffffffff7fffffffffffffffe8ffffffff",
            INIT_64 => X"ffffffd7ffffffffffffff8dffffffff0000008300000000ffffffccffffffff",
            INIT_65 => X"0000003800000000ffffffabfffffffffffffff2ffffffffffffffc4ffffffff",
            INIT_66 => X"ffffff9cffffffff0000000900000000ffffff4fffffffffffffffc8ffffffff",
            INIT_67 => X"ffffffe3fffffffffffffff7ffffffffffffff9fffffffffffffff04ffffffff",
            INIT_68 => X"000000150000000000000019000000000000000200000000fffffff9ffffffff",
            INIT_69 => X"ffffffdbffffffffffffffecffffffff0000000b000000000000001200000000",
            INIT_6A => X"ffffffa3ffffffffffffff29fffffffffffffff5ffffffffffffff88ffffffff",
            INIT_6B => X"00000094000000000000006200000000ffffff8affffffff0000007d00000000",
            INIT_6C => X"ffffffa0ffffffff0000002e0000000000000005000000000000011b00000000",
            INIT_6D => X"ffffffdfffffffff0000005f00000000000000b5000000000000008e00000000",
            INIT_6E => X"ffffffdaffffffff000000ad0000000000000051000000000000001900000000",
            INIT_6F => X"0000003200000000ffffffbeffffffff000001a9000000000000002300000000",
            INIT_70 => X"ffffffc8ffffffff00000024000000000000009c00000000fffffef9ffffffff",
            INIT_71 => X"ffffff29ffffffffffffff56ffffffffffffff31ffffffffffffffe6ffffffff",
            INIT_72 => X"ffffff7affffffff000000a400000000ffffffd3ffffffff0000003000000000",
            INIT_73 => X"fffffedfffffffff000000eb00000000ffffff3affffffffffffffa0ffffffff",
            INIT_74 => X"0000004a000000000000008000000000ffffffedffffffffffffff2bffffffff",
            INIT_75 => X"0000002f00000000ffffff77ffffffffffffffbcffffffff0000003700000000",
            INIT_76 => X"ffffffeeffffffff0000000600000000ffffff51ffffffffffffffd7ffffffff",
            INIT_77 => X"fffffec2ffffffffffffffa6ffffffffffffffd2fffffffffffffeebffffffff",
            INIT_78 => X"0000007d000000000000001f00000000ffffff95ffffffffffffff52ffffffff",
            INIT_79 => X"0000001100000000ffffff94ffffffff00000017000000000000003b00000000",
            INIT_7A => X"0000009b00000000ffffff75fffffffffffffff3ffffffff000000a400000000",
            INIT_7B => X"ffffff50ffffffff000000de00000000fffffe96ffffffffffffff4affffffff",
            INIT_7C => X"fffffe46ffffffffffffff67fffffffffffffec9fffffffffffffffbffffffff",
            INIT_7D => X"000000d200000000ffffff0bffffffff0000000700000000ffffff9dffffffff",
            INIT_7E => X"ffffff9dffffffff0000000900000000ffffff97fffffffffffffefbffffffff",
            INIT_7F => X"0000009b00000000ffffff20ffffffff0000002100000000ffffffebffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE4;


    MEM_IWGHT_LAYER1_INSTANCE5 : if BRAM_NAME = "iwght_layer1_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000aa0000000000000076000000000000005500000000ffffff99ffffffff",
            INIT_01 => X"ffffffe6ffffffff0000004a00000000ffffffe9ffffffff0000007400000000",
            INIT_02 => X"000000490000000000000035000000000000003700000000000000a200000000",
            INIT_03 => X"000000280000000000000072000000000000002500000000ffffff55ffffffff",
            INIT_04 => X"ffffff07ffffffffffffffb7ffffffff000000b5000000000000009500000000",
            INIT_05 => X"fffffd30fffffffffffffcf6ffffffffffffff80fffffffffffffdf2ffffffff",
            INIT_06 => X"fffffe2afffffffffffffff0ffffffff000000e600000000fffffc6effffffff",
            INIT_07 => X"000000ce00000000ffffffb7ffffffffffffffb1ffffffff000000d600000000",
            INIT_08 => X"0000010900000000000000690000000000000051000000000000008900000000",
            INIT_09 => X"0000000c00000000ffffffe2ffffffffffffff37ffffffff000000c100000000",
            INIT_0A => X"ffffffefffffffffffffffbeffffffffffffff15ffffffffffffff18ffffffff",
            INIT_0B => X"fffffff1fffffffffffffff2fffffffffffffeaefffffffffffffd98ffffffff",
            INIT_0C => X"0000001500000000ffffffe1ffffffffffffffecfffffffffffffffbffffffff",
            INIT_0D => X"00000073000000000000000d00000000ffffffecffffffff0000001300000000",
            INIT_0E => X"fffffff9ffffffffffffffc5ffffffff0000003600000000fffffed6ffffffff",
            INIT_0F => X"fffffdfdffffffff000000d4000000000000003600000000ffffffa6ffffffff",
            INIT_10 => X"0000007300000000ffffffd2ffffffff0000002e000000000000007b00000000",
            INIT_11 => X"ffffffbeffffffff0000006b000000000000007a000000000000003c00000000",
            INIT_12 => X"00000035000000000000001c000000000000002300000000ffffffb5ffffffff",
            INIT_13 => X"0000004c000000000000001e000000000000006200000000ffffffa5ffffffff",
            INIT_14 => X"ffffffbbffffffffffffffaeffffffffffffff5dfffffffffffffff3ffffffff",
            INIT_15 => X"0000004300000000ffffffb9ffffffff00000075000000000000002a00000000",
            INIT_16 => X"0000007400000000ffffffa0ffffffff0000000600000000ffffff50ffffffff",
            INIT_17 => X"ffffff57ffffffff00000001000000000000005800000000ffffffbeffffffff",
            INIT_18 => X"ffffff91ffffffff0000003a000000000000001800000000ffffffecffffffff",
            INIT_19 => X"00000060000000000000004f000000000000005100000000ffffffbdffffffff",
            INIT_1A => X"ffffffcbffffffff0000008c00000000ffffffe7ffffffff0000004800000000",
            INIT_1B => X"ffffff5affffffffffffff60ffffffffffffff64fffffffffffffea5ffffffff",
            INIT_1C => X"ffffffbaffffffff000000aa00000000000000a500000000ffffffc8ffffffff",
            INIT_1D => X"ffffff5bffffffff0000008a00000000ffffff4bffffffffffffffb0ffffffff",
            INIT_1E => X"ffffffd8ffffffff0000005100000000ffffff83ffffffff0000000500000000",
            INIT_1F => X"0000005500000000ffffff96ffffffff00000029000000000000001f00000000",
            INIT_20 => X"0000001600000000ffffff99ffffffff00000001000000000000009200000000",
            INIT_21 => X"ffffffe2ffffffff0000000c0000000000000028000000000000000300000000",
            INIT_22 => X"0000007500000000ffffff93ffffffffffffffcbffffffffffffffddffffffff",
            INIT_23 => X"ffffffd5ffffffff00000043000000000000000e00000000000000be00000000",
            INIT_24 => X"ffffff89ffffffffffffffc1ffffffff0000005a00000000ffffff77ffffffff",
            INIT_25 => X"ffffff92ffffffff0000001d00000000ffffff92ffffffff0000002d00000000",
            INIT_26 => X"0000002600000000fffffe6dffffffff0000008600000000fffffff2ffffffff",
            INIT_27 => X"000000390000000000000036000000000000006400000000fffffeabffffffff",
            INIT_28 => X"0000004a00000000ffffff9cffffffffffffff89ffffffff0000008600000000",
            INIT_29 => X"0000005900000000000000470000000000000086000000000000002000000000",
            INIT_2A => X"0000000700000000fffffff5ffffffff0000006b000000000000000800000000",
            INIT_2B => X"0000006400000000ffffff4effffffff0000005500000000ffffffdbffffffff",
            INIT_2C => X"0000009700000000ffffff64ffffffffffffffc6ffffffff0000008b00000000",
            INIT_2D => X"ffffffc1ffffffffffffffc2ffffffffffffffceffffffff0000001d00000000",
            INIT_2E => X"ffffff94ffffffff0000003e00000000ffffff64ffffffffffffff19ffffffff",
            INIT_2F => X"0000000700000000ffffffe6ffffffffffffffe1ffffffffffffffe5ffffffff",
            INIT_30 => X"0000000d00000000ffffffd9ffffffff0000000d000000000000001a00000000",
            INIT_31 => X"0000002c00000000fffffff2fffffffffffffff6ffffffffffffffefffffffff",
            INIT_32 => X"ffffffdfffffffffffffff68ffffffffffffffffffffffffffffffd9ffffffff",
            INIT_33 => X"000000800000000000000029000000000000004400000000fffffff0ffffffff",
            INIT_34 => X"0000000300000000ffffffe8ffffffffffffff0affffffffffffffe3ffffffff",
            INIT_35 => X"0000008f000000000000008b0000000000000058000000000000011d00000000",
            INIT_36 => X"0000004000000000fffffffcffffffff00000078000000000000005700000000",
            INIT_37 => X"0000005d0000000000000027000000000000000200000000ffffffd6ffffffff",
            INIT_38 => X"ffffffe2ffffffffffffffc8ffffffff0000004700000000ffffffdeffffffff",
            INIT_39 => X"0000004c00000000fffffffcffffffff0000001c00000000ffffffecffffffff",
            INIT_3A => X"ffffff4cffffffff000000ab000000000000000400000000000000af00000000",
            INIT_3B => X"ffffffd7ffffffffffffffa6ffffffff0000003c00000000ffffffe0ffffffff",
            INIT_3C => X"0000001b00000000000000c50000000000000003000000000000001800000000",
            INIT_3D => X"ffffffebffffffff0000005b00000000ffffffd9ffffffff0000001700000000",
            INIT_3E => X"ffffffcdffffffff000000070000000000000099000000000000000200000000",
            INIT_3F => X"ffffffedffffffffffffff8dffffffffffffff3afffffffffffffffaffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffff3dfffffffffffffffdffffffffffffffe6ffffffffffffff76ffffffff",
            INIT_41 => X"000000620000000000000020000000000000004600000000ffffffe7ffffffff",
            INIT_42 => X"0000001300000000ffffffc7ffffffff0000001900000000ffffffa0ffffffff",
            INIT_43 => X"0000007f00000000ffffffeaffffffff0000000500000000ffffffd5ffffffff",
            INIT_44 => X"fffffff4ffffffff000000b700000000ffffffb4ffffffff0000005200000000",
            INIT_45 => X"ffffff8bffffffff00000011000000000000007c00000000ffffffbaffffffff",
            INIT_46 => X"ffffff86ffffffffffffffc6ffffffffffffff37fffffffffffffee4ffffffff",
            INIT_47 => X"000000c1000000000000006e000000000000010500000000fffffffeffffffff",
            INIT_48 => X"ffffff32ffffffffffffffc9ffffffffffffffc5ffffffff0000002000000000",
            INIT_49 => X"ffffffbaffffffffffffff92ffffffff000000ba00000000ffffff66ffffffff",
            INIT_4A => X"ffffffe5ffffffffffffffe0ffffffff0000007a00000000000000bd00000000",
            INIT_4B => X"ffffffa9ffffffff00000008000000000000001a000000000000001d00000000",
            INIT_4C => X"ffffff5cffffffff000000e500000000ffffffc7ffffffffffffff95ffffffff",
            INIT_4D => X"ffffff2dffffffff0000002600000000ffffff80ffffffffffffff5effffffff",
            INIT_4E => X"000000f60000000000000054000000000000005f00000000fffffff8ffffffff",
            INIT_4F => X"0000002b00000000ffffff5fffffffffffffff57ffffffff0000002a00000000",
            INIT_50 => X"ffffffd9fffffffffffffffdffffffffffffff73ffffffffffffff99ffffffff",
            INIT_51 => X"ffffffd6ffffffff0000001a0000000000000054000000000000002f00000000",
            INIT_52 => X"fffffff9ffffffffffffffb5ffffffff0000002b000000000000001f00000000",
            INIT_53 => X"fffffff5fffffffffffffffeffffffff0000002200000000ffffffbdffffffff",
            INIT_54 => X"0000001600000000fffffffbffffffff00000009000000000000000b00000000",
            INIT_55 => X"0000003800000000ffffffeaffffffff0000001d00000000ffffffe2ffffffff",
            INIT_56 => X"ffffff1cffffffff0000001a0000000000000037000000000000001400000000",
            INIT_57 => X"ffffffc7ffffffffffffff94ffffffffffffff80ffffffffffffffbcffffffff",
            INIT_58 => X"ffffffe9ffffffffffffff77ffffffffffffffdeffffffffffffffe1ffffffff",
            INIT_59 => X"fffffee9ffffffffffffffd7ffffffffffffff85fffffffffffffe96ffffffff",
            INIT_5A => X"00000000000000000000004b00000000fffffff8ffffffffffffff97ffffffff",
            INIT_5B => X"00000028000000000000001f0000000000000009000000000000003400000000",
            INIT_5C => X"ffffff95ffffffff0000008300000000ffffffaeffffffffffffffd2ffffffff",
            INIT_5D => X"0000005000000000ffffffa9ffffffffffffff28ffffffffffffffe7ffffffff",
            INIT_5E => X"fffffff9ffffffff00000017000000000000002b00000000ffffffe2ffffffff",
            INIT_5F => X"ffffffadffffffff0000001200000000fffffffeffffffffffffffdfffffffff",
            INIT_60 => X"000000450000000000000037000000000000001c000000000000004200000000",
            INIT_61 => X"0000001f000000000000004a0000000000000049000000000000003e00000000",
            INIT_62 => X"0000002a00000000ffffff99ffffffff0000004a00000000000000ae00000000",
            INIT_63 => X"0000004100000000ffffffacfffffffffffffffdffffffffffffffecffffffff",
            INIT_64 => X"ffffffb8ffffffff00000000000000000000004900000000fffffffeffffffff",
            INIT_65 => X"ffffffc9ffffffff00000034000000000000006f00000000ffffffcbffffffff",
            INIT_66 => X"ffffffb2ffffffffffffffe9fffffffffffffffafffffffffffffff5ffffffff",
            INIT_67 => X"0000002400000000ffffff48ffffffff00000013000000000000001900000000",
            INIT_68 => X"ffffff0effffffffffffff6fffffffff00000052000000000000008c00000000",
            INIT_69 => X"ffffff61ffffffffffffffd9ffffffff0000004000000000ffffff27ffffffff",
            INIT_6A => X"00000002000000000000004b00000000fffffff0ffffffff0000000e00000000",
            INIT_6B => X"ffffffd0ffffffffffffffd5ffffffff00000057000000000000008300000000",
            INIT_6C => X"0000004600000000ffffffe0ffffffffffffffb0ffffffffffffff69ffffffff",
            INIT_6D => X"0000001f00000000000000110000000000000031000000000000004900000000",
            INIT_6E => X"ffffff9fffffffff0000005900000000ffffffddffffffffffffffa9ffffffff",
            INIT_6F => X"000000cd000000000000009400000000fffffff4ffffffffffffffb0ffffffff",
            INIT_70 => X"0000001900000000fffffff4ffffffff000000a6000000000000001c00000000",
            INIT_71 => X"ffffffe5ffffffffffffffdeffffffffffffffc9ffffffffffffffe0ffffffff",
            INIT_72 => X"ffffff74ffffffffffffffe7ffffffff0000003a000000000000005a00000000",
            INIT_73 => X"ffffffcdffffffff0000000100000000fffffff8ffffffffffffff95ffffffff",
            INIT_74 => X"000000210000000000000009000000000000005400000000ffffffdfffffffff",
            INIT_75 => X"00000007000000000000003500000000fffffffeffffffff0000004900000000",
            INIT_76 => X"0000007b00000000ffffffb5ffffffffffffff9cffffffffffffffdbffffffff",
            INIT_77 => X"0000001100000000fffffff1ffffffff00000016000000000000002600000000",
            INIT_78 => X"0000000600000000ffffffecffffffff00000000000000000000001500000000",
            INIT_79 => X"ffffffdfffffffff0000000c000000000000000500000000ffffffedffffffff",
            INIT_7A => X"00000055000000000000002a00000000ffffffbaffffffff0000006500000000",
            INIT_7B => X"fffffff7ffffffff0000004700000000ffffffb2ffffffff0000000f00000000",
            INIT_7C => X"000000ec000000000000005200000000ffffffefffffffff0000003200000000",
            INIT_7D => X"0000007700000000fffffff6ffffffffffffffd1ffffffff0000007800000000",
            INIT_7E => X"000000020000000000000079000000000000001800000000ffffff73ffffffff",
            INIT_7F => X"ffffffa7fffffffffffffffdffffffffffffffe5ffffffff000000a000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE5;


    MEM_IWGHT_LAYER1_INSTANCE6 : if BRAM_NAME = "iwght_layer1_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b7000000000000004100000000ffffff1dffffffffffffff74ffffffff",
            INIT_01 => X"ffffffa6ffffffffffffffe7ffffffff000000d700000000000000a200000000",
            INIT_02 => X"ffffff38ffffffff00000056000000000000001400000000ffffffa5ffffffff",
            INIT_03 => X"0000002600000000ffffffbbffffffffffffffe1ffffffffffffffe1ffffffff",
            INIT_04 => X"fffffff1ffffffffffffff9fffffffffffffff4bffffffffffffffe2ffffffff",
            INIT_05 => X"ffffffadffffffffffffff3dffffffffffffff9fffffffff0000001600000000",
            INIT_06 => X"fffffef9ffffffff0000003a00000000fffffec2ffffffffffffff40ffffffff",
            INIT_07 => X"0000000500000000ffffffafffffffffffffffa6ffffffffffffff58ffffffff",
            INIT_08 => X"0000000000000000fffffffcffffffff0000001d00000000ffffffe2ffffffff",
            INIT_09 => X"000000100000000000000007000000000000008700000000ffffffa5ffffffff",
            INIT_0A => X"0000000000000000ffffff48fffffffffffffff3ffffffffffffff9bffffffff",
            INIT_0B => X"ffffffc0ffffffffffffff8bffffffffffffff76fffffffffffffe95ffffffff",
            INIT_0C => X"000000ba00000000ffffff40ffffffff0000007300000000000000e300000000",
            INIT_0D => X"000000aa00000000fffffe78ffffffffffffff8cfffffffffffffffeffffffff",
            INIT_0E => X"0000005700000000000000280000000000000046000000000000006100000000",
            INIT_0F => X"ffffffe7ffffffffffffffd4ffffffff00000088000000000000001400000000",
            INIT_10 => X"0000005600000000ffffff5fffffffff0000008f00000000fffffff4ffffffff",
            INIT_11 => X"00000017000000000000004d000000000000006400000000ffffff8affffffff",
            INIT_12 => X"ffffff93ffffffff0000000100000000ffffffe5fffffffffffffee7ffffffff",
            INIT_13 => X"0000002900000000ffffff7dffffffffffffffa6ffffffff0000005d00000000",
            INIT_14 => X"ffffffcbffffffffffffffdfffffffff0000008400000000ffffffaaffffffff",
            INIT_15 => X"ffffff70ffffffffffffffdcffffffff00000043000000000000003b00000000",
            INIT_16 => X"fffffefcffffffffffffff16ffffffffffffff5effffffff0000000800000000",
            INIT_17 => X"0000003b00000000ffffffefffffffff00000017000000000000001500000000",
            INIT_18 => X"0000008c000000000000002f00000000ffffffa4ffffffff0000003500000000",
            INIT_19 => X"0000002b000000000000007500000000ffffffddffffffffffffff90ffffffff",
            INIT_1A => X"000000a9000000000000003c000000000000005700000000ffffff8dffffffff",
            INIT_1B => X"0000001d00000000ffffffe1ffffffff0000008800000000fffffff0ffffffff",
            INIT_1C => X"00000002000000000000000000000000fffffff4ffffffffffffffe5ffffffff",
            INIT_1D => X"0000005a0000000000000019000000000000000900000000fffffff2ffffffff",
            INIT_1E => X"0000008700000000ffffffadffffffffffffff2affffffff0000002b00000000",
            INIT_1F => X"fffffff9ffffffff00000010000000000000001c000000000000003c00000000",
            INIT_20 => X"ffffffd8ffffffff0000003600000000ffffff95ffffffffffffff3dffffffff",
            INIT_21 => X"000000c5000000000000002c000000000000006b00000000000000ae00000000",
            INIT_22 => X"00000014000000000000005c000000000000004800000000fffffee3ffffffff",
            INIT_23 => X"fffffc9effffffff0000000800000000ffffffa5ffffffffffffff64ffffffff",
            INIT_24 => X"ffffffd5ffffffff0000006b00000000fffffeacffffffffffffffd0ffffffff",
            INIT_25 => X"00000031000000000000002800000000ffffff60ffffffff0000003600000000",
            INIT_26 => X"0000006f00000000000000cb0000000000000006000000000000004900000000",
            INIT_27 => X"0000003700000000000000af00000000000000a700000000fffffffcffffffff",
            INIT_28 => X"fffffeeaffffffffffffff65ffffffffffffff78ffffffff0000003e00000000",
            INIT_29 => X"ffffffecffffffffffffffb9ffffffffffffff67ffffffff0000001800000000",
            INIT_2A => X"0000006800000000000000610000000000000035000000000000003b00000000",
            INIT_2B => X"fffffff2ffffffffffffffc7ffffffffffffffc4ffffffff0000004300000000",
            INIT_2C => X"ffffffedffffffffffffff9effffffffffffff8dffffffffffffffcbffffffff",
            INIT_2D => X"00000050000000000000006e00000000ffffff01ffffffffffffff75ffffffff",
            INIT_2E => X"ffffffa1ffffffff0000008800000000ffffff7dffffffff0000005900000000",
            INIT_2F => X"0000001b00000000fffffedafffffffffffffea7fffffffffffffeeaffffffff",
            INIT_30 => X"fffffffdffffffffffffffd8ffffffffffffffeefffffffffffffff7ffffffff",
            INIT_31 => X"0000009e00000000ffffffc2ffffffffffffffb1ffffffff0000008300000000",
            INIT_32 => X"ffffffb0ffffffff0000003000000000000000a600000000ffffffd4ffffffff",
            INIT_33 => X"ffffff13ffffffffffffffabffffffff0000002700000000fffffff2ffffffff",
            INIT_34 => X"0000004d00000000ffffffe5ffffffff000000c9000000000000007900000000",
            INIT_35 => X"000000c300000000ffffff3bffffffffffffffacffffffff0000005a00000000",
            INIT_36 => X"000000bd000000000000003d00000000fffffef8fffffffffffffc0affffffff",
            INIT_37 => X"ffffff86ffffffffffffffc7ffffffffffffffe4ffffffff0000000500000000",
            INIT_38 => X"0000004800000000000000720000000000000002000000000000003f00000000",
            INIT_39 => X"ffffff97ffffffffffffff6dffffffff000000dd000000000000000d00000000",
            INIT_3A => X"0000000100000000ffffff73fffffffffffffea1fffffffffffffff9ffffffff",
            INIT_3B => X"ffffffb6ffffffff00000024000000000000007600000000fffffffaffffffff",
            INIT_3C => X"ffffffb8ffffffffffffffc5ffffffff0000008d000000000000001a00000000",
            INIT_3D => X"ffffffddffffffffffffffd9ffffffffffffffcfffffffff0000002d00000000",
            INIT_3E => X"0000005000000000ffffffd5ffffffffffffffc2ffffffff000000b100000000",
            INIT_3F => X"0000000d000000000000001b0000000000000006000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000d00000000fffffff5ffffffff0000000000000000ffffffdeffffffff",
            INIT_41 => X"ffffff94ffffffff0000002100000000ffffffffffffffffffffffefffffffff",
            INIT_42 => X"ffffff82ffffffffffffff38ffffffffffffffdbffffffff0000004800000000",
            INIT_43 => X"fffffffdfffffffffffffff2ffffffffffffffb8ffffffff0000000700000000",
            INIT_44 => X"000000d500000000ffffffa3ffffffffffffff69ffffffffffffff98ffffffff",
            INIT_45 => X"0000000a000000000000001f00000000ffffffd4ffffffffffffff36ffffffff",
            INIT_46 => X"ffffffe4ffffffffffffff4dffffffffffffff89ffffffff0000005700000000",
            INIT_47 => X"ffffff72ffffffff0000007200000000ffffffd5fffffffffffffff9ffffffff",
            INIT_48 => X"0000002e00000000000000390000000000000044000000000000005b00000000",
            INIT_49 => X"ffffffdcffffffffffffffbeffffffffffffff68ffffffff0000002400000000",
            INIT_4A => X"0000004d00000000ffffffc7ffffffffffffffa3ffffffff0000006500000000",
            INIT_4B => X"000000b9000000000000005f00000000ffffffcbffffffff0000006200000000",
            INIT_4C => X"00000058000000000000000f000000000000001700000000ffffff8affffffff",
            INIT_4D => X"ffffffe9ffffffffffffffd6ffffffff0000001600000000ffffffe3ffffffff",
            INIT_4E => X"ffffff41ffffffffffffff8affffffffffffffeeffffffff0000009400000000",
            INIT_4F => X"0000004900000000ffffffdbfffffffffffffff5ffffffff0000000b00000000",
            INIT_50 => X"0000002400000000ffffffdfffffffffffffffcdffffffff0000007c00000000",
            INIT_51 => X"0000004900000000ffffffe7ffffffffffffff83ffffffff0000005300000000",
            INIT_52 => X"0000003c00000000000000850000000000000076000000000000000f00000000",
            INIT_53 => X"ffffffe8ffffffff00000089000000000000003b000000000000003300000000",
            INIT_54 => X"0000009b00000000fffffff1ffffffffffffffe6ffffffffffffffa5ffffffff",
            INIT_55 => X"ffffffa8ffffffffffffff41ffffffffffffffb9ffffffff000000c700000000",
            INIT_56 => X"ffffffb9ffffffffffffffa9fffffffffffffff2ffffffff0000003f00000000",
            INIT_57 => X"0000005200000000000000320000000000000000000000000000000200000000",
            INIT_58 => X"ffffff5affffffffffffffbeffffffffffffff9effffffff0000004c00000000",
            INIT_59 => X"ffffffebffffffffffffff26ffffffffffffff85ffffffffffffff07ffffffff",
            INIT_5A => X"0000003e00000000ffffff8fffffffff000000c100000000ffffff78ffffffff",
            INIT_5B => X"ffffffbdffffffff00000065000000000000002d000000000000002900000000",
            INIT_5C => X"ffffffd5ffffffffffffffcdffffffffffffffe6ffffffffffffff2effffffff",
            INIT_5D => X"ffffff85ffffffff0000006a000000000000001700000000ffffffa6ffffffff",
            INIT_5E => X"0000001600000000ffffffb3ffffffffffffffe8ffffffff0000000200000000",
            INIT_5F => X"00000068000000000000004900000000ffffffd6ffffffffffffffd0ffffffff",
            INIT_60 => X"ffffffa9ffffffff0000000d000000000000001900000000ffffffa8ffffffff",
            INIT_61 => X"00000060000000000000008300000000000000e8000000000000003e00000000",
            INIT_62 => X"000000e4000000000000007a000000000000000d00000000000000a100000000",
            INIT_63 => X"ffffffffffffffff0000001200000000ffffff71ffffffffffffffc6ffffffff",
            INIT_64 => X"0000000100000000fffffff1fffffffffffffffdffffffff0000000500000000",
            INIT_65 => X"ffffffa1ffffffff0000000b00000000ffffffe7ffffffffffffffdeffffffff",
            INIT_66 => X"ffffffd6ffffffff00000019000000000000001d00000000ffffffedffffffff",
            INIT_67 => X"00000010000000000000009d00000000ffffffd8ffffffffffffffc8ffffffff",
            INIT_68 => X"ffffffb3ffffffff0000002e000000000000007700000000ffffff58ffffffff",
            INIT_69 => X"fffffffdfffffffffffffffaffffffff000000e6000000000000000f00000000",
            INIT_6A => X"0000000300000000ffffffd4ffffffff0000000f000000000000001800000000",
            INIT_6B => X"ffffffebfffffffffffffff7ffffffff0000000100000000fffffe6dffffffff",
            INIT_6C => X"0000005600000000ffffffbaffffffffffffff91fffffffffffffe7fffffffff",
            INIT_6D => X"ffffffcdfffffffffffffeaafffffffffffffeb2ffffffff0000007300000000",
            INIT_6E => X"fffffffcffffffffffffff18fffffffffffffed9ffffffffffffff7dffffffff",
            INIT_6F => X"ffffffabfffffffffffffff0ffffffff0000007300000000000000cc00000000",
            INIT_70 => X"ffffffcdfffffffffffffe62ffffffffffffff82ffffffff0000003400000000",
            INIT_71 => X"fffffeaeffffffff0000002600000000000000b9000000000000002e00000000",
            INIT_72 => X"fffffeebffffffffffffff22ffffffffffffffe1ffffffffffffff73ffffffff",
            INIT_73 => X"0000000100000000fffffff0ffffffff0000000200000000fffffe80ffffffff",
            INIT_74 => X"ffffffccffffffff0000009e000000000000004200000000ffffffc7ffffffff",
            INIT_75 => X"00000051000000000000007c0000000000000045000000000000000100000000",
            INIT_76 => X"ffffff4cffffffffffffff2dfffffffffffffe64ffffffff0000003700000000",
            INIT_77 => X"ffffffd8fffffffffffffd8cfffffffffffffe21fffffffffffffe63ffffffff",
            INIT_78 => X"ffffffbdffffffff0000003e000000000000008300000000ffffffb0ffffffff",
            INIT_79 => X"ffffffe6fffffffffffffff2ffffffffffffffe9ffffffff0000005900000000",
            INIT_7A => X"ffffffebffffffffffffff5fffffffff0000000a00000000ffffffefffffffff",
            INIT_7B => X"00000040000000000000006300000000ffffffecffffffff0000006000000000",
            INIT_7C => X"ffffffb6ffffffffffffff8affffffffffffffd0ffffffff0000001e00000000",
            INIT_7D => X"ffffffb6ffffffff00000047000000000000004d00000000000000bc00000000",
            INIT_7E => X"0000009a000000000000001800000000ffffff54ffffffffffffffa6ffffffff",
            INIT_7F => X"ffffffb3ffffffff0000000600000000ffffffd1ffffffff0000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE6;


    MEM_IWGHT_LAYER1_INSTANCE7 : if BRAM_NAME = "iwght_layer1_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffe7ffffffff00000013000000000000001100000000fffffff4ffffffff",
            INIT_01 => X"ffffffe4ffffffff0000003800000000ffffffd8ffffffff0000001a00000000",
            INIT_02 => X"ffffffafffffffffffffffd1ffffffff0000001d00000000ffffffbcffffffff",
            INIT_03 => X"ffffffe0ffffffff00000058000000000000001f000000000000004d00000000",
            INIT_04 => X"ffffffa1ffffffffffffff77ffffffffffffffdaffffffffffffff7dffffffff",
            INIT_05 => X"0000004900000000ffffffc4ffffffffffffffcaffffffffffffffc9ffffffff",
            INIT_06 => X"fffffcf5ffffffff00000041000000000000006300000000fffffd02ffffffff",
            INIT_07 => X"ffffffe9ffffffff0000001200000000fffffb64fffffffffffffb7cffffffff",
            INIT_08 => X"0000001000000000ffffffe5fffffffffffffff9ffffffff0000001100000000",
            INIT_09 => X"00000044000000000000000c00000000ffffffeefffffffffffffff3ffffffff",
            INIT_0A => X"00000091000000000000005200000000fffffef9ffffffff0000003900000000",
            INIT_0B => X"ffffff8bfffffffffffffff7ffffffff00000054000000000000002300000000",
            INIT_0C => X"0000005b00000000ffffff9dfffffffffffffff5fffffffffffffea9ffffffff",
            INIT_0D => X"ffffff98ffffffff0000007d00000000ffffffdeffffffffffffff75ffffffff",
            INIT_0E => X"ffffffefffffffff0000004100000000000000ab000000000000003e00000000",
            INIT_0F => X"ffffff90ffffffff00000054000000000000000f00000000ffffffd3ffffffff",
            INIT_10 => X"ffffffebffffffffffffff97ffffffff00000057000000000000003e00000000",
            INIT_11 => X"ffffff3cffffffff00000088000000000000009e00000000ffffff10ffffffff",
            INIT_12 => X"00000034000000000000000200000000ffffffbaffffffff0000003a00000000",
            INIT_13 => X"ffffff7fffffffffffffff98ffffffff0000000700000000ffffffcbffffffff",
            INIT_14 => X"ffffff43ffffffff0000003000000000ffffffd8ffffffffffffff5cffffffff",
            INIT_15 => X"ffffffc5ffffffff00000004000000000000009f00000000ffffff85ffffffff",
            INIT_16 => X"0000004d00000000ffffffb8ffffffff00000033000000000000002e00000000",
            INIT_17 => X"0000002c00000000ffffff86ffffffffffffff56ffffffff0000004c00000000",
            INIT_18 => X"00000054000000000000004b0000000000000012000000000000004200000000",
            INIT_19 => X"fffffff6ffffffff000000230000000000000048000000000000002f00000000",
            INIT_1A => X"ffffffb4fffffffffffffffcffffffffffffffd9ffffffffffffffc1ffffffff",
            INIT_1B => X"00000072000000000000004200000000ffffff7fffffffff0000002300000000",
            INIT_1C => X"0000004f00000000ffffff99ffffffff0000005000000000000000bf00000000",
            INIT_1D => X"ffffffb2ffffffffffffff66ffffffffffffff09ffffffff0000006700000000",
            INIT_1E => X"00000079000000000000003700000000ffffffc8ffffffffffffff87ffffffff",
            INIT_1F => X"ffffff7bffffffff000000c300000000ffffffeaffffffffffffff63ffffffff",
            INIT_20 => X"0000005b00000000ffffff9bffffffffffffffd4ffffffff0000004100000000",
            INIT_21 => X"fffffffcffffffff0000001000000000ffffffdeffffffff0000001b00000000",
            INIT_22 => X"ffffffd5ffffffffffffff02ffffffff0000007700000000ffffffd8ffffffff",
            INIT_23 => X"ffffff90ffffffff00000060000000000000002400000000ffffffdeffffffff",
            INIT_24 => X"000000ad00000000ffffffaeffffffff0000001100000000fffffffbffffffff",
            INIT_25 => X"0000004b00000000000000b700000000fffffffeffffffff0000003700000000",
            INIT_26 => X"ffffffddffffffffffffff94ffffffffffffffe2fffffffffffffff4ffffffff",
            INIT_27 => X"ffffff7bffffffff0000007d000000000000008c000000000000004800000000",
            INIT_28 => X"ffffffcdffffffffffffffbdffffffffffffff5efffffffffffffebeffffffff",
            INIT_29 => X"0000001900000000fffffff5ffffffff0000002100000000ffffffebffffffff",
            INIT_2A => X"0000000900000000ffffffdcffffffff00000018000000000000000700000000",
            INIT_2B => X"00000014000000000000000500000000ffffffa8ffffffff0000005900000000",
            INIT_2C => X"fffffffdffffffff000000180000000000000019000000000000000100000000",
            INIT_2D => X"00000070000000000000000100000000ffffffe3ffffffff0000000200000000",
            INIT_2E => X"ffffff62ffffffff0000003800000000ffffffd2ffffffffffffff34ffffffff",
            INIT_2F => X"00000084000000000000002d000000000000007e000000000000000a00000000",
            INIT_30 => X"ffffffc1ffffffffffffffe1ffffffffffffffc0ffffffffffffffc8ffffffff",
            INIT_31 => X"00000001000000000000014b00000000fffffffaffffffffffffff95ffffffff",
            INIT_32 => X"ffffffe9ffffffff0000005400000000ffffffc3ffffffffffffff8dffffffff",
            INIT_33 => X"fffffff1ffffffffffffff7affffffff00000057000000000000000900000000",
            INIT_34 => X"0000001b00000000ffffffffffffffff0000004100000000ffffffc6ffffffff",
            INIT_35 => X"ffffff5affffffff00000042000000000000002b000000000000003000000000",
            INIT_36 => X"00000024000000000000004f000000000000001e00000000fffffffaffffffff",
            INIT_37 => X"ffffffe1ffffffff00000042000000000000002900000000000000c500000000",
            INIT_38 => X"0000005800000000ffffffefffffffffffffffa4ffffffff0000005300000000",
            INIT_39 => X"ffffffacffffffffffffffacffffffff00000013000000000000006f00000000",
            INIT_3A => X"000000ca00000000fffffffbffffffff0000000f00000000ffffffd8ffffffff",
            INIT_3B => X"00000057000000000000000e0000000000000003000000000000007800000000",
            INIT_3C => X"ffffff66ffffffffffffffd4ffffffffffffff86ffffffffffffff31ffffffff",
            INIT_3D => X"0000000c00000000ffffffeffffffffffffffffaffffffff0000002100000000",
            INIT_3E => X"000000a300000000ffffffd3ffffffff00000030000000000000005e00000000",
            INIT_3F => X"fffffffdffffffff00000056000000000000002000000000ffffffbeffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000056000000000000002000000000ffffff90ffffffff0000005d00000000",
            INIT_41 => X"0000002d00000000000000890000000000000068000000000000001400000000",
            INIT_42 => X"ffffff50ffffffff0000004b00000000000000c700000000fffffecaffffffff",
            INIT_43 => X"fffffff6ffffffffffffff5affffffffffffff61fffffffffffffff5ffffffff",
            INIT_44 => X"fffffff4ffffffff0000006d00000000ffffffb6ffffffff0000002e00000000",
            INIT_45 => X"ffffff09fffffffffffffe84ffffffffffffff15ffffffff0000000600000000",
            INIT_46 => X"fffffffcffffffffffffff5effffffff0000000200000000ffffff7dffffffff",
            INIT_47 => X"ffffffc9ffffffffffffffc5ffffffff0000000500000000ffffff85ffffffff",
            INIT_48 => X"ffffffc8ffffffff0000001500000000ffffffaaffffffff0000003700000000",
            INIT_49 => X"0000000100000000ffffffebffffffff0000006d000000000000001b00000000",
            INIT_4A => X"0000006900000000fffffff2ffffffffffffffa3ffffffff0000005500000000",
            INIT_4B => X"000000200000000000000053000000000000004a000000000000008200000000",
            INIT_4C => X"ffffffd1ffffffffffffff9fffffffff00000019000000000000003300000000",
            INIT_4D => X"00000024000000000000002d000000000000000800000000fffffffbffffffff",
            INIT_4E => X"0000000300000000000000050000000000000017000000000000002e00000000",
            INIT_4F => X"ffffffedffffffff0000001200000000ffffffa5fffffffffffffffeffffffff",
            INIT_50 => X"fffffff5ffffffff0000001200000000ffffffe6ffffffffffffffeaffffffff",
            INIT_51 => X"ffffff77ffffffff0000001b000000000000000f00000000fffffff9ffffffff",
            INIT_52 => X"0000000800000000ffffffe0ffffffff0000000000000000fffffffcffffffff",
            INIT_53 => X"0000006a000000000000004800000000fffffea0fffffffffffffe20ffffffff",
            INIT_54 => X"ffffff73ffffffffffffffe1ffffffff0000009a00000000ffffffd4ffffffff",
            INIT_55 => X"ffffff23ffffffff0000002500000000000000ca000000000000005200000000",
            INIT_56 => X"000000080000000000000051000000000000003700000000ffffffe0ffffffff",
            INIT_57 => X"000000ac00000000ffffff94ffffffffffffffa4ffffffff0000006100000000",
            INIT_58 => X"fffffffdffffffff00000017000000000000003c00000000fffffff6ffffffff",
            INIT_59 => X"0000006b000000000000000c000000000000003800000000fffffffeffffffff",
            INIT_5A => X"ffffffccffffffff00000063000000000000002000000000ffffff8dffffffff",
            INIT_5B => X"fffffff9ffffffff0000003c00000000ffffff43fffffffffffffff0ffffffff",
            INIT_5C => X"ffffffe3ffffffff000000aa0000000000000049000000000000000000000000",
            INIT_5D => X"ffffffb9fffffffffffffffaffffffff0000002700000000ffffffeeffffffff",
            INIT_5E => X"ffffff88ffffffffffffffd8ffffffff0000000a00000000ffffff82ffffffff",
            INIT_5F => X"00000017000000000000004600000000ffffffbfffffffffffffffa3ffffffff",
            INIT_60 => X"00000011000000000000001400000000ffffff61ffffffffffffffdfffffffff",
            INIT_61 => X"0000006b000000000000002800000000ffffffd9ffffffff0000005c00000000",
            INIT_62 => X"0000000f000000000000002d000000000000003200000000ffffff8effffffff",
            INIT_63 => X"00000070000000000000007b00000000000000ad00000000ffffff6affffffff",
            INIT_64 => X"0000000f00000000fffffff8ffffffffffffff92ffffffff0000001100000000",
            INIT_65 => X"ffffffdeffffffffffffffa2ffffffffffffffc9ffffffff0000003400000000",
            INIT_66 => X"ffffffabffffffff00000078000000000000002f00000000ffffff6cffffffff",
            INIT_67 => X"ffffff73ffffffffffffffcaffffffff00000094000000000000003500000000",
            INIT_68 => X"ffffff84ffffffff000000460000000000000044000000000000000d00000000",
            INIT_69 => X"ffffff1fffffffff00000075000000000000007e00000000ffffff3cffffffff",
            INIT_6A => X"ffffffc4ffffffff00000014000000000000005000000000ffffffa1ffffffff",
            INIT_6B => X"ffffffdeffffffffffffffc2ffffffffffffffecffffffff0000000a00000000",
            INIT_6C => X"ffffff70ffffffff0000004900000000ffffff8fffffffff0000003a00000000",
            INIT_6D => X"00000019000000000000004d000000000000005600000000ffffffd9ffffffff",
            INIT_6E => X"ffffffcfffffffffffffff60ffffffffffffffc5ffffffff0000000800000000",
            INIT_6F => X"0000001d00000000ffffff5affffffffffffff52ffffffffffffff04ffffffff",
            INIT_70 => X"0000001c000000000000006200000000fffffffdffffffffffffffe2ffffffff",
            INIT_71 => X"ffffffbcffffffff000000000000000000000028000000000000001a00000000",
            INIT_72 => X"ffffffb0ffffffff0000008200000000000000ce000000000000006d00000000",
            INIT_73 => X"0000000900000000ffffffebffffffff0000000500000000000000c600000000",
            INIT_74 => X"00000000000000000000001d000000000000001500000000fffffff3ffffffff",
            INIT_75 => X"0000007600000000fffffff6fffffffffffffff8ffffffff0000000200000000",
            INIT_76 => X"000000a000000000ffffff6fffffffffffffffbbffffffff0000002e00000000",
            INIT_77 => X"0000007c000000000000003400000000ffffffb2ffffffff0000001600000000",
            INIT_78 => X"000000e200000000fffffff4ffffffff0000002c00000000ffffffbfffffffff",
            INIT_79 => X"ffffff57ffffffffffffffd4ffffffffffffffeeffffffff0000003a00000000",
            INIT_7A => X"ffffffdaffffffffffffff8effffffff0000002300000000ffffffd6ffffffff",
            INIT_7B => X"ffffff61fffffffffffffffeffffffffffffff7affffffffffffffd4ffffffff",
            INIT_7C => X"0000002f000000000000002b0000000000000028000000000000009b00000000",
            INIT_7D => X"ffffffafffffffff0000001b000000000000001700000000ffffff84ffffffff",
            INIT_7E => X"ffffffdaffffffff0000002d000000000000003200000000ffffffd3ffffffff",
            INIT_7F => X"ffffff29ffffffffffffffdfffffffffffffffecffffffffffffff2bffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE7;


    MEM_IWGHT_LAYER1_INSTANCE8 : if BRAM_NAME = "iwght_layer1_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000038000000000000005d00000000ffffffa8ffffffffffffff90ffffffff",
            INIT_01 => X"0000000b000000000000001600000000ffffffffffffffffffffffd9ffffffff",
            INIT_02 => X"0000004700000000000000000000000000000043000000000000004f00000000",
            INIT_03 => X"ffffffe7ffffffff0000007b000000000000002600000000000000cc00000000",
            INIT_04 => X"0000007500000000ffffffc2ffffffff0000007000000000ffffffd7ffffffff",
            INIT_05 => X"ffffff14ffffffffffffff33ffffffffffffffc9ffffffff0000005c00000000",
            INIT_06 => X"ffffff9dffffffffffffffd9ffffffffffffffdeffffffffffffffcdffffffff",
            INIT_07 => X"ffffffabffffffff0000000100000000ffffff7cffffffffffffffd8ffffffff",
            INIT_08 => X"0000000c00000000000000b7000000000000002200000000ffffffe4ffffffff",
            INIT_09 => X"ffffff75ffffffffffffff23ffffffffffffff24fffffffffffffed1ffffffff",
            INIT_0A => X"0000006300000000ffffff93ffffffffffffffedffffffff0000000000000000",
            INIT_0B => X"0000009a000000000000000e0000000000000010000000000000008900000000",
            INIT_0C => X"ffffffedffffffffffffffdcffffffff00000020000000000000004c00000000",
            INIT_0D => X"0000008b00000000ffffff54ffffffff0000000000000000fffffff4ffffffff",
            INIT_0E => X"ffffffe0ffffffffffffffebffffffffffffffdfffffffffffffffe1ffffffff",
            INIT_0F => X"ffffffd3ffffffffffffffbcffffffffffffffc8ffffffffffffffebffffffff",
            INIT_10 => X"000000d100000000000000a4000000000000007e00000000ffffff35ffffffff",
            INIT_11 => X"ffffffc9ffffffffffffffc9ffffffff0000007a000000000000003700000000",
            INIT_12 => X"ffffffb6ffffffffffffff75ffffffffffffffcaffffffffffffff1dffffffff",
            INIT_13 => X"ffffffc1ffffffff0000000400000000ffffffe0fffffffffffffff4ffffffff",
            INIT_14 => X"0000004d000000000000002f00000000ffffffcaffffffff0000004e00000000",
            INIT_15 => X"ffffffb4ffffffff00000015000000000000006b000000000000004900000000",
            INIT_16 => X"0000008b000000000000008a000000000000000f00000000ffffffbfffffffff",
            INIT_17 => X"ffffffe0ffffffff0000001100000000ffffff96ffffffffffffffa7ffffffff",
            INIT_18 => X"00000007000000000000001c00000000ffffffe9ffffffff0000001700000000",
            INIT_19 => X"fffffff7ffffffff00000000000000000000001e000000000000000f00000000",
            INIT_1A => X"0000004e000000000000006a000000000000003d00000000ffffffc1ffffffff",
            INIT_1B => X"ffffffdbffffffff00000072000000000000000700000000ffffffabffffffff",
            INIT_1C => X"0000004c00000000ffffffceffffffffffffffc9ffffffff000000a100000000",
            INIT_1D => X"ffffff90ffffffffffffffb9ffffffffffffffceffffffff000000a100000000",
            INIT_1E => X"ffffffb2ffffffff00000026000000000000002e00000000ffffffefffffffff",
            INIT_1F => X"0000008b0000000000000045000000000000007e00000000ffffffbaffffffff",
            INIT_20 => X"ffffffecffffffffffffffe9ffffffffffffff85ffffffff0000000000000000",
            INIT_21 => X"00000011000000000000006100000000ffffffd0ffffffff0000001f00000000",
            INIT_22 => X"ffffffecffffffffffffffcaffffffff0000000000000000ffffffceffffffff",
            INIT_23 => X"0000002e000000000000001a0000000000000064000000000000000000000000",
            INIT_24 => X"0000003f000000000000001800000000ffffffbbffffffff0000002600000000",
            INIT_25 => X"ffffffffffffffff0000003100000000ffffff9fffffffffffffffccffffffff",
            INIT_26 => X"0000002400000000fffffffdffffffffffffffd2ffffffffffffffb5ffffffff",
            INIT_27 => X"ffffff0effffffffffffff97ffffffff0000007e00000000ffffffbbffffffff",
            INIT_28 => X"ffffffb7ffffffffffffffebffffffff00000056000000000000004900000000",
            INIT_29 => X"ffffffd6ffffffff0000005d00000000000000a9000000000000000d00000000",
            INIT_2A => X"ffffffc1ffffffff000000a00000000000000055000000000000003600000000",
            INIT_2B => X"00000019000000000000000600000000fffffffdfffffffffffffffeffffffff",
            INIT_2C => X"ffffffa2ffffffffffffff49ffffffff00000022000000000000003300000000",
            INIT_2D => X"ffffffbaffffffff00000015000000000000004d00000000000000a400000000",
            INIT_2E => X"0000007300000000ffffff16ffffffffffffffd8ffffffff000000bf00000000",
            INIT_2F => X"0000008000000000ffffffbffffffffffffffff3ffffffff0000006200000000",
            INIT_30 => X"00000046000000000000000900000000ffffffaeffffffffffffff97ffffffff",
            INIT_31 => X"ffffffeeffffffff0000000500000000fffffffdffffffff0000001100000000",
            INIT_32 => X"fffffefaffffffff0000004500000000ffffffb4ffffffff000000be00000000",
            INIT_33 => X"ffffffa2ffffffff0000006b00000000ffffffc4ffffffff000000a200000000",
            INIT_34 => X"ffffff47ffffffff00000042000000000000003700000000ffffffdaffffffff",
            INIT_35 => X"ffffffe2ffffffff000000f500000000ffffffbfffffffffffffff48ffffffff",
            INIT_36 => X"ffffffcdffffffff000000b6000000000000008400000000ffffff6fffffffff",
            INIT_37 => X"00000031000000000000000900000000ffffffc5ffffffff0000009900000000",
            INIT_38 => X"ffffffc2ffffffff0000003600000000ffffffe1ffffffffffffffbaffffffff",
            INIT_39 => X"00000007000000000000007400000000ffffffd5ffffffff0000001200000000",
            INIT_3A => X"000000470000000000000091000000000000003400000000ffffff86ffffffff",
            INIT_3B => X"0000000a00000000ffffffddffffffff0000004f000000000000007500000000",
            INIT_3C => X"ffffffeffffffffffffffffcffffffff0000000700000000ffffffe5ffffffff",
            INIT_3D => X"ffffffb6ffffffffffffffe3fffffffffffffff3ffffffffffffffdbffffffff",
            INIT_3E => X"0000006f000000000000010b00000000ffffff44fffffffffffffeb7ffffffff",
            INIT_3F => X"fffffff0ffffffff00000083000000000000001d00000000ffffff77ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffa2ffffffff0000002900000000ffffff9effffffff0000000900000000",
            INIT_41 => X"ffffffe0ffffffff0000003c000000000000009d00000000ffffffa0ffffffff",
            INIT_42 => X"ffffffc7ffffffff00000024000000000000000b00000000ffffffc0ffffffff",
            INIT_43 => X"fffffff3ffffffff0000007a00000000ffffffeaffffffffffffffc0ffffffff",
            INIT_44 => X"ffffff55ffffffffffffff96ffffffff00000063000000000000004500000000",
            INIT_45 => X"000000470000000000000037000000000000000200000000ffffffa1ffffffff",
            INIT_46 => X"000000f400000000000000050000000000000076000000000000005900000000",
            INIT_47 => X"fffffffcffffffff0000004b000000000000003300000000000000c600000000",
            INIT_48 => X"fffffe52ffffffff0000007200000000ffffffacffffffffffffffbaffffffff",
            INIT_49 => X"ffffff1cffffffff0000008a000000000000003b000000000000005a00000000",
            INIT_4A => X"ffffffa6ffffffffffffff52ffffffffffffffc8ffffffffffffffd4ffffffff",
            INIT_4B => X"ffffffd6ffffffff0000003500000000ffffffe3ffffffffffffffd8ffffffff",
            INIT_4C => X"000000000000000000000025000000000000000600000000ffffffc4ffffffff",
            INIT_4D => X"ffffff9fffffffffffffffe8ffffffffffffffc1ffffffff0000000200000000",
            INIT_4E => X"fffffff5ffffffffffffffbffffffffffffffef4ffffffffffffff78ffffffff",
            INIT_4F => X"ffffff77ffffffffffffff60ffffffff00000047000000000000000c00000000",
            INIT_50 => X"ffffff96ffffffffffffffc9ffffffffffffff95ffffffffffffff79ffffffff",
            INIT_51 => X"ffffffd6ffffffff0000010f00000000ffffff6cffffffff0000004b00000000",
            INIT_52 => X"0000000100000000ffffffbbffffffffffffffd5ffffffffffffff0affffffff",
            INIT_53 => X"0000008b000000000000007c0000000000000091000000000000003200000000",
            INIT_54 => X"ffffff3dffffffff000000020000000000000049000000000000002900000000",
            INIT_55 => X"ffffff8cffffffff000000510000000000000089000000000000004700000000",
            INIT_56 => X"0000008800000000fffffff9ffffffff0000009100000000ffffffdfffffffff",
            INIT_57 => X"00000027000000000000008800000000000000d1000000000000004d00000000",
            INIT_58 => X"ffffff87ffffffffffffff64ffffffffffffff9fffffffff0000002100000000",
            INIT_59 => X"000000a9000000000000003200000000fffffff4ffffffffffffffc3ffffffff",
            INIT_5A => X"0000002b000000000000001d00000000ffffffc0ffffffff000000c400000000",
            INIT_5B => X"0000006a000000000000003a0000000000000053000000000000001000000000",
            INIT_5C => X"00000026000000000000006d0000000000000026000000000000008a00000000",
            INIT_5D => X"fffffe97ffffffffffffff70ffffffffffffff36ffffffffffffff83ffffffff",
            INIT_5E => X"ffffffdbffffffffffffff5bffffffffffffff05fffffffffffffff6ffffffff",
            INIT_5F => X"0000000a000000000000001d000000000000003e00000000ffffff80ffffffff",
            INIT_60 => X"0000000200000000fffffffbffffffff00000002000000000000001000000000",
            INIT_61 => X"ffffffc8ffffffff0000001a000000000000001500000000ffffffe9ffffffff",
            INIT_62 => X"0000005f0000000000000056000000000000003600000000ffffffc4ffffffff",
            INIT_63 => X"ffffffe6ffffffffffffffd5ffffffff0000004f000000000000002b00000000",
            INIT_64 => X"0000000b000000000000008200000000ffffff75ffffffffffffffe6ffffffff",
            INIT_65 => X"0000004000000000000000110000000000000047000000000000004500000000",
            INIT_66 => X"fffffffaffffffff0000004400000000fffffffaffffffff0000002d00000000",
            INIT_67 => X"ffffffa5ffffffff00000034000000000000007a000000000000004c00000000",
            INIT_68 => X"ffffffafffffffff0000000b0000000000000044000000000000009000000000",
            INIT_69 => X"ffffffe2ffffffff0000001900000000ffffff90ffffffff0000002c00000000",
            INIT_6A => X"0000001b00000000000000310000000000000008000000000000006b00000000",
            INIT_6B => X"ffffff5effffffff0000001e00000000fffffff3ffffffff0000007000000000",
            INIT_6C => X"fffffffeffffffff0000002000000000fffffff4ffffffff0000003200000000",
            INIT_6D => X"ffffffc6ffffffffffffffe4ffffffff00000005000000000000002200000000",
            INIT_6E => X"ffffffeaffffffff000000120000000000000014000000000000000900000000",
            INIT_6F => X"fffffff7ffffffff000000c6000000000000008400000000ffffffe1ffffffff",
            INIT_70 => X"ffffffb5ffffffffffffffa3ffffffffffffffdaffffffff0000000b00000000",
            INIT_71 => X"0000007d0000000000000025000000000000003200000000ffffffd2ffffffff",
            INIT_72 => X"0000006000000000ffffffb3ffffffffffffffd7ffffffff0000005300000000",
            INIT_73 => X"ffffffa3fffffffffffffffdffffffff0000002300000000ffffffcbffffffff",
            INIT_74 => X"ffffff7bffffffffffffffe0ffffffffffffffd2ffffffff0000000d00000000",
            INIT_75 => X"0000004000000000ffffff83ffffffff00000036000000000000006800000000",
            INIT_76 => X"0000002f00000000000000150000000000000000000000000000003c00000000",
            INIT_77 => X"0000008f00000000ffffffebffffffff0000000d000000000000008300000000",
            INIT_78 => X"ffffffd9ffffffffffffffceffffffffffffffd4ffffffffffffffd6ffffffff",
            INIT_79 => X"0000005600000000ffffffc1ffffffffffffffaaffffffffffffffd8ffffffff",
            INIT_7A => X"0000006e00000000ffffffe4ffffffffffffffc4ffffffffffffff98ffffffff",
            INIT_7B => X"fffffec6fffffffffffffe9dffffffffffffff7affffffffffffff68ffffffff",
            INIT_7C => X"fffffff4ffffffffffffffa3ffffffffffffff04ffffffffffffffbbffffffff",
            INIT_7D => X"ffffffe3ffffffffffffffc9ffffffff0000002200000000fffffff4ffffffff",
            INIT_7E => X"0000005d000000000000006600000000ffffffbaffffffff0000001f00000000",
            INIT_7F => X"ffffffb8ffffffff00000013000000000000006a000000000000000b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE8;


    MEM_IWGHT_LAYER1_INSTANCE9 : if BRAM_NAME = "iwght_layer1_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002d00000000fffffff8ffffffff00000017000000000000000d00000000",
            INIT_01 => X"0000001100000000ffffffd9ffffffff00000046000000000000000a00000000",
            INIT_02 => X"0000000600000000ffffffbeffffffffffffff82ffffffffffffff7dffffffff",
            INIT_03 => X"ffffffe9ffffffffffffffffffffffffffffffb9ffffffff0000004600000000",
            INIT_04 => X"0000000c000000000000001c00000000fffffff7ffffffff0000001500000000",
            INIT_05 => X"0000003300000000ffffffebfffffffffffffff0ffffffffffffffedffffffff",
            INIT_06 => X"ffffffcaffffffffffffff6affffffffffffffafffffffff0000008d00000000",
            INIT_07 => X"ffffff9effffffff0000004e00000000ffffff88ffffffff0000005f00000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE9;


    MEM_IWGHT_LAYER2_INSTANCE0 : if BRAM_NAME = "iwght_layer2_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000a69d00000000ffff468bffffffff000014a900000000fffff36fffffffff",
            INIT_01 => X"000094ea00000000fffff2d6ffffffffffffafeaffffffff00001aaf00000000",
            INIT_02 => X"0001b05000000000ffffa509ffffffff00005aef00000000ffff088bffffffff",
            INIT_03 => X"000015b700000000fffff3b1ffffffff00003a6200000000fffff194ffffffff",
            INIT_04 => X"00009f08000000000000f52c000000000000bd8d0000000000002b9900000000",
            INIT_05 => X"ffffb8c1ffffffff000037fa00000000fffff730fffffffffffef5aaffffffff",
            INIT_06 => X"00002a4c00000000ffff6bc1ffffffffffff2bf8ffffffffffffbe26ffffffff",
            INIT_07 => X"00002cd700000000ffff7f5affffffff000063f4000000000001defc00000000",
            INIT_08 => X"fffff550ffffffffffffa7d9ffffffffffffe9a3fffffffffffeafc6ffffffff",
            INIT_09 => X"0000497f00000000ffffdcd6ffffffff0000553f00000000000044d000000000",
            INIT_0A => X"0000a6d90000000000005bef00000000ffffd7c1ffffffff0002878000000000",
            INIT_0B => X"ffff8540ffffffff00003068000000000000be8f00000000ffffe07bffffffff",
            INIT_0C => X"0000f0a800000000000106840000000000006e5300000000ffffea8fffffffff",
            INIT_0D => X"0000dc4000000000fffff064ffffffff000076850000000000013e4100000000",
            INIT_0E => X"0000a0c900000000000008ba00000000ffff7409ffffffff000031f000000000",
            INIT_0F => X"ffffcdf9ffffffff000125b800000000000027e600000000fffff041ffffffff",
            INIT_10 => X"fffffff7fffffffffffffffdffffffff0000000000000000fffffff5ffffffff",
            INIT_11 => X"000000030000000000000009000000000000000200000000ffffffe7ffffffff",
            INIT_12 => X"ffffffebfffffffffffffffaffffffff0000000700000000ffffffeeffffffff",
            INIT_13 => X"fffffff1ffffffff00000003000000000000000900000000fffffffbffffffff",
            INIT_14 => X"0000000600000000fffffff5fffffffffffffff3ffffffff0000000200000000",
            INIT_15 => X"fffffff2ffffffff0000000000000000fffffffcfffffffffffffff4ffffffff",
            INIT_16 => X"fffffffcffffffff0000000200000000fffffffaffffffff0000000800000000",
            INIT_17 => X"fffffff6fffffffffffffffefffffffffffffffbfffffffffffffff7ffffffff",
            INIT_18 => X"fffffff0ffffffffffffffe7fffffffffffffff3fffffffffffffffcffffffff",
            INIT_19 => X"000000020000000000000003000000000000000600000000fffffff1ffffffff",
            INIT_1A => X"0000000500000000ffffffe9ffffffff0000000600000000fffffffcffffffff",
            INIT_1B => X"ffffffedffffffff00000001000000000000000500000000ffffffeaffffffff",
            INIT_1C => X"ffffffe5fffffffffffffff8ffffffff00000006000000000000000100000000",
            INIT_1D => X"ffffffe7ffffffffffffffe5fffffffffffffffeffffffff0000000400000000",
            INIT_1E => X"0000001100000000fffffffdffffffff0000000400000000ffffffe8ffffffff",
            INIT_1F => X"fffffff5fffffffffffffff5ffffffff00000005000000000000000100000000",
            INIT_20 => X"fffffffffffffffffffffffaffffffff0000000500000000ffffffedffffffff",
            INIT_21 => X"0000000a00000000fffffff7ffffffffffffffefffffffffffffffefffffffff",
            INIT_22 => X"fffffff1ffffffff00000007000000000000000000000000ffffffefffffffff",
            INIT_23 => X"ffffffffffffffffffffffeffffffffffffffff9fffffffffffffff8ffffffff",
            INIT_24 => X"ffffffffffffffff000000050000000000000006000000000000000000000000",
            INIT_25 => X"fffffff5ffffffff0000000e000000000000000f000000000000000900000000",
            INIT_26 => X"ffffffebffffffffffffffecffffffff0000000a000000000000000000000000",
            INIT_27 => X"0000000500000000ffffffffffffffffffffffedffffffffffffffecffffffff",
            INIT_28 => X"ffffffe2ffffffffffffffeeffffffffffffffffffffffff0000000000000000",
            INIT_29 => X"ffffffe1ffffffffffffffe5ffffffffffffffe6ffffffffffffffe2ffffffff",
            INIT_2A => X"0000000000000000fffffff7ffffffff0000000200000000fffffff0ffffffff",
            INIT_2B => X"ffffffe5fffffffffffffff9ffffffff0000000900000000fffffffbffffffff",
            INIT_2C => X"fffffff5ffffffff0000000100000000ffffffebfffffffffffffff2ffffffff",
            INIT_2D => X"0000000500000000fffffff7ffffffffffffffecffffffff0000000b00000000",
            INIT_2E => X"000000120000000000000005000000000000000000000000fffffff3ffffffff",
            INIT_2F => X"fffffff1fffffffffffffffffffffffffffffff5ffffffffffffffedffffffff",
            INIT_30 => X"fffffffaffffffffffffffebfffffffffffffff1ffffffffffffffffffffffff",
            INIT_31 => X"ffffffedffffffff00000001000000000000000000000000fffffff5ffffffff",
            INIT_32 => X"ffffffffffffffffffffffedffffffffffffffecfffffffffffffffcffffffff",
            INIT_33 => X"fffffffcfffffffffffffff7fffffffffffffff1ffffffffffffffedffffffff",
            INIT_34 => X"ffffffe1ffffffff0000000200000000ffffffedffffffffffffffecffffffff",
            INIT_35 => X"ffffffffffffffff0000000000000000fffffffefffffffffffffff2ffffffff",
            INIT_36 => X"fffffff9ffffffff0000001300000000fffffff1ffffffffffffffebffffffff",
            INIT_37 => X"fffffff5ffffffff00000005000000000000001200000000ffffffffffffffff",
            INIT_38 => X"ffffffe9fffffffffffffffaffffffff0000000300000000ffffffedffffffff",
            INIT_39 => X"fffffffcfffffffffffffffefffffffffffffffbffffffff0000000800000000",
            INIT_3A => X"ffffffe4ffffffffffffffeeffffffff0000000300000000fffffff4ffffffff",
            INIT_3B => X"00000000000000000000000300000000ffffffe3ffffffffffffffeeffffffff",
            INIT_3C => X"ffffffeaffffffffffffffe9ffffffffffffffeffffffffffffffff5ffffffff",
            INIT_3D => X"ffffffefffffffff00000000000000000000000000000000ffffffecffffffff",
            INIT_3E => X"ffffffe7ffffffff0000000b000000000000000f000000000000001000000000",
            INIT_3F => X"ffffffe0ffffffffffffffe8ffffffff00000009000000000000000300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000f00000000fffffff9ffffffffffffffe8fffffffffffffffeffffffff",
            INIT_41 => X"0000001100000000fffffff5ffffffff0000000800000000fffffffaffffffff",
            INIT_42 => X"000000070000000000000013000000000000000200000000ffffffe6ffffffff",
            INIT_43 => X"ffffffe8fffffffffffffffaffffffff0000000e00000000fffffffcffffffff",
            INIT_44 => X"0000000500000000ffffffe9fffffffffffffff5fffffffffffffff7ffffffff",
            INIT_45 => X"ffffffe5fffffffffffffffcffffffffffffffffffffffff0000000400000000",
            INIT_46 => X"fffffffeffffffff0000000500000000fffffff2ffffffff0000000700000000",
            INIT_47 => X"00000000000000000000000200000000fffffff7ffffffff0000000000000000",
            INIT_48 => X"fffffff6ffffffffffffffecffffffff0000000200000000ffffffeaffffffff",
            INIT_49 => X"fffffff3fffffffffffffff2fffffffffffffff9ffffffff0000000600000000",
            INIT_4A => X"0000000800000000ffffffdfffffffff0000000700000000fffffff8ffffffff",
            INIT_4B => X"fffffffdfffffffffffffff6ffffffff0000000100000000ffffffefffffffff",
            INIT_4C => X"ffffffe9ffffffff0000000400000000fffffff5fffffffffffffff5ffffffff",
            INIT_4D => X"ffffffe6fffffffffffffff1ffffffffffffffeafffffffffffffff1ffffffff",
            INIT_4E => X"0000000000000000fffffffffffffffffffffffcffffffffffffffecffffffff",
            INIT_4F => X"ffffffecffffffffffffffe2ffffffff0000000600000000fffffff1ffffffff",
            INIT_50 => X"fffffff2fffffffffffffff8ffffffff0000000100000000fffffff5ffffffff",
            INIT_51 => X"0000000200000000ffffffeffffffffffffffffdffffffffffffffe6ffffffff",
            INIT_52 => X"fffffff6ffffffff0000000500000000ffffffe3ffffffff0000000800000000",
            INIT_53 => X"0000000100000000fffffff9fffffffffffffff2fffffffffffffffeffffffff",
            INIT_54 => X"ffffffedffffffff00000007000000000000001300000000ffffffebffffffff",
            INIT_55 => X"ffffffeafffffffffffffffeffffffffffffffeaffffffffffffffefffffffff",
            INIT_56 => X"ffffffedffffffffffffffe2ffffffffffffffeafffffffffffffff6ffffffff",
            INIT_57 => X"fffffffbffffffff0000000700000000fffffff2ffffffffffffffe6ffffffff",
            INIT_58 => X"ffffffd0ffffffffffffff9fffffffff00000017000000000000004a00000000",
            INIT_59 => X"0000008500000000ffffff17ffffffffffffffadffffffff0000003000000000",
            INIT_5A => X"ffffffe8ffffffffffffff58fffffffffffffe9affffffff0000001500000000",
            INIT_5B => X"0000001600000000ffffff3dffffffff0000005a00000000ffffffdeffffffff",
            INIT_5C => X"00000095000000000000002800000000fffffff4ffffffff000000a000000000",
            INIT_5D => X"0000008000000000fffffff3ffffffffffffff9fffffffff0000002100000000",
            INIT_5E => X"0000004700000000ffffffb3ffffffff0000001b000000000000006300000000",
            INIT_5F => X"0000003b0000000000000042000000000000003c000000000000004700000000",
            INIT_60 => X"00000045000000000000004700000000ffffffd6ffffffff0000004200000000",
            INIT_61 => X"ffffffd0ffffffff0000002000000000ffffff89ffffffffffffff85ffffffff",
            INIT_62 => X"00000142000000000000002d00000000ffffffbeffffffff0000000200000000",
            INIT_63 => X"ffffffd4ffffffff00000059000000000000000b000000000000008400000000",
            INIT_64 => X"ffffff61ffffffff000000cf00000000ffffffa4ffffffffffffffc2ffffffff",
            INIT_65 => X"0000000a00000000ffffff46ffffffff0000000000000000ffffff81ffffffff",
            INIT_66 => X"00000043000000000000005500000000000000e1000000000000001100000000",
            INIT_67 => X"ffffffb0ffffffff0000001e00000000ffffffb4ffffffffffffffcaffffffff",
            INIT_68 => X"fffffe82ffffffffffffff42ffffffffffffff78ffffffff0000001200000000",
            INIT_69 => X"ffffff71ffffffffffffffadffffffffffffffe5ffffffff0000002900000000",
            INIT_6A => X"fffffefaffffffff00000041000000000000006800000000ffffff54ffffffff",
            INIT_6B => X"ffffffa1ffffffffffffffe0ffffffff0000006300000000ffffff6affffffff",
            INIT_6C => X"ffffff90ffffffffffffff9effffffffffffffd4ffffffffffffff0effffffff",
            INIT_6D => X"ffffffd1fffffffffffffef6ffffffff0000002400000000ffffff0cffffffff",
            INIT_6E => X"ffffff9fffffffff000000b800000000ffffffb2ffffffff0000002300000000",
            INIT_6F => X"ffffff79ffffffffffffff7effffffffffffffa4fffffffffffffff6ffffffff",
            INIT_70 => X"ffffffa8ffffffffffffff80ffffffff0000007900000000ffffffdcffffffff",
            INIT_71 => X"ffffffcbffffffffffffff93ffffffffffffff8bffffffff0000006f00000000",
            INIT_72 => X"00000036000000000000008f000000000000009800000000ffffffe6ffffffff",
            INIT_73 => X"ffffff52ffffffffffffffaaffffffff0000007d000000000000005000000000",
            INIT_74 => X"ffffff96fffffffffffffff7ffffffffffffff96ffffffff000000c200000000",
            INIT_75 => X"0000000200000000fffffffdffffffffffffffffffffffffffffff95ffffffff",
            INIT_76 => X"fffffff4ffffffffffffffffffffffffffffffeffffffffffffffff9ffffffff",
            INIT_77 => X"0000004900000000ffffff8bffffffff0000000f00000000ffffffffffffffff",
            INIT_78 => X"0000008c00000000ffffff5fffffffff00000009000000000000001400000000",
            INIT_79 => X"0000002300000000fffffefeffffffff0000001d00000000ffffffe9ffffffff",
            INIT_7A => X"ffffff7dffffffff00000067000000000000001500000000ffffffe4ffffffff",
            INIT_7B => X"0000007f00000000ffffffbbffffffff00000066000000000000006e00000000",
            INIT_7C => X"ffffffa8ffffffff0000002300000000fffffff5ffffffffffffffedffffffff",
            INIT_7D => X"ffffff35ffffffff0000007c000000000000003a00000000ffffffceffffffff",
            INIT_7E => X"fffffffdffffffffffffffc5ffffffffffffffccffffffff0000000200000000",
            INIT_7F => X"0000005900000000ffffff0afffffffffffffffffffffffffffffffcffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE0;


    MEM_IWGHT_LAYER2_INSTANCE1 : if BRAM_NAME = "iwght_layer2_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffeeffffffff0000001e0000000000000058000000000000004d00000000",
            INIT_01 => X"00000069000000000000002700000000ffffffeeffffffff0000009800000000",
            INIT_02 => X"00000070000000000000000100000000ffffff66ffffffff0000006300000000",
            INIT_03 => X"ffffffc0ffffffff000000e700000000ffffffb6ffffffff0000001e00000000",
            INIT_04 => X"00000070000000000000002c000000000000000b00000000ffffff67ffffffff",
            INIT_05 => X"0000002000000000ffffffa2ffffffff0000001c00000000ffffffbfffffffff",
            INIT_06 => X"00000067000000000000001300000000ffffffecffffffff0000004600000000",
            INIT_07 => X"ffffff54ffffffff0000006b00000000000000a2000000000000003b00000000",
            INIT_08 => X"ffffff4bffffffffffffffe7ffffffffffffff59ffffffffffffffbcffffffff",
            INIT_09 => X"ffffff22fffffffffffffe70ffffffffffffffaeffffffff0000008000000000",
            INIT_0A => X"0000012500000000ffffffd1ffffffff000000e600000000fffffef7ffffffff",
            INIT_0B => X"fffffff7ffffffffffffff6affffffff00000056000000000000003900000000",
            INIT_0C => X"ffffff37ffffffffffffffcefffffffffffffea0ffffffff0000000a00000000",
            INIT_0D => X"ffffff9effffffffffffff25ffffffff0000001b00000000000000b400000000",
            INIT_0E => X"0000005e000000000000002c00000000fffffffcffffffff0000004b00000000",
            INIT_0F => X"fffffff1ffffffff0000003100000000ffffffe8ffffffff0000005700000000",
            INIT_10 => X"000000390000000000000058000000000000000d000000000000009000000000",
            INIT_11 => X"0000002b00000000ffffffb4ffffffff00000051000000000000008000000000",
            INIT_12 => X"0000002100000000ffffff51ffffffffffffffdcffffffffffffff2bffffffff",
            INIT_13 => X"fffffe6effffffff0000006900000000ffffffe2ffffffffffffffd0ffffffff",
            INIT_14 => X"00000078000000000000007a00000000ffffffaeffffffffffffffd9ffffffff",
            INIT_15 => X"0000007100000000fffffffbffffffff0000001500000000ffffff44ffffffff",
            INIT_16 => X"ffffff92ffffffff000000020000000000000059000000000000005b00000000",
            INIT_17 => X"000000a0000000000000007000000000ffffffa8ffffffff0000002b00000000",
            INIT_18 => X"ffffff50ffffffffffffff45ffffffff000000de000000000000008d00000000",
            INIT_19 => X"ffffff1bffffffffffffff76ffffffffffffffe6ffffffffffffff68ffffffff",
            INIT_1A => X"0000001000000000ffffff6bfffffffffffffe77ffffffffffffff6bffffffff",
            INIT_1B => X"0000002000000000ffffffefffffffff0000001600000000ffffff35ffffffff",
            INIT_1C => X"ffffffa5ffffffff000000c200000000ffffff9cffffffff0000008e00000000",
            INIT_1D => X"000000de000000000000001f000000000000007900000000ffffff2bffffffff",
            INIT_1E => X"ffffffc2ffffffffffffffc5ffffffff00000000000000000000001f00000000",
            INIT_1F => X"ffffffc7ffffffffffffff57fffffffffffffff8ffffffff0000007700000000",
            INIT_20 => X"0000003700000000ffffffc8ffffffff0000002f00000000fffffffaffffffff",
            INIT_21 => X"0000005800000000ffffff57ffffffff00000062000000000000007b00000000",
            INIT_22 => X"000000ab00000000fffffff4ffffffff0000005b000000000000002600000000",
            INIT_23 => X"0000002e000000000000006a0000000000000108000000000000005100000000",
            INIT_24 => X"ffffff3cffffffff00000070000000000000008400000000ffffff57ffffffff",
            INIT_25 => X"ffffff32fffffffffffffe9cffffffffffffffd2ffffffffffffff2bffffffff",
            INIT_26 => X"00000072000000000000009b00000000ffffffd6ffffffff0000005300000000",
            INIT_27 => X"ffffff31ffffffff0000001c000000000000013a00000000ffffffa4ffffffff",
            INIT_28 => X"ffffff67ffffffffffffff9fffffffff000000a400000000ffffffdaffffffff",
            INIT_29 => X"0000005200000000000000b8000000000000008700000000ffffff53ffffffff",
            INIT_2A => X"0000005800000000ffffffd7ffffffffffffffa9ffffffff0000003300000000",
            INIT_2B => X"ffffffc4ffffffff0000002d00000000fffffde0ffffffff0000004e00000000",
            INIT_2C => X"ffffff61ffffffffffffffe5ffffffff0000001e000000000000008b00000000",
            INIT_2D => X"fffffffaffffffff0000005c00000000ffffffc1ffffffff0000003400000000",
            INIT_2E => X"0000004100000000ffffffc2ffffffffffffff9effffffff0000002600000000",
            INIT_2F => X"0000006300000000ffffff45ffffffff0000000f00000000ffffffbfffffffff",
            INIT_30 => X"ffffff31ffffffffffffff03ffffffff00000067000000000000000100000000",
            INIT_31 => X"00000055000000000000004500000000ffffffc0ffffffffffffffc0ffffffff",
            INIT_32 => X"0000000f00000000ffffffceffffffff0000006800000000ffffff9bffffffff",
            INIT_33 => X"000000d900000000ffffff42ffffffffffffffb1ffffffffffffffa4ffffffff",
            INIT_34 => X"000000d800000000ffffff31fffffffffffffff2ffffffff0000002100000000",
            INIT_35 => X"ffffffd8ffffffff0000001400000000ffffff60ffffffff0000004300000000",
            INIT_36 => X"0000003a00000000ffffffecffffffff0000002a000000000000004e00000000",
            INIT_37 => X"ffffff7effffffffffffff7dffffffffffffff84ffffffffffffffa4ffffffff",
            INIT_38 => X"000000d100000000fffffffbffffffff00000073000000000000000b00000000",
            INIT_39 => X"fffffeb9ffffffffffffffcbffffffff0000004900000000ffffff05ffffffff",
            INIT_3A => X"ffffff99fffffffffffffffcffffffff0000001400000000ffffff06ffffffff",
            INIT_3B => X"000000e1000000000000001900000000ffffffebffffffffffffffb4ffffffff",
            INIT_3C => X"0000001300000000ffffff31ffffffff00000026000000000000006700000000",
            INIT_3D => X"fffffff6ffffffffffffffffffffffff00000019000000000000002100000000",
            INIT_3E => X"fffffff4ffffffff0000000c00000000ffffffedfffffffffffffff3ffffffff",
            INIT_3F => X"0000008e00000000000000800000000000000007000000000000000800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000009000000000000004700000000ffffffb0ffffffff0000002500000000",
            INIT_41 => X"fffffff8ffffffffffffffdeffffffffffffffdaffffffffffffffbeffffffff",
            INIT_42 => X"0000002a00000000fffffef3ffffffffffffffdcfffffffffffffe77ffffffff",
            INIT_43 => X"ffffff99ffffffffffffff80ffffffffffffff75ffffffffffffffc7ffffffff",
            INIT_44 => X"0000007b0000000000000085000000000000009100000000000000a900000000",
            INIT_45 => X"fffffff3ffffffff0000001c00000000fffffe96ffffffffffffffe0ffffffff",
            INIT_46 => X"0000008200000000fffffca5ffffffff0000002700000000000000ab00000000",
            INIT_47 => X"ffffff2bffffffff000000e400000000ffffff53ffffffff0000002600000000",
            INIT_48 => X"ffffff84ffffffffffffff7bffffffff00000092000000000000013200000000",
            INIT_49 => X"000000cc000000000000010100000000ffffff60ffffffffffffff40ffffffff",
            INIT_4A => X"ffffffc6ffffffffffffffe1ffffffff000000cc00000000ffffffd0ffffffff",
            INIT_4B => X"ffffffc9ffffffffffffffe1ffffffff0000001b00000000000000a800000000",
            INIT_4C => X"ffffff09ffffffffffffffe1ffffffff000000a3000000000000005600000000",
            INIT_4D => X"ffffffbcffffffff00000025000000000000005b000000000000001000000000",
            INIT_4E => X"ffffff51fffffffffffffe87ffffffffffffff0cffffffff000000c700000000",
            INIT_4F => X"ffffff49fffffffffffffd67ffffffff000000a000000000ffffff3affffffff",
            INIT_50 => X"ffffffdbffffffffffffff76fffffffffffffe41ffffffffffffff53ffffffff",
            INIT_51 => X"ffffff02ffffffffffffff8dffffffff00000083000000000000009500000000",
            INIT_52 => X"0000000800000000ffffff2ffffffffffffffeebffffffffffffffdcffffffff",
            INIT_53 => X"000000630000000000000105000000000000000300000000ffffff6effffffff",
            INIT_54 => X"0000005e000000000000003d000000000000001000000000ffffff1affffffff",
            INIT_55 => X"ffffff99ffffffff0000008c00000000ffffff21ffffffff0000009e00000000",
            INIT_56 => X"ffffff7bffffffffffffffb2ffffffff0000008f000000000000007f00000000",
            INIT_57 => X"ffffff88ffffffff000000660000000000000153000000000000000f00000000",
            INIT_58 => X"fffffef4ffffffffffffffdaffffffff0000006d00000000ffffffc9ffffffff",
            INIT_59 => X"ffffffb7ffffffffffffff37ffffffff0000002500000000ffffff54ffffffff",
            INIT_5A => X"00000074000000000000003f00000000ffffffc9fffffffffffffff6ffffffff",
            INIT_5B => X"0000002e0000000000000043000000000000006900000000fffffe8cffffffff",
            INIT_5C => X"fffffec8ffffffffffffffe6ffffffff000000f400000000fffffec8ffffffff",
            INIT_5D => X"ffffff10ffffffffffffffd8ffffffff0000003b000000000000004600000000",
            INIT_5E => X"0000008900000000000000e500000000ffffffbdffffffff0000001100000000",
            INIT_5F => X"0000006600000000fffffff7fffffffffffffef5ffffffffffffff45ffffffff",
            INIT_60 => X"000000bc000000000000008e000000000000006500000000fffffee0ffffffff",
            INIT_61 => X"0000006c0000000000000094000000000000009200000000ffffff4dffffffff",
            INIT_62 => X"ffffff86ffffffff00000002000000000000006100000000ffffffebffffffff",
            INIT_63 => X"0000001f000000000000001800000000fffffef9ffffffff0000005a00000000",
            INIT_64 => X"000000c800000000ffffffa0ffffffff0000005200000000ffffff64ffffffff",
            INIT_65 => X"0000005f00000000ffffffe7ffffffff0000000c00000000ffffff4bffffffff",
            INIT_66 => X"ffffffdcffffffff0000001400000000ffffff8cfffffffffffffed9ffffffff",
            INIT_67 => X"0000003a00000000ffffff9cffffffff000000bb000000000000001700000000",
            INIT_68 => X"ffffffffffffffffffffff88ffffffff0000003d000000000000007000000000",
            INIT_69 => X"fffffebcffffffffffffff2ffffffffffffffeddfffffffffffffe67ffffffff",
            INIT_6A => X"000000890000000000000015000000000000000700000000ffffffa7ffffffff",
            INIT_6B => X"000000a0000000000000005600000000000000bf000000000000001000000000",
            INIT_6C => X"0000005500000000ffffffc3ffffffff00000027000000000000006c00000000",
            INIT_6D => X"ffffff6cffffffffffffffaaffffffff0000007a000000000000004300000000",
            INIT_6E => X"0000004f00000000ffffffdfffffffff0000005e000000000000005800000000",
            INIT_6F => X"0000006600000000ffffffdbffffffffffffffe2ffffffffffffffb2ffffffff",
            INIT_70 => X"ffffffcfffffffffffffff8affffffff0000002e000000000000001800000000",
            INIT_71 => X"000000a600000000fffffff8ffffffff00000053000000000000003d00000000",
            INIT_72 => X"ffffff9effffffff0000006700000000ffffff4cffffffff0000008500000000",
            INIT_73 => X"ffffffdaffffffffffffffe6ffffffffffffff90ffffffffffffffacffffffff",
            INIT_74 => X"fffffed9ffffffffffffff52ffffffffffffffb6ffffffffffffff3affffffff",
            INIT_75 => X"ffffff88ffffffffffffffebffffffffffffffd4ffffffffffffff10ffffffff",
            INIT_76 => X"0000005200000000ffffff4affffffffffffffdfffffffff000000e000000000",
            INIT_77 => X"0000000000000000ffffff28fffffffffffffe9affffffffffffff50ffffffff",
            INIT_78 => X"ffffff8fffffffffffffff34ffffffffffffffc5ffffffffffffff86ffffffff",
            INIT_79 => X"ffffff4dfffffffffffffe96ffffffffffffff31ffffffffffffff48ffffffff",
            INIT_7A => X"ffffffe0ffffffffffffffd7ffffffffffffffd5ffffffff0000000400000000",
            INIT_7B => X"ffffff5cffffffffffffffc2ffffffffffffffa4ffffffff0000004b00000000",
            INIT_7C => X"ffffffb7ffffffff000000350000000000000005000000000000006700000000",
            INIT_7D => X"ffffff8effffffffffffff3fffffffffffffff11ffffffffffffffdeffffffff",
            INIT_7E => X"ffffffebffffffff0000002d00000000fffffdafffffffffffffff32ffffffff",
            INIT_7F => X"fffffeb7fffffffffffffeefffffffffffffffd1ffffffffffffffffffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE1;


    MEM_IWGHT_LAYER2_INSTANCE2 : if BRAM_NAME = "iwght_layer2_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000004000000000000002100000000ffffff6dffffffffffffff4effffffff",
            INIT_01 => X"0000003c00000000ffffffffffffffff0000002100000000ffffffefffffffff",
            INIT_02 => X"0000008700000000ffffffa6fffffffffffffff0ffffffff000000aa00000000",
            INIT_03 => X"fffffffaffffffff0000008c000000000000001c00000000ffffffc4ffffffff",
            INIT_04 => X"000000a300000000000000d200000000fffffff0ffffffff000000b700000000",
            INIT_05 => X"0000000f00000000000000100000000000000000000000000000004500000000",
            INIT_06 => X"0000000000000000ffffffe5ffffffffffffffeffffffffffffffff6ffffffff",
            INIT_07 => X"fffffffdffffffff0000001f00000000fffffffffffffffffffffff1ffffffff",
            INIT_08 => X"ffffff46ffffffffffffffdaffffffff0000004700000000ffffff71ffffffff",
            INIT_09 => X"ffffff7cffffffff0000001900000000ffffffd4ffffffff0000001100000000",
            INIT_0A => X"ffffffe0ffffffff0000005c000000000000004900000000ffffffafffffffff",
            INIT_0B => X"ffffff62ffffffff0000001200000000000000b8000000000000005200000000",
            INIT_0C => X"ffffff16ffffffff0000006100000000fffffffdffffffff0000005600000000",
            INIT_0D => X"fffffff1ffffffff0000001700000000ffffffd3ffffffffffffff5cffffffff",
            INIT_0E => X"0000003000000000ffffff64ffffffffffffffa4ffffffffffffff27ffffffff",
            INIT_0F => X"ffffff8fffffffff000000f800000000000000d100000000ffffffdcffffffff",
            INIT_10 => X"ffffff87ffffffff000000730000000000000034000000000000011b00000000",
            INIT_11 => X"ffffffeafffffffffffffffcffffffff0000000000000000ffffffebffffffff",
            INIT_12 => X"ffffff6effffffffffffffd1ffffffff0000006300000000ffffff21ffffffff",
            INIT_13 => X"000000a600000000ffffff9dfffffffffffffff6ffffffff0000006a00000000",
            INIT_14 => X"0000003f00000000ffffffbbffffffff0000005700000000fffffff9ffffffff",
            INIT_15 => X"0000001100000000ffffffebffffffff00000009000000000000001500000000",
            INIT_16 => X"0000003d000000000000001a00000000ffffffb1ffffffff0000000400000000",
            INIT_17 => X"0000009800000000ffffffeeffffffff0000003900000000ffffffb1ffffffff",
            INIT_18 => X"0000003200000000fffffff0ffffffff0000000d00000000ffffffd4ffffffff",
            INIT_19 => X"00000013000000000000001700000000ffffffc3ffffffffffffff8affffffff",
            INIT_1A => X"ffffff56ffffffffffffff0affffffff0000006a00000000ffffffa1ffffffff",
            INIT_1B => X"000000c6000000000000002a00000000ffffffa7ffffffff0000000700000000",
            INIT_1C => X"00000009000000000000002200000000ffffff2fffffffffffffff58ffffffff",
            INIT_1D => X"000000af00000000000000e700000000ffffffdaffffffff0000005f00000000",
            INIT_1E => X"0000001d00000000ffffff9bfffffffffffffff3ffffffff0000007b00000000",
            INIT_1F => X"00000044000000000000002d0000000000000021000000000000007800000000",
            INIT_20 => X"0000008300000000000000290000000000000031000000000000003b00000000",
            INIT_21 => X"0000000a000000000000003800000000ffffffbbffffffff0000000100000000",
            INIT_22 => X"ffffffd9ffffffffffffffd8ffffffffffffff4affffffffffffffddffffffff",
            INIT_23 => X"ffffffb5ffffffffffffffdfffffffff0000007400000000ffffffe1ffffffff",
            INIT_24 => X"0000004d000000000000002e00000000ffffffdeffffffff0000009300000000",
            INIT_25 => X"0000011d000000000000002600000000fffffffeffffffff0000007500000000",
            INIT_26 => X"0000004600000000000000e8000000000000007c00000000000000cb00000000",
            INIT_27 => X"ffffffc6ffffffff0000006a0000000000000011000000000000003400000000",
            INIT_28 => X"ffffffbfffffffffffffffa9ffffffffffffffb8ffffffff0000001500000000",
            INIT_29 => X"0000003b0000000000000070000000000000000a000000000000007c00000000",
            INIT_2A => X"0000013300000000000000bd00000000000000a5000000000000006000000000",
            INIT_2B => X"fffffff7ffffffff00000066000000000000001a000000000000010800000000",
            INIT_2C => X"ffffffcaffffffffffffffcfffffffff00000005000000000000003000000000",
            INIT_2D => X"ffffff8effffffffffffffabfffffffffffffff5ffffffffffffff8dffffffff",
            INIT_2E => X"000000cf00000000ffffff99ffffffff0000005200000000fffffffcffffffff",
            INIT_2F => X"ffffff50ffffffffffffffb9ffffffff000000b900000000ffffffc1ffffffff",
            INIT_30 => X"ffffff69ffffffff00000028000000000000007400000000ffffffc5ffffffff",
            INIT_31 => X"000000ae00000000000000a300000000ffffff25ffffffff0000008400000000",
            INIT_32 => X"ffffffcbffffffffffffff52ffffffff00000043000000000000006700000000",
            INIT_33 => X"ffffff81ffffffffffffff86ffffffffffffff6effffffff0000000300000000",
            INIT_34 => X"ffffff0fffffffff000000da00000000ffffffbdffffffff0000004a00000000",
            INIT_35 => X"0000008600000000ffffff2affffffffffffff63ffffffff0000004000000000",
            INIT_36 => X"fffffedeffffffffffffffabffffffffffffff5effffffffffffffdbffffffff",
            INIT_37 => X"00000032000000000000001300000000fffffec7ffffffff0000002a00000000",
            INIT_38 => X"0000002b00000000ffffff36ffffffffffffffd5ffffffffffffff5dffffffff",
            INIT_39 => X"ffffffd6fffffffffffffef0fffffffffffffffaffffffffffffffcaffffffff",
            INIT_3A => X"fffffeeeffffffff00000035000000000000004f000000000000003500000000",
            INIT_3B => X"ffffff01fffffffffffffff5ffffffff0000010d000000000000002400000000",
            INIT_3C => X"ffffffffffffffff00000075000000000000000400000000ffffff38ffffffff",
            INIT_3D => X"fffffe6efffffffffffffefcffffffffffffff34ffffffffffffff71ffffffff",
            INIT_3E => X"ffffff6affffffffffffffb1fffffffffffffe5dfffffffffffffdd1ffffffff",
            INIT_3F => X"ffffffc9ffffffffffffff47ffffffff0000005e00000000ffffffeaffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffff60fffffffffffffef9ffffffff000000b6000000000000004600000000",
            INIT_41 => X"0000000d00000000ffffffddffffffff0000001000000000ffffffadffffffff",
            INIT_42 => X"ffffff6dffffffffffffffa1ffffffff0000008a00000000ffffff74ffffffff",
            INIT_43 => X"ffffff7effffffff0000006f00000000000000e2000000000000007c00000000",
            INIT_44 => X"fffffeb0ffffffffffffffa4ffffffff0000002000000000ffffff9fffffffff",
            INIT_45 => X"0000008f000000000000005c00000000ffffffeaffffffff0000001700000000",
            INIT_46 => X"0000000d00000000ffffffa6ffffffff0000005500000000fffffffdffffffff",
            INIT_47 => X"0000003d000000000000006400000000000000a900000000ffffffc3ffffffff",
            INIT_48 => X"ffffff84ffffffff0000001300000000fffffff9ffffffff0000001b00000000",
            INIT_49 => X"ffffff37ffffffffffffff4dffffffff00000000000000000000002800000000",
            INIT_4A => X"0000008000000000ffffff7fffffffff000000b500000000ffffffefffffffff",
            INIT_4B => X"ffffff03ffffffff000000530000000000000048000000000000009100000000",
            INIT_4C => X"0000009400000000000000f9000000000000005d00000000ffffffebffffffff",
            INIT_4D => X"0000000000000000fffffffaffffffff00000005000000000000007200000000",
            INIT_4E => X"ffffffebffffffff00000005000000000000000400000000ffffffeeffffffff",
            INIT_4F => X"000000df000000000000002700000000fffffff9ffffffff0000000200000000",
            INIT_50 => X"00000037000000000000000e00000000fffffffeffffffffffffffc5ffffffff",
            INIT_51 => X"ffffff5fffffffff0000005e000000000000003600000000ffffff9cffffffff",
            INIT_52 => X"0000001700000000ffffff6cffffffffffffffd8ffffffff0000005700000000",
            INIT_53 => X"ffffff4bfffffffffffffff1ffffffff0000005300000000ffffffbbffffffff",
            INIT_54 => X"ffffffeafffffffffffffefaffffffffffffff34ffffffffffffffb2ffffffff",
            INIT_55 => X"ffffffa9ffffffff00000032000000000000009400000000ffffffd5ffffffff",
            INIT_56 => X"0000002c00000000ffffffd9ffffffff000000f6000000000000001a00000000",
            INIT_57 => X"000000eb000000000000005a000000000000006b000000000000003600000000",
            INIT_58 => X"0000009100000000ffffffdfffffffffffffffa4ffffffff0000005200000000",
            INIT_59 => X"00000109000000000000012f00000000ffffff3affffffffffffffefffffffff",
            INIT_5A => X"000000cf000000000000015a00000000ffffffdfffffffff0000005a00000000",
            INIT_5B => X"0000001d00000000ffffff2ffffffffffffffc7cffffffffffffffe1ffffffff",
            INIT_5C => X"ffffff8dffffffff000000c9000000000000008100000000fffffe9cffffffff",
            INIT_5D => X"ffffff39ffffffffffffffa1ffffffffffffffd9ffffffff0000006c00000000",
            INIT_5E => X"ffffff4fffffffffffffffa6ffffffff0000007b00000000000000da00000000",
            INIT_5F => X"0000000300000000fffffff9ffffffff0000008d00000000ffffffc6ffffffff",
            INIT_60 => X"ffffff98ffffffff00000061000000000000003b000000000000004b00000000",
            INIT_61 => X"0000005e00000000ffffffa9fffffffffffffeb7fffffffffffffee6ffffffff",
            INIT_62 => X"0000016f00000000000000be000000000000001400000000ffffff9bffffffff",
            INIT_63 => X"ffffff7ffffffffffffffe9cffffffffffffff86ffffffff000000e700000000",
            INIT_64 => X"ffffff1effffffff0000004200000000000000aa00000000ffffffb1ffffffff",
            INIT_65 => X"000000480000000000000000000000000000005c000000000000002100000000",
            INIT_66 => X"ffffff78fffffffffffffffeffffffff0000000e000000000000006400000000",
            INIT_67 => X"ffffff5fffffffff00000028000000000000002a00000000ffffff48ffffffff",
            INIT_68 => X"fffffc9effffffffffffffe5ffffffffffffffaeffffffff0000001900000000",
            INIT_69 => X"0000001700000000fffffea7ffffffff00000042000000000000006000000000",
            INIT_6A => X"fffffefaffffffff0000009d00000000fffffe23ffffffff0000002f00000000",
            INIT_6B => X"00000011000000000000002d00000000ffffff3cfffffffffffffef9ffffffff",
            INIT_6C => X"000000e600000000ffffffe4fffffffffffffe07ffffffff000001b800000000",
            INIT_6D => X"fffffef1ffffffffffffff44fffffffffffffeb9ffffffffffffffa4ffffffff",
            INIT_6E => X"00000055000000000000003f00000000ffffff90fffffffffffffef4ffffffff",
            INIT_6F => X"ffffff66ffffffff000000c5000000000000003d000000000000007b00000000",
            INIT_70 => X"ffffffc3ffffffff0000005900000000fffffffeffffffff000000b900000000",
            INIT_71 => X"0000005800000000ffffffa0ffffffffffffff30ffffffff0000005200000000",
            INIT_72 => X"00000038000000000000006c0000000000000096000000000000007600000000",
            INIT_73 => X"ffffffcdffffffff0000005d00000000ffffffb2ffffffffffffff57ffffffff",
            INIT_74 => X"ffffff29ffffffff00000043000000000000005400000000ffffff23ffffffff",
            INIT_75 => X"ffffffddffffffffffffff51ffffffff0000001200000000ffffff3dffffffff",
            INIT_76 => X"0000009100000000ffffff99fffffffffffffeb1ffffffffffffff84ffffffff",
            INIT_77 => X"ffffff5fffffffff0000000800000000ffffffbdfffffffffffffefeffffffff",
            INIT_78 => X"00000047000000000000000b0000000000000012000000000000002b00000000",
            INIT_79 => X"000000760000000000000032000000000000007a00000000000000ed00000000",
            INIT_7A => X"fffffff6ffffffff000000410000000000000018000000000000001a00000000",
            INIT_7B => X"0000007e00000000ffffffe1ffffffff00000057000000000000008a00000000",
            INIT_7C => X"000000360000000000000026000000000000001f000000000000000d00000000",
            INIT_7D => X"fffffef9ffffffff0000005d00000000ffffffceffffffff0000008b00000000",
            INIT_7E => X"0000000000000000ffffffe6ffffffff00000010000000000000008600000000",
            INIT_7F => X"fffffe6fffffffff00000018000000000000006f00000000ffffff51ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE2;


    MEM_IWGHT_LAYER2_INSTANCE3 : if BRAM_NAME = "iwght_layer2_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffd9ffffffffffffff44ffffffff0000008300000000ffffff14ffffffff",
            INIT_01 => X"0000003100000000fffffff5ffffffffffffff7effffffff0000000900000000",
            INIT_02 => X"0000002c00000000ffffffe3ffffffff00000042000000000000001400000000",
            INIT_03 => X"ffffffd5ffffffff00000019000000000000001f000000000000005f00000000",
            INIT_04 => X"0000008500000000ffffffc1ffffffff0000008c00000000ffffffe9ffffffff",
            INIT_05 => X"00000032000000000000003f00000000fffffffcffffffff0000000c00000000",
            INIT_06 => X"0000005900000000ffffffedffffffffffffff51ffffffff0000002400000000",
            INIT_07 => X"00000044000000000000008800000000fffffffdffffffffffffff4cffffffff",
            INIT_08 => X"ffffff1fffffffffffffffbeffffffffffffffe5ffffffff0000007000000000",
            INIT_09 => X"0000004600000000fffffffbffffffff0000003400000000ffffffaeffffffff",
            INIT_0A => X"0000000600000000ffffffcdffffffff0000008000000000ffffffe3ffffffff",
            INIT_0B => X"ffffff81fffffffffffffff9fffffffffffffee9ffffffff0000004700000000",
            INIT_0C => X"ffffffd2ffffffffffffff86ffffffff00000034000000000000001400000000",
            INIT_0D => X"ffffffe6ffffffff0000000600000000ffffff5fffffffff0000006a00000000",
            INIT_0E => X"ffffff74ffffffff000000d800000000ffffffe6ffffffff0000000e00000000",
            INIT_0F => X"ffffff48ffffffff00000081000000000000007300000000fffffec5ffffffff",
            INIT_10 => X"ffffffa0ffffffff000000280000000000000035000000000000002f00000000",
            INIT_11 => X"ffffff65ffffffffffffff88ffffffff000000be00000000ffffff94ffffffff",
            INIT_12 => X"0000003500000000ffffff82ffffffff00000060000000000000003400000000",
            INIT_13 => X"ffffff45ffffffff000000df00000000ffffffcdffffffffffffffbbffffffff",
            INIT_14 => X"00000038000000000000000200000000ffffffd0ffffffffffffff23ffffffff",
            INIT_15 => X"0000000c00000000fffffffaffffffff0000000200000000ffffffa5ffffffff",
            INIT_16 => X"fffffff2ffffffffffffffe3ffffffff0000001b000000000000001700000000",
            INIT_17 => X"ffffff21ffffffffffffffeafffffffffffffffbffffffff0000000700000000",
            INIT_18 => X"0000009d00000000000000aa00000000ffffffc9fffffffffffffff2ffffffff",
            INIT_19 => X"ffffff78ffffffff0000004a000000000000006b000000000000002800000000",
            INIT_1A => X"fffffe6dffffffffffffffdeffffffff000000cd00000000fffffee9ffffffff",
            INIT_1B => X"ffffff4fffffffffffffff4bffffffff0000000700000000fffffee3ffffffff",
            INIT_1C => X"0000009a000000000000003a000000000000002c00000000000000dc00000000",
            INIT_1D => X"fffffea7ffffffffffffff90ffffffffffffffebffffffffffffffafffffffff",
            INIT_1E => X"00000082000000000000000a00000000ffffffb5ffffffff0000001200000000",
            INIT_1F => X"ffffffadffffffffffffff05ffffffffffffff99ffffffff0000005600000000",
            INIT_20 => X"ffffffe7ffffffffffffffdaffffffffffffff18ffffffff0000000a00000000",
            INIT_21 => X"000000500000000000000003000000000000004400000000ffffff97ffffffff",
            INIT_22 => X"0000006700000000000000c8000000000000006b00000000ffffffffffffffff",
            INIT_23 => X"0000001700000000ffffffecffffffffffffffacffffffffffffffa2ffffffff",
            INIT_24 => X"0000002d00000000000000e7000000000000006400000000ffffff0effffffff",
            INIT_25 => X"0000002b00000000ffffff3bffffffff00000081000000000000001f00000000",
            INIT_26 => X"ffffffe1ffffffff0000009300000000ffffff84ffffffffffffffadffffffff",
            INIT_27 => X"00000017000000000000004f000000000000005100000000ffffffe3ffffffff",
            INIT_28 => X"000000cc00000000fffffff7ffffffff0000004200000000ffffff90ffffffff",
            INIT_29 => X"ffffff9dffffffffffffff1effffffffffffff4afffffffffffffffcffffffff",
            INIT_2A => X"00000031000000000000003d00000000ffffffd6ffffffffffffffe5ffffffff",
            INIT_2B => X"ffffff90ffffffff0000007800000000fffffed2ffffffffffffff40ffffffff",
            INIT_2C => X"ffffffdaffffffff0000006b00000000ffffffefffffffffffffff69ffffffff",
            INIT_2D => X"000000ce00000000000000aa000000000000002300000000fffffffdffffffff",
            INIT_2E => X"ffffff70ffffffff0000001500000000ffffff98ffffffffffffff74ffffffff",
            INIT_2F => X"0000004d00000000000000e3000000000000001300000000ffffff2bffffffff",
            INIT_30 => X"fffffff6ffffffff0000000300000000ffffffcfffffffffffffff92ffffffff",
            INIT_31 => X"ffffff88ffffffffffffffd7ffffffff0000004400000000fffffff9ffffffff",
            INIT_32 => X"ffffffe0ffffffffffffffddffffffffffffffcdffffffffffffffbeffffffff",
            INIT_33 => X"000000d900000000ffffffebffffffffffffffadffffffffffffffd5ffffffff",
            INIT_34 => X"0000000800000000ffffffcfffffffff0000004b000000000000002600000000",
            INIT_35 => X"ffffffabffffffff0000005a00000000ffffffd3ffffffff0000001200000000",
            INIT_36 => X"000000bf00000000000000090000000000000014000000000000003f00000000",
            INIT_37 => X"ffffff8effffffff000000180000000000000018000000000000004900000000",
            INIT_38 => X"ffffff92ffffffff0000001500000000000000cc000000000000000000000000",
            INIT_39 => X"0000006400000000ffffff79ffffffffffffffddffffffff0000007900000000",
            INIT_3A => X"ffffffc6ffffffff000000100000000000000039000000000000000000000000",
            INIT_3B => X"00000021000000000000009e000000000000004100000000fffffffbffffffff",
            INIT_3C => X"ffffff02ffffffffffffffb8ffffffff0000002e00000000ffffff78ffffffff",
            INIT_3D => X"ffffff8efffffffffffffff1ffffffff0000000a00000000ffffffcaffffffff",
            INIT_3E => X"ffffffefffffffffffffffd1ffffffff0000005600000000ffffffa5ffffffff",
            INIT_3F => X"000000d4000000000000002b000000000000000f000000000000001000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffffffffffffffffffff3ffffffffffffffebffffffff0000000400000000",
            INIT_41 => X"fffffff7fffffffffffffffaffffffff0000000a00000000fffffff6ffffffff",
            INIT_42 => X"ffffffebffffffffffffffefffffffff0000000e00000000ffffffdfffffffff",
            INIT_43 => X"00000003000000000000000600000000ffffffe9ffffffffffffffefffffffff",
            INIT_44 => X"ffffffebffffffff0000000700000000fffffff3ffffffffffffffe7ffffffff",
            INIT_45 => X"fffffff7ffffffffffffffe2ffffffffffffffe7fffffffffffffff4ffffffff",
            INIT_46 => X"0000000800000000fffffff3fffffffffffffff2fffffffffffffff5ffffffff",
            INIT_47 => X"ffffffe7fffffffffffffffafffffffffffffff6ffffffffffffffedffffffff",
            INIT_48 => X"ffffffe8fffffffffffffffdfffffffffffffff6ffffffffffffffeeffffffff",
            INIT_49 => X"0000000300000000fffffff9ffffffff0000000500000000ffffffedffffffff",
            INIT_4A => X"00000005000000000000000b0000000000000008000000000000000800000000",
            INIT_4B => X"0000000500000000fffffff3ffffffff0000000b00000000ffffffeaffffffff",
            INIT_4C => X"fffffffefffffffffffffff3ffffffff00000005000000000000000600000000",
            INIT_4D => X"0000000400000000ffffffebffffffff00000005000000000000000500000000",
            INIT_4E => X"0000000000000000fffffff5fffffffffffffff0ffffffff0000000300000000",
            INIT_4F => X"fffffff0ffffffffffffffefffffffff0000000400000000fffffff3ffffffff",
            INIT_50 => X"fffffffefffffffffffffffcffffffff0000000a000000000000000b00000000",
            INIT_51 => X"0000000300000000fffffffbffffffff0000000a00000000fffffff5ffffffff",
            INIT_52 => X"0000000200000000fffffffefffffffffffffff2fffffffffffffff2ffffffff",
            INIT_53 => X"fffffff1ffffffff0000000c00000000ffffffefffffffffffffffffffffffff",
            INIT_54 => X"0000000d00000000fffffff2ffffffffffffffeaffffffffffffffe6ffffffff",
            INIT_55 => X"fffffff9fffffffffffffff3fffffffffffffff8ffffffff0000000800000000",
            INIT_56 => X"ffffffe2ffffffffffffffe4ffffffff0000000000000000fffffff1ffffffff",
            INIT_57 => X"00000011000000000000000300000000fffffffafffffffffffffff8ffffffff",
            INIT_58 => X"ffffffe7ffffffff0000000300000000fffffff7fffffffffffffff2ffffffff",
            INIT_59 => X"fffffff8fffffffffffffff9fffffffffffffff9fffffffffffffff2ffffffff",
            INIT_5A => X"ffffffdeffffffffffffffffffffffffffffffe0fffffffffffffff0ffffffff",
            INIT_5B => X"fffffff1fffffffffffffffdffffffffffffffe8fffffffffffffffeffffffff",
            INIT_5C => X"0000000a00000000fffffff8ffffffffffffffe8fffffffffffffff3ffffffff",
            INIT_5D => X"0000000200000000fffffff5fffffffffffffff0ffffffff0000000a00000000",
            INIT_5E => X"fffffffeffffffff0000000f00000000fffffffbffffffffffffffecffffffff",
            INIT_5F => X"0000000000000000ffffffe9ffffffffffffffedffffffff0000000f00000000",
            INIT_60 => X"fffffff6ffffffffffffffe4ffffffff0000000d000000000000000a00000000",
            INIT_61 => X"0000000500000000ffffffebffffffffffffffeefffffffffffffffaffffffff",
            INIT_62 => X"00000004000000000000000100000000fffffff0ffffffffffffffe8ffffffff",
            INIT_63 => X"fffffffeffffffffffffffe8fffffffffffffffafffffffffffffff9ffffffff",
            INIT_64 => X"ffffffebffffffffffffffeaffffffffffffffeeffffffffffffffe6ffffffff",
            INIT_65 => X"ffffffecfffffffffffffffcfffffffffffffffaffffffff0000000100000000",
            INIT_66 => X"fffffffdffffffffffffffebffffffff00000000000000000000000700000000",
            INIT_67 => X"0000000f000000000000000800000000fffffffffffffffffffffff7ffffffff",
            INIT_68 => X"fffffff6ffffffff00000002000000000000000d000000000000000300000000",
            INIT_69 => X"fffffff7ffffffffffffffe5ffffffff0000000000000000ffffffecffffffff",
            INIT_6A => X"fffffffbffffffff0000000000000000ffffffefffffffff0000000a00000000",
            INIT_6B => X"fffffff2fffffffffffffff3ffffffff0000000400000000fffffffeffffffff",
            INIT_6C => X"00000007000000000000000b000000000000000700000000fffffff4ffffffff",
            INIT_6D => X"ffffffe7ffffffffffffffe9ffffffffffffffffffffffff0000000100000000",
            INIT_6E => X"0000000900000000fffffff7fffffffffffffffaffffffff0000000d00000000",
            INIT_6F => X"0000000800000000fffffff0ffffffffffffffefffffffffffffffe7ffffffff",
            INIT_70 => X"fffffffbffffffff00000000000000000000000700000000ffffffeaffffffff",
            INIT_71 => X"0000000500000000fffffff5fffffffffffffff2fffffffffffffff8ffffffff",
            INIT_72 => X"ffffffebfffffffffffffff7fffffffffffffff3ffffffffffffffeaffffffff",
            INIT_73 => X"fffffff0fffffffffffffffaffffffff0000000a000000000000000800000000",
            INIT_74 => X"ffffffeaffffffffffffffebffffffff0000000900000000fffffff9ffffffff",
            INIT_75 => X"ffffffecffffffff0000000a00000000fffffff5fffffffffffffff0ffffffff",
            INIT_76 => X"00000007000000000000000300000000ffffffe3fffffffffffffffcffffffff",
            INIT_77 => X"0000000000000000fffffff0ffffffff0000000500000000fffffff9ffffffff",
            INIT_78 => X"fffffffefffffffffffffff1fffffffffffffff6fffffffffffffffcffffffff",
            INIT_79 => X"fffffffeffffffffffffffeefffffffffffffff7ffffffff0000000700000000",
            INIT_7A => X"0000000200000000fffffffaffffffff0000000800000000fffffffdffffffff",
            INIT_7B => X"000000020000000000000002000000000000000c000000000000000400000000",
            INIT_7C => X"ffffffe8ffffffffffffffe1ffffffff0000000a00000000ffffffeaffffffff",
            INIT_7D => X"ffffffe6ffffffffffffffe6ffffffffffffffe9ffffffff0000000700000000",
            INIT_7E => X"00000005000000000000000000000000ffffffe5fffffffffffffff6ffffffff",
            INIT_7F => X"0000000600000000fffffff4ffffffffffffffe9ffffffff0000000300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE3;


    MEM_IWGHT_LAYER2_INSTANCE4 : if BRAM_NAME = "iwght_layer2_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff4ffffffff0000000700000000fffffff5fffffffffffffff7ffffffff",
            INIT_01 => X"fffffff5fffffffffffffff9ffffffff0000000400000000ffffffe2ffffffff",
            INIT_02 => X"0000000100000000fffffff0ffffffff0000000800000000fffffffcffffffff",
            INIT_03 => X"fffffff1fffffffffffffff5ffffffffffffffe7ffffffff0000000700000000",
            INIT_04 => X"ffffffecffffffff0000000d00000000ffffffebfffffffffffffff6ffffffff",
            INIT_05 => X"fffffffbffffffffffffffeeffffffff0000000600000000ffffffeaffffffff",
            INIT_06 => X"ffffffecfffffffffffffff4fffffffffffffff5ffffffffffffffffffffffff",
            INIT_07 => X"fffffffafffffffffffffffdffffffffffffffedfffffffffffffff9ffffffff",
            INIT_08 => X"ffffff66ffffffffffffff83ffffffffffffff78ffffffffffffffcbffffffff",
            INIT_09 => X"fffffeb0fffffffffffffef7ffffffffffffff8bfffffffffffffec5ffffffff",
            INIT_0A => X"ffffffb1fffffffffffffff6ffffffffffffffc0ffffffffffffff7bffffffff",
            INIT_0B => X"0000003000000000fffffff7ffffffff00000020000000000000000200000000",
            INIT_0C => X"0000004200000000ffffff71ffffffff00000017000000000000007e00000000",
            INIT_0D => X"0000005400000000000000d700000000ffffff50ffffffffffffffa7ffffffff",
            INIT_0E => X"ffffff57ffffffff0000006400000000ffffffe5ffffffff000000c400000000",
            INIT_0F => X"0000001000000000ffffff4effffffff0000007d00000000ffffff1cffffffff",
            INIT_10 => X"0000002800000000ffffff6fffffffff000000a1000000000000003f00000000",
            INIT_11 => X"0000008800000000fffffff1ffffffffffffff68ffffffffffffffbfffffffff",
            INIT_12 => X"000000160000000000000093000000000000000c000000000000002b00000000",
            INIT_13 => X"ffffff7cffffffffffffffbdffffffff00000012000000000000005c00000000",
            INIT_14 => X"ffffffdcffffffffffffff8fffffffffffffff7efffffffffffffff3ffffffff",
            INIT_15 => X"ffffff84ffffffff0000006200000000ffffffc0ffffffff0000000400000000",
            INIT_16 => X"ffffff1fffffffff00000096000000000000007f000000000000000100000000",
            INIT_17 => X"000000a30000000000000074000000000000005300000000ffffffbdffffffff",
            INIT_18 => X"000000350000000000000060000000000000008600000000ffffffcbffffffff",
            INIT_19 => X"fffffffcfffffffffffffff8ffffffff00000051000000000000005100000000",
            INIT_1A => X"ffffffc6ffffffff0000000800000000ffffffccffffffff0000005f00000000",
            INIT_1B => X"ffffff9fffffffff0000005c000000000000006600000000ffffffc4ffffffff",
            INIT_1C => X"ffffff92fffffffffffffef1ffffffffffffff87ffffffffffffff66ffffffff",
            INIT_1D => X"ffffff7dfffffffffffffedcfffffffffffffe7cffffffffffffff4dffffffff",
            INIT_1E => X"ffffffe0ffffffffffffff93ffffffffffffff77ffffffff0000006c00000000",
            INIT_1F => X"ffffff71ffffffffffffff98ffffffff00000012000000000000003100000000",
            INIT_20 => X"00000068000000000000003900000000ffffff72ffffffff0000002200000000",
            INIT_21 => X"0000004c000000000000001500000000000000a4000000000000004a00000000",
            INIT_22 => X"0000003600000000ffffffcdffffffffffffff90fffffffffffffff8ffffffff",
            INIT_23 => X"ffffffb0ffffffff00000038000000000000005b00000000fffffff9ffffffff",
            INIT_24 => X"0000007000000000ffffffbfffffffffffffffd6ffffffffffffffe3ffffffff",
            INIT_25 => X"00000013000000000000000500000000fffffff0ffffffff0000004800000000",
            INIT_26 => X"fffffff3ffffffff0000000f0000000000000002000000000000000c00000000",
            INIT_27 => X"ffffff94ffffffffffffffcafffffffffffffff1ffffffffffffffe0ffffffff",
            INIT_28 => X"00000026000000000000000f00000000ffffffe1ffffffffffffffa7ffffffff",
            INIT_29 => X"ffffff81ffffffff0000002f00000000ffffffd8ffffffffffffff29ffffffff",
            INIT_2A => X"ffffff1fffffffff00000045000000000000003c00000000fffffec2ffffffff",
            INIT_2B => X"0000006c0000000000000008000000000000008600000000ffffff22ffffffff",
            INIT_2C => X"0000009b00000000ffffffb2ffffffff0000003300000000000000a500000000",
            INIT_2D => X"0000000700000000000000a00000000000000009000000000000002e00000000",
            INIT_2E => X"000000fd00000000ffffff48ffffffffffffff5efffffffffffffe2affffffff",
            INIT_2F => X"ffffffb2ffffffffffffff78ffffffff000000bc000000000000003f00000000",
            INIT_30 => X"ffffffb9ffffffffffffffbcffffffff0000003800000000000000ec00000000",
            INIT_31 => X"00000012000000000000000d00000000ffffffd9ffffffffffffffd2ffffffff",
            INIT_32 => X"00000020000000000000009600000000ffffffceffffffffffffffcbffffffff",
            INIT_33 => X"ffffffe9ffffffff00000078000000000000001800000000ffffff0effffffff",
            INIT_34 => X"0000008b0000000000000019000000000000003800000000fffffff0ffffffff",
            INIT_35 => X"ffffffb3ffffffff000000ac000000000000003d00000000ffffffdfffffffff",
            INIT_36 => X"ffffff88ffffffff00000059000000000000000500000000ffffffe0ffffffff",
            INIT_37 => X"ffffff52fffffffffffffee6ffffffff0000006900000000ffffff2dffffffff",
            INIT_38 => X"0000011000000000ffffffcaffffffff0000008c00000000ffffff8cffffffff",
            INIT_39 => X"0000002200000000ffffff69ffffffffffffffbfffffffffffffffc6ffffffff",
            INIT_3A => X"fffffffaffffffffffffffd6ffffffffffffffc7ffffffffffffff26ffffffff",
            INIT_3B => X"ffffffdcffffffffffffffc3ffffffffffffffa9ffffffff0000008d00000000",
            INIT_3C => X"0000002b000000000000003300000000ffffff9cfffffffffffffff6ffffffff",
            INIT_3D => X"000000800000000000000047000000000000004e00000000ffffffd4ffffffff",
            INIT_3E => X"0000006f00000000ffffffa8ffffffffffffffe2ffffffff0000007800000000",
            INIT_3F => X"fffffff1ffffffff0000005b00000000ffffffc0fffffffffffffff5ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffffffffffff0000002900000000ffffffc5ffffffff0000008500000000",
            INIT_41 => X"fffffefcffffffffffffff75ffffffff0000005d00000000ffffff5fffffffff",
            INIT_42 => X"ffffffd5ffffffffffffff9cffffffffffffffbdffffffff000000fe00000000",
            INIT_43 => X"00000091000000000000005600000000ffffff76ffffffff0000002c00000000",
            INIT_44 => X"00000088000000000000001a00000000ffffff83ffffffff0000004c00000000",
            INIT_45 => X"0000004d00000000ffffffe7fffffffffffffff5ffffffff0000003e00000000",
            INIT_46 => X"0000010a000000000000008e00000000ffffff7affffffff0000008a00000000",
            INIT_47 => X"ffffffeaffffffffffffffd3fffffffffffffff7ffffffff0000005000000000",
            INIT_48 => X"ffffffbeffffffff0000001000000000ffffffa9ffffffffffffffc0ffffffff",
            INIT_49 => X"ffffffeaffffffff0000004b000000000000001900000000ffffff8dffffffff",
            INIT_4A => X"0000008400000000000000470000000000000124000000000000000300000000",
            INIT_4B => X"ffffffbbffffffffffffffa6ffffffff00000030000000000000004d00000000",
            INIT_4C => X"ffffffceffffffffffffff9bffffffff0000005a00000000ffffff6affffffff",
            INIT_4D => X"000000cb00000000ffffff97ffffffff00000043000000000000006e00000000",
            INIT_4E => X"00000014000000000000003100000000ffffffdaffffffff0000001e00000000",
            INIT_4F => X"0000001200000000ffffff81ffffffff0000001800000000fffffff7ffffffff",
            INIT_50 => X"ffffffdcffffffff0000002d00000000000000a3000000000000000f00000000",
            INIT_51 => X"0000008100000000000000130000000000000067000000000000006b00000000",
            INIT_52 => X"ffffff63ffffffff0000001e00000000ffffff4cffffffff0000007000000000",
            INIT_53 => X"ffffffe6ffffffff0000006200000000ffffffb2ffffffff0000004d00000000",
            INIT_54 => X"0000000b0000000000000090000000000000001200000000ffffff7bffffffff",
            INIT_55 => X"0000001e0000000000000081000000000000003300000000ffffff79ffffffff",
            INIT_56 => X"0000000f00000000fffffff1fffffffffffffff5fffffffffffffff8ffffffff",
            INIT_57 => X"0000011d000000000000001800000000ffffff95ffffffff000000b600000000",
            INIT_58 => X"ffffffc6ffffffff0000006d000000000000000c000000000000002500000000",
            INIT_59 => X"000000060000000000000015000000000000005000000000fffffff6ffffffff",
            INIT_5A => X"ffffffe2ffffffffffffff91ffffffff0000006f000000000000005000000000",
            INIT_5B => X"ffffffd3ffffffff000000af00000000fffffffcffffffff0000007400000000",
            INIT_5C => X"0000002700000000ffffff68ffffffffffffffd2ffffffff0000006d00000000",
            INIT_5D => X"ffffff97ffffffff0000000b00000000ffffff97ffffffff0000003800000000",
            INIT_5E => X"0000008f00000000ffffff69ffffffff00000061000000000000006500000000",
            INIT_5F => X"ffffff4effffffffffffff8effffffff0000004a00000000ffffffa6ffffffff",
            INIT_60 => X"ffffffe8ffffffff00000076000000000000001800000000ffffffe9ffffffff",
            INIT_61 => X"ffffffebffffffff000000a3000000000000008000000000ffffffe6ffffffff",
            INIT_62 => X"ffffff09ffffffff0000005700000000ffffffd6ffffffffffffff39ffffffff",
            INIT_63 => X"ffffffc6ffffffff00000046000000000000004b00000000ffffff6affffffff",
            INIT_64 => X"0000000a0000000000000070000000000000002c000000000000003200000000",
            INIT_65 => X"0000003d0000000000000055000000000000000800000000ffffffe8ffffffff",
            INIT_66 => X"ffffff8affffffff00000006000000000000003f000000000000006900000000",
            INIT_67 => X"ffffff75ffffffffffffffc4ffffffff0000007b000000000000001000000000",
            INIT_68 => X"ffffff39ffffffff0000004900000000000000d1000000000000000900000000",
            INIT_69 => X"00000048000000000000000500000000ffffff37ffffffffffffffe9ffffffff",
            INIT_6A => X"0000008f000000000000000500000000ffffff86ffffffff0000008800000000",
            INIT_6B => X"ffffffefffffffffffffff66ffffffffffffffe8ffffffff0000006400000000",
            INIT_6C => X"0000003100000000ffffff97ffffffffffffffdcffffffff0000005c00000000",
            INIT_6D => X"fffffff3ffffffff00000006000000000000000000000000fffffffbffffffff",
            INIT_6E => X"fffffff2fffffffffffffff4fffffffffffffff3ffffffff0000000700000000",
            INIT_6F => X"ffffffe4ffffffff00000015000000000000001300000000fffffff7ffffffff",
            INIT_70 => X"0000000d0000000000000023000000000000006500000000fffffff5ffffffff",
            INIT_71 => X"0000004400000000ffffffddffffffff0000006600000000ffffffb7ffffffff",
            INIT_72 => X"ffffffd6ffffffffffffffa0ffffffff0000006500000000ffffff91ffffffff",
            INIT_73 => X"ffffffeaffffffffffffff38ffffffffffffff4bffffffff0000005a00000000",
            INIT_74 => X"ffffff78ffffffff000000000000000000000039000000000000008600000000",
            INIT_75 => X"0000008d00000000ffffffefffffffffffffffdfffffffff0000000900000000",
            INIT_76 => X"0000001f00000000ffffff21fffffffffffffca5ffffffff0000009d00000000",
            INIT_77 => X"ffffffa4ffffffff0000007100000000ffffffffffffffff0000006e00000000",
            INIT_78 => X"0000000000000000ffffffbbffffffffffffffa7ffffffff0000012a00000000",
            INIT_79 => X"0000006400000000ffffff8bffffffffffffff8cffffffff0000000b00000000",
            INIT_7A => X"ffffff9dffffffffffffffebffffffffffffffb3ffffffff0000009700000000",
            INIT_7B => X"ffffff50ffffffffffffffe6ffffffff000000cc000000000000002e00000000",
            INIT_7C => X"ffffffb3ffffffff0000002800000000ffffff65ffffffff0000007d00000000",
            INIT_7D => X"ffffffd4ffffffffffffffe9ffffffffffffffe0ffffffff0000006500000000",
            INIT_7E => X"ffffffe3ffffffffffffffbeffffffff0000000f000000000000002f00000000",
            INIT_7F => X"ffffff45ffffffffffffff58ffffffff000000ec000000000000008e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE4;


    MEM_IWGHT_LAYER2_INSTANCE5 : if BRAM_NAME = "iwght_layer2_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffee4ffffffffffffffabffffffff0000003100000000ffffff40ffffffff",
            INIT_01 => X"000000cd00000000ffffff38ffffffffffffff77ffffffff0000002b00000000",
            INIT_02 => X"ffffffd3ffffffff0000002b000000000000006400000000fffffffeffffffff",
            INIT_03 => X"ffffffa9ffffffffffffffa4ffffffffffffffdfffffffff0000007500000000",
            INIT_04 => X"0000000c000000000000007c00000000ffffff50ffffffffffffff74ffffffff",
            INIT_05 => X"00000080000000000000007300000000ffffffd4ffffffff0000004100000000",
            INIT_06 => X"000000aa000000000000000f00000000ffffffb0ffffffff000000c400000000",
            INIT_07 => X"0000001d000000000000002100000000ffffffc7ffffffff0000001400000000",
            INIT_08 => X"ffffffeeffffffff0000008100000000ffffffabffffffff0000006d00000000",
            INIT_09 => X"ffffff24ffffffffffffff4dffffffff00000039000000000000002600000000",
            INIT_0A => X"00000016000000000000004b00000000fffffff0ffffffffffffffe2ffffffff",
            INIT_0B => X"ffffff92ffffffffffffffeeffffffff0000005f000000000000004500000000",
            INIT_0C => X"ffffffd4ffffffffffffff2affffffff0000000b000000000000008600000000",
            INIT_0D => X"00000025000000000000002200000000ffffffa7fffffffffffffff4ffffffff",
            INIT_0E => X"000000d700000000000000ce00000000000000a3000000000000001f00000000",
            INIT_0F => X"fffffef5ffffffff0000004100000000ffffff2bffffffff0000010400000000",
            INIT_10 => X"ffffffb3ffffffffffffff93ffffffff0000000f000000000000002c00000000",
            INIT_11 => X"ffffff96fffffffffffffedcffffffffffffff6dffffffff0000002500000000",
            INIT_12 => X"ffffff56ffffffffffffff69ffffffff00000008000000000000003000000000",
            INIT_13 => X"00000006000000000000000d000000000000000c00000000ffffffe2ffffffff",
            INIT_14 => X"ffffffedfffffffffffffff0fffffffffffffe1affffffff0000001600000000",
            INIT_15 => X"ffffffbeffffffff0000002600000000ffffff05ffffffffffffffb4ffffffff",
            INIT_16 => X"ffffffa4ffffffffffffff3dffffffffffffffd4ffffffffffffff48ffffffff",
            INIT_17 => X"000000e3000000000000002200000000ffffff39ffffffff000000ed00000000",
            INIT_18 => X"0000007000000000ffffffe2ffffffffffffffefffffffff000000a500000000",
            INIT_19 => X"0000003b0000000000000088000000000000001100000000fffffff4ffffffff",
            INIT_1A => X"ffffffe9ffffffffffffffaaffffffffffffff72ffffffff0000002900000000",
            INIT_1B => X"ffffff60ffffffff0000006000000000ffffffc9ffffffff0000006300000000",
            INIT_1C => X"0000006600000000ffffff82ffffffff00000081000000000000006400000000",
            INIT_1D => X"ffffffa0ffffffff0000003c000000000000005a00000000000000b800000000",
            INIT_1E => X"ffffffa9ffffffffffffffaeffffffff0000007b00000000ffffff1cffffffff",
            INIT_1F => X"ffffffd0fffffffffffffe6dffffffff0000001100000000ffffff78ffffffff",
            INIT_20 => X"000000b000000000ffffffbcffffffffffffffc2ffffffff0000001b00000000",
            INIT_21 => X"0000004e00000000ffffffe6ffffffff0000005900000000ffffff88ffffffff",
            INIT_22 => X"ffffffaaffffffff0000002900000000fffffff6ffffffffffffffc7ffffffff",
            INIT_23 => X"ffffffc2ffffffffffffffcbffffffff000000a800000000ffffff24ffffffff",
            INIT_24 => X"00000017000000000000005400000000ffffffefffffffffffffffeeffffffff",
            INIT_25 => X"ffffffbcffffffffffffffe5ffffffff000000c000000000ffffffb3ffffffff",
            INIT_26 => X"000000aa00000000ffffff6effffffff0000004400000000ffffffd9ffffffff",
            INIT_27 => X"ffffff74ffffffffffffff9afffffffffffffff2ffffffff0000000b00000000",
            INIT_28 => X"ffffff8bfffffffffffffeceffffffffffffffbcffffffffffffffc4ffffffff",
            INIT_29 => X"000000e2000000000000003e00000000ffffff4bffffffffffffff82ffffffff",
            INIT_2A => X"0000008a00000000ffffff94ffffffff0000000000000000000000b200000000",
            INIT_2B => X"0000001500000000ffffffb0ffffffff0000001f000000000000004600000000",
            INIT_2C => X"fffffee8ffffffff0000006a000000000000007e00000000ffffff9fffffffff",
            INIT_2D => X"0000002a00000000ffffffc9fffffffffffffffdffffffffffffff8fffffffff",
            INIT_2E => X"000000400000000000000008000000000000004c000000000000001a00000000",
            INIT_2F => X"ffffff76ffffffffffffff6cffffffffffffff65ffffffff0000004c00000000",
            INIT_30 => X"ffffff93fffffffffffffffbffffffffffffff8effffffffffffff89ffffffff",
            INIT_31 => X"ffffff20ffffffffffffff0cffffffff0000001d00000000ffffff96ffffffff",
            INIT_32 => X"00000004000000000000006500000000ffffff40ffffffff0000008000000000",
            INIT_33 => X"0000007800000000fffffff2ffffffff000000bb000000000000003d00000000",
            INIT_34 => X"ffffffaeffffffffffffff36ffffffffffffff91ffffffffffffffbdffffffff",
            INIT_35 => X"ffffffeffffffffffffffff9ffffffff0000000400000000ffffffd7ffffffff",
            INIT_36 => X"fffffff1fffffffffffffff1fffffffffffffff9ffffffff0000000100000000",
            INIT_37 => X"0000003200000000000000340000000000000000000000000000000900000000",
            INIT_38 => X"0000000700000000ffffff7dffffffff0000005300000000fffffff5ffffffff",
            INIT_39 => X"ffffff8dffffffffffffffa0ffffffff00000027000000000000006100000000",
            INIT_3A => X"ffffffe0fffffffffffffff6ffffffffffffff20ffffffffffffff49ffffffff",
            INIT_3B => X"00000029000000000000001a00000000ffffff4cffffffffffffffafffffffff",
            INIT_3C => X"00000035000000000000005600000000000000b700000000ffffffbfffffffff",
            INIT_3D => X"ffffffdeffffffff00000001000000000000004b00000000ffffff56ffffffff",
            INIT_3E => X"ffffff69fffffffffffffffafffffffffffffdd3ffffffff0000002700000000",
            INIT_3F => X"fffffecdffffffff0000003200000000000000aa00000000ffffff6cffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a1000000000000005200000000000000d2000000000000004f00000000",
            INIT_41 => X"ffffffd9ffffffff0000003e000000000000001d00000000000000b800000000",
            INIT_42 => X"ffffffbbffffffff0000003d00000000ffffff46ffffffffffffffbbffffffff",
            INIT_43 => X"0000008d00000000ffffff69ffffffffffffffceffffffffffffffd7ffffffff",
            INIT_44 => X"ffffff55ffffffffffffffaaffffffffffffff0bffffffff0000000d00000000",
            INIT_45 => X"000000c8000000000000005800000000ffffffddffffffffffffff70ffffffff",
            INIT_46 => X"0000003a00000000ffffff9affffffffffffffe3ffffffff0000006300000000",
            INIT_47 => X"000000ff00000000ffffff8fffffffffffffff9dffffffffffffffabffffffff",
            INIT_48 => X"ffffffbdffffffff0000004100000000ffffff62ffffffff000000a400000000",
            INIT_49 => X"00000095000000000000003a0000000000000026000000000000006d00000000",
            INIT_4A => X"00000010000000000000000e00000000ffffff68ffffffff0000009900000000",
            INIT_4B => X"000000bf00000000ffffff3fffffffff0000004c00000000fffffef2ffffffff",
            INIT_4C => X"ffffffd7ffffffffffffffa0ffffffffffffffd4ffffffff0000004700000000",
            INIT_4D => X"000000a8000000000000007d0000000000000048000000000000003200000000",
            INIT_4E => X"ffffffc5ffffffffffffff2fffffffffffffff05ffffffff0000001d00000000",
            INIT_4F => X"ffffff9bffffffff00000062000000000000000100000000ffffff78ffffffff",
            INIT_50 => X"000000110000000000000073000000000000001600000000000000a300000000",
            INIT_51 => X"ffffff4bffffffff0000000500000000000000a0000000000000007000000000",
            INIT_52 => X"0000008100000000000000dd0000000000000095000000000000005b00000000",
            INIT_53 => X"0000001d000000000000006d00000000ffffffdfffffffff0000001e00000000",
            INIT_54 => X"0000007b00000000ffffffeeffffffffffffffc7fffffffffffffff0ffffffff",
            INIT_55 => X"ffffffa4ffffffff0000000c00000000ffffffb2fffffffffffffff9ffffffff",
            INIT_56 => X"0000005a000000000000001a0000000000000030000000000000001900000000",
            INIT_57 => X"ffffff5fffffffffffffff53ffffffffffffff25ffffffffffffffe9ffffffff",
            INIT_58 => X"fffffff9ffffffff000000740000000000000032000000000000006300000000",
            INIT_59 => X"0000004900000000ffffffe9ffffffff0000006e00000000ffffffe2ffffffff",
            INIT_5A => X"0000003e0000000000000099000000000000006700000000ffffff8effffffff",
            INIT_5B => X"ffffffc7ffffffffffffff60ffffffffffffffc4ffffffffffffff40ffffffff",
            INIT_5C => X"0000000500000000ffffff47ffffffff000000a9000000000000008100000000",
            INIT_5D => X"0000004c0000000000000008000000000000014700000000ffffffb0ffffffff",
            INIT_5E => X"ffffffb9ffffffff00000007000000000000002b00000000ffffffb1ffffffff",
            INIT_5F => X"000000220000000000000020000000000000003000000000ffffffb7ffffffff",
            INIT_60 => X"0000004c00000000ffffffdfffffffffffffff26ffffffff0000004500000000",
            INIT_61 => X"000000b5000000000000004400000000ffffffe2ffffffffffffff9cffffffff",
            INIT_62 => X"0000005d00000000ffffff8dffffffffffffff84ffffffffffffff69ffffffff",
            INIT_63 => X"ffffffc3ffffffff0000002800000000ffffffeaffffffffffffffe3ffffffff",
            INIT_64 => X"ffffffb7ffffffff0000003800000000ffffffe5ffffffffffffff86ffffffff",
            INIT_65 => X"00000140000000000000008900000000ffffff03ffffffff0000006100000000",
            INIT_66 => X"0000003000000000fffffd5fffffffff0000007900000000000000c800000000",
            INIT_67 => X"0000009100000000ffffffa0ffffffffffffffeaffffffff0000009400000000",
            INIT_68 => X"ffffff75ffffffffffffff7bffffffffffffffa7ffffffff0000005600000000",
            INIT_69 => X"0000001600000000ffffffe0ffffffff0000005400000000ffffff47ffffffff",
            INIT_6A => X"0000005a00000000fffffff3ffffffff0000001a00000000ffffff23ffffffff",
            INIT_6B => X"000000c00000000000000099000000000000005e00000000ffffff86ffffffff",
            INIT_6C => X"fffffeeaffffffff00000058000000000000003600000000ffffff49ffffffff",
            INIT_6D => X"0000002e000000000000005500000000fffffe8ffffffffffffffef4ffffffff",
            INIT_6E => X"ffffff1affffffffffffffc8ffffffffffffffedffffffff0000005c00000000",
            INIT_6F => X"ffffff95ffffffffffffff6dffffffffffffff88ffffffff0000009100000000",
            INIT_70 => X"ffffffe1ffffffffffffff4cfffffffffffffec5ffffffff000000b000000000",
            INIT_71 => X"0000003900000000ffffffe4ffffffffffffff8affffffff0000008400000000",
            INIT_72 => X"ffffffc0ffffffffffffffc6ffffffff0000008300000000ffffff81ffffffff",
            INIT_73 => X"ffffff1cffffffffffffff69ffffffffffffffbbffffffff0000002b00000000",
            INIT_74 => X"0000001900000000fffffff9fffffffffffffed4ffffffff0000002900000000",
            INIT_75 => X"ffffffc5ffffffff00000009000000000000006500000000ffffffefffffffff",
            INIT_76 => X"ffffff96ffffffffffffffd7ffffffff0000006b00000000000000be00000000",
            INIT_77 => X"ffffff59ffffffffffffffffffffffff0000009f00000000ffffff2dffffffff",
            INIT_78 => X"0000002c00000000ffffffdeffffffff0000001b000000000000000400000000",
            INIT_79 => X"ffffffe3ffffffffffffff7effffffffffffffd2ffffffff0000004f00000000",
            INIT_7A => X"0000006400000000ffffffa3ffffffffffffff87ffffffffffffffadffffffff",
            INIT_7B => X"000000b100000000fffffff3ffffffff0000000700000000ffffff87ffffffff",
            INIT_7C => X"00000044000000000000004100000000ffffff9affffffff0000008200000000",
            INIT_7D => X"0000000000000000fffffff6fffffffffffffffbffffffffffffff2bffffffff",
            INIT_7E => X"ffffffedfffffffffffffff1ffffffff00000001000000000000000400000000",
            INIT_7F => X"fffffef5fffffffffffffff3fffffffffffffff5ffffffff0000001300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE5;


    MEM_IWGHT_LAYER2_INSTANCE6 : if BRAM_NAME = "iwght_layer2_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffcdffffffffffffffa5ffffffff0000007e00000000fffffff9ffffffff",
            INIT_01 => X"0000002b00000000ffffff98ffffffff000000a500000000ffffff1effffffff",
            INIT_02 => X"ffffff2fffffffffffffffa9ffffffff0000006400000000ffffff58ffffffff",
            INIT_03 => X"fffffff3ffffffff00000047000000000000003e000000000000008300000000",
            INIT_04 => X"ffffffcbffffffff000000220000000000000040000000000000002d00000000",
            INIT_05 => X"ffffff4bffffffffffffff16ffffffffffffff0effffffffffffffa3ffffffff",
            INIT_06 => X"00000104000000000000007000000000ffffff87ffffffff000000bd00000000",
            INIT_07 => X"0000003d000000000000004200000000ffffffa7ffffffff0000015200000000",
            INIT_08 => X"fffffff8ffffffffffffffd6fffffffffffffeeafffffffffffffffbffffffff",
            INIT_09 => X"000000db0000000000000039000000000000018200000000fffffefcffffffff",
            INIT_0A => X"ffffff8bfffffffffffffebafffffffffffffe1fffffffff000000b500000000",
            INIT_0B => X"ffffffa6ffffffffffffffadfffffffffffffff0ffffffff0000001100000000",
            INIT_0C => X"ffffff52fffffffffffffeb2ffffffff000000cf00000000ffffffb6ffffffff",
            INIT_0D => X"ffffffd3ffffffff000000020000000000000077000000000000003400000000",
            INIT_0E => X"ffffff57ffffffff0000004f00000000ffffffedffffffff0000001b00000000",
            INIT_0F => X"fffffff2ffffffffffffffcffffffffffffffed5ffffffff0000006700000000",
            INIT_10 => X"fffffe1dffffffff00000051000000000000007100000000fffffffaffffffff",
            INIT_11 => X"0000009b0000000000000121000000000000000200000000ffffffdbffffffff",
            INIT_12 => X"0000004c000000000000007100000000000000b6000000000000008000000000",
            INIT_13 => X"0000002d000000000000004100000000ffffff8cffffffff000000be00000000",
            INIT_14 => X"fffffecbffffffff0000004d000000000000012500000000ffffff94ffffffff",
            INIT_15 => X"fffffeb1ffffffff000000c000000000ffffff9fffffffffffffffc4ffffffff",
            INIT_16 => X"ffffffa6ffffffffffffff92ffffffffffffffe0ffffffffffffff5affffffff",
            INIT_17 => X"fffffe74ffffffff000000c200000000fffffee2ffffffffffffff1effffffff",
            INIT_18 => X"ffffff73ffffffff0000005e000000000000002000000000ffffffb5ffffffff",
            INIT_19 => X"00000029000000000000004f00000000ffffff9affffffff0000007b00000000",
            INIT_1A => X"ffffff19fffffffffffffff0ffffffffffffff1efffffffffffffc89ffffffff",
            INIT_1B => X"00000068000000000000000d00000000ffffffd2ffffffff0000000000000000",
            INIT_1C => X"0000003500000000ffffffcbffffffff00000003000000000000005700000000",
            INIT_1D => X"0000000200000000ffffff8effffffff0000009f000000000000003900000000",
            INIT_1E => X"0000002900000000ffffffe1ffffffff000000ac00000000ffffffe4ffffffff",
            INIT_1F => X"000000c0000000000000009800000000ffffffd4fffffffffffffe89ffffffff",
            INIT_20 => X"ffffff60ffffffff000000630000000000000117000000000000007900000000",
            INIT_21 => X"0000002400000000ffffffa2ffffffff000000d1000000000000003f00000000",
            INIT_22 => X"ffffff70ffffffffffffffb7fffffffffffffff8ffffffffffffffe3ffffffff",
            INIT_23 => X"ffffffb6ffffffff000000d0000000000000002b000000000000004a00000000",
            INIT_24 => X"ffffff67ffffffffffffffbeffffffff0000001200000000ffffffd3ffffffff",
            INIT_25 => X"ffffffc8ffffffff0000003b00000000ffffffe8ffffffffffffffe6ffffffff",
            INIT_26 => X"000000de000000000000000000000000ffffffc5ffffffff0000001f00000000",
            INIT_27 => X"0000005a00000000ffffff9affffffffffffffd6ffffffffffffff7cffffffff",
            INIT_28 => X"0000008f000000000000001100000000ffffffdfffffffff0000005e00000000",
            INIT_29 => X"ffffff7bffffffff0000001a0000000000000028000000000000006d00000000",
            INIT_2A => X"ffffffbdfffffffffffffffcffffffff00000001000000000000000100000000",
            INIT_2B => X"000000fe000000000000001e00000000fffffff3ffffffffffffffc0ffffffff",
            INIT_2C => X"000000b60000000000000024000000000000007100000000ffffff37ffffffff",
            INIT_2D => X"0000004f00000000ffffff1fffffffffffffff34ffffffff0000002600000000",
            INIT_2E => X"ffffff54ffffffff0000003400000000ffffff02ffffffffffffff82ffffffff",
            INIT_2F => X"ffffffcbffffffff0000006b00000000fffffff5ffffffffffffffc1ffffffff",
            INIT_30 => X"0000003900000000ffffffedffffffffffffffc1ffffffffffffff93ffffffff",
            INIT_31 => X"0000000200000000ffffffffffffffffffffffb0ffffffffffffffecffffffff",
            INIT_32 => X"0000004200000000fffffffbffffffff00000024000000000000001200000000",
            INIT_33 => X"ffffffd9ffffffff0000007d000000000000000e00000000ffffff9cffffffff",
            INIT_34 => X"ffffffcbffffffff0000001e000000000000003500000000ffffffcbffffffff",
            INIT_35 => X"ffffffb4ffffffffffffff63ffffffff0000005600000000ffffff9affffffff",
            INIT_36 => X"ffffffe7ffffffffffffff9cffffffffffffffcbffffffffffffffa5ffffffff",
            INIT_37 => X"ffffffe3ffffffffffffffc3ffffffffffffff93ffffffff0000000b00000000",
            INIT_38 => X"00000096000000000000001d00000000ffffff9ffffffffffffffff0ffffffff",
            INIT_39 => X"ffffffd9ffffffff0000003d00000000ffffff54ffffffff0000000e00000000",
            INIT_3A => X"fffffff1fffffffffffffffdffffffff00000020000000000000006f00000000",
            INIT_3B => X"fffffffeffffffff000000130000000000000039000000000000003100000000",
            INIT_3C => X"0000003c0000000000000048000000000000002d000000000000001900000000",
            INIT_3D => X"ffffffbbffffffffffffff6bffffffff0000005d000000000000003100000000",
            INIT_3E => X"000000e2000000000000004300000000ffffffcdffffffffffffffd2ffffffff",
            INIT_3F => X"ffffffe3ffffffff000000ae0000000000000046000000000000005b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d4000000000000002700000000ffffff8cffffffffffffff5affffffff",
            INIT_41 => X"fffffff9ffffffff0000004400000000fffffff3ffffffffffffff5affffffff",
            INIT_42 => X"ffffff8bffffffffffffffe1fffffffffffffff2ffffffffffffffa5ffffffff",
            INIT_43 => X"ffffffc9ffffffff00000016000000000000004b00000000ffffffc6ffffffff",
            INIT_44 => X"fffffff8ffffffff00000008000000000000001500000000ffffffa8ffffffff",
            INIT_45 => X"00000000000000000000000b00000000fffffffaffffffff0000005200000000",
            INIT_46 => X"fffffff3fffffffffffffff2ffffffff00000012000000000000000900000000",
            INIT_47 => X"0000009a000000000000004b00000000fffffff7ffffffff0000000c00000000",
            INIT_48 => X"00000003000000000000000a0000000000000009000000000000001100000000",
            INIT_49 => X"ffffff89ffffffffffffff7fffffffff0000001700000000ffffff9bffffffff",
            INIT_4A => X"ffffffd7ffffffff0000004900000000000000ad00000000ffffffceffffffff",
            INIT_4B => X"ffffff75ffffffff00000060000000000000002300000000ffffffb3ffffffff",
            INIT_4C => X"ffffffadffffffff0000002e000000000000005500000000ffffffb4ffffffff",
            INIT_4D => X"fffffedbffffffffffffff0bfffffffffffffeefffffffffffffffaeffffffff",
            INIT_4E => X"0000001800000000fffffff3ffffffff0000003200000000ffffff9dffffffff",
            INIT_4F => X"00000018000000000000013d000000000000000700000000ffffffd9ffffffff",
            INIT_50 => X"0000003600000000ffffffc7ffffffff0000005300000000ffffffcfffffffff",
            INIT_51 => X"ffffffe1ffffffff0000001c00000000ffffffd4ffffffffffffffdaffffffff",
            INIT_52 => X"ffffff5cffffffff000000440000000000000045000000000000002400000000",
            INIT_53 => X"ffffffb0ffffffffffffff2cffffffffffffff75ffffffff0000003d00000000",
            INIT_54 => X"0000000100000000ffffff41ffffffffffffff7bffffffffffffff1fffffffff",
            INIT_55 => X"ffffffdaffffffffffffff9effffffffffffffc3ffffffffffffff96ffffffff",
            INIT_56 => X"000000070000000000000045000000000000007800000000ffffffb0ffffffff",
            INIT_57 => X"0000006300000000ffffff79ffffffff0000003400000000ffffff49ffffffff",
            INIT_58 => X"0000004e000000000000003700000000ffffff84ffffffff0000002500000000",
            INIT_59 => X"0000002e000000000000000c00000000ffffffc7ffffffffffffffadffffffff",
            INIT_5A => X"fffffff4ffffffffffffffb3ffffffff0000005d000000000000000300000000",
            INIT_5B => X"0000008a000000000000002c00000000000000c700000000000000a000000000",
            INIT_5C => X"00000032000000000000000e000000000000001100000000ffffffa0ffffffff",
            INIT_5D => X"ffffffbcffffffff0000002f0000000000000060000000000000001b00000000",
            INIT_5E => X"0000005900000000ffffff8effffffffffffffeeffffffffffffffcaffffffff",
            INIT_5F => X"0000001800000000ffffffccffffffffffffffdcffffffff000000c400000000",
            INIT_60 => X"ffffffe1ffffffff000000210000000000000022000000000000005f00000000",
            INIT_61 => X"000000a300000000ffffffebffffffffffffffa2ffffffffffffff84ffffffff",
            INIT_62 => X"0000008e00000000ffffffadfffffffffffffff5ffffffffffffff49ffffffff",
            INIT_63 => X"ffffffadffffffffffffff33ffffffffffffffe7ffffffff0000001700000000",
            INIT_64 => X"0000001c00000000ffffffd7ffffffffffffffb4ffffffffffffffaeffffffff",
            INIT_65 => X"0000006600000000000000250000000000000076000000000000006e00000000",
            INIT_66 => X"ffffffc3ffffffff0000000000000000fffffff2ffffffff000000ba00000000",
            INIT_67 => X"fffffff6ffffffffffffffe0ffffffffffffffc6ffffffffffffff7affffffff",
            INIT_68 => X"ffffff81ffffffff000000120000000000000046000000000000005000000000",
            INIT_69 => X"0000001a000000000000002b00000000ffffffd6ffffffff0000003100000000",
            INIT_6A => X"ffffffc7ffffffffffffffe9ffffffffffffffa3fffffffffffffefdffffffff",
            INIT_6B => X"ffffffa7ffffffff0000008200000000ffffffe6ffffffff0000005e00000000",
            INIT_6C => X"00000042000000000000005b000000000000003c00000000fffffff6ffffffff",
            INIT_6D => X"ffffffd9ffffffffffffffd8ffffffffffffffdeffffffff0000004500000000",
            INIT_6E => X"ffffffbeffffffffffffffe5ffffffffffffffa7ffffffffffffffb2ffffffff",
            INIT_6F => X"fffffff1ffffffff00000054000000000000006b000000000000008800000000",
            INIT_70 => X"0000004000000000ffffffaaffffffff00000026000000000000008300000000",
            INIT_71 => X"00000070000000000000000b00000000ffffffd8ffffffff0000004600000000",
            INIT_72 => X"000000a6000000000000004100000000ffffff38ffffffff0000009400000000",
            INIT_73 => X"0000001200000000fffffff5fffffffffffffffeffffffffffffff78ffffffff",
            INIT_74 => X"ffffff99ffffffffffffff6affffffffffffffb7ffffffff0000003c00000000",
            INIT_75 => X"ffffff96ffffffffffffff90ffffffff00000068000000000000004d00000000",
            INIT_76 => X"0000002c00000000ffffffa0ffffffffffffff97ffffffffffffffd7ffffffff",
            INIT_77 => X"ffffffe7ffffffff0000002100000000ffffffe3ffffffff0000005400000000",
            INIT_78 => X"0000005f00000000fffffff2ffffffffffffff35ffffffffffffffadffffffff",
            INIT_79 => X"00000025000000000000001c0000000000000065000000000000000200000000",
            INIT_7A => X"0000002f0000000000000070000000000000001f00000000ffffffd1ffffffff",
            INIT_7B => X"ffffffe8ffffffffffffffc6ffffffff00000019000000000000007000000000",
            INIT_7C => X"fffffff2ffffffff000000aa00000000fffffffeffffffffffffffc2ffffffff",
            INIT_7D => X"ffffffe6fffffffffffffef6ffffffff0000007a00000000ffffff87ffffffff",
            INIT_7E => X"ffffff79fffffffffffffeffffffffffffffff9cffffffff0000001e00000000",
            INIT_7F => X"ffffffcbffffffffffffff20ffffffffffffff9affffffffffffffbbffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE6;


    MEM_IWGHT_LAYER2_INSTANCE7 : if BRAM_NAME = "iwght_layer2_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000c200000000ffffffa9ffffffff0000002d000000000000006500000000",
            INIT_01 => X"fffffff8ffffffffffffffebffffffff0000006200000000fffffff2ffffffff",
            INIT_02 => X"0000004e00000000ffffffa1ffffffffffffffbfffffffffffffffe5ffffffff",
            INIT_03 => X"ffffffd8ffffffff0000000a00000000ffffff37ffffffffffffffc9ffffffff",
            INIT_04 => X"ffffffd3ffffffff0000002f00000000000000de000000000000007900000000",
            INIT_05 => X"0000001f0000000000000003000000000000006b00000000000000a400000000",
            INIT_06 => X"00000017000000000000006800000000ffffffb2ffffffffffffffeaffffffff",
            INIT_07 => X"ffffff8ffffffffffffffffaffffffffffffffa6ffffffffffffffddffffffff",
            INIT_08 => X"ffffffa8ffffffffffffffecffffffffffffffe5ffffffff0000001700000000",
            INIT_09 => X"ffffff74ffffffff00000055000000000000005600000000ffffff0dffffffff",
            INIT_0A => X"00000001000000000000004200000000fffffff0ffffffffffffff5dffffffff",
            INIT_0B => X"ffffffcfffffffffffffffdffffffffffffffee5ffffffffffffffcbffffffff",
            INIT_0C => X"000000400000000000000024000000000000004500000000000000a400000000",
            INIT_0D => X"0000000300000000fffffff8ffffffff00000003000000000000007f00000000",
            INIT_0E => X"00000006000000000000001000000000fffffffdffffffff0000001a00000000",
            INIT_0F => X"0000006f000000000000000900000000fffffffaffffffffffffffebffffffff",
            INIT_10 => X"0000000c00000000fffffff6ffffffff0000008200000000ffffffc2ffffffff",
            INIT_11 => X"00000054000000000000007b000000000000003700000000ffffffb8ffffffff",
            INIT_12 => X"ffffffccffffffff0000004700000000ffffff92ffffffffffffffffffffffff",
            INIT_13 => X"0000006800000000ffffffb5ffffffff00000085000000000000007600000000",
            INIT_14 => X"0000004a00000000ffffffc8ffffffff0000000e00000000ffffffd8ffffffff",
            INIT_15 => X"0000004c000000000000000a000000000000003400000000ffffffffffffffff",
            INIT_16 => X"000000b600000000ffffffaaffffffffffffff7affffffffffffffddffffffff",
            INIT_17 => X"000000b6000000000000001500000000ffffffe0ffffffffffffff26ffffffff",
            INIT_18 => X"ffffff82ffffffff0000002700000000000000e900000000ffffff67ffffffff",
            INIT_19 => X"ffffffd0ffffffffffffffe2ffffffffffffffd1ffffffff0000004500000000",
            INIT_1A => X"ffffffc9ffffffff000000a600000000ffffffecffffffff0000004600000000",
            INIT_1B => X"ffffffd5ffffffff0000001c000000000000003c00000000fffffffdffffffff",
            INIT_1C => X"ffffff51ffffffffffffffebffffffff0000001c000000000000006700000000",
            INIT_1D => X"ffffffc6ffffffff00000036000000000000001700000000000000e900000000",
            INIT_1E => X"ffffff11ffffffffffffffa0ffffffffffffff95ffffffffffffffcbffffffff",
            INIT_1F => X"0000003600000000ffffff9dffffffff00000033000000000000008000000000",
            INIT_20 => X"00000091000000000000003c000000000000000000000000fffffffcffffffff",
            INIT_21 => X"0000001d00000000ffffffccffffffff0000000c00000000ffffffc4ffffffff",
            INIT_22 => X"0000006200000000ffffffdcffffffff0000004600000000ffffffeaffffffff",
            INIT_23 => X"0000009f00000000ffffff50ffffffff0000004f000000000000005500000000",
            INIT_24 => X"ffffffedffffffffffffff9cffffffff0000000400000000ffffffa9ffffffff",
            INIT_25 => X"00000109000000000000003f000000000000004200000000ffffffefffffffff",
            INIT_26 => X"ffffff3fffffffff0000008f00000000ffffff63fffffffffffffffcffffffff",
            INIT_27 => X"ffffff84ffffffffffffff65ffffffff0000003300000000ffffffd7ffffffff",
            INIT_28 => X"00000059000000000000002e000000000000009200000000ffffffc4ffffffff",
            INIT_29 => X"0000006400000000000000050000000000000077000000000000001800000000",
            INIT_2A => X"0000001f00000000ffffff86ffffffffffffffcdffffffff0000002600000000",
            INIT_2B => X"0000004900000000fffffff0ffffffffffffff36ffffffff000000f900000000",
            INIT_2C => X"ffffffd4ffffffffffffffb2fffffffffffffff3ffffffff0000005c00000000",
            INIT_2D => X"0000004000000000ffffff77ffffffffffffff85ffffffffffffffc2ffffffff",
            INIT_2E => X"0000005c00000000ffffffb3ffffffffffffff40ffffffff0000004e00000000",
            INIT_2F => X"ffffffbfffffffff000000aa00000000ffffff52ffffffffffffff6cffffffff",
            INIT_30 => X"00000029000000000000002e0000000000000043000000000000003b00000000",
            INIT_31 => X"00000082000000000000004c00000000ffffff69ffffffffffffff3fffffffff",
            INIT_32 => X"000000cf000000000000001400000000fffffffcffffffffffffffc9ffffffff",
            INIT_33 => X"ffffff8dffffffff000000360000000000000026000000000000008700000000",
            INIT_34 => X"00000071000000000000000900000000ffffffe4ffffffffffffffc7ffffffff",
            INIT_35 => X"0000003400000000ffffff7effffffff0000001300000000ffffff41ffffffff",
            INIT_36 => X"fffffff2ffffffffffffffe2ffffffff0000006800000000ffffff4bffffffff",
            INIT_37 => X"000000180000000000000087000000000000008700000000ffffff9bffffffff",
            INIT_38 => X"000000c800000000ffffffe1ffffffff0000001300000000ffffffceffffffff",
            INIT_39 => X"fffffff3ffffffff0000000000000000ffffffadfffffffffffffff7ffffffff",
            INIT_3A => X"0000000400000000fffffe57ffffffffffffffb5ffffffff0000002a00000000",
            INIT_3B => X"ffffff6dfffffffffffffff9ffffffff0000003e00000000ffffffbaffffffff",
            INIT_3C => X"fffffed4ffffffff000000520000000000000084000000000000013200000000",
            INIT_3D => X"fffffd8affffffffffffffe8fffffffffffffffeffffffffffffff67ffffffff",
            INIT_3E => X"0000002700000000ffffff0efffffffffffffefcffffffffffffff5fffffffff",
            INIT_3F => X"ffffff9dffffffffffffffc5ffffffff0000003300000000fffffffcffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000db000000000000002a000000000000006c000000000000003f00000000",
            INIT_41 => X"0000009a000000000000001400000000ffffffafffffffffffffff40ffffffff",
            INIT_42 => X"ffffffdeffffffff0000009c00000000ffffffb1ffffffff0000007800000000",
            INIT_43 => X"ffffffd0ffffffffffffffcfffffffff0000005000000000ffffffabffffffff",
            INIT_44 => X"ffffffb8ffffffffffffffeaffffffff000000ed00000000000000b600000000",
            INIT_45 => X"00000047000000000000002c00000000ffffffc0ffffffffffffffdcffffffff",
            INIT_46 => X"0000004b00000000ffffff74ffffffff00000015000000000000007c00000000",
            INIT_47 => X"ffffff4effffffff0000003800000000ffffff7dffffffff0000002d00000000",
            INIT_48 => X"ffffff80ffffffff0000004e00000000ffffff6bffffffff0000001600000000",
            INIT_49 => X"ffffffe4ffffffff0000008e000000000000001100000000ffffff68ffffffff",
            INIT_4A => X"ffffffa7ffffffff0000002e00000000000000b8000000000000005700000000",
            INIT_4B => X"ffffffb3ffffffff00000003000000000000006500000000ffffffeaffffffff",
            INIT_4C => X"0000002700000000000000270000000000000074000000000000006700000000",
            INIT_4D => X"00000032000000000000001d0000000000000023000000000000007000000000",
            INIT_4E => X"ffffffe8ffffffffffffffa2ffffffff00000008000000000000003000000000",
            INIT_4F => X"0000002b00000000fffffff8ffffffff0000002f00000000ffffff6dffffffff",
            INIT_50 => X"0000001500000000ffffff3cffffffff0000004e00000000ffffffb4ffffffff",
            INIT_51 => X"ffffff2cffffffffffffffccffffffff0000004400000000000000d500000000",
            INIT_52 => X"0000006400000000ffffff0affffffff0000002e00000000ffffffffffffffff",
            INIT_53 => X"fffffff0ffffffffffffffcdffffffffffffff8fffffffff0000000400000000",
            INIT_54 => X"ffffffd7ffffffffffffffffffffffff0000001c000000000000008800000000",
            INIT_55 => X"0000000a00000000fffffffffffffffffffffff4ffffffffffffffcaffffffff",
            INIT_56 => X"fffffff6ffffffff0000000000000000fffffff5ffffffff0000000d00000000",
            INIT_57 => X"ffffffc4ffffffffffffff84ffffffff0000000c00000000ffffffefffffffff",
            INIT_58 => X"ffffff9dffffffff00000017000000000000005400000000fffffff8ffffffff",
            INIT_59 => X"000000ee00000000ffffff86ffffffff00000032000000000000001200000000",
            INIT_5A => X"0000004c00000000fffffefcffffffffffffffbeffffffffffffffcbffffffff",
            INIT_5B => X"ffffff1fffffffffffffffb2ffffffff0000006300000000ffffffb7ffffffff",
            INIT_5C => X"0000001000000000ffffff2afffffffffffffeddffffffffffffffd0ffffffff",
            INIT_5D => X"ffffff70ffffffff0000007a0000000000000034000000000000005f00000000",
            INIT_5E => X"ffffff6affffffff0000019f000000000000013f00000000ffffff3affffffff",
            INIT_5F => X"ffffff9effffffff000000180000000000000063000000000000000b00000000",
            INIT_60 => X"00000021000000000000001d00000000ffffff8bffffffffffffffecffffffff",
            INIT_61 => X"fffffebafffffffffffffeb1ffffffffffffffb7ffffffff0000000900000000",
            INIT_62 => X"000000a5000000000000009c000000000000004d00000000000000ba00000000",
            INIT_63 => X"fffffeedffffffffffffffefffffffff0000008e00000000000000ae00000000",
            INIT_64 => X"00000004000000000000014300000000ffffff71ffffffffffffffafffffffff",
            INIT_65 => X"fffffff8ffffffff0000008b000000000000007d000000000000006e00000000",
            INIT_66 => X"ffffff33fffffffffffffe2dffffffff0000006800000000ffffffd9ffffffff",
            INIT_67 => X"fffffff9ffffffff00000022000000000000003000000000000000bf00000000",
            INIT_68 => X"ffffff5dffffffffffffffebffffffff0000005000000000ffffff6affffffff",
            INIT_69 => X"0000006500000000fffffffcffffffffffffff68ffffffff0000003400000000",
            INIT_6A => X"0000003100000000ffffff76ffffffffffffff9affffffffffffff5cffffffff",
            INIT_6B => X"00000022000000000000000500000000000000ea000000000000003500000000",
            INIT_6C => X"ffffffd9ffffffffffffffaaffffffffffffffdeffffffffffffff3bffffffff",
            INIT_6D => X"0000001500000000ffffff1cffffffff0000002600000000fffffee6ffffffff",
            INIT_6E => X"0000006400000000000000220000000000000026000000000000001e00000000",
            INIT_6F => X"0000006600000000fffffff5ffffffffffffff69ffffffff0000009d00000000",
            INIT_70 => X"fffffffffffffffffffffe4affffffffffffff74fffffffffffffff4ffffffff",
            INIT_71 => X"0000001f00000000ffffff45ffffffffffffffb2ffffffffffffff82ffffffff",
            INIT_72 => X"0000005200000000fffffeddffffffff0000002a00000000ffffffd5ffffffff",
            INIT_73 => X"0000005100000000ffffff9dffffffffffffff75ffffffffffffffdcffffffff",
            INIT_74 => X"0000005b00000000000000fa00000000ffffffb9ffffffff000000d600000000",
            INIT_75 => X"000000b70000000000000032000000000000004b000000000000005b00000000",
            INIT_76 => X"0000006500000000ffffff90ffffffff0000001c000000000000003e00000000",
            INIT_77 => X"ffffff3fffffffff0000001b00000000000000af000000000000001100000000",
            INIT_78 => X"ffffff91ffffffffffffff57ffffffff00000014000000000000003000000000",
            INIT_79 => X"ffffff9dfffffffffffffff2ffffffffffffffa8fffffffffffffffcffffffff",
            INIT_7A => X"0000002600000000ffffff4affffffffffffff3dffffffffffffff0fffffffff",
            INIT_7B => X"0000000200000000000000c3000000000000003600000000ffffff47ffffffff",
            INIT_7C => X"ffffffc8ffffffff000000eb00000000ffffffd2ffffffffffffffe2ffffffff",
            INIT_7D => X"0000009900000000ffffff8bffffffff000000a100000000fffffdc4ffffffff",
            INIT_7E => X"000000a2000000000000002b000000000000000300000000ffffffe2ffffffff",
            INIT_7F => X"0000001e00000000ffffff9affffffffffffff7cffffffffffffff12ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE7;


    MEM_IWGHT_LAYER2_INSTANCE8 : if BRAM_NAME = "iwght_layer2_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffffcffffffff0000000200000000ffffffe6fffffffffffffff3ffffffff",
            INIT_01 => X"0000000d00000000ffffffddffffffff0000000c00000000fffffff2ffffffff",
            INIT_02 => X"fffffff3fffffffffffffffffffffffffffffff1fffffffffffffff9ffffffff",
            INIT_03 => X"fffffff7ffffffffffffffe3ffffffffffffffeafffffffffffffff1ffffffff",
            INIT_04 => X"ffffffe8ffffffffffffffe0ffffffff0000000e000000000000000300000000",
            INIT_05 => X"fffffff1fffffffffffffffdffffffffffffffe5ffffffffffffffdbffffffff",
            INIT_06 => X"fffffffcfffffffffffffff6fffffffffffffffcfffffffffffffff2ffffffff",
            INIT_07 => X"ffffffecffffffffffffffe2ffffffffffffffe8ffffffffffffffe4ffffffff",
            INIT_08 => X"fffffffaffffffffffffffe8ffffffff0000000d00000000fffffff6ffffffff",
            INIT_09 => X"ffffffe3fffffffffffffff8ffffffffffffffe7ffffffffffffffe5ffffffff",
            INIT_0A => X"fffffff8ffffffff0000000400000000fffffff3ffffffffffffffebffffffff",
            INIT_0B => X"fffffffefffffffffffffff5ffffffff00000002000000000000000700000000",
            INIT_0C => X"0000000500000000fffffff3ffffffffffffffeaffffffffffffffdeffffffff",
            INIT_0D => X"ffffffedfffffffffffffffdffffffffffffffe8ffffffffffffffefffffffff",
            INIT_0E => X"fffffffefffffffffffffffeffffffffffffffdfffffffff0000001200000000",
            INIT_0F => X"fffffff3fffffffffffffff5ffffffff00000000000000000000000500000000",
            INIT_10 => X"ffffffffffffffff0000000400000000fffffff9fffffffffffffff1ffffffff",
            INIT_11 => X"000000030000000000000004000000000000001100000000fffffff6ffffffff",
            INIT_12 => X"fffffff6fffffffffffffffdffffffff0000000100000000fffffffdffffffff",
            INIT_13 => X"ffffffdfffffffffffffffe6fffffffffffffffffffffffffffffffcffffffff",
            INIT_14 => X"ffffffe8fffffffffffffff0fffffffffffffff5ffffffffffffffffffffffff",
            INIT_15 => X"ffffffeeffffffffffffffe4ffffffff0000000300000000ffffffebffffffff",
            INIT_16 => X"0000000800000000ffffffecffffffff0000001600000000fffffff6ffffffff",
            INIT_17 => X"fffffff8fffffffffffffff1fffffffffffffff2ffffffff0000000a00000000",
            INIT_18 => X"fffffffcffffffffffffffe8ffffffffffffffe2ffffffffffffffecffffffff",
            INIT_19 => X"fffffff4ffffffff0000000300000000ffffffeffffffffffffffff5ffffffff",
            INIT_1A => X"0000000600000000ffffffdffffffffffffffff3fffffffffffffff1ffffffff",
            INIT_1B => X"fffffff4fffffffffffffff3fffffffffffffffaffffffffffffffd9ffffffff",
            INIT_1C => X"ffffffdaffffffffffffffecffffffffffffffebffffffff0000000300000000",
            INIT_1D => X"fffffffaffffffff0000000e000000000000000700000000fffffffcffffffff",
            INIT_1E => X"0000000500000000fffffff5ffffffffffffffefffffffff0000000600000000",
            INIT_1F => X"fffffff0ffffffff000000000000000000000000000000000000000300000000",
            INIT_20 => X"0000000400000000fffffffaffffffff0000000a000000000000000f00000000",
            INIT_21 => X"ffffffedfffffffffffffff9fffffffffffffff5ffffffff0000001600000000",
            INIT_22 => X"0000000500000000fffffff9ffffffffffffffe7ffffffffffffffe6ffffffff",
            INIT_23 => X"0000000200000000fffffff4ffffffff0000000400000000ffffffe5ffffffff",
            INIT_24 => X"fffffff7ffffffff0000000a00000000fffffff0fffffffffffffffbffffffff",
            INIT_25 => X"fffffffefffffffffffffff2ffffffff0000000a00000000fffffff4ffffffff",
            INIT_26 => X"fffffff5fffffffffffffff3ffffffff0000001100000000fffffff6ffffffff",
            INIT_27 => X"ffffffebfffffffffffffff1ffffffff0000001100000000fffffff8ffffffff",
            INIT_28 => X"0000000800000000ffffffeafffffffffffffff3ffffffff0000000400000000",
            INIT_29 => X"fffffffbffffffff0000000a000000000000000100000000ffffffeeffffffff",
            INIT_2A => X"ffffffeaffffffffffffffebfffffffffffffff7fffffffffffffffeffffffff",
            INIT_2B => X"ffffffffffffffff0000000c00000000ffffffe5fffffffffffffffdffffffff",
            INIT_2C => X"0000000100000000fffffff5ffffffff0000001400000000fffffffaffffffff",
            INIT_2D => X"fffffff1ffffffff0000000000000000ffffffefffffffffffffffe2ffffffff",
            INIT_2E => X"ffffffe4ffffffffffffffffffffffff0000000300000000fffffffaffffffff",
            INIT_2F => X"0000000000000000fffffffdfffffffffffffffeffffffff0000000000000000",
            INIT_30 => X"ffffffeaffffffffffffffebfffffffffffffff0ffffffff0000000000000000",
            INIT_31 => X"fffffffbffffffffffffffeeffffffff0000000000000000fffffff2ffffffff",
            INIT_32 => X"fffffff3ffffffffffffffe8fffffffffffffff5ffffffff0000000a00000000",
            INIT_33 => X"fffffff7ffffffff0000000b0000000000000013000000000000000000000000",
            INIT_34 => X"00000002000000000000000600000000fffffff0ffffffffffffffeaffffffff",
            INIT_35 => X"ffffffe5fffffffffffffffbfffffffffffffff9fffffffffffffff2ffffffff",
            INIT_36 => X"fffffffeffffffff0000000b00000000fffffff0fffffffffffffff5ffffffff",
            INIT_37 => X"0000000b00000000fffffffefffffffffffffff7ffffffffffffffe8ffffffff",
            INIT_38 => X"fffffff3ffffffffffffffedffffffff0000000900000000fffffffaffffffff",
            INIT_39 => X"fffffff3ffffffff00000006000000000000000c00000000fffffffaffffffff",
            INIT_3A => X"0000000000000000fffffff7fffffffffffffff3fffffffffffffffeffffffff",
            INIT_3B => X"00000004000000000000000d000000000000000000000000fffffffaffffffff",
            INIT_3C => X"ffffffdfffffffff0000000d00000000fffffff3ffffffff0000000400000000",
            INIT_3D => X"ffffffffffffffffffffffedfffffffffffffff1fffffffffffffff6ffffffff",
            INIT_3E => X"00000001000000000000000400000000ffffffe1fffffffffffffffbffffffff",
            INIT_3F => X"ffffffe8ffffffff0000000400000000fffffff3fffffffffffffffeffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000400000000fffffffcfffffffffffffff5ffffffffffffffe6ffffffff",
            INIT_41 => X"0000000300000000ffffffebffffffff0000000800000000ffffffffffffffff",
            INIT_42 => X"fffffff0ffffffff0000000400000000fffffff1fffffffffffffff6ffffffff",
            INIT_43 => X"0000000400000000fffffff8ffffffffffffffefffffffff0000000b00000000",
            INIT_44 => X"fffffff4fffffffffffffff9ffffffff00000001000000000000000a00000000",
            INIT_45 => X"ffffffebffffffff0000000c000000000000000200000000fffffff4ffffffff",
            INIT_46 => X"ffffffe4fffffffffffffff9ffffffff0000000700000000ffffffedffffffff",
            INIT_47 => X"ffffffedffffffff0000000400000000ffffffe7ffffffffffffffe1ffffffff",
            INIT_48 => X"ffffffaeffffffff0000001f00000000ffffffb7ffffffff0000006000000000",
            INIT_49 => X"ffffff81ffffffffffffffd9ffffffff00000042000000000000002100000000",
            INIT_4A => X"000000d600000000ffffffb0ffffffffffffffaefffffffffffffff3ffffffff",
            INIT_4B => X"ffffff9affffffff0000000d000000000000003300000000ffffff81ffffffff",
            INIT_4C => X"000000a300000000ffffff70ffffffffffffff5bffffffffffffff9cffffffff",
            INIT_4D => X"ffffff95ffffffff000000bc000000000000002500000000ffffffdbffffffff",
            INIT_4E => X"fffffffcffffffffffffffc5ffffffff0000001300000000fffffff2ffffffff",
            INIT_4F => X"000000190000000000000082000000000000003200000000ffffff91ffffffff",
            INIT_50 => X"0000008500000000000000050000000000000048000000000000001500000000",
            INIT_51 => X"0000002700000000fffffffeffffffffffffff47ffffffffffffffcdffffffff",
            INIT_52 => X"ffffffe2ffffffff0000007100000000ffffff75ffffffffffffffccffffffff",
            INIT_53 => X"0000001a0000000000000025000000000000003c000000000000003100000000",
            INIT_54 => X"ffffffdaffffffff000000ee00000000000000dc00000000ffffffbeffffffff",
            INIT_55 => X"0000004400000000ffffff8dffffffff0000008000000000ffffffa3ffffffff",
            INIT_56 => X"00000051000000000000003500000000ffffffe7ffffffffffffff42ffffffff",
            INIT_57 => X"ffffffa7ffffffff000000bc00000000ffffffa5ffffffff0000003f00000000",
            INIT_58 => X"ffffffedffffffff0000005d00000000fffffff8ffffffffffffff81ffffffff",
            INIT_59 => X"000000f6000000000000006200000000ffffff99ffffffff0000002500000000",
            INIT_5A => X"ffffff93ffffffffffffffd7ffffffff000000c700000000fffffff8ffffffff",
            INIT_5B => X"ffffff74ffffffff0000000a00000000ffffffc5ffffffff000000a700000000",
            INIT_5C => X"fffffff6ffffffff0000001f00000000ffffffd1ffffffffffffff3dffffffff",
            INIT_5D => X"000000840000000000000081000000000000005e00000000ffffffdeffffffff",
            INIT_5E => X"fffffffcffffffff000000a900000000ffffffe3ffffffffffffffadffffffff",
            INIT_5F => X"0000005200000000000000460000000000000046000000000000009d00000000",
            INIT_60 => X"0000004500000000000000410000000000000091000000000000000400000000",
            INIT_61 => X"ffffffacffffffff0000001900000000ffffff9bffffffff0000003e00000000",
            INIT_62 => X"ffffff20ffffffff0000002a000000000000000300000000ffffffeeffffffff",
            INIT_63 => X"00000014000000000000005700000000ffffffc0ffffffffffffffdfffffffff",
            INIT_64 => X"ffffffffffffffff00000065000000000000003800000000ffffffddffffffff",
            INIT_65 => X"0000000000000000fffffffbffffffff0000001a000000000000003000000000",
            INIT_66 => X"00000006000000000000000f000000000000000b000000000000000a00000000",
            INIT_67 => X"0000003d00000000ffffffcafffffffffffffffdfffffffffffffff3ffffffff",
            INIT_68 => X"ffffffe6ffffffffffffffcaffffffff0000002d000000000000006400000000",
            INIT_69 => X"ffffff8affffffff0000002200000000ffffffd1ffffffffffffffa6ffffffff",
            INIT_6A => X"fffffff4ffffffff00000028000000000000002b00000000ffffffbdffffffff",
            INIT_6B => X"0000005f00000000ffffffc4ffffffffffffffb6ffffffffffffffe9ffffffff",
            INIT_6C => X"ffffff6dffffffffffffffd4ffffffff0000002300000000ffffff23ffffffff",
            INIT_6D => X"ffffffa4ffffffff000000c100000000ffffff76ffffffffffffff73ffffffff",
            INIT_6E => X"fffffe44ffffffff000000f500000000000000a600000000ffffff90ffffffff",
            INIT_6F => X"0000007000000000ffffffbdffffffffffffffa4ffffffff0000008500000000",
            INIT_70 => X"00000087000000000000000a000000000000001d00000000fffffeb2ffffffff",
            INIT_71 => X"00000086000000000000002000000000ffffffcdffffffff0000003300000000",
            INIT_72 => X"0000000d0000000000000015000000000000006700000000ffffff1effffffff",
            INIT_73 => X"0000004600000000fffffe01ffffffff0000011700000000ffffff5bffffffff",
            INIT_74 => X"0000007a00000000ffffffefffffffffffffffe4fffffffffffffee9ffffffff",
            INIT_75 => X"ffffffcdfffffffffffffedbffffffffffffff64ffffffff0000008900000000",
            INIT_76 => X"ffffffa2ffffffff0000008800000000ffffffadffffffffffffffc1ffffffff",
            INIT_77 => X"000000030000000000000076000000000000002100000000fffffe0fffffffff",
            INIT_78 => X"ffffffcfffffffffffffff04ffffffffffffffe7ffffffffffffffa6ffffffff",
            INIT_79 => X"00000005000000000000009e00000000ffffffc2ffffffffffffffedffffffff",
            INIT_7A => X"000000b600000000ffffffeaffffffffffffffe0ffffffff0000002700000000",
            INIT_7B => X"00000043000000000000009b0000000000000072000000000000007700000000",
            INIT_7C => X"0000004600000000ffffff95ffffffff0000002000000000ffffff97ffffffff",
            INIT_7D => X"ffffff9effffffffffffff73ffffffff00000049000000000000006d00000000",
            INIT_7E => X"0000009000000000ffffffceffffffffffffffa1ffffffffffffffd5ffffffff",
            INIT_7F => X"0000003800000000000000390000000000000033000000000000009200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE8;


    MEM_IWGHT_LAYER2_INSTANCE9 : if BRAM_NAME = "iwght_layer2_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffc2ffffffffffffffcdffffffffffffff51ffffffff0000013200000000",
            INIT_01 => X"ffffffdbffffffffffffffe9ffffffff0000005b00000000ffffff29ffffffff",
            INIT_02 => X"0000005700000000ffffff76ffffffffffffffb3ffffffff0000003800000000",
            INIT_03 => X"ffffffb4ffffffffffffffffffffffffffffff98ffffffff0000006400000000",
            INIT_04 => X"0000003c00000000ffffffe7ffffffffffffff77ffffffffffffffe6ffffffff",
            INIT_05 => X"ffffffb8fffffffffffffff1ffffffff00000023000000000000002000000000",
            INIT_06 => X"0000007c000000000000004900000000fffffff4ffffffff0000002600000000",
            INIT_07 => X"0000003100000000ffffff47ffffffff000000d8000000000000003600000000",
            INIT_08 => X"ffffff4cffffffffffffffe8ffffffffffffff86ffffffffffffffb4ffffffff",
            INIT_09 => X"0000001500000000ffffffc9ffffffff000000a6000000000000002200000000",
            INIT_0A => X"ffffffd1ffffffff000000d200000000ffffffafffffffffffffff79ffffffff",
            INIT_0B => X"0000002b00000000000000a700000000ffffffd1ffffffffffffffcfffffffff",
            INIT_0C => X"0000002800000000ffffffdaffffffff0000003200000000ffffffaeffffffff",
            INIT_0D => X"0000002300000000ffffffb6ffffffff0000003f00000000ffffff9dffffffff",
            INIT_0E => X"ffffff83ffffffffffffff6fffffffffffffffffffffffff000000a100000000",
            INIT_0F => X"ffffff25ffffffff0000006300000000ffffff90ffffffffffffffb5ffffffff",
            INIT_10 => X"fffffeedffffffff0000002f00000000ffffff9dffffffffffffff7bffffffff",
            INIT_11 => X"ffffffeefffffffffffffeedfffffffffffffff3ffffffff0000000100000000",
            INIT_12 => X"ffffffd2ffffffff00000070000000000000003b00000000fffffff8ffffffff",
            INIT_13 => X"ffffffa6ffffffff0000008200000000000000a000000000ffffff63ffffffff",
            INIT_14 => X"0000003200000000000000ef000000000000006300000000ffffff9fffffffff",
            INIT_15 => X"ffffffedffffffffffffffd6fffffffffffffffaffffffffffffff84ffffffff",
            INIT_16 => X"ffffff9dffffffff00000073000000000000003000000000fffffff7ffffffff",
            INIT_17 => X"0000004800000000ffffffd4ffffffffffffff9bffffffffffffff72ffffffff",
            INIT_18 => X"0000004b00000000fffffff5ffffffff0000002d00000000ffffffcdffffffff",
            INIT_19 => X"ffffff20ffffffffffffff25ffffffffffffffbfffffffff0000002f00000000",
            INIT_1A => X"ffffffc4fffffffffffffd09ffffffffffffffb4fffffffffffffebdffffffff",
            INIT_1B => X"0000002f0000000000000093000000000000004e00000000fffffffeffffffff",
            INIT_1C => X"ffffff68ffffffff0000005f000000000000000d00000000000000af00000000",
            INIT_1D => X"ffffffb3ffffffff0000002a00000000fffffeb5ffffffff0000009500000000",
            INIT_1E => X"ffffffd6fffffffffffffffcffffffffffffffc2ffffffff0000003600000000",
            INIT_1F => X"000000530000000000000065000000000000002400000000ffffffb6ffffffff",
            INIT_20 => X"0000000300000000ffffffa0ffffffff00000079000000000000002400000000",
            INIT_21 => X"ffffff7bffffffff0000009c00000000ffffff12ffffffff0000002100000000",
            INIT_22 => X"0000001a00000000ffffffe3ffffffffffffffe8ffffffffffffff91ffffffff",
            INIT_23 => X"000000f800000000ffffff9bffffffff0000001000000000ffffff62ffffffff",
            INIT_24 => X"ffffff1fffffffffffffffdcffffffff0000004800000000ffffff5affffffff",
            INIT_25 => X"ffffff16ffffffffffffff47ffffffffffffff7effffffffffffff01ffffffff",
            INIT_26 => X"ffffffecffffffff00000064000000000000006300000000fffffddbffffffff",
            INIT_27 => X"ffffff6affffffff00000094000000000000000a00000000ffffff99ffffffff",
            INIT_28 => X"00000037000000000000002f000000000000006a00000000ffffffb5ffffffff",
            INIT_29 => X"0000004700000000fffffffbffffffffffffffd7ffffffff0000003900000000",
            INIT_2A => X"ffffff9effffffff0000000c000000000000004300000000000000cf00000000",
            INIT_2B => X"ffffffaaffffffff00000052000000000000008800000000ffffffddffffffff",
            INIT_2C => X"ffffff22ffffffffffffffc3ffffffffffffffccffffffffffffffc4ffffffff",
            INIT_2D => X"fffffff7fffffffffffffff9fffffffffffffff8ffffffffffffff3dffffffff",
            INIT_2E => X"fffffff3ffffffff00000014000000000000001300000000fffffff6ffffffff",
            INIT_2F => X"ffffffc1ffffffffffffff4dfffffffffffffff4fffffffffffffff0ffffffff",
            INIT_30 => X"ffffff4fffffffffffffffddfffffffffffffedcffffffffffffffc3ffffffff",
            INIT_31 => X"00000004000000000000006800000000ffffff41fffffffffffffedfffffffff",
            INIT_32 => X"ffffffd0fffffffffffffffcffffffffffffff64ffffffff0000004700000000",
            INIT_33 => X"ffffff36ffffffff000000ba000000000000008300000000ffffff93ffffffff",
            INIT_34 => X"ffffff9effffffff0000008400000000ffffffbcffffffffffffffaaffffffff",
            INIT_35 => X"ffffff37ffffffff00000038000000000000002f00000000ffffff78ffffffff",
            INIT_36 => X"0000008f0000000000000112000000000000003000000000ffffff29ffffffff",
            INIT_37 => X"0000013c00000000fffffee6ffffffffffffff91ffffffff000000a900000000",
            INIT_38 => X"ffffffcaffffffffffffffbbfffffffffffffff2ffffffffffffffa6ffffffff",
            INIT_39 => X"0000006b0000000000000051000000000000004e00000000ffffffe1ffffffff",
            INIT_3A => X"0000000000000000fffffff9ffffffff0000002000000000000000fe00000000",
            INIT_3B => X"ffffffd8ffffffff000000de00000000ffffff7dffffffffffffffe1ffffffff",
            INIT_3C => X"00000036000000000000008f00000000ffffffc1ffffffff0000009200000000",
            INIT_3D => X"fffffff5ffffffffffffff59ffffffff0000002600000000ffffff2cffffffff",
            INIT_3E => X"0000002a00000000ffffff56ffffffff0000007a000000000000004e00000000",
            INIT_3F => X"0000004a000000000000005700000000ffffffbaffffffff0000004500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffff23ffffffffffffff63ffffffffffffffbdffffffffffffff72ffffffff",
            INIT_41 => X"0000008500000000ffffff56ffffffffffffffbfffffffff0000001c00000000",
            INIT_42 => X"ffffffb7ffffffff0000002a00000000ffffff60ffffffffffffff9cffffffff",
            INIT_43 => X"ffffffb4ffffffff0000006a000000000000003100000000fffffffcffffffff",
            INIT_44 => X"ffffff84ffffffff000000790000000000000064000000000000005300000000",
            INIT_45 => X"ffffffe8ffffffffffffff03ffffffff0000003a000000000000015000000000",
            INIT_46 => X"0000001a000000000000009500000000ffffffe3ffffffffffffffe7ffffffff",
            INIT_47 => X"fffffff8ffffffff0000003f000000000000000e00000000ffffffc9ffffffff",
            INIT_48 => X"000000a800000000ffffff5affffffffffffffcfffffffff0000006600000000",
            INIT_49 => X"00000000000000000000003100000000ffffff4effffffff000000cd00000000",
            INIT_4A => X"ffffffbafffffffffffffff2ffffffff0000002300000000ffffffd3ffffffff",
            INIT_4B => X"00000049000000000000005100000000ffffff8effffffff0000003a00000000",
            INIT_4C => X"0000003b000000000000003700000000ffffff77ffffffff0000004c00000000",
            INIT_4D => X"ffffff65ffffffff0000006500000000fffffff4ffffffff0000002d00000000",
            INIT_4E => X"0000002300000000ffffffddffffffff000000cd00000000ffffffdfffffffff",
            INIT_4F => X"ffffffcdfffffffffffffffdffffffff0000004100000000fffffff7ffffffff",
            INIT_50 => X"fffffff8ffffffff0000003a00000000ffffff86ffffffffffffffd5ffffffff",
            INIT_51 => X"00000056000000000000005900000000ffffffc2ffffffff0000002100000000",
            INIT_52 => X"0000001700000000000000c500000000fffffff8ffffffff0000004700000000",
            INIT_53 => X"0000005900000000ffffffa5ffffffff0000006400000000ffffff87ffffffff",
            INIT_54 => X"ffffffdeffffffffffffffdfffffffff0000002f00000000fffffff7ffffffff",
            INIT_55 => X"0000007e00000000ffffff4bffffffff0000001500000000000000b900000000",
            INIT_56 => X"ffffff71ffffffff000000740000000000000044000000000000001d00000000",
            INIT_57 => X"0000003000000000fffffff4ffffffff0000007200000000ffffffe4ffffffff",
            INIT_58 => X"ffffff4dffffffffffffffd1ffffffffffffff95ffffffffffffff01ffffffff",
            INIT_59 => X"fffffff5ffffffffffffff89ffffffffffffff0effffffffffffffd1ffffffff",
            INIT_5A => X"ffffff83ffffffffffffffbcffffffffffffffcdffffffffffffffecffffffff",
            INIT_5B => X"0000004b00000000ffffff8effffffff0000001400000000000000ef00000000",
            INIT_5C => X"fffffffbfffffffffffffff5ffffffff0000006c00000000ffffffbbffffffff",
            INIT_5D => X"ffffffccffffffffffffff5affffffff0000006800000000ffffff2dffffffff",
            INIT_5E => X"0000008000000000ffffff75ffffffffffffff8affffffff0000000c00000000",
            INIT_5F => X"ffffff87ffffffff0000006a0000000000000042000000000000005100000000",
            INIT_60 => X"0000008300000000ffffff93ffffffffffffff93ffffffffffffff48ffffffff",
            INIT_61 => X"000000ce000000000000007d00000000000000b7000000000000000c00000000",
            INIT_62 => X"ffffffd9ffffffff0000004200000000ffffffd8ffffffff0000002300000000",
            INIT_63 => X"0000009000000000ffffff82ffffffffffffff27ffffffffffffff8cffffffff",
            INIT_64 => X"0000006c000000000000001000000000ffffffd2ffffffffffffffebffffffff",
            INIT_65 => X"fffffffaffffffff0000004b00000000ffffffd1ffffffff0000002f00000000",
            INIT_66 => X"ffffff4bfffffffffffffe9bffffffffffffffe7ffffffff0000002e00000000",
            INIT_67 => X"ffffffadffffffffffffffc8ffffffffffffffe5ffffffffffffffeeffffffff",
            INIT_68 => X"ffffff9dffffffff0000001c00000000ffffff27ffffffffffffff50ffffffff",
            INIT_69 => X"ffffff75ffffffff00000011000000000000005500000000ffffff61ffffffff",
            INIT_6A => X"ffffff83ffffffffffffff42fffffffffffffffeffffffff0000006200000000",
            INIT_6B => X"ffffff9affffffff000000130000000000000045000000000000002c00000000",
            INIT_6C => X"ffffffe2ffffffffffffff86ffffffffffffffb2ffffffff000000df00000000",
            INIT_6D => X"000000b3000000000000001c000000000000006c000000000000002f00000000",
            INIT_6E => X"ffffff8effffffffffffff4fffffffffffffff9fffffffff0000005c00000000",
            INIT_6F => X"fffffff0ffffffff0000001800000000ffffff4cffffffffffffffddffffffff",
            INIT_70 => X"0000004e000000000000004700000000ffffffd2ffffffffffffffcfffffffff",
            INIT_71 => X"ffffffc7ffffffff000000b000000000ffffffb4ffffffffffffff97ffffffff",
            INIT_72 => X"0000002300000000ffffffaeffffffff0000002c00000000ffffff34ffffffff",
            INIT_73 => X"ffffff85ffffffff000000030000000000000052000000000000001d00000000",
            INIT_74 => X"00000027000000000000008200000000ffffffd9ffffffff0000003400000000",
            INIT_75 => X"fffffffbffffffff0000000f00000000fffffff4ffffffff0000001600000000",
            INIT_76 => X"fffffff9ffffffff0000000d00000000fffffff5fffffffffffffff1ffffffff",
            INIT_77 => X"0000005a000000000000002700000000fffffff9ffffffff0000000600000000",
            INIT_78 => X"fffffffbffffffff0000000000000000fffffff8ffffffff0000000b00000000",
            INIT_79 => X"00000054000000000000003b000000000000006600000000ffffffccffffffff",
            INIT_7A => X"0000001e00000000fffffff3ffffffffffffffc9ffffffff0000001200000000",
            INIT_7B => X"ffffffc1ffffffffffffffd0ffffffff0000005e000000000000003e00000000",
            INIT_7C => X"0000001400000000fffffff2ffffffffffffff94ffffffff0000001f00000000",
            INIT_7D => X"ffffffc2ffffffff000000300000000000000045000000000000001c00000000",
            INIT_7E => X"0000002d00000000ffffffc0ffffffff0000010e000000000000004000000000",
            INIT_7F => X"000000b900000000ffffff51ffffffff0000003700000000ffffffb9ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE9;


    MEM_IWGHT_LAYER2_INSTANCE10 : if BRAM_NAME = "iwght_layer2_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffff90ffffffff00000054000000000000006d00000000fffffff5ffffffff",
            INIT_01 => X"0000001900000000ffffffaaffffffff0000007e00000000ffffff89ffffffff",
            INIT_02 => X"0000002e000000000000000300000000ffffff27ffffffff0000002a00000000",
            INIT_03 => X"ffffff41ffffffff0000002300000000fffffffaffffffff0000007300000000",
            INIT_04 => X"ffffff80ffffffff0000008000000000000000a300000000ffffff80ffffffff",
            INIT_05 => X"00000047000000000000006b0000000000000047000000000000001f00000000",
            INIT_06 => X"ffffffeaffffffff00000080000000000000001600000000ffffff3bffffffff",
            INIT_07 => X"0000003f000000000000007800000000ffffffb0ffffffff0000008100000000",
            INIT_08 => X"ffffff83ffffffff0000002c00000000ffffff8fffffffff0000000300000000",
            INIT_09 => X"000000e500000000000000f7000000000000006400000000ffffff6fffffffff",
            INIT_0A => X"0000005900000000ffffffc5ffffffff0000001300000000ffffff91ffffffff",
            INIT_0B => X"ffffffd2ffffffffffffff2cffffffff00000061000000000000009700000000",
            INIT_0C => X"ffffff7fffffffff00000027000000000000007f00000000ffffffbdffffffff",
            INIT_0D => X"0000000000000000fffffff9ffffffffffffff70fffffffffffffff6ffffffff",
            INIT_0E => X"00000083000000000000004d00000000ffffff32ffffffff0000007900000000",
            INIT_0F => X"ffffff16ffffffff0000000800000000000000a600000000ffffffb5ffffffff",
            INIT_10 => X"000000230000000000000012000000000000001100000000ffffffd5ffffffff",
            INIT_11 => X"0000004b00000000000000540000000000000036000000000000003400000000",
            INIT_12 => X"0000003b00000000ffffff8afffffffffffffff0ffffffffffffffccffffffff",
            INIT_13 => X"0000007000000000ffffff32ffffffffffffffefffffffff0000000500000000",
            INIT_14 => X"00000042000000000000000f00000000fffffffdffffffff000000f000000000",
            INIT_15 => X"ffffffe6ffffffff0000003e00000000ffffffe8fffffffffffffff5ffffffff",
            INIT_16 => X"ffffffe4ffffffff000000b80000000000000029000000000000000000000000",
            INIT_17 => X"ffffffdfffffffff0000003200000000ffffff9affffffffffffffedffffffff",
            INIT_18 => X"00000023000000000000002a000000000000006600000000ffffffe7ffffffff",
            INIT_19 => X"ffffffb4ffffffff0000005e000000000000009f00000000ffffffacffffffff",
            INIT_1A => X"000000fd0000000000000003000000000000008a000000000000002800000000",
            INIT_1B => X"ffffff7cffffffffffffff41ffffffffffffff9fffffffff000000ae00000000",
            INIT_1C => X"0000000700000000ffffff4effffffff00000023000000000000008d00000000",
            INIT_1D => X"0000000a000000000000000700000000fffffff9ffffffffffffffe9ffffffff",
            INIT_1E => X"0000008f00000000fffffff1fffffffffffffff2ffffffffffffffceffffffff",
            INIT_1F => X"000000f700000000ffffffeeffffffffffffff54ffffffffffffffe9ffffffff",
            INIT_20 => X"0000006f00000000ffffff9bfffffffffffffffbffffffffffffff4dffffffff",
            INIT_21 => X"00000033000000000000005d0000000000000000000000000000005200000000",
            INIT_22 => X"00000014000000000000000f000000000000002500000000ffffffb9ffffffff",
            INIT_23 => X"0000006e00000000000000000000000000000095000000000000005000000000",
            INIT_24 => X"ffffffe0ffffffff0000002500000000ffffff8bffffffff0000007000000000",
            INIT_25 => X"0000005d000000000000003900000000ffffffa2ffffffff000000ba00000000",
            INIT_26 => X"0000001f00000000fffffebdfffffffffffffed8ffffffffffffffaeffffffff",
            INIT_27 => X"ffffff35ffffffff0000009800000000ffffffd1ffffffff0000007c00000000",
            INIT_28 => X"ffffffbcffffffff0000002600000000ffffff60ffffffffffffff97ffffffff",
            INIT_29 => X"ffffff7cfffffffffffffeb1fffffffffffffeb7ffffffffffffff76ffffffff",
            INIT_2A => X"ffffff4cffffffffffffff74ffffffffffffff7dffffffffffffff6affffffff",
            INIT_2B => X"0000004400000000ffffffa8ffffffffffffff4effffffffffffffeeffffffff",
            INIT_2C => X"ffffffc3ffffffff0000005c0000000000000092000000000000004b00000000",
            INIT_2D => X"ffffffb3ffffffff00000090000000000000003f000000000000008200000000",
            INIT_2E => X"ffffff76ffffffff0000006000000000000000c000000000ffffffdbffffffff",
            INIT_2F => X"0000003700000000ffffffe9ffffffff0000000f000000000000002f00000000",
            INIT_30 => X"0000001700000000ffffffe6ffffffff0000003f00000000ffffff4bffffffff",
            INIT_31 => X"ffffffbbffffffff000000460000000000000055000000000000001000000000",
            INIT_32 => X"ffffffa3ffffffffffffff79fffffffffffffff6ffffffffffffffdaffffffff",
            INIT_33 => X"ffffff1effffffffffffffbcffffffffffffff57fffffffffffffffaffffffff",
            INIT_34 => X"0000001000000000ffffffa1ffffffffffffff8affffffff0000005100000000",
            INIT_35 => X"ffffff8cffffffffffffff44ffffffffffffff78ffffffffffffffa9ffffffff",
            INIT_36 => X"000000c100000000ffffff5dffffffff0000007a00000000ffffffccffffffff",
            INIT_37 => X"ffffffc2ffffffff0000005500000000000000ed000000000000006600000000",
            INIT_38 => X"ffffffe8ffffffff00000041000000000000000c00000000ffffff73ffffffff",
            INIT_39 => X"ffffffafffffffff0000003f0000000000000056000000000000003600000000",
            INIT_3A => X"000000a800000000ffffffc7ffffffffffffffc0ffffffff0000007500000000",
            INIT_3B => X"ffffff2effffffff00000033000000000000003100000000ffffff96ffffffff",
            INIT_3C => X"ffffff52ffffffffffffffa1ffffffffffffff0dffffffffffffff78ffffffff",
            INIT_3D => X"0000000100000000ffffffe9ffffffff0000000b00000000000000f500000000",
            INIT_3E => X"fffffffafffffffffffffff3fffffffffffffffdfffffffffffffff3ffffffff",
            INIT_3F => X"ffffffd4ffffffffffffff7effffffff0000001f000000000000000d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002400000000ffffffc0ffffffff0000006f00000000fffffed8ffffffff",
            INIT_41 => X"ffffffd9ffffffffffffff5effffffff0000006200000000ffffffefffffffff",
            INIT_42 => X"0000008900000000ffffff66ffffffffffffff12ffffffff0000001600000000",
            INIT_43 => X"0000002100000000fffffffaffffffff0000000300000000ffffff03ffffffff",
            INIT_44 => X"000000b10000000000000173000000000000007d00000000ffffffc2ffffffff",
            INIT_45 => X"fffffffeffffffffffffffe1ffffffff00000007000000000000001c00000000",
            INIT_46 => X"ffffff45ffffffff0000000200000000ffffff6dffffffff0000002200000000",
            INIT_47 => X"ffffff91ffffffff0000007300000000ffffff68ffffffff0000000000000000",
            INIT_48 => X"0000002f00000000ffffff3fffffffffffffff77ffffffffffffff65ffffffff",
            INIT_49 => X"ffffff6effffffff00000060000000000000002c000000000000000800000000",
            INIT_4A => X"ffffffd6ffffffffffffff91ffffffffffffff4effffffff0000013300000000",
            INIT_4B => X"ffffff84ffffffffffffffc3ffffffffffffffb6ffffffff0000014600000000",
            INIT_4C => X"000000da00000000ffffff3effffffffffffff73fffffffffffffed5ffffffff",
            INIT_4D => X"ffffff9bffffffffffffff94ffffffffffffff7affffffffffffff8dffffffff",
            INIT_4E => X"ffffffe1fffffffffffffffcffffffff0000008400000000000000b900000000",
            INIT_4F => X"ffffffb6ffffffff0000004300000000ffffffdfffffffff0000001400000000",
            INIT_50 => X"ffffffdaffffffff000000f600000000ffffffb2ffffffffffffff88ffffffff",
            INIT_51 => X"ffffffdcffffffff0000000000000000fffffef6ffffffffffffffdaffffffff",
            INIT_52 => X"ffffff9bffffffffffffffb4ffffffff00000052000000000000008500000000",
            INIT_53 => X"ffffffdcffffffffffffffe9ffffffff0000005400000000ffffffe6ffffffff",
            INIT_54 => X"0000000600000000ffffffcaffffffffffffff9dffffffff0000009800000000",
            INIT_55 => X"0000005600000000ffffff52ffffffff0000002900000000ffffffb3ffffffff",
            INIT_56 => X"fffffffeffffffffffffff49fffffffffffffec0ffffffff000000af00000000",
            INIT_57 => X"0000001a000000000000009600000000ffffff07ffffffff0000006d00000000",
            INIT_58 => X"000000ad00000000ffffff1affffffffffffffc5ffffffff0000004200000000",
            INIT_59 => X"0000000000000000ffffff2effffffff0000000c00000000ffffffe8ffffffff",
            INIT_5A => X"0000002800000000ffffff9dffffffff0000002d000000000000001b00000000",
            INIT_5B => X"ffffff6fffffffff0000003e00000000ffffffb3ffffffffffffffecffffffff",
            INIT_5C => X"0000000f000000000000001f00000000ffffff52fffffffffffffff6ffffffff",
            INIT_5D => X"0000006f0000000000000022000000000000004b000000000000000a00000000",
            INIT_5E => X"ffffffa0ffffffffffffff55ffffffff0000007c000000000000002300000000",
            INIT_5F => X"0000007d000000000000005000000000ffffff52ffffffff0000003e00000000",
            INIT_60 => X"ffffff85ffffffff0000005600000000ffffffeeffffffff0000006800000000",
            INIT_61 => X"ffffffeeffffffff0000001c000000000000004400000000ffffff94ffffffff",
            INIT_62 => X"0000004e00000000ffffff95ffffffffffffffd4ffffffff0000009b00000000",
            INIT_63 => X"0000000f00000000ffffff42ffffffff0000002300000000ffffff60ffffffff",
            INIT_64 => X"0000002a000000000000008e00000000ffffffc2fffffffffffffff2ffffffff",
            INIT_65 => X"0000008000000000ffffffe6ffffffffffffffd0ffffffff0000006800000000",
            INIT_66 => X"000000240000000000000025000000000000003c00000000ffffffa4ffffffff",
            INIT_67 => X"ffffffd2ffffffffffffff33fffffffffffffffffffffffffffffffaffffffff",
            INIT_68 => X"00000001000000000000002700000000ffffff81ffffffffffffff8cffffffff",
            INIT_69 => X"00000076000000000000000500000000000000c6000000000000005600000000",
            INIT_6A => X"0000002e00000000ffffff85ffffffff00000004000000000000005b00000000",
            INIT_6B => X"fffffff1ffffffffffffffd4ffffffffffffff69ffffffff0000003300000000",
            INIT_6C => X"ffffff9dffffffff0000008800000000ffffffddffffffffffffff66ffffffff",
            INIT_6D => X"ffffff8affffffff0000010a0000000000000009000000000000003e00000000",
            INIT_6E => X"ffffff8effffffff0000000000000000ffffffe4ffffffffffffff9cffffffff",
            INIT_6F => X"ffffffb4ffffffffffffff81ffffffff0000005b000000000000008a00000000",
            INIT_70 => X"ffffffe3ffffffffffffff91ffffffff00000006000000000000002000000000",
            INIT_71 => X"0000005500000000ffffff7cffffffffffffff9affffffffffffffd3ffffffff",
            INIT_72 => X"fffffed8ffffffffffffffbeffffffffffffff53fffffffffffffff4ffffffff",
            INIT_73 => X"0000005a0000000000000024000000000000001e000000000000006f00000000",
            INIT_74 => X"ffffffd5ffffffffffffffb3ffffffff0000004a00000000fffffee4ffffffff",
            INIT_75 => X"fffffe9affffffffffffff71ffffffffffffffa9ffffffff0000008800000000",
            INIT_76 => X"fffffff5ffffffffffffff85ffffffff0000003900000000ffffff31ffffffff",
            INIT_77 => X"ffffffefffffffffffffff77ffffffffffffff4cffffffff0000008300000000",
            INIT_78 => X"0000003800000000ffffff51ffffffff0000002500000000ffffff70ffffffff",
            INIT_79 => X"0000006100000000ffffff6fffffffffffffffbffffffffffffffffdffffffff",
            INIT_7A => X"fffffea3ffffffff0000008100000000ffffff5bffffffffffffff8dffffffff",
            INIT_7B => X"0000003f00000000ffffff8cffffffff00000076000000000000004a00000000",
            INIT_7C => X"0000003c000000000000001e00000000ffffff97ffffffffffffffe2ffffffff",
            INIT_7D => X"ffffffe8ffffffff000000080000000000000076000000000000002200000000",
            INIT_7E => X"ffffffabffffffff0000001c00000000ffffffddffffffffffffffa4ffffffff",
            INIT_7F => X"000000c0000000000000001800000000ffffff92ffffffff0000008b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE10;


    MEM_IWGHT_LAYER2_INSTANCE11 : if BRAM_NAME = "iwght_layer2_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000049000000000000002f000000000000009700000000fffffffaffffffff",
            INIT_01 => X"ffffff86ffffffff000000cc00000000ffffffb9ffffffffffffffa2ffffffff",
            INIT_02 => X"0000006600000000ffffffe6ffffffffffffff86fffffffffffffff5ffffffff",
            INIT_03 => X"00000001000000000000003f00000000ffffffc6ffffffffffffff57ffffffff",
            INIT_04 => X"0000003700000000ffffff26ffffffff000000d700000000000000bb00000000",
            INIT_05 => X"fffffffdffffffff0000000000000000ffffffffffffffff0000003d00000000",
            INIT_06 => X"fffffff2fffffffffffffffffffffffffffffffbffffffff0000001300000000",
            INIT_07 => X"ffffff69ffffffff0000000500000000ffffffedfffffffffffffffbffffffff",
            INIT_08 => X"ffffffb5ffffffffffffffd9ffffffffffffffc6ffffffff0000005700000000",
            INIT_09 => X"ffffffdcffffffff0000000700000000fffffffbffffffff0000005600000000",
            INIT_0A => X"ffffffc9ffffffff0000008000000000ffffffeaffffffffffffff33ffffffff",
            INIT_0B => X"ffffffeaffffffffffffffceffffffffffffffbdffffffff0000005000000000",
            INIT_0C => X"ffffff08ffffffff0000001f000000000000009d000000000000005600000000",
            INIT_0D => X"0000004900000000ffffffabffffffff000000c200000000000000a900000000",
            INIT_0E => X"0000002f00000000ffffffeeffffffff0000007c00000000000000cb00000000",
            INIT_0F => X"0000004100000000ffffff3dffffffff0000004100000000000000ec00000000",
            INIT_10 => X"ffffff97ffffffffffffff45ffffffffffffffacffffffff0000007b00000000",
            INIT_11 => X"000000a90000000000000013000000000000009a00000000ffffffc9ffffffff",
            INIT_12 => X"ffffffa2ffffffffffffffbcffffffffffffffd4ffffffffffffffadffffffff",
            INIT_13 => X"0000003a00000000fffffff0ffffffff0000001c000000000000001f00000000",
            INIT_14 => X"000000090000000000000016000000000000003500000000fffffffdffffffff",
            INIT_15 => X"0000003400000000ffffff33ffffffff0000003400000000ffffff88ffffffff",
            INIT_16 => X"0000004f00000000ffffffbeffffffffffffffa7ffffffffffffffafffffffff",
            INIT_17 => X"000000670000000000000084000000000000000800000000ffffffd9ffffffff",
            INIT_18 => X"0000002800000000ffffffa8ffffffff00000062000000000000008500000000",
            INIT_19 => X"ffffffecffffffff0000009a00000000ffffff71ffffffffffffff93ffffffff",
            INIT_1A => X"000000890000000000000033000000000000007e000000000000008200000000",
            INIT_1B => X"ffffffe3fffffffffffffff8ffffffff00000015000000000000000d00000000",
            INIT_1C => X"fffffffbffffffff0000005a00000000ffffff88ffffffff0000004f00000000",
            INIT_1D => X"0000002000000000ffffff91ffffffffffffff73ffffffff0000000f00000000",
            INIT_1E => X"0000002e00000000fffffff8ffffffff000000b9000000000000003000000000",
            INIT_1F => X"00000018000000000000003100000000ffffffd0ffffffffffffffafffffffff",
            INIT_20 => X"0000001f00000000ffffff3dffffffffffffffbaffffffffffffff5bffffffff",
            INIT_21 => X"ffffffc1ffffffff000000060000000000000026000000000000006400000000",
            INIT_22 => X"ffffffe0ffffffffffffffd9ffffffffffffffeaffffffff0000004700000000",
            INIT_23 => X"0000007e00000000ffffffaeffffffff0000004200000000ffffff5fffffffff",
            INIT_24 => X"fffffecaffffffff0000001c000000000000001a000000000000007500000000",
            INIT_25 => X"ffffff25ffffffff00000053000000000000001a00000000ffffff5cffffffff",
            INIT_26 => X"ffffff64ffffffffffffffe4ffffffffffffffa0ffffffffffffff33ffffffff",
            INIT_27 => X"ffffffaeffffffff0000003300000000000000cf000000000000002400000000",
            INIT_28 => X"0000002b000000000000000800000000ffffffdfffffffffffffffc4ffffffff",
            INIT_29 => X"0000005f00000000ffffffa0ffffffffffffffe0ffffffff0000003c00000000",
            INIT_2A => X"ffffffadffffffffffffffa2ffffffffffffffacffffffffffffff87ffffffff",
            INIT_2B => X"00000010000000000000004a000000000000008700000000ffffffb0ffffffff",
            INIT_2C => X"0000005600000000000000160000000000000035000000000000003600000000",
            INIT_2D => X"ffffffdfffffffffffffffe3ffffffff0000009b000000000000001100000000",
            INIT_2E => X"0000008100000000ffffffa8ffffffff0000002300000000ffffffd4ffffffff",
            INIT_2F => X"ffffffddffffffff0000007f0000000000000002000000000000006f00000000",
            INIT_30 => X"00000055000000000000002d0000000000000074000000000000003e00000000",
            INIT_31 => X"0000005600000000ffffffa5ffffffff0000008a000000000000006600000000",
            INIT_32 => X"fffffff2ffffffff0000001c000000000000008300000000ffffffceffffffff",
            INIT_33 => X"000000a800000000000000870000000000000092000000000000008a00000000",
            INIT_34 => X"0000001f000000000000002f000000000000002800000000000000a200000000",
            INIT_35 => X"ffffff9affffffff0000000800000000ffffff99ffffffffffffff46ffffffff",
            INIT_36 => X"ffffffabfffffffffffffed9ffffffff000000d2000000000000007a00000000",
            INIT_37 => X"000000da000000000000001800000000ffffff3cffffffffffffff94ffffffff",
            INIT_38 => X"0000008600000000ffffffebffffffff00000079000000000000008b00000000",
            INIT_39 => X"ffffffceffffffff00000073000000000000007b00000000ffffffacffffffff",
            INIT_3A => X"ffffff3effffffff0000003c000000000000002f000000000000009800000000",
            INIT_3B => X"fffffff9ffffffff000000020000000000000087000000000000009500000000",
            INIT_3C => X"ffffff4bffffffffffffffbeffffffffffffffb0ffffffff0000004300000000",
            INIT_3D => X"fffffff7ffffffffffffffdcfffffffffffffe76ffffffffffffffeeffffffff",
            INIT_3E => X"ffffff72fffffffffffffffaffffffff0000001200000000ffffffe7ffffffff",
            INIT_3F => X"fffffe97ffffffff0000002900000000fffffed1ffffffff0000006300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008f00000000ffffff46ffffffff0000000200000000ffffff05ffffffff",
            INIT_41 => X"0000008f0000000000000019000000000000000f000000000000005c00000000",
            INIT_42 => X"ffffffa2ffffffff0000001a0000000000000061000000000000004d00000000",
            INIT_43 => X"0000004d00000000fffffef0ffffffffffffffa1ffffffffffffffb4ffffffff",
            INIT_44 => X"0000001c000000000000002e00000000000000b200000000ffffffb2ffffffff",
            INIT_45 => X"ffffff90ffffffff00000005000000000000005000000000ffffffceffffffff",
            INIT_46 => X"ffffffa9ffffffff0000001800000000ffffffacffffffffffffff36ffffffff",
            INIT_47 => X"0000007e00000000ffffffa4ffffffff0000005700000000ffffffe9ffffffff",
            INIT_48 => X"fffffff5ffffffff000000a9000000000000003000000000ffffff97ffffffff",
            INIT_49 => X"00000000000000000000005700000000ffffffedffffffffffffff9dffffffff",
            INIT_4A => X"0000000b000000000000000900000000ffffffa6ffffffffffffffedffffffff",
            INIT_4B => X"000000000000000000000049000000000000007400000000ffffffe2ffffffff",
            INIT_4C => X"ffffff89ffffffffffffff4cffffffffffffff2cffffffff0000000400000000",
            INIT_4D => X"00000000000000000000000c0000000000000011000000000000006000000000",
            INIT_4E => X"fffffff8ffffffff0000000900000000fffffff1ffffffff0000000400000000",
            INIT_4F => X"000000d4000000000000000a00000000fffffffaffffffffffffffedffffffff",
            INIT_50 => X"ffffffabffffffffffffffe0ffffffff0000008c000000000000005b00000000",
            INIT_51 => X"ffffff7effffffffffffff53ffffffffffffff1fffffffffffffff7effffffff",
            INIT_52 => X"0000000a00000000fffffffeffffffffffffffebfffffffffffffeb1ffffffff",
            INIT_53 => X"0000007b00000000000000560000000000000095000000000000007900000000",
            INIT_54 => X"ffffff00ffffffffffffffcaffffffffffffffd0ffffffff0000005800000000",
            INIT_55 => X"00000033000000000000003200000000ffffffd9ffffffffffffff92ffffffff",
            INIT_56 => X"ffffff76ffffffffffffff96ffffffff0000007700000000ffffffc9ffffffff",
            INIT_57 => X"ffffffa6ffffffffffffffa0ffffffffffffffb1ffffffff0000002c00000000",
            INIT_58 => X"0000004200000000ffffffe6ffffffff00000056000000000000008000000000",
            INIT_59 => X"0000007100000000ffffffebffffffffffffff94ffffffffffffff5dffffffff",
            INIT_5A => X"0000000a000000000000003f00000000ffffff9fffffffff0000001f00000000",
            INIT_5B => X"0000004100000000ffffffa6ffffffff0000003a00000000ffffff58ffffffff",
            INIT_5C => X"ffffffecffffffff0000008100000000ffffff4effffffff0000008800000000",
            INIT_5D => X"ffffffa9fffffffffffffffbffffffff0000006200000000ffffff7affffffff",
            INIT_5E => X"ffffff9bffffffff00000042000000000000004200000000ffffff05ffffffff",
            INIT_5F => X"0000004300000000ffffff50fffffffffffffff1ffffffff0000007000000000",
            INIT_60 => X"ffffff55ffffffff000000830000000000000009000000000000001200000000",
            INIT_61 => X"ffffffa0ffffffff00000077000000000000007400000000ffffffecffffffff",
            INIT_62 => X"ffffff62ffffffffffffff74ffffffffffffffd8fffffffffffffffaffffffff",
            INIT_63 => X"ffffff78ffffffffffffffb9ffffffffffffffddffffffff0000004500000000",
            INIT_64 => X"000000ba000000000000004400000000ffffffe0ffffffffffffffa7ffffffff",
            INIT_65 => X"ffffffe4ffffffff0000001400000000fffffff6ffffffffffffffd9ffffffff",
            INIT_66 => X"ffffffedffffffffffffffdaffffffffffffff9cffffffffffffff70ffffffff",
            INIT_67 => X"000000ff00000000000000c70000000000000068000000000000001e00000000",
            INIT_68 => X"ffffff3effffffff0000004e0000000000000004000000000000011000000000",
            INIT_69 => X"000000da000000000000000700000000ffffff6effffffffffffff32ffffffff",
            INIT_6A => X"00000070000000000000005f0000000000000011000000000000002b00000000",
            INIT_6B => X"ffffffd2ffffffffffffffefffffffffffffffb5ffffffff0000004500000000",
            INIT_6C => X"00000080000000000000008e00000000ffffffb4ffffffffffffffe4ffffffff",
            INIT_6D => X"000000a500000000ffffffc1ffffffff00000062000000000000009500000000",
            INIT_6E => X"0000000400000000ffffff73ffffffffffffffe4ffffffffffffffe5ffffffff",
            INIT_6F => X"0000004200000000fffffffaffffffff00000007000000000000008200000000",
            INIT_70 => X"0000006100000000ffffffa7ffffffffffffffbfffffffffffffff66ffffffff",
            INIT_71 => X"0000000c000000000000005900000000000000b0000000000000000500000000",
            INIT_72 => X"0000001c00000000ffffff6bffffffff0000000b000000000000003a00000000",
            INIT_73 => X"fffffeedffffffffffffff9bffffffff00000019000000000000002e00000000",
            INIT_74 => X"00000012000000000000000d000000000000001000000000ffffff84ffffffff",
            INIT_75 => X"ffffffefffffffff000000c300000000ffffff86ffffffffffffffe1ffffffff",
            INIT_76 => X"ffffffa7fffffffffffffff0fffffffffffffff4ffffffffffffffe7ffffffff",
            INIT_77 => X"000000220000000000000024000000000000006f000000000000002500000000",
            INIT_78 => X"fffffff5fffffffffffffffeffffffff0000001100000000fffffff9ffffffff",
            INIT_79 => X"ffffffe6fffffffffffffffeffffffff0000000300000000ffffffefffffffff",
            INIT_7A => X"ffffffeaffffffff0000000700000000ffffffe6fffffffffffffffeffffffff",
            INIT_7B => X"0000000200000000ffffffebfffffffffffffff5ffffffff0000000b00000000",
            INIT_7C => X"0000000100000000fffffffeffffffffffffffffffffffffffffffe0ffffffff",
            INIT_7D => X"00000003000000000000000d00000000fffffffbfffffffffffffffeffffffff",
            INIT_7E => X"ffffffe4ffffffff0000000200000000fffffff7fffffffffffffff8ffffffff",
            INIT_7F => X"fffffff6ffffffff0000000700000000fffffffaffffffff0000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE11;


    MEM_IWGHT_LAYER2_INSTANCE12 : if BRAM_NAME = "iwght_layer2_instance12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff4ffffffff00000004000000000000000200000000fffffff9ffffffff",
            INIT_01 => X"fffffff2ffffffffffffffe8ffffffffffffffffffffffff0000000e00000000",
            INIT_02 => X"0000000b00000000fffffff8ffffffffffffffefffffffffffffffffffffffff",
            INIT_03 => X"ffffffefffffffffffffffecffffffffffffffe7ffffffff0000000e00000000",
            INIT_04 => X"ffffffecffffffff0000000000000000fffffffdfffffffffffffffeffffffff",
            INIT_05 => X"fffffff6fffffffffffffffdffffffff0000000200000000ffffffe4ffffffff",
            INIT_06 => X"ffffffeafffffffffffffff5ffffffffffffffe1ffffffff0000000200000000",
            INIT_07 => X"0000000600000000ffffffe7ffffffff00000012000000000000000000000000",
            INIT_08 => X"0000000300000000fffffff8ffffffff0000000a00000000ffffffeaffffffff",
            INIT_09 => X"0000000200000000ffffffeeffffffff00000003000000000000001100000000",
            INIT_0A => X"fffffffcffffffff0000000d0000000000000005000000000000000300000000",
            INIT_0B => X"fffffffdffffffffffffffe9fffffffffffffff9fffffffffffffff8ffffffff",
            INIT_0C => X"fffffff3fffffffffffffff4ffffffffffffffebffffffffffffffebffffffff",
            INIT_0D => X"fffffff5ffffffffffffffeeffffffff0000000000000000fffffffaffffffff",
            INIT_0E => X"fffffffcfffffffffffffffaffffffff0000000000000000ffffffe8ffffffff",
            INIT_0F => X"0000000700000000ffffffebfffffffffffffff1fffffffffffffff2ffffffff",
            INIT_10 => X"0000000300000000ffffffe9ffffffff0000000b00000000fffffff4ffffffff",
            INIT_11 => X"ffffffeaffffffffffffffeffffffffffffffff6ffffffff0000000000000000",
            INIT_12 => X"fffffff3ffffffff0000000b00000000fffffff4fffffffffffffff6ffffffff",
            INIT_13 => X"fffffff1fffffffffffffff7fffffffffffffff9ffffffff0000000400000000",
            INIT_14 => X"0000000c00000000ffffffddffffffff0000000900000000fffffff0ffffffff",
            INIT_15 => X"00000004000000000000000e00000000fffffffdfffffffffffffff2ffffffff",
            INIT_16 => X"ffffffefffffffff0000000800000000fffffff9ffffffff0000000e00000000",
            INIT_17 => X"fffffff5ffffffff0000000000000000ffffffedffffffff0000000f00000000",
            INIT_18 => X"fffffffcffffffff0000000500000000fffffff9fffffffffffffffbffffffff",
            INIT_19 => X"ffffffe5fffffffffffffffbffffffffffffffefffffffff0000000e00000000",
            INIT_1A => X"0000000000000000ffffffe7fffffffffffffffdfffffffffffffff6ffffffff",
            INIT_1B => X"ffffffebfffffffffffffff3ffffffffffffffe6ffffffff0000000700000000",
            INIT_1C => X"fffffff9fffffffffffffff2ffffffffffffffffffffffffffffffeaffffffff",
            INIT_1D => X"fffffffcffffffff0000000000000000fffffffdfffffffffffffffcffffffff",
            INIT_1E => X"fffffffdffffffffffffffebffffffff00000005000000000000000000000000",
            INIT_1F => X"0000001300000000ffffffffffffffff0000000f000000000000000000000000",
            INIT_20 => X"0000000000000000fffffffdffffffff0000000b000000000000000600000000",
            INIT_21 => X"ffffffedffffffffffffffe8fffffffffffffff2fffffffffffffff6ffffffff",
            INIT_22 => X"0000000000000000fffffffdfffffffffffffff9ffffffff0000000100000000",
            INIT_23 => X"fffffff5fffffffffffffff4ffffffff00000000000000000000000700000000",
            INIT_24 => X"fffffffbffffffff0000000100000000ffffffeffffffffffffffff7ffffffff",
            INIT_25 => X"0000000000000000fffffffbffffffff0000000000000000fffffff8ffffffff",
            INIT_26 => X"ffffffedffffffffffffffe8fffffffffffffff2ffffffff0000000700000000",
            INIT_27 => X"fffffff5fffffffffffffffaffffffff00000003000000000000000a00000000",
            INIT_28 => X"0000000a00000000ffffffeefffffffffffffff8fffffffffffffff6ffffffff",
            INIT_29 => X"0000000a00000000ffffffe8ffffffffffffffe7ffffffffffffffefffffffff",
            INIT_2A => X"fffffffefffffffffffffffefffffffffffffffafffffffffffffffaffffffff",
            INIT_2B => X"ffffffeaffffffffffffffeefffffffffffffff5ffffffffffffffffffffffff",
            INIT_2C => X"fffffff3ffffffffffffffe8fffffffffffffff1ffffffffffffffecffffffff",
            INIT_2D => X"fffffffcffffffff0000000100000000fffffff7fffffffffffffffeffffffff",
            INIT_2E => X"fffffff5fffffffffffffff7ffffffffffffffecffffffff0000000300000000",
            INIT_2F => X"fffffff9ffffffff0000000200000000ffffffffffffffff0000001300000000",
            INIT_30 => X"00000008000000000000000100000000fffffff2ffffffffffffffeaffffffff",
            INIT_31 => X"ffffffe6ffffffff000000050000000000000008000000000000000c00000000",
            INIT_32 => X"00000000000000000000000000000000fffffff9ffffffff0000000a00000000",
            INIT_33 => X"ffffffe4fffffffffffffffdffffffffffffffe4ffffffffffffffe9ffffffff",
            INIT_34 => X"00000003000000000000000100000000fffffff4ffffffff0000000000000000",
            INIT_35 => X"fffffffcfffffffffffffffaffffffff0000000700000000fffffff1ffffffff",
            INIT_36 => X"fffffffefffffffffffffff6ffffffffffffffecffffffff0000000000000000",
            INIT_37 => X"00000000000000000000000600000000fffffff5ffffffffffffffffffffffff",
            INIT_38 => X"ffffffeeffffffff00000002000000000000000800000000fffffff4ffffffff",
            INIT_39 => X"0000000700000000000000030000000000000006000000000000000000000000",
            INIT_3A => X"ffffffedffffffff0000000a0000000000000001000000000000000100000000",
            INIT_3B => X"000000140000000000000011000000000000000000000000ffffffe5ffffffff",
            INIT_3C => X"0000000500000000fffffffdfffffffffffffff2ffffffffffffffeaffffffff",
            INIT_3D => X"00000007000000000000000000000000fffffff1ffffffffffffffefffffffff",
            INIT_3E => X"ffffffe0ffffffff0000000900000000ffffffe3fffffffffffffff3ffffffff",
            INIT_3F => X"fffffff8fffffffffffffff6ffffffffffffffdfffffffff0000000400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffffffffffffffffff9dffffffffffffff84ffffffff0000002100000000",
            INIT_41 => X"ffffff92ffffffffffffffe2ffffffff0000000100000000ffffffbaffffffff",
            INIT_42 => X"fffffff2ffffffff000000ab00000000fffffff2ffffffffffffffdcffffffff",
            INIT_43 => X"ffffffefffffffff0000002e000000000000003a00000000ffffff75ffffffff",
            INIT_44 => X"0000004e000000000000004c00000000ffffff3affffffffffffffa6ffffffff",
            INIT_45 => X"0000004b000000000000002c000000000000000f00000000ffffffd6ffffffff",
            INIT_46 => X"ffffff7effffffff0000006100000000ffffff85ffffffff0000000000000000",
            INIT_47 => X"00000064000000000000002f00000000ffffffb5ffffffff0000008600000000",
            INIT_48 => X"ffffff45ffffffffffffffe1ffffffff0000000d000000000000002600000000",
            INIT_49 => X"ffffffd3ffffffffffffffefffffffff00000001000000000000001000000000",
            INIT_4A => X"0000008e00000000ffffffa4ffffffffffffff8fffffffff0000002000000000",
            INIT_4B => X"ffffff81ffffffff000000070000000000000000000000000000007500000000",
            INIT_4C => X"fffffff2ffffffffffffffe6ffffffff00000007000000000000008a00000000",
            INIT_4D => X"ffffffb9ffffffffffffffd1ffffffff00000051000000000000000800000000",
            INIT_4E => X"0000001b000000000000001100000000fffffeddffffffff0000005300000000",
            INIT_4F => X"0000002e000000000000005400000000000000c900000000ffffff40ffffffff",
            INIT_50 => X"000000dd000000000000006600000000ffffffefffffffff0000005a00000000",
            INIT_51 => X"ffffffc9ffffffffffffffb8ffffffffffffffd0ffffffff0000000700000000",
            INIT_52 => X"ffffff71ffffffffffffff24ffffffff0000001000000000ffffff9bffffffff",
            INIT_53 => X"ffffff75ffffffffffffffd3ffffffff00000048000000000000000900000000",
            INIT_54 => X"ffffffaefffffffffffffed2ffffffffffffffddffffffff0000008200000000",
            INIT_55 => X"fffffff0ffffffffffffff52ffffffffffffffaaffffffff0000002900000000",
            INIT_56 => X"ffffffe1ffffffffffffffc2ffffffff000000a5000000000000007500000000",
            INIT_57 => X"ffffffcafffffffffffffffdffffffff0000000a00000000000000c800000000",
            INIT_58 => X"ffffffafffffffff0000000b0000000000000038000000000000001300000000",
            INIT_59 => X"00000083000000000000009800000000ffffffcaffffffff0000007e00000000",
            INIT_5A => X"0000001100000000ffffff57ffffffffffffff30ffffffff0000001600000000",
            INIT_5B => X"0000001400000000ffffff4cfffffffffffffecaffffffff0000002900000000",
            INIT_5C => X"0000010000000000000000a000000000ffffffa7ffffffff0000000800000000",
            INIT_5D => X"fffffff9fffffffffffffffaffffffff0000000c000000000000001200000000",
            INIT_5E => X"00000014000000000000000900000000ffffffebffffffff0000000d00000000",
            INIT_5F => X"ffffff6affffffffffffffa2ffffffffffffffffffffffff0000000600000000",
            INIT_60 => X"00000056000000000000002600000000ffffffc0ffffffffffffff98ffffffff",
            INIT_61 => X"ffffffafffffffffffffffb9ffffffffffffff97fffffffffffffffeffffffff",
            INIT_62 => X"0000000000000000ffffff90ffffffffffffff5dffffffff000000fc00000000",
            INIT_63 => X"ffffff46fffffffffffffed8ffffffff0000002000000000ffffffe8ffffffff",
            INIT_64 => X"0000002900000000fffffff9ffffffff0000005d000000000000003f00000000",
            INIT_65 => X"0000003900000000000000050000000000000085000000000000003b00000000",
            INIT_66 => X"ffffff48ffffffffffffff3bffffffffffffffceffffffffffffffe7ffffffff",
            INIT_67 => X"0000003800000000ffffff93ffffffff0000016e00000000ffffff7fffffffff",
            INIT_68 => X"0000003a00000000ffffff71ffffffff000000b300000000ffffff7dffffffff",
            INIT_69 => X"ffffff5affffffff0000000d00000000ffffff41ffffffffffffffe8ffffffff",
            INIT_6A => X"ffffffb2ffffffffffffff2fffffffff0000003f00000000ffffffe8ffffffff",
            INIT_6B => X"0000003400000000ffffffc5fffffffffffffff5ffffffff0000004300000000",
            INIT_6C => X"ffffffe8ffffffff0000004200000000ffffff5dffffffff0000005400000000",
            INIT_6D => X"00000073000000000000003b00000000000000af000000000000003400000000",
            INIT_6E => X"ffffff5cffffffffffffffc3ffffffff00000003000000000000003d00000000",
            INIT_6F => X"ffffff26ffffffffffffff5fffffffffffffff25ffffffffffffff85ffffffff",
            INIT_70 => X"0000000500000000ffffffa4ffffffff000000dc00000000ffffffc9ffffffff",
            INIT_71 => X"ffffffcaffffffff0000005700000000ffffffe2ffffffff0000000b00000000",
            INIT_72 => X"ffffffaaffffffff00000029000000000000003600000000000000d200000000",
            INIT_73 => X"ffffffddffffffff0000005a000000000000004300000000ffffffb3ffffffff",
            INIT_74 => X"00000065000000000000007600000000ffffff04ffffffffffffffabffffffff",
            INIT_75 => X"000000120000000000000008000000000000005400000000ffffffd7ffffffff",
            INIT_76 => X"ffffff84ffffffff0000005c000000000000002e00000000ffffff51ffffffff",
            INIT_77 => X"000000360000000000000045000000000000007a000000000000004e00000000",
            INIT_78 => X"ffffffecffffffff0000005c00000000fffffff3ffffffff0000002a00000000",
            INIT_79 => X"ffffffc5ffffffff0000004100000000ffffff79fffffffffffffff5ffffffff",
            INIT_7A => X"000000f90000000000000011000000000000008400000000ffffffcfffffffff",
            INIT_7B => X"0000006d000000000000004800000000ffffffc5ffffffff0000002000000000",
            INIT_7C => X"0000005e00000000ffffff52fffffffffffffe6affffffffffffffa9ffffffff",
            INIT_7D => X"ffffffe1ffffffff0000006f00000000ffffff89ffffffffffffff11ffffffff",
            INIT_7E => X"0000006900000000ffffffe1ffffffff0000007700000000ffffff74ffffffff",
            INIT_7F => X"0000000600000000fffffec6ffffffffffffff39ffffffffffffff20ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE12;


    MEM_IWGHT_LAYER2_INSTANCE13 : if BRAM_NAME = "iwght_layer2_instance13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007f00000000000000ec00000000ffffffd4ffffffffffffff28ffffffff",
            INIT_01 => X"ffffffc1ffffffffffffff1bffffffff0000004c000000000000005c00000000",
            INIT_02 => X"00000008000000000000003f0000000000000079000000000000005300000000",
            INIT_03 => X"ffffff86fffffffffffffff3ffffffff0000004500000000ffffff7dffffffff",
            INIT_04 => X"ffffff9fffffffff0000009600000000000000be00000000fffffe99ffffffff",
            INIT_05 => X"0000005f0000000000000007000000000000008600000000ffffff9affffffff",
            INIT_06 => X"000000df00000000ffffff64ffffffffffffffaffffffffffffffeb3ffffffff",
            INIT_07 => X"0000005a00000000000000fd00000000ffffff7fffffffff0000000a00000000",
            INIT_08 => X"00000043000000000000002b00000000ffffffb6ffffffff0000003e00000000",
            INIT_09 => X"ffffffc5ffffffffffffffbdffffffff000000c3000000000000002000000000",
            INIT_0A => X"0000004400000000ffffffd4ffffffff0000003b000000000000009900000000",
            INIT_0B => X"ffffffb6ffffffffffffffc3ffffffff00000031000000000000002900000000",
            INIT_0C => X"ffffffe8ffffffff0000002e000000000000008200000000ffffffecffffffff",
            INIT_0D => X"ffffff19ffffffff00000037000000000000003600000000ffffffd9ffffffff",
            INIT_0E => X"00000127000000000000003a00000000ffffff80ffffffffffffff57ffffffff",
            INIT_0F => X"0000004a00000000fffffee8ffffffffffffffbcffffffffffffff73ffffffff",
            INIT_10 => X"ffffff85ffffffff00000069000000000000007600000000ffffffbbffffffff",
            INIT_11 => X"ffffffc0fffffffffffffffeffffffffffffff57ffffffff0000007400000000",
            INIT_12 => X"000000040000000000000010000000000000000900000000ffffff56ffffffff",
            INIT_13 => X"ffffff68fffffffffffffe97ffffffffffffff98fffffffffffffff8ffffffff",
            INIT_14 => X"0000007200000000ffffffdcffffffffffffff8bffffffff0000007d00000000",
            INIT_15 => X"ffffff95ffffffffffffff80ffffffffffffffa1ffffffffffffffc4ffffffff",
            INIT_16 => X"ffffff91ffffffff0000002a00000000ffffff0bffffffff0000004800000000",
            INIT_17 => X"0000011500000000ffffff6fffffffffffffffc2ffffffff0000005400000000",
            INIT_18 => X"0000002700000000000000a000000000ffffffb0ffffffffffffffdfffffffff",
            INIT_19 => X"0000003700000000ffffffe2ffffffff00000099000000000000007a00000000",
            INIT_1A => X"ffffffd0ffffffffffffffc3ffffffffffffffa6ffffffff0000003f00000000",
            INIT_1B => X"ffffffcfffffffffffffff70ffffffffffffffbeffffffffffffff89ffffffff",
            INIT_1C => X"000000430000000000000028000000000000005900000000ffffffb7ffffffff",
            INIT_1D => X"ffffff8affffffff000000630000000000000043000000000000000600000000",
            INIT_1E => X"0000001900000000000000b000000000ffffff8dffffffff0000004400000000",
            INIT_1F => X"fffffff9ffffffff0000006d000000000000000300000000000000b400000000",
            INIT_20 => X"ffffffcfffffffff000000450000000000000019000000000000001900000000",
            INIT_21 => X"ffffff5bfffffffffffffff1ffffffff0000000000000000ffffffe7ffffffff",
            INIT_22 => X"fffffffcffffffff00000017000000000000003c00000000000000c500000000",
            INIT_23 => X"ffffffecffffffff0000003b0000000000000024000000000000002b00000000",
            INIT_24 => X"000000b900000000000000a5000000000000009600000000000000f500000000",
            INIT_25 => X"0000000400000000ffffffecffffffff0000000300000000ffffffdfffffffff",
            INIT_26 => X"fffffff7ffffffff00000017000000000000000000000000ffffffe2ffffffff",
            INIT_27 => X"ffffffc9ffffffff0000009b00000000ffffffe8fffffffffffffffaffffffff",
            INIT_28 => X"ffffffc5ffffffffffffff8affffffffffffff7effffffff0000007d00000000",
            INIT_29 => X"fffffff1ffffffff0000004b00000000ffffff54ffffffffffffff8dffffffff",
            INIT_2A => X"0000005e00000000ffffffe1ffffffffffffff42ffffffff0000007c00000000",
            INIT_2B => X"ffffffddffffffff0000008200000000ffffff7dffffffff0000002a00000000",
            INIT_2C => X"ffffff5fffffffffffffffaaffffffffffffff82fffffffffffffeb5ffffffff",
            INIT_2D => X"0000003400000000ffffff1fffffffffffffffaeffffffffffffff70ffffffff",
            INIT_2E => X"fffffff7ffffffff0000007a00000000ffffff79ffffffff0000001500000000",
            INIT_2F => X"0000005900000000ffffff6cffffffff0000007f00000000ffffffbeffffffff",
            INIT_30 => X"0000002c00000000ffffff84ffffffff000000b7000000000000000700000000",
            INIT_31 => X"000000c30000000000000067000000000000000200000000ffffff20ffffffff",
            INIT_32 => X"ffffffe7ffffffff0000003100000000ffffffe8ffffffff0000006c00000000",
            INIT_33 => X"000000cf00000000ffffffc9ffffffffffffffeaffffffff000000a800000000",
            INIT_34 => X"0000004100000000fffffef8ffffffff000000d9000000000000007800000000",
            INIT_35 => X"ffffff2effffffff0000001e00000000ffffff02ffffffffffffff90ffffffff",
            INIT_36 => X"0000003600000000fffffffcffffffffffffffe8ffffffff0000011000000000",
            INIT_37 => X"ffffffc2ffffffffffffff72ffffffff0000010e00000000ffffffcaffffffff",
            INIT_38 => X"000000730000000000000095000000000000001000000000fffffeedffffffff",
            INIT_39 => X"ffffff91ffffffff000000b900000000000000c100000000ffffff38ffffffff",
            INIT_3A => X"ffffffb8ffffffffffffff7dffffffffffffffd9ffffffff0000000400000000",
            INIT_3B => X"0000006100000000fffffd61ffffffff0000007500000000ffffff6fffffffff",
            INIT_3C => X"0000006000000000ffffffe1ffffffffffffff95fffffffffffffffbffffffff",
            INIT_3D => X"0000005500000000ffffff99ffffffff0000008200000000ffffffc1ffffffff",
            INIT_3E => X"ffffffe9ffffffffffffffe9ffffffffffffff21ffffffffffffffafffffffff",
            INIT_3F => X"ffffffaeffffffff000000c80000000000000095000000000000001a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffdf8fffffffffffffff7fffffffffffffed7ffffffffffffffb1ffffffff",
            INIT_41 => X"00000023000000000000008600000000ffffffbbffffffffffffff68ffffffff",
            INIT_42 => X"ffffffb0ffffffff00000002000000000000006e00000000ffffff60ffffffff",
            INIT_43 => X"ffffffd0ffffffff0000004d00000000ffffff5fffffffffffffff72ffffffff",
            INIT_44 => X"0000001000000000000000a300000000000000c2000000000000003d00000000",
            INIT_45 => X"ffffff3fffffffffffffffe6ffffffffffffff0bffffffff0000000600000000",
            INIT_46 => X"fffffffeffffffffffffffdbffffffff0000002c00000000fffffecfffffffff",
            INIT_47 => X"ffffff8bffffffffffffff5ffffffffffffffff6ffffffffffffff05ffffffff",
            INIT_48 => X"000000b100000000ffffffb6ffffffffffffffe2fffffffffffffee3ffffffff",
            INIT_49 => X"0000005600000000000000c6000000000000006400000000fffffe8affffffff",
            INIT_4A => X"0000002d0000000000000050000000000000001f000000000000003a00000000",
            INIT_4B => X"ffffff93fffffffffffffeb0ffffffff00000042000000000000001600000000",
            INIT_4C => X"0000003700000000fffffef1ffffffffffffff0effffffff0000004b00000000",
            INIT_4D => X"ffffff5fffffffff0000005a00000000fffffff9ffffffffffffffc4ffffffff",
            INIT_4E => X"fffffffbffffffffffffffe4ffffffff000000a2000000000000005e00000000",
            INIT_4F => X"0000000100000000ffffff6cffffffffffffffcbffffffff0000005900000000",
            INIT_50 => X"0000003b000000000000003000000000ffffff53ffffffff0000007000000000",
            INIT_51 => X"0000003700000000ffffff56fffffffffffffff9ffffffffffffff99ffffffff",
            INIT_52 => X"ffffffceffffffff0000003f00000000ffffff66ffffffff0000001100000000",
            INIT_53 => X"0000012e00000000ffffff4bffffffff0000003300000000ffffffc9ffffffff",
            INIT_54 => X"0000001b00000000000000220000000000000076000000000000002b00000000",
            INIT_55 => X"0000002700000000fffffff4ffffffffffffff9bffffffffffffff25ffffffff",
            INIT_56 => X"00000001000000000000001e0000000000000060000000000000008000000000",
            INIT_57 => X"ffffffa6ffffffffffffff78ffffffff0000009b00000000ffffffcdffffffff",
            INIT_58 => X"ffffff85ffffffff0000001800000000ffffffc2ffffffff0000000400000000",
            INIT_59 => X"0000003000000000ffffffacffffffff00000000000000000000007800000000",
            INIT_5A => X"ffffff63ffffffff0000001500000000ffffff4affffffffffffff94ffffffff",
            INIT_5B => X"ffffffc0ffffffffffffffc6ffffffff00000081000000000000002600000000",
            INIT_5C => X"0000008600000000ffffff85ffffffff00000023000000000000000d00000000",
            INIT_5D => X"0000007f000000000000003400000000ffffff7dffffffffffffffaeffffffff",
            INIT_5E => X"ffffffc9ffffffffffffffdcffffffffffffffd8ffffffffffffff45ffffffff",
            INIT_5F => X"0000001000000000ffffffb8ffffffffffffffc9ffffffff0000000100000000",
            INIT_60 => X"ffffffb1ffffffffffffffb5ffffffffffffff8dffffffffffffff40ffffffff",
            INIT_61 => X"0000001500000000ffffffb5fffffffffffffff5ffffffff0000000200000000",
            INIT_62 => X"ffffff7affffffffffffffaaffffffffffffff92ffffffff0000001200000000",
            INIT_63 => X"000000b700000000000000b6000000000000001400000000ffffff8affffffff",
            INIT_64 => X"0000001300000000ffffff78ffffffff0000009200000000ffffffcfffffffff",
            INIT_65 => X"000000b800000000ffffff7fffffffffffffffe4ffffffffffffffaaffffffff",
            INIT_66 => X"fffffff5fffffffffffffff8ffffffff00000044000000000000002500000000",
            INIT_67 => X"000000d600000000000000580000000000000011000000000000004800000000",
            INIT_68 => X"ffffff1dffffffff0000000100000000ffffff98ffffffff0000004000000000",
            INIT_69 => X"fffffff8ffffffffffffffe0fffffffffffffff5fffffffffffffff8ffffffff",
            INIT_6A => X"0000002800000000000000900000000000000072000000000000002b00000000",
            INIT_6B => X"000000810000000000000033000000000000008100000000fffffff7ffffffff",
            INIT_6C => X"0000004100000000ffffffe5ffffffff0000002d000000000000004500000000",
            INIT_6D => X"fffffff9fffffffffffffffcfffffffffffffff6ffffffffffffffcfffffffff",
            INIT_6E => X"fffffff2ffffffff0000001100000000fffffffaffffffff0000000000000000",
            INIT_6F => X"ffffff8affffffffffffff77ffffffff00000000000000000000000000000000",
            INIT_70 => X"ffffff9effffffffffffffe5ffffffff0000004700000000ffffffd1ffffffff",
            INIT_71 => X"ffffffb0ffffffff0000003d000000000000000e000000000000004e00000000",
            INIT_72 => X"ffffff64ffffffffffffff95ffffffff0000006f00000000ffffff9bffffffff",
            INIT_73 => X"000000500000000000000033000000000000006400000000ffffffdeffffffff",
            INIT_74 => X"fffffff5ffffffff0000002900000000ffffff9affffffff0000004400000000",
            INIT_75 => X"00000039000000000000006f000000000000001f00000000ffffffb7ffffffff",
            INIT_76 => X"ffffff42ffffffff000000d200000000ffffff79fffffffffffffff1ffffffff",
            INIT_77 => X"000000ce00000000000000320000000000000048000000000000006800000000",
            INIT_78 => X"0000005b00000000000000a9000000000000005000000000000000be00000000",
            INIT_79 => X"0000004100000000ffffff01ffffffff0000006200000000ffffffd7ffffffff",
            INIT_7A => X"00000069000000000000000a00000000ffffffe9ffffffffffffffd3ffffffff",
            INIT_7B => X"0000002100000000ffffffd6ffffffff00000064000000000000001300000000",
            INIT_7C => X"0000001600000000ffffff17ffffffff0000004300000000ffffffdaffffffff",
            INIT_7D => X"ffffff5affffffffffffffcdffffffffffffff38ffffffffffffff7effffffff",
            INIT_7E => X"000000fa00000000000000350000000000000018000000000000005b00000000",
            INIT_7F => X"ffffff1bffffffffffffff87ffffffff00000036000000000000006300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE13;


    MEM_IWGHT_LAYER2_INSTANCE14 : if BRAM_NAME = "iwght_layer2_instance14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffff86ffffffff0000001600000000000000ad000000000000000b00000000",
            INIT_01 => X"ffffff49ffffffff00000053000000000000009400000000ffffffc1ffffffff",
            INIT_02 => X"0000004b000000000000000700000000ffffffc1fffffffffffffffdffffffff",
            INIT_03 => X"ffffff11ffffffffffffff37ffffffffffffff72ffffffff0000006e00000000",
            INIT_04 => X"0000000700000000fffffff8ffffffff0000007e000000000000000b00000000",
            INIT_05 => X"ffffffb6ffffffffffffff9dffffffff00000033000000000000007400000000",
            INIT_06 => X"00000025000000000000001f000000000000016600000000ffffff94ffffffff",
            INIT_07 => X"0000006a00000000fffffedeffffffffffffffe8ffffffff0000006c00000000",
            INIT_08 => X"0000000900000000ffffff60ffffffffffffffd3ffffffff000000a300000000",
            INIT_09 => X"000000630000000000000030000000000000004d000000000000008d00000000",
            INIT_0A => X"0000003800000000ffffff50ffffffff0000005a00000000ffffff52ffffffff",
            INIT_0B => X"ffffffe1ffffffff00000098000000000000009200000000000000a600000000",
            INIT_0C => X"0000001600000000ffffff23fffffffffffffffffffffffffffffffaffffffff",
            INIT_0D => X"00000061000000000000000c000000000000002f000000000000003800000000",
            INIT_0E => X"0000000d00000000ffffff97ffffffffffffffc8ffffffffffffff78ffffffff",
            INIT_0F => X"ffffff55ffffffffffffff8affffffff0000005800000000000000c500000000",
            INIT_10 => X"ffffff4bffffffffffffff7effffffff0000008d000000000000008700000000",
            INIT_11 => X"00000024000000000000003700000000ffffffcfffffffff0000000300000000",
            INIT_12 => X"ffffff0cffffffff0000008e00000000ffffffe0ffffffffffffff54ffffffff",
            INIT_13 => X"0000004700000000fffffe96ffffffff0000001c00000000ffffff91ffffffff",
            INIT_14 => X"fffffff0ffffffff0000006f00000000fffffeaaffffffffffffff9fffffffff",
            INIT_15 => X"00000089000000000000001f000000000000003d00000000ffffffedffffffff",
            INIT_16 => X"00000069000000000000003b0000000000000103000000000000005c00000000",
            INIT_17 => X"ffffffc0fffffffffffffddaffffffffffffff0fffffffffffffffa8ffffffff",
            INIT_18 => X"0000001c00000000ffffffd0ffffffff000000b3000000000000009800000000",
            INIT_19 => X"0000000000000000ffffffa3ffffffff0000005b000000000000007100000000",
            INIT_1A => X"0000007d0000000000000052000000000000003a00000000ffffffc6ffffffff",
            INIT_1B => X"fffffe80ffffffffffffffd1ffffffff0000001000000000ffffff5cffffffff",
            INIT_1C => X"ffffffd5ffffffffffffff99ffffffffffffff0dffffffff0000001800000000",
            INIT_1D => X"00000042000000000000009c000000000000011e00000000000000a100000000",
            INIT_1E => X"00000014000000000000002700000000ffffffe1ffffffff0000000d00000000",
            INIT_1F => X"0000004600000000ffffffcfffffffff0000002500000000000000bc00000000",
            INIT_20 => X"ffffffddffffffffffffffa8fffffffffffffff6ffffffff0000006200000000",
            INIT_21 => X"000000460000000000000023000000000000009300000000fffffff4ffffffff",
            INIT_22 => X"ffffffe7ffffffff000000d100000000ffffffffffffffff000000a200000000",
            INIT_23 => X"ffffffebffffffffffffff5affffffffffffffffffffffff0000006700000000",
            INIT_24 => X"ffffff01ffffffff0000006200000000ffffffd5ffffffffffffff16ffffffff",
            INIT_25 => X"ffffff7affffffffffffffb2ffffffffffffffedffffffffffffffcaffffffff",
            INIT_26 => X"0000002300000000fffffff4ffffffffffffffb2ffffffff0000005f00000000",
            INIT_27 => X"fffffff4ffffffff0000004a00000000fffffff9ffffffff0000009d00000000",
            INIT_28 => X"00000070000000000000004e00000000ffffff80ffffffffffffff9cffffffff",
            INIT_29 => X"ffffff72ffffffff00000046000000000000006c00000000ffffffe9ffffffff",
            INIT_2A => X"0000000a00000000ffffff16ffffffffffffff63ffffffff0000004500000000",
            INIT_2B => X"ffffffb0ffffffffffffffd2ffffffff00000008000000000000004500000000",
            INIT_2C => X"000000a6000000000000007a0000000000000062000000000000004500000000",
            INIT_2D => X"00000004000000000000000b00000000000000e000000000000000fc00000000",
            INIT_2E => X"0000005f00000000fffffff0ffffffffffffffa2ffffffff0000001000000000",
            INIT_2F => X"fffffffbffffffff00000031000000000000005900000000ffffffefffffffff",
            INIT_30 => X"fffffff2ffffffffffffffc2ffffffff0000000e00000000ffffffbdffffffff",
            INIT_31 => X"00000053000000000000005200000000ffffff9dffffffffffffff5fffffffff",
            INIT_32 => X"ffffffe7ffffffff0000005800000000000000a500000000ffffff7affffffff",
            INIT_33 => X"0000001000000000000000a70000000000000043000000000000000c00000000",
            INIT_34 => X"ffffff7dffffffffffffff7bffffffffffffffb6ffffffff0000003d00000000",
            INIT_35 => X"000000100000000000000014000000000000001500000000fffffffaffffffff",
            INIT_36 => X"fffffff9fffffffffffffff8fffffffffffffff1ffffffff0000000d00000000",
            INIT_37 => X"00000098000000000000001b00000000fffffff8ffffffffffffffffffffffff",
            INIT_38 => X"000000ce00000000000000700000000000000043000000000000003500000000",
            INIT_39 => X"ffffffd7ffffffffffffffd0ffffffffffffff52ffffffffffffff20ffffffff",
            INIT_3A => X"00000031000000000000005e00000000ffffff43ffffffff0000004800000000",
            INIT_3B => X"ffffffcfffffffff0000000e000000000000009900000000ffffffddffffffff",
            INIT_3C => X"00000026000000000000009700000000ffffff9fffffffff0000001700000000",
            INIT_3D => X"fffffff0ffffffff0000007400000000ffffffcfffffffffffffffe4ffffffff",
            INIT_3E => X"0000006e000000000000008300000000ffffff14ffffffff0000000b00000000",
            INIT_3F => X"ffffffc7ffffffff000000df00000000ffffffa0ffffffff0000006100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffeb4ffffffffffffffd3ffffffff00000164000000000000006400000000",
            INIT_41 => X"00000000000000000000003b00000000ffffff8cffffffffffffffabffffffff",
            INIT_42 => X"0000007b000000000000005000000000ffffffe7ffffffff0000001200000000",
            INIT_43 => X"0000004e000000000000007100000000ffffff4affffffff0000005400000000",
            INIT_44 => X"00000055000000000000004a0000000000000037000000000000005b00000000",
            INIT_45 => X"0000004400000000ffffffcaffffffff0000001500000000ffffff90ffffffff",
            INIT_46 => X"ffffffb7ffffffffffffffceffffffff00000019000000000000004500000000",
            INIT_47 => X"0000002b00000000000000500000000000000010000000000000005900000000",
            INIT_48 => X"0000006000000000000000340000000000000098000000000000003b00000000",
            INIT_49 => X"ffffff31ffffffff0000001c00000000ffffff1cffffffffffffffbeffffffff",
            INIT_4A => X"00000019000000000000001d00000000ffffff92ffffffffffffffb6ffffffff",
            INIT_4B => X"ffffff7affffffff0000001d00000000ffffff13ffffffffffffffd0ffffffff",
            INIT_4C => X"0000008000000000000000a500000000ffffffa8ffffffff0000000800000000",
            INIT_4D => X"000000000000000000000026000000000000002600000000fffffff8ffffffff",
            INIT_4E => X"000000a800000000ffffff5bffffffff0000003c00000000ffffffbfffffffff",
            INIT_4F => X"0000008e00000000ffffffe7ffffffffffffffe0ffffffff0000005900000000",
            INIT_50 => X"fffffff2ffffffff0000002900000000fffffff1fffffffffffffffdffffffff",
            INIT_51 => X"0000007500000000ffffff12ffffffffffffff45ffffffffffffff7fffffffff",
            INIT_52 => X"00000014000000000000000300000000ffffffc7ffffffff0000008200000000",
            INIT_53 => X"0000001b00000000fffffffdffffffffffffffffffffffffffffffd9ffffffff",
            INIT_54 => X"ffffff39ffffffffffffff6affffffff0000005200000000ffffff85ffffffff",
            INIT_55 => X"ffffff58ffffffffffffffd2ffffffffffffffefffffffff0000004a00000000",
            INIT_56 => X"0000000d00000000fffffe6bffffffffffffff61ffffffffffffff15ffffffff",
            INIT_57 => X"0000002700000000ffffffa5ffffffffffffffabffffffff0000004900000000",
            INIT_58 => X"0000000600000000fffffffeffffffff00000062000000000000002400000000",
            INIT_59 => X"fffffff1ffffffff000000420000000000000035000000000000003c00000000",
            INIT_5A => X"ffffffe3ffffffff0000003300000000ffffffb8ffffffffffffffc4ffffffff",
            INIT_5B => X"0000006800000000ffffffffffffffffffffffe9ffffffffffffff06ffffffff",
            INIT_5C => X"000000520000000000000068000000000000008500000000ffffffe1ffffffff",
            INIT_5D => X"0000001600000000ffffffadfffffffffffffffdffffffff0000003500000000",
            INIT_5E => X"ffffff68ffffffffffffff8cffffffff0000006d000000000000000700000000",
            INIT_5F => X"ffffff57ffffffffffffffd8ffffffff0000009900000000ffffff68ffffffff",
            INIT_60 => X"0000008e00000000fffffff2ffffffffffffffe8ffffffffffffffeaffffffff",
            INIT_61 => X"0000003d000000000000000400000000ffffff5dfffffffffffffff0ffffffff",
            INIT_62 => X"ffffffd7ffffffffffffff7effffffff000000b200000000ffffffdfffffffff",
            INIT_63 => X"ffffff5cfffffffffffffffdffffffff0000005b000000000000003a00000000",
            INIT_64 => X"0000002c00000000ffffffa7ffffffff000000b1000000000000001000000000",
            INIT_65 => X"0000001100000000ffffffefffffffffffffff8fffffffff0000008800000000",
            INIT_66 => X"ffffff61ffffffff00000086000000000000000500000000ffffff8dffffffff",
            INIT_67 => X"000000b800000000ffffffdfffffffffffffffd9ffffffff0000005700000000",
            INIT_68 => X"fffffffbffffffff00000050000000000000007300000000ffffff41ffffffff",
            INIT_69 => X"fffffffdffffffffffffff8effffffff0000006d00000000ffffff25ffffffff",
            INIT_6A => X"ffffffe3fffffffffffffff6ffffffffffffffbcffffffffffffffc3ffffffff",
            INIT_6B => X"ffffff63ffffffffffffffefffffffff00000044000000000000009e00000000",
            INIT_6C => X"0000001e000000000000005300000000ffffffbeffffffff000000ac00000000",
            INIT_6D => X"0000001300000000000000650000000000000017000000000000006700000000",
            INIT_6E => X"ffffffcbffffffff00000026000000000000006b00000000ffffff8cffffffff",
            INIT_6F => X"0000000700000000ffffffedffffffff0000005c000000000000009c00000000",
            INIT_70 => X"ffffffc6ffffffff0000003f00000000ffffffa8ffffffff0000005100000000",
            INIT_71 => X"ffffff84ffffffff0000001c00000000ffffffccffffffff0000002500000000",
            INIT_72 => X"0000007400000000ffffff83ffffffffffffff41ffffffffffffffa0ffffffff",
            INIT_73 => X"ffffff51ffffffff0000006500000000ffffffbdffffffffffffff96ffffffff",
            INIT_74 => X"0000000e0000000000000057000000000000000a00000000ffffffe5ffffffff",
            INIT_75 => X"ffffff9fffffffff0000000f000000000000009d00000000fffffffeffffffff",
            INIT_76 => X"0000005300000000ffffffdfffffffffffffffdeffffffffffffffb0ffffffff",
            INIT_77 => X"0000000d000000000000003c000000000000000c000000000000006100000000",
            INIT_78 => X"0000007500000000ffffff42ffffffff0000003100000000ffffffe1ffffffff",
            INIT_79 => X"ffffff37ffffffffffffffc0ffffffffffffff27ffffffffffffffeeffffffff",
            INIT_7A => X"000000580000000000000004000000000000002000000000ffffffbaffffffff",
            INIT_7B => X"ffffffc0ffffffff00000087000000000000005500000000ffffffe7ffffffff",
            INIT_7C => X"0000009f00000000000000160000000000000048000000000000000100000000",
            INIT_7D => X"0000000800000000fffffffcfffffffffffffffdffffffff0000004700000000",
            INIT_7E => X"00000000000000000000000700000000fffffff2ffffffffffffffffffffffff",
            INIT_7F => X"0000000900000000ffffffb6ffffffff00000002000000000000000100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE14;


    MEM_IWGHT_LAYER2_INSTANCE15 : if BRAM_NAME = "iwght_layer2_instance15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffff91ffffffffffffffcdffffffffffffffa9ffffffffffffff7dffffffff",
            INIT_01 => X"ffffffdbffffffff000000340000000000000062000000000000004a00000000",
            INIT_02 => X"0000000f00000000ffffffeeffffffff0000009c00000000ffffffb9ffffffff",
            INIT_03 => X"ffffff0effffffff00000053000000000000007d00000000fffffff1ffffffff",
            INIT_04 => X"ffffff9cffffffffffffffe3ffffffffffffffa3ffffffff0000005b00000000",
            INIT_05 => X"ffffff1effffffff0000000e00000000ffffff70ffffffff000000a100000000",
            INIT_06 => X"ffffff94ffffffff00000037000000000000007900000000ffffffd5ffffffff",
            INIT_07 => X"ffffff3bffffffffffffffcbffffffff000000b6000000000000003900000000",
            INIT_08 => X"0000004300000000ffffffb4ffffffff0000006d000000000000000500000000",
            INIT_09 => X"00000023000000000000003e000000000000001f00000000ffffffefffffffff",
            INIT_0A => X"fffffffdffffffff0000000d00000000fffffffbffffffffffffff65ffffffff",
            INIT_0B => X"0000008c00000000ffffffd9ffffffff0000006700000000ffffff7effffffff",
            INIT_0C => X"0000005a00000000000000180000000000000045000000000000002600000000",
            INIT_0D => X"fffffeb2ffffffff0000007200000000000000ba00000000ffffffe2ffffffff",
            INIT_0E => X"0000003d000000000000008f00000000000000d700000000ffffff85ffffffff",
            INIT_0F => X"ffffff72ffffffffffffff82ffffffff000000f600000000ffffffc2ffffffff",
            INIT_10 => X"0000000400000000ffffff33ffffffffffffffdaffffffff0000001500000000",
            INIT_11 => X"0000000800000000ffffff59ffffffffffffff41ffffffffffffff4fffffffff",
            INIT_12 => X"ffffffdefffffffffffffff4ffffffff0000004400000000000000d500000000",
            INIT_13 => X"000000ac000000000000001900000000ffffffebffffffffffffffd3ffffffff",
            INIT_14 => X"00000022000000000000008a00000000ffffffd4ffffffff0000006400000000",
            INIT_15 => X"0000003700000000ffffffd5ffffffff0000008900000000ffffffa4ffffffff",
            INIT_16 => X"000000ad00000000ffffffb5ffffffff0000008e00000000ffffffc5ffffffff",
            INIT_17 => X"ffffff6bffffffff0000003b00000000fffffebeffffffff0000003800000000",
            INIT_18 => X"0000006300000000fffffff0ffffffff000000a100000000fffffff8ffffffff",
            INIT_19 => X"fffffef6ffffffffffffffc6ffffffff0000004800000000ffffff47ffffffff",
            INIT_1A => X"ffffffcfffffffffffffffa7ffffffffffffffb2ffffffff0000003f00000000",
            INIT_1B => X"000000d8000000000000001e00000000ffffff24ffffffff0000005c00000000",
            INIT_1C => X"fffffff9ffffffff000000f000000000ffffff17ffffffffffffff48ffffffff",
            INIT_1D => X"ffffffefffffffffffffffe9ffffffffffffffdaffffffff0000006600000000",
            INIT_1E => X"0000007600000000ffffff6efffffffffffffef2ffffffffffffffafffffffff",
            INIT_1F => X"0000004f0000000000000041000000000000000c00000000ffffffebffffffff",
            INIT_20 => X"fffffffdffffffff0000008b00000000fffffe2affffffff0000007600000000",
            INIT_21 => X"ffffffeeffffffff0000004d00000000000000d3000000000000007d00000000",
            INIT_22 => X"0000003e00000000ffffffbffffffffffffffff9ffffffffffffffeaffffffff",
            INIT_23 => X"ffffff00ffffffff000000af00000000ffffffb9ffffffffffffffadffffffff",
            INIT_24 => X"ffffffadffffffffffffff99ffffffff00000008000000000000003000000000",
            INIT_25 => X"00000071000000000000008900000000000000a400000000ffffffdcffffffff",
            INIT_26 => X"000000cd000000000000009d00000000ffffff4dffffffff0000003600000000",
            INIT_27 => X"ffffff50ffffffff00000005000000000000004600000000ffffff17ffffffff",
            INIT_28 => X"00000099000000000000001100000000ffffff82ffffffffffffff68ffffffff",
            INIT_29 => X"0000006c000000000000002b000000000000000500000000ffffff9dffffffff",
            INIT_2A => X"ffffff2cfffffffffffffffaffffffffffffff76ffffffff0000008600000000",
            INIT_2B => X"0000006b00000000ffffff8dffffffff0000004b00000000ffffffabffffffff",
            INIT_2C => X"000000a400000000000000220000000000000057000000000000009300000000",
            INIT_2D => X"000000190000000000000103000000000000008f00000000ffffff0bffffffff",
            INIT_2E => X"0000000d000000000000004600000000fffffff1fffffffffffffe4affffffff",
            INIT_2F => X"0000000600000000ffffffb9ffffffffffffff32ffffffffffffffa8ffffffff",
            INIT_30 => X"ffffffd6ffffffffffffffc5ffffffffffffff93ffffffffffffff24ffffffff",
            INIT_31 => X"ffffff0affffffffffffffd1ffffffff00000002000000000000000400000000",
            INIT_32 => X"00000068000000000000001f00000000ffffff96ffffffff0000003700000000",
            INIT_33 => X"0000001b00000000ffffff63ffffffffffffffc1ffffffff0000007200000000",
            INIT_34 => X"0000001b00000000ffffff99ffffffffffffffc2ffffffff0000008700000000",
            INIT_35 => X"ffffffcfffffffff0000003400000000000000b7000000000000008d00000000",
            INIT_36 => X"0000001e00000000000000a500000000ffffffd3ffffffff0000006100000000",
            INIT_37 => X"00000000000000000000005300000000000000aa000000000000000500000000",
            INIT_38 => X"ffffff25ffffffffffffff99ffffffffffffffc3ffffffffffffff58ffffffff",
            INIT_39 => X"000000bb00000000ffffff6cffffffffffffff33ffffffffffffff80ffffffff",
            INIT_3A => X"0000007200000000ffffff75ffffffff00000050000000000000004f00000000",
            INIT_3B => X"0000000900000000000000d0000000000000000e000000000000002b00000000",
            INIT_3C => X"0000006c000000000000003100000000ffffffe2ffffffff0000008100000000",
            INIT_3D => X"0000000b00000000ffffff96ffffffff00000037000000000000007a00000000",
            INIT_3E => X"0000002600000000ffffffccffffffffffffffc4ffffffff0000002c00000000",
            INIT_3F => X"ffffffb1fffffffffffffffcffffffff0000004900000000ffffffd4ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffff92ffffffffffffff3affffffffffffffb4ffffffff0000001600000000",
            INIT_41 => X"0000001100000000fffffffdffffffff00000025000000000000006100000000",
            INIT_42 => X"ffffffd2ffffffffffffff6affffffff0000003c000000000000006300000000",
            INIT_43 => X"0000008c00000000fffffff3ffffffff0000008b00000000ffffffb7ffffffff",
            INIT_44 => X"000000000000000000000001000000000000004300000000ffffff6fffffffff",
            INIT_45 => X"0000000f0000000000000005000000000000000c00000000ffffff47ffffffff",
            INIT_46 => X"fffffff5ffffffffffffffebfffffffffffffff5ffffffff0000000300000000",
            INIT_47 => X"00000038000000000000000400000000ffffffedfffffffffffffff0ffffffff",
            INIT_48 => X"ffffffe7ffffffff000000bb00000000fffffff9ffffffff0000005200000000",
            INIT_49 => X"ffffffc4ffffffff000000f600000000000000cc00000000fffffff3ffffffff",
            INIT_4A => X"0000005100000000ffffff92ffffffff00000084000000000000006d00000000",
            INIT_4B => X"ffffffa6ffffffffffffff1effffffffffffff81ffffffff0000006200000000",
            INIT_4C => X"ffffffe7ffffffffffffffbaffffffff00000149000000000000002800000000",
            INIT_4D => X"fffffee5ffffffffffffff18ffffffff0000009600000000000000b000000000",
            INIT_4E => X"000000c1000000000000004f00000000ffffffdeffffffffffffffc1ffffffff",
            INIT_4F => X"0000000300000000ffffffa2ffffffffffffff49ffffffff0000009600000000",
            INIT_50 => X"ffffffcfffffffffffffff73ffffffffffffffaeffffffffffffff79ffffffff",
            INIT_51 => X"0000006d00000000ffffffe3ffffffffffffff87ffffffffffffff66ffffffff",
            INIT_52 => X"ffffffdbffffffffffffff3dffffffffffffff84ffffffffffffffb9ffffffff",
            INIT_53 => X"0000006e00000000ffffffb5ffffffff0000001600000000000000bd00000000",
            INIT_54 => X"0000008c00000000ffffff8dffffffffffffff8bffffffff0000009200000000",
            INIT_55 => X"ffffff9bffffffff00000033000000000000003e000000000000008200000000",
            INIT_56 => X"ffffffdefffffffffffffe9fffffffff0000008d000000000000002600000000",
            INIT_57 => X"0000008a000000000000008100000000fffffffcffffffffffffff99ffffffff",
            INIT_58 => X"ffffff33ffffffff00000025000000000000005900000000ffffff81ffffffff",
            INIT_59 => X"000000c4000000000000001a00000000ffffffa0ffffffffffffff44ffffffff",
            INIT_5A => X"fffffffcffffffff000000ce000000000000003600000000ffffffd2ffffffff",
            INIT_5B => X"0000006600000000fffffff6ffffffff0000009000000000ffffff12ffffffff",
            INIT_5C => X"ffffff40ffffffff0000007c000000000000004600000000ffffff9dffffffff",
            INIT_5D => X"000000510000000000000037000000000000000a00000000ffffff31ffffffff",
            INIT_5E => X"ffffff65ffffffffffffffa7ffffffffffffffceffffffffffffffdcffffffff",
            INIT_5F => X"0000002f000000000000007e000000000000007500000000fffffef0ffffffff",
            INIT_60 => X"0000009d00000000ffffff3fffffffff0000006100000000fffffe8bffffffff",
            INIT_61 => X"000000a6000000000000002d00000000ffffff32ffffffffffffff89ffffffff",
            INIT_62 => X"ffffffadffffffffffffff93ffffffffffffff73ffffffffffffffd2ffffffff",
            INIT_63 => X"fffffffaffffffff0000005b000000000000004e00000000fffffff7ffffffff",
            INIT_64 => X"ffffffcbffffffff00000019000000000000000000000000ffffff29ffffffff",
            INIT_65 => X"0000004600000000ffffffd5fffffffffffffffdffffffffffffff81ffffffff",
            INIT_66 => X"00000085000000000000003000000000ffffff73ffffffff0000002000000000",
            INIT_67 => X"fffffff4ffffffff0000000200000000fffffffcffffffffffffff6bffffffff",
            INIT_68 => X"0000002b00000000ffffff4bffffffffffffffe5ffffffff0000005d00000000",
            INIT_69 => X"0000002b000000000000004f000000000000008900000000000000f600000000",
            INIT_6A => X"0000001700000000ffffff6effffffff00000035000000000000001600000000",
            INIT_6B => X"ffffffecffffffffffffffafffffffff0000001c000000000000005500000000",
            INIT_6C => X"0000001500000000ffffff6affffffffffffffc5ffffffffffffff7effffffff",
            INIT_6D => X"0000008f00000000fffffeb7ffffffffffffff5efffffffffffffe93ffffffff",
            INIT_6E => X"ffffffa6ffffffffffffffc1fffffffffffffff9ffffffff0000005300000000",
            INIT_6F => X"0000004100000000ffffff98ffffffff0000005500000000ffffffdcffffffff",
            INIT_70 => X"ffffff79ffffffff0000007700000000ffffffd4ffffffff0000004100000000",
            INIT_71 => X"ffffffecfffffffffffffff9ffffffff00000066000000000000004000000000",
            INIT_72 => X"fffffff5ffffffff0000010900000000fffffffdffffffff0000001700000000",
            INIT_73 => X"fffffff5ffffffffffffff85ffffffffffffffacffffffff0000002200000000",
            INIT_74 => X"0000003100000000fffffff8ffffffff0000000600000000ffffffd5ffffffff",
            INIT_75 => X"000000b0000000000000002d00000000fffffffbffffffff0000001200000000",
            INIT_76 => X"0000000200000000ffffffb7ffffffffffffffe8fffffffffffffff8ffffffff",
            INIT_77 => X"ffffff7effffffff0000001800000000ffffffbdffffffffffffff1dffffffff",
            INIT_78 => X"ffffffe0ffffffffffffffb4ffffffff0000003700000000ffffff7bffffffff",
            INIT_79 => X"0000005700000000ffffff8dffffffffffffffbdffffffff0000006d00000000",
            INIT_7A => X"00000030000000000000004300000000fffffff7ffffffff0000004e00000000",
            INIT_7B => X"ffffffbeffffffff0000004a000000000000006100000000ffffff9affffffff",
            INIT_7C => X"0000005500000000fffffff3ffffffff0000005e00000000ffffff09ffffffff",
            INIT_7D => X"ffffff15ffffffff0000004f0000000000000066000000000000004a00000000",
            INIT_7E => X"ffffffebffffffff0000001400000000ffffff0dffffffffffffff73ffffffff",
            INIT_7F => X"0000005900000000ffffffe2ffffffffffffffe8ffffffff0000002000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE15;


    MEM_IWGHT_LAYER2_INSTANCE16 : if BRAM_NAME = "iwght_layer2_instance16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffafffffffffffffff7bffffffff00000019000000000000002800000000",
            INIT_01 => X"ffffff72ffffffffffffff26ffffffffffffff8cffffffffffffff86ffffffff",
            INIT_02 => X"000000140000000000000020000000000000005b00000000ffffff8cffffffff",
            INIT_03 => X"0000006d00000000ffffffb8ffffffff0000002300000000ffffff0cffffffff",
            INIT_04 => X"0000001a00000000ffffffa9ffffffff0000007900000000ffffffb4ffffffff",
            INIT_05 => X"00000009000000000000003a00000000ffffffefffffffffffffffa1ffffffff",
            INIT_06 => X"0000007b00000000ffffffbbffffffff0000003a00000000ffffffbaffffffff",
            INIT_07 => X"000000ce00000000ffffffaaffffffffffffffc1ffffffff000000d900000000",
            INIT_08 => X"ffffffebffffffff00000058000000000000002f000000000000004d00000000",
            INIT_09 => X"00000052000000000000005600000000ffffff43fffffffffffffff3ffffffff",
            INIT_0A => X"0000001a000000000000000300000000000000d500000000ffffff7fffffffff",
            INIT_0B => X"0000003a000000000000003a00000000ffffffe9ffffffffffffffe9ffffffff",
            INIT_0C => X"000000900000000000000034000000000000004600000000ffffffc9ffffffff",
            INIT_0D => X"fffffff8ffffffff0000000a0000000000000001000000000000003800000000",
            INIT_0E => X"000000150000000000000010000000000000001500000000fffffff8ffffffff",
            INIT_0F => X"ffffff67ffffffff0000002d000000000000000900000000fffffff9ffffffff",
            INIT_10 => X"0000000f000000000000002200000000ffffffdaffffffffffffff9affffffff",
            INIT_11 => X"ffffffe9ffffffff0000006f00000000fffffffdffffffff0000001200000000",
            INIT_12 => X"0000000e00000000ffffffcaffffffff00000040000000000000001700000000",
            INIT_13 => X"0000002d000000000000004100000000ffffff8dffffffff0000004100000000",
            INIT_14 => X"ffffffb2fffffffffffffe10ffffffffffffff92ffffffff0000000500000000",
            INIT_15 => X"ffffffa1ffffffffffffffdfffffffffffffff56ffffffffffffff7cffffffff",
            INIT_16 => X"ffffff1fffffffffffffffdeffffffffffffffd8fffffffffffffef5ffffffff",
            INIT_17 => X"ffffffccffffffffffffff47fffffffffffffee3ffffffffffffffffffffffff",
            INIT_18 => X"ffffffc5ffffffffffffff98ffffffffffffff19ffffffffffffffdeffffffff",
            INIT_19 => X"0000001900000000ffffffacffffffff000000c100000000ffffffbfffffffff",
            INIT_1A => X"00000105000000000000000200000000ffffffc4ffffffff0000003700000000",
            INIT_1B => X"ffffff11ffffffffffffff44ffffffffffffff8dffffffffffffffbcffffffff",
            INIT_1C => X"0000000600000000ffffffa1ffffffff000000c2000000000000003600000000",
            INIT_1D => X"ffffffe2ffffffff0000003800000000ffffffe6ffffffffffffffbfffffffff",
            INIT_1E => X"000000130000000000000059000000000000007000000000ffffff37ffffffff",
            INIT_1F => X"ffffffecffffffff0000001a00000000fffffec0ffffffff0000002b00000000",
            INIT_20 => X"ffffffd2fffffffffffffedeffffffff0000000c000000000000004600000000",
            INIT_21 => X"ffffff59ffffffff0000003900000000ffffff3cffffffffffffffd4ffffffff",
            INIT_22 => X"ffffffc3fffffffffffffff1ffffffff000000e5000000000000006100000000",
            INIT_23 => X"0000004200000000ffffffcaffffffff0000001100000000ffffffa5ffffffff",
            INIT_24 => X"0000003300000000ffffffecffffffff0000001200000000ffffffd9ffffffff",
            INIT_25 => X"0000000e00000000ffffff6fffffffffffffffefffffffffffffff66ffffffff",
            INIT_26 => X"ffffff62ffffffff000000660000000000000013000000000000006900000000",
            INIT_27 => X"ffffffc8ffffffffffffff48fffffffffffffff3ffffffffffffff83ffffffff",
            INIT_28 => X"ffffffb4fffffffffffffefafffffffffffffee5ffffffffffffff62ffffffff",
            INIT_29 => X"ffffffffffffffffffffffa6ffffffffffffff21fffffffffffffefbffffffff",
            INIT_2A => X"fffffebaffffffff0000002a00000000fffffeebffffffffffffff53ffffffff",
            INIT_2B => X"ffffffd6ffffffffffffff68ffffffffffffff62ffffffffffffffe3ffffffff",
            INIT_2C => X"0000004600000000fffffed9ffffffff0000000700000000ffffffccffffffff",
            INIT_2D => X"0000004b000000000000000400000000000000f100000000ffffffcfffffffff",
            INIT_2E => X"0000004400000000ffffff91ffffffffffffffcaffffffff0000009600000000",
            INIT_2F => X"0000006a00000000ffffff98ffffffffffffffecffffffff0000007900000000",
            INIT_30 => X"ffffffb8ffffffff0000004300000000ffffffd8ffffffffffffffacffffffff",
            INIT_31 => X"0000000c00000000000000330000000000000046000000000000004700000000",
            INIT_32 => X"ffffffadfffffffffffffff0ffffffffffffffdfffffffffffffff94ffffffff",
            INIT_33 => X"000000e200000000ffffff78ffffffffffffff94ffffffffffffffd3ffffffff",
            INIT_34 => X"ffffff77ffffffffffffffd5ffffffff000000ae000000000000001c00000000",
            INIT_35 => X"ffffffb0ffffffff0000002700000000ffffffe5ffffffffffffffedffffffff",
            INIT_36 => X"000000050000000000000003000000000000001c000000000000006100000000",
            INIT_37 => X"ffffffecffffffff000000120000000000000020000000000000008b00000000",
            INIT_38 => X"0000003f000000000000000600000000ffffffeeffffffff0000000f00000000",
            INIT_39 => X"0000007c00000000ffffff33ffffffff0000008700000000ffffffa6ffffffff",
            INIT_3A => X"ffffffb4ffffffff0000005100000000ffffffe2ffffffff000000d100000000",
            INIT_3B => X"0000005b00000000ffffff66ffffffff000000e100000000fffffec7ffffffff",
            INIT_3C => X"ffffff8bffffffff0000004c00000000ffffff61ffffffff000000b000000000",
            INIT_3D => X"0000000700000000fffffffeffffffff0000002300000000ffffff65ffffffff",
            INIT_3E => X"000000ab00000000ffffffbaffffffff000000a300000000ffffff9cffffffff",
            INIT_3F => X"00000066000000000000000000000000ffffff6cffffffff0000001d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffeeffffffff000000bd00000000fffffff2ffffffffffffffe9ffffffff",
            INIT_41 => X"ffffffe3ffffffff0000000a00000000fffffffdffffffff0000001900000000",
            INIT_42 => X"0000001e000000000000002f0000000000000001000000000000003700000000",
            INIT_43 => X"0000006c00000000ffffffeeffffffffffffffc4ffffffff0000008300000000",
            INIT_44 => X"ffffff2bffffffff0000006100000000ffffff2effffffffffffff2cffffffff",
            INIT_45 => X"0000003200000000ffffff40ffffffffffffffbcffffffffffffff95ffffffff",
            INIT_46 => X"ffffff94ffffffffffffff0dffffffffffffff7dffffffff0000006c00000000",
            INIT_47 => X"0000000600000000ffffffb3ffffffffffffffceffffffffffffffbbffffffff",
            INIT_48 => X"ffffff70ffffffffffffff28ffffffff0000002c00000000ffffff0dffffffff",
            INIT_49 => X"ffffff6cffffffffffffffa0fffffffffffffeb1fffffffffffffeceffffffff",
            INIT_4A => X"0000004a000000000000007000000000fffffeffffffffff0000007000000000",
            INIT_4B => X"ffffffe9ffffffff0000000a00000000ffffff00ffffffffffffffc8ffffffff",
            INIT_4C => X"fffffff5ffffffff000000f800000000000000e300000000ffffffd9ffffffff",
            INIT_4D => X"ffffffc6ffffffff0000002900000000000000f0000000000000000d00000000",
            INIT_4E => X"0000009400000000ffffffb6fffffffffffffff5ffffffffffffffdeffffffff",
            INIT_4F => X"000000db000000000000002900000000ffffff91ffffffff0000006600000000",
            INIT_50 => X"ffffff1effffffff00000004000000000000004200000000ffffff7fffffffff",
            INIT_51 => X"0000002b0000000000000011000000000000009600000000ffffffd7ffffffff",
            INIT_52 => X"ffffffd5ffffffffffffffe6ffffffff0000000f000000000000003600000000",
            INIT_53 => X"0000003f00000000ffffff60ffffffff0000000000000000ffffffd0ffffffff",
            INIT_54 => X"0000000f00000000ffffffefffffffffffffffe6ffffffffffffffe4ffffffff",
            INIT_55 => X"0000000400000000fffffffbffffffff0000000c00000000ffffff31ffffffff",
            INIT_56 => X"fffffff7fffffffffffffff0ffffffff00000004000000000000000800000000",
            INIT_57 => X"ffffffbdffffffffffffffdfffffffff00000006000000000000000600000000",
            INIT_58 => X"0000004700000000000000b50000000000000041000000000000005c00000000",
            INIT_59 => X"0000005900000000000000ad00000000ffffffc7ffffffffffffffaeffffffff",
            INIT_5A => X"00000032000000000000002100000000ffffff91ffffffffffffffacffffffff",
            INIT_5B => X"ffffff83ffffffff00000052000000000000001a000000000000003900000000",
            INIT_5C => X"ffffff79ffffffff000000000000000000000013000000000000000100000000",
            INIT_5D => X"ffffffacffffffffffffffcfffffffff0000001800000000ffffffaeffffffff",
            INIT_5E => X"ffffff0dffffffffffffffc7ffffffff0000000000000000ffffffccffffffff",
            INIT_5F => X"0000014300000000ffffff5cfffffffffffffe9effffffffffffffd7ffffffff",
            INIT_60 => X"ffffff98ffffffff00000025000000000000000a00000000000000c200000000",
            INIT_61 => X"ffffff68ffffffffffffffe5ffffffff00000035000000000000007400000000",
            INIT_62 => X"000000c6000000000000004d000000000000007f00000000ffffff4fffffffff",
            INIT_63 => X"0000004400000000fffffff6ffffffffffffff47ffffffff0000002300000000",
            INIT_64 => X"ffffffccffffffff00000058000000000000003600000000ffffff95ffffffff",
            INIT_65 => X"000000b800000000fffffff9ffffffff00000033000000000000002200000000",
            INIT_66 => X"0000003700000000ffffffe4ffffffffffffff91ffffffff0000003200000000",
            INIT_67 => X"ffffff9dffffffffffffff8fffffffff00000065000000000000000000000000",
            INIT_68 => X"fffffff7ffffffffffffffb9ffffffff00000070000000000000000000000000",
            INIT_69 => X"ffffffa7ffffffff0000002800000000ffffffa6ffffffffffffff96ffffffff",
            INIT_6A => X"ffffff63ffffffff00000050000000000000006b00000000ffffffecffffffff",
            INIT_6B => X"ffffff5fffffffff0000000500000000fffffed6ffffffffffffff45ffffffff",
            INIT_6C => X"0000000d0000000000000063000000000000007b00000000ffffffcdffffffff",
            INIT_6D => X"0000005a000000000000004100000000ffffffecffffffffffffffe7ffffffff",
            INIT_6E => X"0000003900000000ffffff9cffffffff0000006300000000ffffffbaffffffff",
            INIT_6F => X"0000001f000000000000000b00000000ffffff65ffffffffffffffc8ffffffff",
            INIT_70 => X"ffffffdeffffffff0000000800000000fffffffcffffffff0000004a00000000",
            INIT_71 => X"0000000000000000ffffff47ffffffffffffffa8ffffffffffffffb7ffffffff",
            INIT_72 => X"0000000000000000ffffffcdfffffffffffffffaffffffff0000000e00000000",
            INIT_73 => X"ffffff98ffffffffffffffebffffffff000000db000000000000007c00000000",
            INIT_74 => X"ffffffd2ffffffff000000f600000000000000b800000000ffffff94ffffffff",
            INIT_75 => X"ffffff7affffffffffffff5effffffff0000007400000000ffffffd6ffffffff",
            INIT_76 => X"00000010000000000000005e000000000000000b000000000000003000000000",
            INIT_77 => X"ffffff31ffffffff00000021000000000000006a000000000000006400000000",
            INIT_78 => X"00000018000000000000001e00000000fffffffaffffffff0000004500000000",
            INIT_79 => X"0000001200000000ffffff65ffffffffffffffe1ffffffff000000ae00000000",
            INIT_7A => X"0000008900000000ffffffd7ffffffff00000062000000000000002400000000",
            INIT_7B => X"ffffff8bffffffffffffff74ffffffff0000003d00000000ffffffd9ffffffff",
            INIT_7C => X"0000008e000000000000011400000000ffffff1effffffffffffffc9ffffffff",
            INIT_7D => X"ffffffc0ffffffffffffff86fffffffffffffff9ffffffffffffff62ffffffff",
            INIT_7E => X"0000000400000000ffffffc8ffffffff0000000800000000ffffff8bffffffff",
            INIT_7F => X"000000c100000000ffffff4fffffffffffffff6fffffffff0000006a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE16;


    MEM_IWGHT_LAYER2_INSTANCE17 : if BRAM_NAME = "iwght_layer2_instance17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffffffffffff000000ad000000000000008c00000000ffffffb5ffffffff",
            INIT_01 => X"ffffff6bfffffffffffffe31ffffffff00000052000000000000006d00000000",
            INIT_02 => X"0000002f00000000ffffffeeffffffffffffff97ffffffffffffffcfffffffff",
            INIT_03 => X"ffffff6fffffffff0000003f00000000ffffffacffffffff0000005900000000",
            INIT_04 => X"0000003000000000ffffff6dffffffffffffff9fffffffff0000000000000000",
            INIT_05 => X"ffffff90ffffffff0000009f000000000000003c000000000000005100000000",
            INIT_06 => X"0000005800000000ffffff00ffffffff0000004f00000000fffffff5ffffffff",
            INIT_07 => X"ffffffd0ffffffff0000006300000000ffffffceffffffffffffff81ffffffff",
            INIT_08 => X"0000007f00000000ffffff2affffffffffffffecffffffffffffff93ffffffff",
            INIT_09 => X"fffffff4ffffffff000000620000000000000022000000000000000e00000000",
            INIT_0A => X"0000002b00000000ffffff6afffffffffffffec1fffffffffffffffaffffffff",
            INIT_0B => X"ffffffbfffffffffffffffb1ffffffffffffff88ffffffff000000a000000000",
            INIT_0C => X"0000002600000000ffffffe9ffffffffffffffc6ffffffffffffff56ffffffff",
            INIT_0D => X"ffffffa5ffffffffffffffcbffffffffffffff5affffffffffffff9dffffffff",
            INIT_0E => X"0000007200000000ffffffaaffffffff00000049000000000000000e00000000",
            INIT_0F => X"ffffffefffffffff000000c300000000ffffffa1ffffffff0000001800000000",
            INIT_10 => X"fffffec0fffffffffffffff2ffffffff00000002000000000000001b00000000",
            INIT_11 => X"0000006c00000000ffffffebffffffffffffff7dfffffffffffffff2ffffffff",
            INIT_12 => X"0000000100000000000000fd00000000fffffff0fffffffffffffff8ffffffff",
            INIT_13 => X"0000006e00000000fffffe75ffffffffffffffa4fffffffffffffec7ffffffff",
            INIT_14 => X"ffffff48ffffffff0000005000000000000000a1000000000000008700000000",
            INIT_15 => X"fffffeaaffffffff00000017000000000000007e00000000ffffffcaffffffff",
            INIT_16 => X"000000cf00000000ffffff01ffffffff0000003d00000000ffffff84ffffffff",
            INIT_17 => X"fffffff3ffffffffffffff2cfffffffffffffe7bffffffff0000004500000000",
            INIT_18 => X"ffffffadffffffff0000001f00000000fffffebfffffffffffffff58ffffffff",
            INIT_19 => X"00000042000000000000001800000000ffffffdaffffffffffffff16ffffffff",
            INIT_1A => X"00000065000000000000001200000000ffffffc9ffffffff000000d800000000",
            INIT_1B => X"ffffff8efffffffffffffec6ffffffffffffff85ffffffff0000006100000000",
            INIT_1C => X"0000000e00000000ffffffeaffffffff00000002000000000000001f00000000",
            INIT_1D => X"0000000d000000000000000b000000000000000c00000000ffffffd5ffffffff",
            INIT_1E => X"fffffff9ffffffff00000006000000000000000a000000000000000700000000",
            INIT_1F => X"0000005300000000fffffffffffffffffffffffdfffffffffffffff7ffffffff",
            INIT_20 => X"0000005500000000000000a000000000ffffffe8ffffffff0000006f00000000",
            INIT_21 => X"ffffff60ffffffff0000002200000000fffffffaffffffffffffff26ffffffff",
            INIT_22 => X"ffffff40ffffffffffffffc4ffffffffffffffa9fffffffffffffeaaffffffff",
            INIT_23 => X"0000008c0000000000000054000000000000004300000000ffffff7fffffffff",
            INIT_24 => X"0000009500000000ffffff9affffffff0000001700000000ffffff1affffffff",
            INIT_25 => X"ffffff97ffffffff000000620000000000000007000000000000003d00000000",
            INIT_26 => X"ffffff2fffffffff0000007400000000fffffeceffffffffffffff17ffffffff",
            INIT_27 => X"00000087000000000000002a00000000fffffe26fffffffffffffd9bffffffff",
            INIT_28 => X"ffffff70ffffffffffffffadffffffff00000068000000000000013200000000",
            INIT_29 => X"0000006a00000000fffffffcffffffff00000041000000000000006300000000",
            INIT_2A => X"00000041000000000000004d00000000ffffff36fffffffffffffeb9ffffffff",
            INIT_2B => X"0000008600000000fffffff1ffffffffffffff8cffffffff0000000900000000",
            INIT_2C => X"000000820000000000000019000000000000007f000000000000006a00000000",
            INIT_2D => X"0000018d00000000000000bc00000000ffffff99ffffffff0000001400000000",
            INIT_2E => X"0000003400000000ffffffb9fffffffffffffff1ffffffffffffff4effffffff",
            INIT_2F => X"000000440000000000000033000000000000003800000000ffffff73ffffffff",
            INIT_30 => X"0000002800000000ffffffa9fffffffffffffff8ffffffff0000002500000000",
            INIT_31 => X"ffffff19ffffffff0000009e000000000000003700000000ffffffc8ffffffff",
            INIT_32 => X"ffffffc9ffffffff0000001100000000fffffefdffffffff0000007b00000000",
            INIT_33 => X"ffffffcbfffffffffffffe22ffffffff000000b000000000ffffffc4ffffffff",
            INIT_34 => X"0000007a00000000ffffffeeffffffffffffffb7ffffffff000000ae00000000",
            INIT_35 => X"ffffff89ffffffffffffffd6ffffffff0000009e00000000fffffff7ffffffff",
            INIT_36 => X"000000e800000000ffffffa2ffffffffffffffafffffffffffffff7fffffffff",
            INIT_37 => X"0000006d00000000000000ef00000000fffffedeffffffffffffffdbffffffff",
            INIT_38 => X"ffffffc0ffffffffffffff4cffffffff0000003000000000ffffffeeffffffff",
            INIT_39 => X"ffffffb0ffffffffffffff2cffffffffffffffb8ffffffffffffffdfffffffff",
            INIT_3A => X"fffffec0ffffffff0000005d000000000000008200000000000000d300000000",
            INIT_3B => X"0000011a00000000ffffff89ffffffffffffff95ffffffffffffffceffffffff",
            INIT_3C => X"00000036000000000000004e00000000ffffffbaffffffff0000004400000000",
            INIT_3D => X"00000079000000000000004b00000000ffffff9cffffffff0000006800000000",
            INIT_3E => X"00000088000000000000007e000000000000010100000000ffffffb1ffffffff",
            INIT_3F => X"ffffff9dffffffff00000037000000000000001c000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004f00000000ffffffc1ffffffffffffffe8ffffffffffffff9dffffffff",
            INIT_41 => X"ffffffc2ffffffffffffffe2ffffffffffffffd8fffffffffffffefcffffffff",
            INIT_42 => X"0000008a00000000000000980000000000000069000000000000005400000000",
            INIT_43 => X"ffffffbbffffffff000000790000000000000001000000000000008200000000",
            INIT_44 => X"ffffffdaffffffffffffffb2ffffffffffffff4cffffffff0000001200000000",
            INIT_45 => X"ffffff4dffffffffffffff51ffffffff0000000d00000000ffffff9cffffffff",
            INIT_46 => X"0000008e00000000ffffff9ffffffffffffffff2ffffffff0000007f00000000",
            INIT_47 => X"000000fb0000000000000065000000000000001c00000000ffffff35ffffffff",
            INIT_48 => X"000000a800000000000000330000000000000061000000000000005100000000",
            INIT_49 => X"ffffffaeffffffff0000002b00000000ffffffa4ffffffffffffffecffffffff",
            INIT_4A => X"0000009f00000000ffffff96ffffffffffffffc5ffffffffffffffe2ffffffff",
            INIT_4B => X"000000c8000000000000008000000000ffffff0effffffff0000004600000000",
            INIT_4C => X"000000690000000000000050000000000000002600000000fffffeefffffffff",
            INIT_4D => X"ffffff83ffffffffffffffb6ffffffff0000005b000000000000006900000000",
            INIT_4E => X"ffffffdffffffffffffffff7ffffffffffffffe1ffffffffffffffe5ffffffff",
            INIT_4F => X"0000002500000000000000eb00000000ffffff47ffffffff000000c800000000",
            INIT_50 => X"ffffff5afffffffffffffe44ffffffffffffff92ffffffffffffff79ffffffff",
            INIT_51 => X"ffffffa8ffffffff00000030000000000000006800000000ffffffebffffffff",
            INIT_52 => X"ffffffb1ffffffffffffff90ffffffff00000048000000000000001200000000",
            INIT_53 => X"ffffffe8ffffffff0000000900000000ffffff72ffffffff0000000900000000",
            INIT_54 => X"000000200000000000000030000000000000005500000000fffffff1ffffffff",
            INIT_55 => X"ffffffe3ffffffffffffff36ffffffff0000003500000000ffffff6dffffffff",
            INIT_56 => X"0000001a00000000ffffff3effffffff0000001900000000ffffffedffffffff",
            INIT_57 => X"fffffed9ffffffff0000008f00000000ffffff8cffffffff0000009500000000",
            INIT_58 => X"ffffff1ffffffffffffffedbfffffffffffffff7ffffffffffffffa1ffffffff",
            INIT_59 => X"0000008b00000000fffffffbffffffffffffff52fffffffffffffff8ffffffff",
            INIT_5A => X"0000000d00000000ffffffbbfffffffffffffebfffffffffffffff78ffffffff",
            INIT_5B => X"0000008b000000000000002000000000ffffffebffffffff0000006400000000",
            INIT_5C => X"fffffeefffffffffffffffe8ffffffff0000008a00000000ffffffbaffffffff",
            INIT_5D => X"000000ca0000000000000102000000000000003f00000000fffffff2ffffffff",
            INIT_5E => X"000000ab00000000fffffff8ffffffff0000000e00000000ffffffccffffffff",
            INIT_5F => X"ffffffb9ffffffffffffffb7ffffffffffffff8dffffffffffffffecffffffff",
            INIT_60 => X"ffffff81ffffffff0000007c000000000000004e00000000ffffffc9ffffffff",
            INIT_61 => X"ffffff6affffffffffffffaaffffffffffffff7cffffffff0000001500000000",
            INIT_62 => X"0000003a00000000000000800000000000000067000000000000000900000000",
            INIT_63 => X"0000003400000000fffffffdffffffff00000069000000000000010400000000",
            INIT_64 => X"fffffff4fffffffffffffff1ffffffffffffffd9ffffffffffffffd4ffffffff",
            INIT_65 => X"fffffffbffffffff0000000900000000fffffff9ffffffffffffffd4ffffffff",
            INIT_66 => X"fffffffeffffffff0000000d00000000fffffffaffffffffffffffedffffffff",
            INIT_67 => X"00000041000000000000005a00000000fffffff4ffffffff0000001400000000",
            INIT_68 => X"ffffffc3ffffffffffffffe0ffffffff00000069000000000000004600000000",
            INIT_69 => X"0000006a000000000000002e00000000ffffffb3ffffffffffffffebffffffff",
            INIT_6A => X"0000003f0000000000000001000000000000009b000000000000001200000000",
            INIT_6B => X"ffffff33ffffffffffffff8cffffffff0000002b00000000ffffffb7ffffffff",
            INIT_6C => X"ffffffd1ffffffff0000000e000000000000004b000000000000004500000000",
            INIT_6D => X"ffffffb8ffffffffffffffa8ffffffff0000004900000000ffffffb7ffffffff",
            INIT_6E => X"000000d100000000000000120000000000000086000000000000001200000000",
            INIT_6F => X"ffffff34ffffffff00000027000000000000012e00000000ffffff4effffffff",
            INIT_70 => X"000000a400000000ffffff73fffffffffffffee8ffffffffffffff4effffffff",
            INIT_71 => X"ffffffb5ffffffff000000b8000000000000000500000000ffffff1fffffffff",
            INIT_72 => X"fffffeaeffffffffffffff71ffffffff0000008c00000000fffffff8ffffffff",
            INIT_73 => X"0000006e00000000fffffee5ffffffffffffff8affffffffffffff62ffffffff",
            INIT_74 => X"000000db00000000ffffff3bffffffffffffff7cffffffffffffff41ffffffff",
            INIT_75 => X"0000006c0000000000000032000000000000007800000000fffffffeffffffff",
            INIT_76 => X"0000003a00000000000000c0000000000000003200000000ffffffffffffffff",
            INIT_77 => X"ffffffc9ffffffff0000003f00000000fffffff6ffffffff0000001700000000",
            INIT_78 => X"fffffe35ffffffffffffffc3ffffffff0000001300000000fffffefdffffffff",
            INIT_79 => X"0000001900000000fffffffdffffffff00000175000000000000004100000000",
            INIT_7A => X"00000086000000000000002400000000ffffffc7ffffffff0000000800000000",
            INIT_7B => X"000000fd00000000ffffffe1ffffffff0000014100000000ffffffa4ffffffff",
            INIT_7C => X"ffffffe5ffffffffffffff03ffffffffffffffb6ffffffff0000004a00000000",
            INIT_7D => X"ffffff23ffffffff0000001e00000000ffffff8cffffffffffffffceffffffff",
            INIT_7E => X"000000370000000000000050000000000000001200000000ffffffb3ffffffff",
            INIT_7F => X"ffffffddffffffffffffffffffffffff00000008000000000000002000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE17;


    MEM_IWGHT_LAYER2_INSTANCE18 : if BRAM_NAME = "iwght_layer2_instance18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005700000000000000ae00000000ffffffdeffffffff0000007d00000000",
            INIT_01 => X"000000c20000000000000057000000000000003d00000000ffffff7effffffff",
            INIT_02 => X"ffffffffffffffff00000001000000000000002600000000ffffffe7ffffffff",
            INIT_03 => X"0000009a000000000000008c00000000fffffff9ffffffff0000004100000000",
            INIT_04 => X"0000003f00000000ffffff01ffffffffffffff8effffffffffffff6cffffffff",
            INIT_05 => X"ffffffebffffffffffffffd4ffffffff0000003e000000000000005c00000000",
            INIT_06 => X"0000007400000000fffffffcffffffffffffffedffffffff0000006600000000",
            INIT_07 => X"0000004a00000000ffffffc4ffffffffffffff8affffffff0000003400000000",
            INIT_08 => X"fffffee2ffffffff000000ad00000000ffffffccffffffff0000000300000000",
            INIT_09 => X"ffffffe9ffffffffffffff33ffffffffffffff12ffffffff0000006a00000000",
            INIT_0A => X"0000000c00000000ffffffb1ffffffffffffff33ffffffff0000004000000000",
            INIT_0B => X"0000009d00000000ffffffaffffffffffffffeedffffffff0000004900000000",
            INIT_0C => X"0000002800000000fffffed8ffffffffffffff70ffffffffffffff8dffffffff",
            INIT_0D => X"ffffff86ffffffffffffffa7fffffffffffffffcffffffffffffffa0ffffffff",
            INIT_0E => X"0000004e000000000000000200000000ffffff8effffffff0000001500000000",
            INIT_0F => X"0000003000000000ffffffbdfffffffffffffeb3ffffffffffffff6affffffff",
            INIT_10 => X"ffffff64ffffffffffffff5ffffffffffffffe8afffffffffffffe9affffffff",
            INIT_11 => X"ffffffe5ffffffff0000001700000000ffffff00fffffffffffffefeffffffff",
            INIT_12 => X"0000016700000000fffffcd6ffffffff0000004400000000ffffff5effffffff",
            INIT_13 => X"0000001200000000ffffff7cffffffff000000ae00000000000000b700000000",
            INIT_14 => X"0000007b00000000000000c000000000000000c700000000000000bd00000000",
            INIT_15 => X"ffffffe2ffffffff0000000100000000fffffff4fffffffffffffeaeffffffff",
            INIT_16 => X"ffffffd0ffffffff00000021000000000000005700000000fffffff7ffffffff",
            INIT_17 => X"0000001c00000000ffffffc8ffffffff00000094000000000000002400000000",
            INIT_18 => X"00000051000000000000002700000000ffffffe7ffffffff000000a200000000",
            INIT_19 => X"00000002000000000000003800000000fffffe61ffffffff000000e800000000",
            INIT_1A => X"00000013000000000000000400000000ffffffc7ffffffff000000f100000000",
            INIT_1B => X"fffffea3ffffffffffffff21fffffffffffffe66ffffffffffffff69ffffffff",
            INIT_1C => X"00000068000000000000001400000000ffffff81ffffffffffffff6effffffff",
            INIT_1D => X"ffffff14fffffffffffffff7ffffffff000000a4000000000000002400000000",
            INIT_1E => X"fffffff0ffffffffffffffbaffffffffffffffeeffffffff0000001d00000000",
            INIT_1F => X"ffffff94fffffffffffffff0ffffffffffffffb7ffffffff0000005a00000000",
            INIT_20 => X"0000006000000000ffffff74ffffffffffffffd2fffffffffffffe6bffffffff",
            INIT_21 => X"0000009700000000ffffffb4ffffffff0000002a000000000000003100000000",
            INIT_22 => X"00000080000000000000000b00000000000000fa00000000ffffffc1ffffffff",
            INIT_23 => X"ffffff81ffffffff0000004600000000ffffff4fffffffffffffffd5ffffffff",
            INIT_24 => X"ffffffdcfffffffffffffdcfffffffff0000000d00000000000000e000000000",
            INIT_25 => X"ffffffb3ffffffff0000011c000000000000004200000000ffffff98ffffffff",
            INIT_26 => X"ffffffc6ffffffffffffffb4ffffffff000000ac00000000ffffff66ffffffff",
            INIT_27 => X"0000008a00000000ffffffa7ffffffffffffff39ffffffff0000007000000000",
            INIT_28 => X"0000003800000000000000f200000000ffffff33ffffffff0000002800000000",
            INIT_29 => X"00000014000000000000000000000000ffffffccffffffffffffff50ffffffff",
            INIT_2A => X"0000002100000000000000350000000000000046000000000000007000000000",
            INIT_2B => X"0000010c00000000fffffe4dffffffffffffff64ffffffffffffffd0ffffffff",
            INIT_2C => X"ffffffbeffffffffffffffb2fffffffffffffe61ffffffff0000010e00000000",
            INIT_2D => X"00000011000000000000000b00000000ffffffedffffffff0000009100000000",
            INIT_2E => X"fffffff6ffffffff0000000d000000000000000400000000fffffff2ffffffff",
            INIT_2F => X"fffffefbffffffffffffff3dfffffffffffffff1ffffffff0000000000000000",
            INIT_30 => X"ffffffb2fffffffffffffef7ffffffff0000003a00000000ffffffc9ffffffff",
            INIT_31 => X"ffffffb6fffffffffffffff4ffffffffffffffafffffffff0000007d00000000",
            INIT_32 => X"00000057000000000000001000000000000000bc000000000000006100000000",
            INIT_33 => X"0000000700000000ffffffeaffffffff00000011000000000000001200000000",
            INIT_34 => X"ffffffc3fffffffffffffff7ffffffffffffff55ffffffff0000007900000000",
            INIT_35 => X"ffffffa2ffffffffffffff32ffffffff0000007300000000fffffff5ffffffff",
            INIT_36 => X"0000001c00000000fffffef3ffffffff0000012a000000000000007900000000",
            INIT_37 => X"ffffff41ffffffff00000037000000000000001c00000000ffffffb8ffffffff",
            INIT_38 => X"ffffffddfffffffffffffff8ffffffff0000008c000000000000006000000000",
            INIT_39 => X"00000053000000000000001200000000ffffffc7ffffffffffffffcbffffffff",
            INIT_3A => X"000000160000000000000000000000000000000e00000000ffffffecffffffff",
            INIT_3B => X"0000009800000000ffffffb6ffffffff000000ab00000000fffffe77ffffffff",
            INIT_3C => X"00000063000000000000003c000000000000000f00000000ffffffdbffffffff",
            INIT_3D => X"ffffff51ffffffffffffff95ffffffff00000036000000000000002000000000",
            INIT_3E => X"fffffff2ffffffffffffffb9ffffffffffffff86ffffffff0000004400000000",
            INIT_3F => X"0000006c00000000000000cd00000000ffffff65ffffffff0000009e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffbcffffffffffffffd0ffffffff00000028000000000000006b00000000",
            INIT_41 => X"ffffff3bffffffff0000004100000000ffffffadffffffff0000000a00000000",
            INIT_42 => X"000001d100000000fffffecaffffffffffffffbeffffffff0000001f00000000",
            INIT_43 => X"00000077000000000000006a00000000ffffffe1ffffffffffffffb4ffffffff",
            INIT_44 => X"00000089000000000000000600000000fffffdaeffffffffffffff4effffffff",
            INIT_45 => X"ffffff4bffffffff000000080000000000000066000000000000006100000000",
            INIT_46 => X"ffffffb6ffffffff000000b200000000000000e000000000ffffff92ffffffff",
            INIT_47 => X"ffffffa2ffffffff00000064000000000000007900000000ffffffe3ffffffff",
            INIT_48 => X"fffffffbfffffffffffffeeaffffffff0000006e00000000ffffff49ffffffff",
            INIT_49 => X"fffffff8ffffffffffffffbeffffffff0000004a00000000000000ae00000000",
            INIT_4A => X"0000001f00000000ffffffe6ffffffff0000000d000000000000002800000000",
            INIT_4B => X"ffffff7dffffffffffffffceffffffff000000a300000000ffffffadffffffff",
            INIT_4C => X"00000067000000000000001b000000000000002c000000000000000b00000000",
            INIT_4D => X"00000037000000000000004b00000000ffffff77ffffffff0000004900000000",
            INIT_4E => X"0000008a00000000ffffffdfffffffff0000003400000000ffffffeaffffffff",
            INIT_4F => X"ffffffb7ffffffffffffffa7ffffffff0000000400000000000000dc00000000",
            INIT_50 => X"fffffff5ffffffff000000400000000000000017000000000000008800000000",
            INIT_51 => X"fffffee7fffffffffffffee7ffffffffffffff0bfffffffffffffffaffffffff",
            INIT_52 => X"00000005000000000000006600000000ffffff90ffffffff000000d700000000",
            INIT_53 => X"0000009500000000fffffee4ffffffffffffffcaffffffff0000006500000000",
            INIT_54 => X"ffffffdeffffffffffffffc2ffffffff00000014000000000000003f00000000",
            INIT_55 => X"ffffffc9ffffffffffffffc9fffffffffffffff8ffffffffffffff7cffffffff",
            INIT_56 => X"00000001000000000000000a000000000000008c00000000ffffffe9ffffffff",
            INIT_57 => X"0000004a00000000ffffff7affffffff0000000b00000000ffffff60ffffffff",
            INIT_58 => X"0000005c0000000000000082000000000000006f000000000000007300000000",
            INIT_59 => X"0000006c00000000000000140000000000000060000000000000009700000000",
            INIT_5A => X"0000004400000000ffffffa5fffffffffffffff0ffffffff0000008200000000",
            INIT_5B => X"ffffffa6ffffffff0000007a00000000ffffff82ffffffffffffffa5ffffffff",
            INIT_5C => X"00000005000000000000002a00000000fffffff9ffffffff0000002600000000",
            INIT_5D => X"000000a7000000000000006900000000ffffff2cffffffffffffff7dffffffff",
            INIT_5E => X"ffffffdeffffffff00000049000000000000008600000000ffffffd7ffffffff",
            INIT_5F => X"00000004000000000000000300000000ffffffc2ffffffffffffffccffffffff",
            INIT_60 => X"0000005900000000ffffffbdffffffff0000005200000000ffffffedffffffff",
            INIT_61 => X"ffffff89ffffffffffffffb7ffffffffffffff67ffffffffffffffaaffffffff",
            INIT_62 => X"ffffff5cffffffffffffffb4fffffffffffffeedffffffffffffff2bffffffff",
            INIT_63 => X"0000008900000000ffffffbdffffffff0000007500000000ffffff01ffffffff",
            INIT_64 => X"000000e100000000fffffffdffffffff00000072000000000000008800000000",
            INIT_65 => X"00000001000000000000000d00000000ffffffe3ffffffff0000009900000000",
            INIT_66 => X"ffffff97ffffffffffffff97ffffffff00000043000000000000003700000000",
            INIT_67 => X"0000002800000000ffffffe2ffffffffffffff96ffffffffffffffe8ffffffff",
            INIT_68 => X"0000008800000000000000780000000000000030000000000000008900000000",
            INIT_69 => X"0000006100000000fffffffdffffffff0000006b000000000000002e00000000",
            INIT_6A => X"fffffff5ffffffff000000590000000000000042000000000000007900000000",
            INIT_6B => X"ffffff6affffffff000000050000000000000047000000000000001400000000",
            INIT_6C => X"0000002e00000000ffffffedffffffff0000002f000000000000004f00000000",
            INIT_6D => X"0000004400000000ffffff82ffffffffffffffffffffffffffffff94ffffffff",
            INIT_6E => X"00000084000000000000003100000000ffffff62ffffffff0000001900000000",
            INIT_6F => X"000000aa000000000000011300000000000000f2000000000000000b00000000",
            INIT_70 => X"ffffff9bffffffff0000008e0000000000000084000000000000009a00000000",
            INIT_71 => X"ffffffc0ffffffffffffff78ffffffff0000001d00000000ffffff8cffffffff",
            INIT_72 => X"ffffffdefffffffffffffff8ffffffffffffffc3ffffffffffffff6affffffff",
            INIT_73 => X"ffffffc0ffffffff0000003400000000fffffff1ffffffff0000002d00000000",
            INIT_74 => X"fffffee5ffffffff0000003400000000ffffff9cffffffffffffffffffffffff",
            INIT_75 => X"ffffffeeffffffff00000004000000000000000100000000ffffff9fffffffff",
            INIT_76 => X"0000000800000000fffffffdfffffffffffffff8ffffffff0000000900000000",
            INIT_77 => X"fffffff7fffffffffffffff7ffffffff00000005000000000000001a00000000",
            INIT_78 => X"ffffff8ffffffffffffffff4ffffffffffffffc9ffffffffffffffe6ffffffff",
            INIT_79 => X"0000004e00000000ffffffd9fffffffffffffff8ffffffffffffffeeffffffff",
            INIT_7A => X"ffffff9dffffffffffffff8bffffffff0000005500000000ffffffcdffffffff",
            INIT_7B => X"0000005c00000000ffffffdeffffffff0000001c000000000000004f00000000",
            INIT_7C => X"0000001400000000000000670000000000000085000000000000000000000000",
            INIT_7D => X"ffffffaeffffffffffffffd6ffffffff0000002200000000000000bf00000000",
            INIT_7E => X"fffffffafffffffffffffea4ffffffffffffffedffffffff0000001c00000000",
            INIT_7F => X"0000009100000000fffffef3ffffffff0000008c000000000000008800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE18;


    MEM_IWGHT_LAYER2_INSTANCE19 : if BRAM_NAME = "iwght_layer2_instance19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a8000000000000000700000000ffffffa9ffffffff000000e100000000",
            INIT_01 => X"ffffffcffffffffffffffffeffffffff0000004500000000ffffff9bffffffff",
            INIT_02 => X"000000c5000000000000009000000000000000a300000000ffffffaeffffffff",
            INIT_03 => X"00000062000000000000003900000000fffffffaffffffff0000004800000000",
            INIT_04 => X"0000002a000000000000008500000000ffffffc6ffffffffffffffe1ffffffff",
            INIT_05 => X"ffffff9affffffffffffffd6ffffffff0000009b00000000ffffff9affffffff",
            INIT_06 => X"0000003900000000ffffffacffffffffffffff99ffffffff0000000c00000000",
            INIT_07 => X"fffffffcffffffff00000005000000000000000400000000ffffffe9ffffffff",
            INIT_08 => X"ffffff68ffffffff00000023000000000000000600000000ffffff59ffffffff",
            INIT_09 => X"0000006c00000000ffffff88fffffffffffffff7ffffffffffffff83ffffffff",
            INIT_0A => X"0000001500000000fffffffeffffffffffffff96ffffffffffffffdaffffffff",
            INIT_0B => X"ffffffe5fffffffffffffff8fffffffffffffed5ffffffff000000d500000000",
            INIT_0C => X"ffffffd0ffffffffffffffc5ffffffff0000002600000000ffffffa3ffffffff",
            INIT_0D => X"ffffff3effffffff00000036000000000000005200000000ffffff10ffffffff",
            INIT_0E => X"0000001f00000000fffffff7ffffffffffffffcbffffffff0000000600000000",
            INIT_0F => X"0000001400000000ffffffbbffffffff00000025000000000000002f00000000",
            INIT_10 => X"ffffff8dffffffffffffff62ffffffff0000000400000000fffffffbffffffff",
            INIT_11 => X"ffffffa9ffffffffffffffdefffffffffffffff6ffffffffffffffccffffffff",
            INIT_12 => X"00000012000000000000008500000000ffffffceffffffffffffff5cffffffff",
            INIT_13 => X"0000005c00000000ffffff7fffffffffffffffe0ffffffff0000004600000000",
            INIT_14 => X"ffffffb0ffffffffffffff99ffffffff0000002d00000000ffffff37ffffffff",
            INIT_15 => X"fffffe4affffffff0000000000000000ffffff6dffffffffffffffbdffffffff",
            INIT_16 => X"ffffff33ffffffffffffffd6ffffffffffffffbbffffffffffffffe1ffffffff",
            INIT_17 => X"ffffffb8ffffffffffffffa4fffffffffffffffeffffffffffffffb6ffffffff",
            INIT_18 => X"0000003c000000000000002e000000000000002900000000fffffff0ffffffff",
            INIT_19 => X"ffffffb6ffffffff0000005400000000ffffff37ffffffff0000007800000000",
            INIT_1A => X"0000000300000000ffffffaeffffffffffffffc9ffffffffffffff61ffffffff",
            INIT_1B => X"ffffff79ffffffffffffffdbffffffffffffff26fffffffffffffef1ffffffff",
            INIT_1C => X"ffffffffffffffff0000000100000000000000a000000000ffffff83ffffffff",
            INIT_1D => X"ffffffbaffffffff00000097000000000000010200000000ffffffdeffffffff",
            INIT_1E => X"0000000800000000fffffff4ffffffff00000048000000000000009f00000000",
            INIT_1F => X"0000006100000000ffffffa3ffffffffffffff4efffffffffffffff1ffffffff",
            INIT_20 => X"ffffffd0ffffffffffffffcfffffffffffffffb1ffffffffffffff5effffffff",
            INIT_21 => X"ffffff79ffffffffffffff90ffffffff0000004b000000000000007f00000000",
            INIT_22 => X"ffffffd5ffffffff000000a100000000ffffff37ffffffff0000006000000000",
            INIT_23 => X"0000004900000000ffffff54ffffffffffffffd8ffffffffffffff92ffffffff",
            INIT_24 => X"0000000f000000000000006700000000ffffffe4ffffffffffffffe8ffffffff",
            INIT_25 => X"ffffffabfffffffffffffffdffffffffffffffedffffffffffffffdcffffffff",
            INIT_26 => X"0000009f00000000fffffff3ffffffffffffff9affffffff0000000a00000000",
            INIT_27 => X"00000068000000000000010800000000ffffffcaffffffffffffff48ffffffff",
            INIT_28 => X"ffffff86ffffffff0000001b00000000ffffffe0ffffffffffffffc8ffffffff",
            INIT_29 => X"0000005f00000000ffffffffffffffffffffffe4ffffffffffffffaaffffffff",
            INIT_2A => X"0000002d000000000000001d000000000000007a000000000000011700000000",
            INIT_2B => X"000000a300000000ffffffb2ffffffffffffffb5fffffffffffffff2ffffffff",
            INIT_2C => X"00000000000000000000000a000000000000001f00000000ffffffa2ffffffff",
            INIT_2D => X"ffffffd4ffffffff00000028000000000000002e000000000000001a00000000",
            INIT_2E => X"0000002400000000000000560000000000000029000000000000000a00000000",
            INIT_2F => X"0000002500000000ffffff8fffffffffffffffefffffffff000000a700000000",
            INIT_30 => X"ffffffedffffffffffffffcbffffffff0000004600000000ffffff88ffffffff",
            INIT_31 => X"ffffffabffffffff0000000a000000000000008000000000ffffff63ffffffff",
            INIT_32 => X"fffffeb6ffffffff00000025000000000000007500000000ffffffecffffffff",
            INIT_33 => X"000000cc0000000000000018000000000000000d00000000ffffff5cffffffff",
            INIT_34 => X"ffffffdffffffffffffffffbffffffffffffff03ffffffffffffffc3ffffffff",
            INIT_35 => X"ffffff21ffffffff000001000000000000000117000000000000001300000000",
            INIT_36 => X"fffffff1fffffffffffffffeffffffff00000062000000000000008600000000",
            INIT_37 => X"ffffffbdffffffffffffff37ffffffff0000001800000000ffffffd4ffffffff",
            INIT_38 => X"0000002900000000000000a30000000000000091000000000000000000000000",
            INIT_39 => X"ffffff26ffffffff00000006000000000000002500000000000000b700000000",
            INIT_3A => X"fffffff3ffffffff00000028000000000000009500000000ffffff61ffffffff",
            INIT_3B => X"0000004100000000ffffffa7ffffffffffffffb1ffffffff0000005b00000000",
            INIT_3C => X"ffffffd7ffffffffffffffdfffffffff0000000f000000000000000000000000",
            INIT_3D => X"ffffffecffffffff0000000f000000000000000800000000fffffff6ffffffff",
            INIT_3E => X"ffffffedffffffffffffffecffffffff00000012000000000000000900000000",
            INIT_3F => X"ffffffe9ffffffffffffffcbffffffff00000007000000000000000a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004f000000000000000f00000000ffffffdfffffffff0000003b00000000",
            INIT_41 => X"0000003000000000000000ef00000000fffffff5ffffffffffffff3fffffffff",
            INIT_42 => X"00000090000000000000006f00000000ffffff9dffffffff0000005600000000",
            INIT_43 => X"000000ae00000000ffffff7fffffffffffffff1cffffffffffffffecffffffff",
            INIT_44 => X"0000000f000000000000006e00000000000000a8000000000000005900000000",
            INIT_45 => X"0000003800000000ffffffaaffffffffffffffaaffffffffffffff8effffffff",
            INIT_46 => X"0000000700000000fffffe45ffffffffffffffeeffffffff0000009100000000",
            INIT_47 => X"ffffffa1ffffffff000000ab00000000ffffff0affffffff0000011c00000000",
            INIT_48 => X"0000001d000000000000002000000000ffffffb6ffffffff0000012b00000000",
            INIT_49 => X"0000001a00000000ffffffd5ffffffff0000001200000000ffffff99ffffffff",
            INIT_4A => X"000000ce00000000ffffff69ffffffffffffff85ffffffffffffffb9ffffffff",
            INIT_4B => X"0000002300000000ffffff61ffffffffffffff81ffffffffffffffd0ffffffff",
            INIT_4C => X"0000007f0000000000000007000000000000001600000000ffffffd5ffffffff",
            INIT_4D => X"0000004200000000ffffff1affffffff0000008a000000000000004000000000",
            INIT_4E => X"0000000c00000000ffffffb9ffffffffffffff34ffffffffffffff42ffffffff",
            INIT_4F => X"0000006c00000000ffffffb6ffffffff0000005b00000000ffffffd4ffffffff",
            INIT_50 => X"0000007b00000000ffffff8bffffffffffffffdcffffffff0000001300000000",
            INIT_51 => X"ffffffbbffffffff00000072000000000000004f00000000fffffeaaffffffff",
            INIT_52 => X"ffffffedffffffff0000006c000000000000005900000000ffffffeaffffffff",
            INIT_53 => X"0000001f00000000000000b2000000000000007900000000ffffff5bffffffff",
            INIT_54 => X"ffffffaeffffffffffffff82ffffffffffffff82ffffffff0000006100000000",
            INIT_55 => X"00000096000000000000001e000000000000004900000000fffffff3ffffffff",
            INIT_56 => X"ffffff3effffffffffffff66ffffffff0000000900000000ffffff74ffffffff",
            INIT_57 => X"000000b800000000ffffffe9fffffffffffffe12ffffffff000000d600000000",
            INIT_58 => X"ffffffdefffffffffffffff1ffffffff000000a500000000ffffff6affffffff",
            INIT_59 => X"0000006900000000ffffffa6ffffffff0000000c000000000000001c00000000",
            INIT_5A => X"00000037000000000000001d00000000ffffffaaffffffffffffffc3ffffffff",
            INIT_5B => X"ffffffd7ffffffff0000005f0000000000000067000000000000003900000000",
            INIT_5C => X"0000003100000000ffffff71fffffffffffffff5ffffffff0000002c00000000",
            INIT_5D => X"ffffff4fffffffff0000007300000000fffffffaffffffffffffffb7ffffffff",
            INIT_5E => X"000000d0000000000000007000000000ffffffe0ffffffffffffff91ffffffff",
            INIT_5F => X"ffffffc6ffffffff0000005500000000ffffff3affffffffffffff78ffffffff",
            INIT_60 => X"ffffffbeffffffff0000003800000000ffffffc4ffffffff0000001a00000000",
            INIT_61 => X"000000a600000000ffffff32ffffffff0000003c000000000000000a00000000",
            INIT_62 => X"ffffffe0ffffffff00000007000000000000000300000000ffffffd0ffffffff",
            INIT_63 => X"0000005f000000000000002e0000000000000018000000000000008b00000000",
            INIT_64 => X"ffffff23ffffffffffffff8bffffffffffffffc2ffffffffffffff8dffffffff",
            INIT_65 => X"fffffff0ffffffff0000008a000000000000008300000000000000b600000000",
            INIT_66 => X"0000006400000000000000a600000000ffffffd7ffffffff0000002100000000",
            INIT_67 => X"ffffff03ffffffffffffffb6ffffffffffffff63fffffffffffffffbffffffff",
            INIT_68 => X"ffffffe7ffffffff0000000c00000000fffffffbffffffff0000000200000000",
            INIT_69 => X"fffffffdffffffffffffffebfffffffffffffff2ffffffff0000000500000000",
            INIT_6A => X"ffffffecffffffff00000006000000000000000100000000ffffffebffffffff",
            INIT_6B => X"ffffffe5fffffffffffffffeffffffffffffffe8ffffffff0000000200000000",
            INIT_6C => X"fffffff0fffffffffffffff2fffffffffffffffeffffffffffffffffffffffff",
            INIT_6D => X"fffffff3fffffffffffffff5ffffffffffffffdeffffffff0000000600000000",
            INIT_6E => X"fffffff6ffffffff0000000000000000ffffffeefffffffffffffff6ffffffff",
            INIT_6F => X"0000000700000000fffffff9fffffffffffffffbffffffff0000000e00000000",
            INIT_70 => X"0000000200000000fffffff6ffffffffffffffedfffffffffffffff7ffffffff",
            INIT_71 => X"ffffffe5ffffffff000000050000000000000000000000000000000800000000",
            INIT_72 => X"0000000400000000ffffffe7ffffffffffffffeaffffffffffffffebffffffff",
            INIT_73 => X"fffffffefffffffffffffff2fffffffffffffff4ffffffffffffffe7ffffffff",
            INIT_74 => X"fffffff3ffffffff00000005000000000000000900000000fffffffbffffffff",
            INIT_75 => X"fffffff0fffffffffffffff0ffffffff0000000c00000000fffffff0ffffffff",
            INIT_76 => X"fffffff0ffffffff0000000c00000000ffffffe8fffffffffffffffcffffffff",
            INIT_77 => X"fffffff3ffffffff0000000900000000fffffff7fffffffffffffffbffffffff",
            INIT_78 => X"ffffffffffffffffffffffefffffffff0000001000000000fffffff4ffffffff",
            INIT_79 => X"fffffff2ffffffffffffffebffffffffffffffe8ffffffff0000000900000000",
            INIT_7A => X"ffffffe5fffffffffffffffbffffffff0000000700000000ffffffe3ffffffff",
            INIT_7B => X"fffffff0fffffffffffffff8fffffffffffffff5fffffffffffffffaffffffff",
            INIT_7C => X"0000000100000000ffffffe5ffffffffffffffefffffffff0000000000000000",
            INIT_7D => X"00000005000000000000000100000000ffffffe6ffffffffffffffefffffffff",
            INIT_7E => X"fffffff8ffffffff00000007000000000000000900000000ffffffecffffffff",
            INIT_7F => X"00000004000000000000000000000000fffffff5ffffffffffffffebffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE19;


    MEM_IWGHT_LAYER2_INSTANCE20 : if BRAM_NAME = "iwght_layer2_instance20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000100000000ffffffffffffffffffffffebffffffffffffffeeffffffff",
            INIT_01 => X"ffffffe8fffffffffffffff1ffffffff0000000100000000ffffffefffffffff",
            INIT_02 => X"ffffffedffffffffffffffe2ffffffffffffffe1fffffffffffffffcffffffff",
            INIT_03 => X"0000000000000000ffffffffffffffffffffffe9ffffffff0000000000000000",
            INIT_04 => X"ffffffeffffffffffffffffbffffffffffffffe4ffffffffffffffefffffffff",
            INIT_05 => X"0000000100000000fffffffdffffffffffffffeffffffffffffffff5ffffffff",
            INIT_06 => X"fffffff0ffffffff00000006000000000000000700000000fffffff4ffffffff",
            INIT_07 => X"fffffff4fffffffffffffffbffffffff00000016000000000000000900000000",
            INIT_08 => X"0000000e00000000ffffffe9ffffffffffffffeafffffffffffffffeffffffff",
            INIT_09 => X"fffffff9ffffffff0000000100000000fffffff3fffffffffffffffbffffffff",
            INIT_0A => X"ffffffe4ffffffffffffffedfffffffffffffff9fffffffffffffff0ffffffff",
            INIT_0B => X"ffffffe8ffffffff00000000000000000000000a00000000fffffff7ffffffff",
            INIT_0C => X"0000000400000000ffffffecffffffff0000000700000000ffffffecffffffff",
            INIT_0D => X"fffffff4ffffffffffffffe9ffffffff0000000000000000ffffffebffffffff",
            INIT_0E => X"fffffffcffffffffffffffe5ffffffff0000000100000000fffffff3ffffffff",
            INIT_0F => X"fffffffdffffffff0000000800000000fffffff6ffffffff0000000b00000000",
            INIT_10 => X"00000009000000000000000200000000ffffffeffffffffffffffffdffffffff",
            INIT_11 => X"fffffff7ffffffff0000000d00000000ffffffe9ffffffff0000000100000000",
            INIT_12 => X"000000020000000000000008000000000000000d00000000fffffffeffffffff",
            INIT_13 => X"ffffffefffffffff0000000200000000fffffff5fffffffffffffff5ffffffff",
            INIT_14 => X"ffffffe8fffffffffffffff2ffffffff0000000900000000fffffffaffffffff",
            INIT_15 => X"00000002000000000000000900000000ffffffeeffffffffffffffe9ffffffff",
            INIT_16 => X"fffffffafffffffffffffff8ffffffffffffffeefffffffffffffff2ffffffff",
            INIT_17 => X"0000000600000000fffffffffffffffffffffff8ffffffffffffffe6ffffffff",
            INIT_18 => X"fffffffcfffffffffffffffaffffffff00000008000000000000000300000000",
            INIT_19 => X"0000000e000000000000000c00000000fffffff4fffffffffffffff6ffffffff",
            INIT_1A => X"00000003000000000000000c00000000ffffffecffffffffffffffffffffffff",
            INIT_1B => X"ffffffe6fffffffffffffffafffffffffffffff6ffffffffffffffe7ffffffff",
            INIT_1C => X"fffffff5fffffffffffffff6ffffffffffffffe7ffffffffffffffedffffffff",
            INIT_1D => X"fffffff4ffffffffffffffefffffffffffffffe4fffffffffffffff8ffffffff",
            INIT_1E => X"fffffff4fffffffffffffffefffffffffffffff3fffffffffffffff9ffffffff",
            INIT_1F => X"ffffffeffffffffffffffff3ffffffff0000000900000000fffffff8ffffffff",
            INIT_20 => X"fffffff0ffffffff00000000000000000000000200000000fffffffbffffffff",
            INIT_21 => X"000000090000000000000007000000000000000b000000000000000000000000",
            INIT_22 => X"00000004000000000000001000000000ffffffedfffffffffffffffcffffffff",
            INIT_23 => X"fffffff3fffffffffffffff5ffffffff0000001200000000ffffffe3ffffffff",
            INIT_24 => X"fffffff7ffffffff0000000c00000000fffffff7fffffffffffffffbffffffff",
            INIT_25 => X"0000000200000000fffffffafffffffffffffff1ffffffff0000000700000000",
            INIT_26 => X"fffffff8ffffffffffffffe8ffffffff0000000500000000fffffff4ffffffff",
            INIT_27 => X"0000000400000000ffffffe9ffffffff00000008000000000000000500000000",
            INIT_28 => X"fffffffefffffffffffffff2ffffffff0000000000000000ffffffedffffffff",
            INIT_29 => X"ffffffe1ffffffff0000000700000000fffffff9ffffffff0000000a00000000",
            INIT_2A => X"fffffff7fffffffffffffff6fffffffffffffffcffffffff0000001000000000",
            INIT_2B => X"ffffffecffffffff00000009000000000000000700000000fffffffbffffffff",
            INIT_2C => X"000000050000000000000001000000000000000400000000ffffffecffffffff",
            INIT_2D => X"fffffffdffffffff0000000b00000000ffffffeafffffffffffffff1ffffffff",
            INIT_2E => X"ffffffe7fffffffffffffff3ffffffffffffffeeffffffffffffffffffffffff",
            INIT_2F => X"ffffffe0ffffffffffffffecffffffffffffffeeffffffffffffffe3ffffffff",
            INIT_30 => X"ffffffeeffffffffffffffaafffffffffffffff5ffffffff0000003e00000000",
            INIT_31 => X"000000890000000000000057000000000000007400000000ffffffd3ffffffff",
            INIT_32 => X"0000003200000000ffffffbfffffffff00000082000000000000006600000000",
            INIT_33 => X"ffffffe3fffffffffffffe56ffffffff0000009700000000ffffffeeffffffff",
            INIT_34 => X"0000009900000000ffffff7fffffffffffffffdfffffffff0000002800000000",
            INIT_35 => X"ffffff78ffffffffffffffa8ffffffff00000071000000000000003800000000",
            INIT_36 => X"ffffffe3fffffffffffffe89ffffffffffffff52ffffffff0000013300000000",
            INIT_37 => X"ffffffa6ffffffffffffff33ffffffff0000009a00000000ffffffe0ffffffff",
            INIT_38 => X"0000001800000000ffffffaefffffffffffffff6ffffffffffffffaaffffffff",
            INIT_39 => X"ffffff10ffffffff00000078000000000000005900000000ffffff52ffffffff",
            INIT_3A => X"0000000a00000000ffffffe0ffffffff00000070000000000000009900000000",
            INIT_3B => X"ffffff3fffffffffffffff53ffffffff00000017000000000000001400000000",
            INIT_3C => X"0000006400000000ffffffeaffffffff00000014000000000000005400000000",
            INIT_3D => X"0000000100000000ffffffd0ffffffff00000096000000000000002600000000",
            INIT_3E => X"ffffffe0ffffffff0000007c00000000fffffff6ffffffffffffff7effffffff",
            INIT_3F => X"0000003600000000ffffffebffffffff0000001700000000ffffffe9ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffa8ffffffff0000002b00000000ffffffffffffffffffffff2fffffffff",
            INIT_41 => X"ffffffdaffffffffffffffcdffffffff000000f000000000ffffffdbffffffff",
            INIT_42 => X"000000430000000000000060000000000000000600000000ffffff75ffffffff",
            INIT_43 => X"0000008d00000000ffffffceffffffff000000ff00000000ffffffbaffffffff",
            INIT_44 => X"ffffff87ffffffffffffffd4ffffffffffffffc8ffffffffffffffc2ffffffff",
            INIT_45 => X"fffffffdffffffff00000056000000000000006f000000000000001a00000000",
            INIT_46 => X"fffffed9ffffffff0000000e00000000fffffff7ffffffffffffffd8ffffffff",
            INIT_47 => X"ffffffb6ffffffffffffffc6ffffffff0000001200000000ffffff0fffffffff",
            INIT_48 => X"000000a30000000000000085000000000000008300000000fffffff6ffffffff",
            INIT_49 => X"00000016000000000000000b00000000ffffffa6ffffffff0000003500000000",
            INIT_4A => X"ffffff50ffffffff00000004000000000000000b000000000000009100000000",
            INIT_4B => X"00000022000000000000000d0000000000000093000000000000001d00000000",
            INIT_4C => X"ffffff97ffffffffffffff67ffffffff00000010000000000000000e00000000",
            INIT_4D => X"00000004000000000000000400000000ffffffe9ffffffffffffffcdffffffff",
            INIT_4E => X"fffffffcfffffffffffffff2fffffffffffffff8fffffffffffffffaffffffff",
            INIT_4F => X"0000008c00000000ffffff9cfffffffffffffff7ffffffff0000000800000000",
            INIT_50 => X"0000002800000000000000a100000000fffffff0ffffffffffffffefffffffff",
            INIT_51 => X"ffffff98ffffffff000000140000000000000030000000000000004000000000",
            INIT_52 => X"0000000300000000ffffffe9ffffffff000000dc000000000000005400000000",
            INIT_53 => X"0000005e000000000000000000000000fffffff3ffffffff000000d500000000",
            INIT_54 => X"ffffff69fffffffffffffed5ffffffffffffff06ffffffffffffff98ffffffff",
            INIT_55 => X"0000000600000000ffffffd6ffffffffffffffdfffffffffffffffadffffffff",
            INIT_56 => X"0000001200000000ffffffdaffffffff000000bf000000000000001800000000",
            INIT_57 => X"0000000600000000000000000000000000000082000000000000009c00000000",
            INIT_58 => X"ffffff35ffffffff0000002500000000ffffff3effffffff0000000400000000",
            INIT_59 => X"0000006b000000000000005c0000000000000084000000000000002a00000000",
            INIT_5A => X"ffffffe9ffffffffffffffdaffffffff0000009a000000000000001a00000000",
            INIT_5B => X"0000006200000000ffffff64ffffffffffffffc9fffffffffffffff1ffffffff",
            INIT_5C => X"0000000b00000000ffffff8cffffffff0000004f000000000000002800000000",
            INIT_5D => X"ffffffe8ffffffffffffff4cffffffffffffff73ffffffff0000009500000000",
            INIT_5E => X"0000004f00000000000000d400000000fffffff5ffffffffffffffa7ffffffff",
            INIT_5F => X"00000089000000000000005600000000ffffffa8ffffffffffffff3effffffff",
            INIT_60 => X"ffffff58ffffffffffffffd8ffffffff00000043000000000000000c00000000",
            INIT_61 => X"ffffff53ffffffff0000007e000000000000007d00000000ffffffafffffffff",
            INIT_62 => X"00000058000000000000002000000000fffffeeafffffffffffffff3ffffffff",
            INIT_63 => X"fffffff8ffffffff00000061000000000000009300000000ffffff28ffffffff",
            INIT_64 => X"ffffffb8ffffffff0000006900000000ffffffe1ffffffffffffffddffffffff",
            INIT_65 => X"0000001b000000000000004800000000ffffffd7ffffffff0000001400000000",
            INIT_66 => X"ffffffbaffffffffffffff72ffffffff0000004900000000ffffff8fffffffff",
            INIT_67 => X"ffffffc1ffffffff0000002700000000fffffed6ffffffffffffffdfffffffff",
            INIT_68 => X"00000011000000000000004d00000000ffffffc7ffffffffffffff9fffffffff",
            INIT_69 => X"0000004d00000000ffffffe3ffffffffffffffcdffffffff0000002700000000",
            INIT_6A => X"ffffffbaffffffff0000003c00000000fffffef6ffffffff0000003f00000000",
            INIT_6B => X"fffffff2ffffffffffffff9bffffffff00000072000000000000002b00000000",
            INIT_6C => X"ffffffc9ffffffffffffffb0ffffffffffffff52ffffffffffffffaaffffffff",
            INIT_6D => X"ffffffe9ffffffffffffffb4ffffffff00000012000000000000002f00000000",
            INIT_6E => X"fffffff4fffffffffffffff6ffffffffffffff2effffffff0000000d00000000",
            INIT_6F => X"ffffffb0ffffffffffffff8bffffffff0000001f000000000000007100000000",
            INIT_70 => X"ffffffe3ffffffff000000330000000000000002000000000000004f00000000",
            INIT_71 => X"0000007f00000000ffffffdaffffffff0000009b000000000000004200000000",
            INIT_72 => X"ffffff98fffffffffffffffcffffffff0000000100000000ffffffcdffffffff",
            INIT_73 => X"fffffff0ffffffff0000006c0000000000000037000000000000009100000000",
            INIT_74 => X"ffffff82ffffffff0000001400000000ffffffecffffffffffffff92ffffffff",
            INIT_75 => X"00000011000000000000008900000000ffffffb8ffffffffffffffa4ffffffff",
            INIT_76 => X"ffffffc2ffffffffffffffa7ffffffffffffffbaffffffff0000006500000000",
            INIT_77 => X"0000008f00000000fffffffcffffffff0000006f00000000ffffffb6ffffffff",
            INIT_78 => X"ffffff1dffffffffffffffedffffffff0000005300000000000000b600000000",
            INIT_79 => X"ffffff14ffffffffffffff5effffffffffffff8ffffffffffffffe8dffffffff",
            INIT_7A => X"00000005000000000000006500000000ffffffd1ffffffffffffff8fffffffff",
            INIT_7B => X"00000027000000000000009d00000000ffffff4fffffffff0000002000000000",
            INIT_7C => X"fffffff3ffffffffffffffb9ffffffffffffffa6ffffffff0000005100000000",
            INIT_7D => X"0000007a00000000ffffffc6ffffffffffffffb8ffffffff0000000500000000",
            INIT_7E => X"0000005400000000ffffffe3ffffffff0000004300000000000000c200000000",
            INIT_7F => X"ffffffdeffffffff0000002b000000000000012a00000000ffffffbdffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE20;


    MEM_IWGHT_LAYER2_INSTANCE21 : if BRAM_NAME = "iwght_layer2_instance21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffff62ffffffffffffff9fffffffff00000021000000000000002c00000000",
            INIT_01 => X"0000000f00000000ffffffe9ffffffffffffffcfffffffffffffff3fffffffff",
            INIT_02 => X"ffffff4effffffff0000007600000000ffffffa4fffffffffffffef2ffffffff",
            INIT_03 => X"0000009b000000000000005e00000000000000a400000000ffffff8effffffff",
            INIT_04 => X"fffffffcffffffff00000019000000000000005200000000ffffffc4ffffffff",
            INIT_05 => X"000000530000000000000068000000000000000c000000000000003900000000",
            INIT_06 => X"ffffffb7ffffffff000000a500000000000000d2000000000000005700000000",
            INIT_07 => X"0000008f0000000000000012000000000000005f00000000ffffffc0ffffffff",
            INIT_08 => X"ffffffe1fffffffffffffff6fffffffffffffff0ffffffffffffffabffffffff",
            INIT_09 => X"ffffffd6ffffffffffffffb1ffffffffffffffc8ffffffff0000007d00000000",
            INIT_0A => X"ffffff90ffffffffffffffbeffffffffffffffc0ffffffff0000005100000000",
            INIT_0B => X"0000002e00000000ffffff18fffffffffffffffaffffffffffffffd8ffffffff",
            INIT_0C => X"ffffffbbffffffff00000006000000000000001300000000ffffffdaffffffff",
            INIT_0D => X"0000000200000000ffffff7affffffffffffff95fffffffffffffe69ffffffff",
            INIT_0E => X"ffffffdcffffffff0000004100000000000000ad00000000ffffff67ffffffff",
            INIT_0F => X"000000450000000000000078000000000000003d00000000ffffffb4ffffffff",
            INIT_10 => X"000000620000000000000000000000000000006a00000000fffffff6ffffffff",
            INIT_11 => X"ffffff43ffffffff0000005600000000fffffffbffffffff0000006200000000",
            INIT_12 => X"ffffffbefffffffffffffff5ffffffff0000000b00000000ffffffbcffffffff",
            INIT_13 => X"0000002e00000000ffffff74ffffffffffffffcdfffffffffffffff4ffffffff",
            INIT_14 => X"000000ad0000000000000018000000000000004c00000000ffffff4bffffffff",
            INIT_15 => X"fffffff5fffffffffffffff8ffffffff00000007000000000000001000000000",
            INIT_16 => X"0000000500000000ffffffefffffffffffffffeefffffffffffffff3ffffffff",
            INIT_17 => X"000000200000000000000051000000000000001b000000000000001000000000",
            INIT_18 => X"fffffeedfffffffffffffed1fffffffffffffff3ffffffff0000009000000000",
            INIT_19 => X"ffffffbfffffffffffffffaaffffffffffffff9effffffffffffff8affffffff",
            INIT_1A => X"ffffffe2ffffffff0000001700000000ffffff17ffffffffffffff81ffffffff",
            INIT_1B => X"0000004800000000ffffffccffffffffffffffd2fffffffffffffffdffffffff",
            INIT_1C => X"00000004000000000000004600000000ffffff86ffffffffffffffb9ffffffff",
            INIT_1D => X"ffffffdcffffffff000000c600000000ffffff2affffffffffffffebffffffff",
            INIT_1E => X"0000003f00000000000000b100000000ffffff95ffffffffffffffb5ffffffff",
            INIT_1F => X"ffffff9fffffffff00000009000000000000005500000000ffffff3bffffffff",
            INIT_20 => X"00000039000000000000000400000000ffffffcdffffffff0000003e00000000",
            INIT_21 => X"0000006d00000000ffffff75ffffffff0000003700000000ffffffb1ffffffff",
            INIT_22 => X"0000004200000000000000ac00000000ffffff92fffffffffffffefcffffffff",
            INIT_23 => X"ffffff8bffffffffffffff47ffffffffffffffaeffffffff0000005800000000",
            INIT_24 => X"ffffff47ffffffff000000f600000000fffffea6ffffffff0000003500000000",
            INIT_25 => X"0000006a000000000000005600000000fffffffcffffffffffffffa2ffffffff",
            INIT_26 => X"ffffff68ffffffffffffff84ffffffff0000000b00000000000000c800000000",
            INIT_27 => X"ffffff90ffffffff0000001100000000ffffff16ffffffff0000002600000000",
            INIT_28 => X"0000009d000000000000003700000000ffffffc9ffffffff0000006400000000",
            INIT_29 => X"ffffffbdffffffff0000011200000000ffffff91ffffffff000000c500000000",
            INIT_2A => X"0000004400000000000000410000000000000080000000000000000900000000",
            INIT_2B => X"00000032000000000000002a00000000fffffffaffffffffffffff75ffffffff",
            INIT_2C => X"0000003400000000000000380000000000000045000000000000005500000000",
            INIT_2D => X"ffffffc6ffffffffffffff66ffffffffffffffd9ffffffffffffffd4ffffffff",
            INIT_2E => X"ffffff6cffffffffffffffc8ffffffffffffff99ffffffff0000008600000000",
            INIT_2F => X"00000045000000000000005b00000000ffffffe3ffffffff000000c800000000",
            INIT_30 => X"0000005f00000000ffffff80ffffffff00000074000000000000004f00000000",
            INIT_31 => X"ffffff7affffffffffffffd1ffffffffffffff7bffffffff0000005f00000000",
            INIT_32 => X"fffffff4ffffffff0000005c00000000ffffff44ffffffffffffff50ffffffff",
            INIT_33 => X"00000044000000000000001b0000000000000077000000000000004300000000",
            INIT_34 => X"0000008800000000ffffffadffffffff00000014000000000000003900000000",
            INIT_35 => X"00000069000000000000003b000000000000002000000000ffffffc1ffffffff",
            INIT_36 => X"0000000700000000ffffffc8fffffffffffffffeffffffffffffffaeffffffff",
            INIT_37 => X"ffffffedffffffffffffff7cffffffff000000bd000000000000004600000000",
            INIT_38 => X"0000000700000000ffffffc0ffffffffffffff07ffffffffffffff6effffffff",
            INIT_39 => X"0000004d00000000ffffffc0ffffffff0000007a000000000000005700000000",
            INIT_3A => X"00000021000000000000002a00000000fffffef3ffffffffffffff80ffffffff",
            INIT_3B => X"000000e100000000ffffff66ffffffff0000004000000000ffffff63ffffffff",
            INIT_3C => X"0000000c00000000ffffffb5ffffffff00000028000000000000001000000000",
            INIT_3D => X"ffffffe4fffffffffffffff9fffffffffffffffbffffffff0000001c00000000",
            INIT_3E => X"ffffffdeffffffff000000e200000000ffffffcfffffffffffffffb8ffffffff",
            INIT_3F => X"0000005600000000ffffffbaffffffffffffffbfffffffff0000009100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff2ffffffffffffff9dffffffffffffff38ffffffffffffffe5ffffffff",
            INIT_41 => X"ffffffe1ffffffff0000004800000000000000ae000000000000005a00000000",
            INIT_42 => X"0000010200000000fffffe79ffffffffffffff0affffffff0000006100000000",
            INIT_43 => X"ffffff76fffffffffffffe36fffffffffffffff9ffffffff0000005300000000",
            INIT_44 => X"0000009200000000ffffffc3ffffffff0000010b000000000000008b00000000",
            INIT_45 => X"ffffffc3ffffffff000000340000000000000008000000000000003700000000",
            INIT_46 => X"ffffff24ffffffff0000005c00000000000000fe00000000ffffff66ffffffff",
            INIT_47 => X"0000008500000000ffffffbfffffffff0000005d00000000ffffff39ffffffff",
            INIT_48 => X"00000070000000000000002e000000000000006400000000ffffffd0ffffffff",
            INIT_49 => X"ffffff54ffffffff0000000200000000ffffff61ffffffff0000004b00000000",
            INIT_4A => X"ffffff67fffffffffffffef3fffffffffffffe64ffffffff0000009200000000",
            INIT_4B => X"ffffffdcffffffff000000ba00000000ffffff90ffffffff0000004600000000",
            INIT_4C => X"ffffffedffffffffffffff83ffffffffffffffc3ffffffffffffffe4ffffffff",
            INIT_4D => X"ffffff99fffffffffffffff7ffffffffffffffedfffffffffffffff1ffffffff",
            INIT_4E => X"fffffe36ffffffffffffffadffffffffffffffc7fffffffffffffe5cffffffff",
            INIT_4F => X"ffffff91ffffffff0000005400000000ffffffb8ffffffffffffffe8ffffffff",
            INIT_50 => X"0000005100000000ffffff89ffffffff0000003300000000ffffffeeffffffff",
            INIT_51 => X"0000008b000000000000004000000000fffffffcffffffffffffff8affffffff",
            INIT_52 => X"ffffffb3ffffffffffffffe2ffffffffffffffa2ffffffffffffffd4ffffffff",
            INIT_53 => X"00000084000000000000005200000000fffffef8ffffffffffffff5fffffffff",
            INIT_54 => X"ffffffc4ffffffff0000002a0000000000000063000000000000000100000000",
            INIT_55 => X"ffffffc7ffffffff000000180000000000000057000000000000005300000000",
            INIT_56 => X"0000006c0000000000000011000000000000004b00000000ffffffa6ffffffff",
            INIT_57 => X"fffffeb4ffffffffffffffb2ffffffffffffffc0ffffffffffffff05ffffffff",
            INIT_58 => X"0000000b000000000000000800000000ffffff1fffffffffffffffb6ffffffff",
            INIT_59 => X"000000170000000000000082000000000000000f000000000000005000000000",
            INIT_5A => X"ffffff37ffffffff0000000d000000000000000a00000000fffffff9ffffffff",
            INIT_5B => X"0000008c00000000ffffff97ffffffff00000026000000000000006b00000000",
            INIT_5C => X"0000006000000000ffffff6effffffffffffffc6ffffffffffffff96ffffffff",
            INIT_5D => X"ffffffffffffffff0000000000000000fffffffcffffffffffffff86ffffffff",
            INIT_5E => X"0000000b000000000000000100000000fffffff2fffffffffffffff8ffffffff",
            INIT_5F => X"0000004c00000000ffffff8efffffffffffffff7fffffffffffffff6ffffffff",
            INIT_60 => X"00000046000000000000005500000000ffffffbfffffffffffffff6cffffffff",
            INIT_61 => X"0000008200000000fffffff3ffffffff0000004f000000000000003d00000000",
            INIT_62 => X"ffffff73ffffffffffffff97ffffffff0000008900000000ffffff7bffffffff",
            INIT_63 => X"00000096000000000000001400000000ffffff5dffffffff0000004600000000",
            INIT_64 => X"ffffffbbffffffffffffffdfffffffff0000003000000000ffffffeaffffffff",
            INIT_65 => X"0000010d00000000ffffffadffffffffffffffeafffffffffffffe97ffffffff",
            INIT_66 => X"0000006f0000000000000058000000000000005300000000fffffff7ffffffff",
            INIT_67 => X"0000002500000000fffffff7ffffffffffffffcfffffffff0000002400000000",
            INIT_68 => X"fffffe8cffffffffffffff5dffffffff000000ba000000000000004c00000000",
            INIT_69 => X"00000069000000000000001800000000fffffffdffffffff0000007500000000",
            INIT_6A => X"00000072000000000000001a00000000ffffffbfffffffff000000b600000000",
            INIT_6B => X"0000004700000000000000c700000000ffffff9bffffffffffffffbfffffffff",
            INIT_6C => X"0000003200000000ffffff49ffffffff00000028000000000000000700000000",
            INIT_6D => X"0000001e00000000ffffffdfffffffff000000f100000000ffffffc6ffffffff",
            INIT_6E => X"0000004200000000ffffff9cffffffff0000005700000000fffffedfffffffff",
            INIT_6F => X"ffffffdbffffffff0000002f000000000000003300000000ffffff6bffffffff",
            INIT_70 => X"00000003000000000000001a000000000000002900000000ffffff76ffffffff",
            INIT_71 => X"ffffff58ffffffff00000097000000000000008500000000ffffff79ffffffff",
            INIT_72 => X"000000df00000000ffffff9fffffffff0000009e00000000ffffffdfffffffff",
            INIT_73 => X"ffffff55ffffffff0000003500000000fffffe69ffffffff0000009300000000",
            INIT_74 => X"0000000800000000ffffff54ffffffffffffff32ffffffff0000000600000000",
            INIT_75 => X"fffffffdffffffffffffffc2ffffffffffffff2cffffffff0000001700000000",
            INIT_76 => X"0000002d000000000000008500000000ffffffd3ffffffff0000001900000000",
            INIT_77 => X"0000004c000000000000008f00000000ffffffb8ffffffffffffffc1ffffffff",
            INIT_78 => X"000000d10000000000000014000000000000001b00000000fffffefcffffffff",
            INIT_79 => X"000000450000000000000014000000000000000600000000ffffffbeffffffff",
            INIT_7A => X"ffffffc3ffffffff000000c300000000fffffe98ffffffffffffffccffffffff",
            INIT_7B => X"000000c1000000000000005400000000ffffff2bffffffff0000002600000000",
            INIT_7C => X"ffffffb7ffffffff0000001f00000000ffffffbcffffffffffffff6bffffffff",
            INIT_7D => X"fffffecdfffffffffffffff4ffffffff00000011000000000000000f00000000",
            INIT_7E => X"0000003b00000000ffffff9dffffffff00000043000000000000002100000000",
            INIT_7F => X"0000004e00000000ffffff38ffffffffffffffa7ffffffffffffffe9ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE21;


    MEM_IWGHT_LAYER2_INSTANCE22 : if BRAM_NAME = "iwght_layer2_instance22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000006300000000000000c0000000000000007700000000ffffffe4ffffffff",
            INIT_01 => X"ffffffa8ffffffffffffffdffffffffffffffef4ffffffffffffffd0ffffffff",
            INIT_02 => X"0000005e00000000ffffffb4ffffffff0000002d000000000000003c00000000",
            INIT_03 => X"0000006200000000000000b3000000000000003e00000000ffffffdcffffffff",
            INIT_04 => X"ffffffa2fffffffffffffee6fffffffffffffff9ffffffff0000002300000000",
            INIT_05 => X"0000005300000000ffffff1cffffffff00000079000000000000000400000000",
            INIT_06 => X"000000b3000000000000002d000000000000007700000000fffffee6ffffffff",
            INIT_07 => X"ffffff9affffffffffffffddffffffffffffff97ffffffff0000001e00000000",
            INIT_08 => X"fffffffaffffffff0000001300000000ffffff21ffffffff0000000900000000",
            INIT_09 => X"0000004700000000ffffffdeffffffff00000024000000000000002800000000",
            INIT_0A => X"ffffff6cffffffff00000056000000000000000a000000000000000600000000",
            INIT_0B => X"ffffff7bffffffff000000be00000000ffffffb1ffffffff0000003f00000000",
            INIT_0C => X"ffffffcfffffffffffffff90ffffffff000000ad00000000000000a000000000",
            INIT_0D => X"ffffff9fffffffffffffffdcffffffff0000000a00000000ffffffffffffffff",
            INIT_0E => X"ffffffcfffffffffffffff85ffffffff00000003000000000000011f00000000",
            INIT_0F => X"ffffffdbffffffffffffffb3ffffffff0000000900000000ffffffd2ffffffff",
            INIT_10 => X"ffffffa7ffffffff0000007200000000ffffffb6ffffffff0000004200000000",
            INIT_11 => X"ffffffc3fffffffffffffffcffffffffffffffbaffffffffffffffd9ffffffff",
            INIT_12 => X"ffffffbbffffffff00000034000000000000000e00000000ffffffdeffffffff",
            INIT_13 => X"00000007000000000000002200000000fffffedaffffffffffffffc3ffffffff",
            INIT_14 => X"00000074000000000000007400000000ffffffe6ffffffffffffff71ffffffff",
            INIT_15 => X"ffffffccffffffff0000005600000000fffffeb5ffffffffffffff28ffffffff",
            INIT_16 => X"0000003400000000ffffff08ffffffffffffffc9ffffffff0000006400000000",
            INIT_17 => X"ffffffa9ffffffff0000004100000000ffffff62ffffffffffffff4bffffffff",
            INIT_18 => X"ffffffcdffffffff0000006200000000ffffffefffffffffffffff11ffffffff",
            INIT_19 => X"ffffffcdffffffff000000d7000000000000008800000000ffffff6dffffffff",
            INIT_1A => X"fffffff3ffffffffffffffa7ffffffffffffffc8ffffffffffffff99ffffffff",
            INIT_1B => X"000000130000000000000043000000000000003600000000ffffff7dffffffff",
            INIT_1C => X"ffffffc0ffffffff000000bf0000000000000080000000000000009c00000000",
            INIT_1D => X"0000005e00000000ffffffbaffffffffffffffbcfffffffffffffff2ffffffff",
            INIT_1E => X"ffffffecffffffff0000003d00000000ffffffd8ffffffffffffffa8ffffffff",
            INIT_1F => X"00000021000000000000005d0000000000000036000000000000003e00000000",
            INIT_20 => X"ffffffb4ffffffffffffff78ffffffff00000050000000000000005c00000000",
            INIT_21 => X"0000007500000000ffffffd4fffffffffffffef2fffffffffffffecbffffffff",
            INIT_22 => X"00000043000000000000007b00000000000000dd00000000000000b300000000",
            INIT_23 => X"0000007e00000000ffffffd6ffffffffffffff8effffffffffffffd8ffffffff",
            INIT_24 => X"0000003a0000000000000094000000000000002f000000000000002d00000000",
            INIT_25 => X"ffffffebfffffffffffffffdffffffffffffffefffffffff0000002300000000",
            INIT_26 => X"0000002000000000fffffff3ffffffffffffffecffffffff0000000c00000000",
            INIT_27 => X"00000036000000000000003700000000ffffffedfffffffffffffff2ffffffff",
            INIT_28 => X"0000002e00000000ffffffc6ffffffff0000005e00000000ffffffd0ffffffff",
            INIT_29 => X"0000000c000000000000004b000000000000005500000000ffffffe3ffffffff",
            INIT_2A => X"0000006800000000ffffffc1ffffffffffffff06ffffffffffffff8bffffffff",
            INIT_2B => X"0000009a00000000000000d600000000000000a500000000ffffffefffffffff",
            INIT_2C => X"0000003900000000ffffff6affffffffffffffceffffffffffffff92ffffffff",
            INIT_2D => X"ffffff42ffffffffffffffa7ffffffffffffff6effffffffffffffd3ffffffff",
            INIT_2E => X"ffffffa2ffffffff0000000800000000ffffffdaffffffffffffffc1ffffffff",
            INIT_2F => X"ffffffaafffffffffffffff5ffffffff0000002b00000000ffffff8affffffff",
            INIT_30 => X"0000004e00000000ffffffc1ffffffff00000119000000000000007500000000",
            INIT_31 => X"fffffec8ffffffffffffffabfffffffffffffeeeffffffffffffffcbffffffff",
            INIT_32 => X"0000003c00000000ffffff26ffffffff0000007b00000000ffffff94ffffffff",
            INIT_33 => X"0000007500000000ffffffdeffffffff0000001000000000ffffffa8ffffffff",
            INIT_34 => X"0000003000000000000000ae000000000000002f00000000ffffffecffffffff",
            INIT_35 => X"ffffffaeffffffffffffff4effffffff00000034000000000000003900000000",
            INIT_36 => X"ffffffd0ffffffff0000002200000000ffffff82ffffffff0000001a00000000",
            INIT_37 => X"0000008700000000000000130000000000000024000000000000000500000000",
            INIT_38 => X"ffffffa1ffffffff00000036000000000000006800000000ffffffb8ffffffff",
            INIT_39 => X"000000d3000000000000000a00000000ffffffbffffffffffffffed2ffffffff",
            INIT_3A => X"000000e800000000ffffffdcffffffffffffffb5ffffffff000000bb00000000",
            INIT_3B => X"ffffffcdfffffffffffffefeffffffff0000006700000000ffffff7affffffff",
            INIT_3C => X"fffffffcffffffffffffff24ffffffff0000001100000000ffffffdfffffffff",
            INIT_3D => X"ffffffffffffffff00000005000000000000007400000000ffffffa5ffffffff",
            INIT_3E => X"0000002900000000ffffff91ffffffffffffff2effffffff0000003d00000000",
            INIT_3F => X"0000001000000000ffffff8effffffffffffffa4ffffffff0000001d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffff5effffffff00000021000000000000010f000000000000006100000000",
            INIT_41 => X"fffffed8fffffffffffffce0ffffffff0000003800000000ffffffccffffffff",
            INIT_42 => X"fffffea5ffffffff0000001500000000ffffffaaffffffff000000b400000000",
            INIT_43 => X"ffffff3dffffffff0000003c00000000ffffffa6ffffffffffffff66ffffffff",
            INIT_44 => X"0000001a00000000ffffffd1ffffffffffffff6bffffffff0000001300000000",
            INIT_45 => X"ffffff2effffffff00000065000000000000000e00000000ffffffb9ffffffff",
            INIT_46 => X"ffffffd8ffffffffffffffcbfffffffffffffff8ffffffffffffffafffffffff",
            INIT_47 => X"ffffffe8ffffffff000000e1000000000000004000000000ffffffebffffffff",
            INIT_48 => X"ffffffb0ffffffff0000000e000000000000006c000000000000001300000000",
            INIT_49 => X"ffffffa5ffffffffffffff60ffffffff0000004500000000ffffff8cffffffff",
            INIT_4A => X"0000002d00000000ffffffc8ffffffffffffff9fffffffff0000003100000000",
            INIT_4B => X"ffffff31ffffffffffffffeeffffffff000000ba000000000000004400000000",
            INIT_4C => X"ffffffbaffffffff000000290000000000000011000000000000005500000000",
            INIT_4D => X"ffffffc7ffffffffffffff93ffffffffffffffb9ffffffff0000001600000000",
            INIT_4E => X"ffffff56ffffffffffffffcfffffffff000000d4000000000000009000000000",
            INIT_4F => X"ffffff6fffffffff0000008c00000000fffffff8ffffffffffffff4bffffffff",
            INIT_50 => X"0000005e00000000ffffffa0ffffffffffffffbcffffffff0000003600000000",
            INIT_51 => X"ffffff9fffffffff0000008b00000000ffffffa3ffffffffffffff72ffffffff",
            INIT_52 => X"ffffffb2ffffffffffffffddffffffff0000007e00000000fffffff7ffffffff",
            INIT_53 => X"0000006500000000ffffffd0ffffffffffffff0cffffffff0000006e00000000",
            INIT_54 => X"ffffff7dffffffff00000049000000000000007a00000000ffffff51ffffffff",
            INIT_55 => X"fffffff8fffffffffffffff9ffffffff00000036000000000000010300000000",
            INIT_56 => X"ffffffbaffffffffffffffc9ffffffffffffff8fffffffffffffff55ffffffff",
            INIT_57 => X"0000001200000000ffffff65fffffffffffffee1ffffffff0000002d00000000",
            INIT_58 => X"ffffffdfffffffff0000001800000000ffffff97ffffffffffffffe8ffffffff",
            INIT_59 => X"ffffff28ffffffffffffff99ffffffffffffffceffffffffffffff88ffffffff",
            INIT_5A => X"ffffffd8ffffffffffffff84ffffffff0000004f00000000fffffef3ffffffff",
            INIT_5B => X"ffffffbbffffffff00000003000000000000007d00000000ffffff78ffffffff",
            INIT_5C => X"0000000300000000ffffff9fffffffffffffffc6ffffffff0000003100000000",
            INIT_5D => X"fffffff7ffffffff0000004100000000ffffffaeffffffff0000001900000000",
            INIT_5E => X"0000003400000000ffffffd9ffffffff0000003c00000000ffffff85ffffffff",
            INIT_5F => X"ffffffd3ffffffff0000001a00000000ffffffdeffffffff0000004800000000",
            INIT_60 => X"ffffffe2ffffffffffffff32ffffffffffffffc7ffffffffffffffb0ffffffff",
            INIT_61 => X"00000054000000000000004a00000000ffffff83ffffffffffffffdfffffffff",
            INIT_62 => X"0000001a00000000ffffffe1ffffffff0000002b000000000000001d00000000",
            INIT_63 => X"0000001d000000000000003500000000fffffff0ffffffffffffffcbffffffff",
            INIT_64 => X"fffffff7ffffffffffffff3fffffffff0000001b000000000000007500000000",
            INIT_65 => X"ffffffcdfffffffffffffee6fffffffffffffed9ffffffffffffffbfffffffff",
            INIT_66 => X"00000000000000000000007b00000000ffffff31ffffffffffffffccffffffff",
            INIT_67 => X"ffffffa4ffffffff00000038000000000000001e00000000ffffffc2ffffffff",
            INIT_68 => X"fffffff8ffffffff0000000000000000ffffffaeffffffffffffffc6ffffffff",
            INIT_69 => X"0000008400000000000000060000000000000014000000000000007200000000",
            INIT_6A => X"0000008000000000ffffffbeffffffff0000006f00000000000000ca00000000",
            INIT_6B => X"fffffe94fffffffffffffffbffffffffffffffd9ffffffffffffffefffffffff",
            INIT_6C => X"ffffffa8ffffffffffffff52ffffffffffffff3affffffffffffff64ffffffff",
            INIT_6D => X"0000000000000000fffffffdffffffff00000008000000000000002700000000",
            INIT_6E => X"fffffff8ffffffff0000000b00000000ffffffecfffffffffffffffbffffffff",
            INIT_6F => X"ffffff88ffffffff0000002e00000000ffffffedffffffff0000000700000000",
            INIT_70 => X"ffffffe8ffffffffffffff6dffffffff0000004d000000000000004100000000",
            INIT_71 => X"ffffffa3ffffffffffffff9effffffff00000035000000000000002900000000",
            INIT_72 => X"ffffffcaffffffffffffffcaffffffffffffffc4ffffffff0000003d00000000",
            INIT_73 => X"ffffff54ffffffffffffff39ffffffff00000021000000000000009000000000",
            INIT_74 => X"ffffff5bffffffff00000001000000000000003400000000ffffff9dffffffff",
            INIT_75 => X"ffffff87ffffffffffffff64ffffffff0000003700000000ffffffb8ffffffff",
            INIT_76 => X"0000002f00000000ffffff3effffffffffffff7effffffffffffff78ffffffff",
            INIT_77 => X"ffffffceffffffff0000004400000000fffffea5ffffffff0000002100000000",
            INIT_78 => X"0000007600000000ffffffeaffffffff0000006700000000fffffe9bffffffff",
            INIT_79 => X"ffffff12fffffffffffffff9ffffffffffffff4cffffffffffffff48ffffffff",
            INIT_7A => X"00000062000000000000003500000000fffffff0ffffffffffffff92ffffffff",
            INIT_7B => X"0000000c000000000000000500000000ffffff56ffffffffffffffcbffffffff",
            INIT_7C => X"0000001400000000ffffff5effffffffffffff8bffffffff0000004100000000",
            INIT_7D => X"ffffff96ffffffffffffffd0ffffffff00000069000000000000003e00000000",
            INIT_7E => X"0000001300000000ffffffc9ffffffff0000005d00000000ffffffb5ffffffff",
            INIT_7F => X"0000003700000000000000680000000000000038000000000000003400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE22;


    MEM_IWGHT_LAYER2_INSTANCE23 : if BRAM_NAME = "iwght_layer2_instance23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffa2ffffffff0000011800000000ffffffbcffffffffffffffc4ffffffff",
            INIT_01 => X"ffffff54ffffffffffffffbcffffffff0000002600000000ffffffcaffffffff",
            INIT_02 => X"000000610000000000000011000000000000003f00000000ffffff8fffffffff",
            INIT_03 => X"fffffff8ffffffffffffff9bffffffff0000000e000000000000000c00000000",
            INIT_04 => X"0000006000000000ffffffb5fffffffffffffff2ffffffffffffffc8ffffffff",
            INIT_05 => X"0000004b00000000000000b5000000000000005300000000ffffffedffffffff",
            INIT_06 => X"ffffff5affffffffffffffc4ffffffffffffffc2ffffffffffffffadffffffff",
            INIT_07 => X"00000066000000000000001c000000000000003b000000000000009400000000",
            INIT_08 => X"ffffffa7ffffffff000000220000000000000021000000000000008300000000",
            INIT_09 => X"0000008b00000000ffffffb5ffffffff0000000900000000ffffff0affffffff",
            INIT_0A => X"0000002c000000000000001e000000000000002f00000000ffffffacffffffff",
            INIT_0B => X"ffffff89ffffffff0000000500000000ffffffd2ffffffffffffffd4ffffffff",
            INIT_0C => X"ffffffd9ffffffff00000048000000000000008a000000000000006b00000000",
            INIT_0D => X"ffffff0effffffffffffffe7fffffffffffffff5fffffffffffffff0ffffffff",
            INIT_0E => X"ffffff46ffffffffffffff6bffffffff0000001800000000ffffffceffffffff",
            INIT_0F => X"ffffff82ffffffff0000001800000000fffffffdffffffffffffff76ffffffff",
            INIT_10 => X"ffffffaeffffffff00000022000000000000004b000000000000000d00000000",
            INIT_11 => X"fffffff6ffffffff00000006000000000000000a000000000000003900000000",
            INIT_12 => X"0000001a000000000000000100000000ffffffc0ffffffffffffff92ffffffff",
            INIT_13 => X"0000000b00000000ffffffafffffffffffffffcaffffffff0000004200000000",
            INIT_14 => X"fffffff8ffffffff0000001000000000ffffffb9ffffffffffffff77ffffffff",
            INIT_15 => X"ffffff5fffffffff0000002500000000ffffffb7ffffffff0000001d00000000",
            INIT_16 => X"0000008f00000000ffffff74ffffffffffffffb6ffffffff0000000900000000",
            INIT_17 => X"000000bf000000000000007b000000000000003a00000000ffffffc3ffffffff",
            INIT_18 => X"0000002100000000ffffffcaffffffffffffff75ffffffff0000004900000000",
            INIT_19 => X"ffffffe7ffffffff0000004900000000ffffffa8ffffffff0000009a00000000",
            INIT_1A => X"ffffffb7ffffffffffffffbfffffffffffffff63ffffffff0000001f00000000",
            INIT_1B => X"ffffffd7ffffffffffffffe9ffffffffffffff20ffffffffffffff8fffffffff",
            INIT_1C => X"ffffffe1ffffffff0000001900000000ffffffe7ffffffffffffffb7ffffffff",
            INIT_1D => X"ffffff28ffffffff0000005b00000000000000ae00000000ffffffacffffffff",
            INIT_1E => X"0000007700000000ffffff40ffffffff0000008e000000000000003600000000",
            INIT_1F => X"0000008e00000000fffffffeffffffff0000002d00000000ffffff80ffffffff",
            INIT_20 => X"ffffff62ffffffffffffffb3ffffffffffffff6ffffffffffffffff7ffffffff",
            INIT_21 => X"00000005000000000000005300000000000000ad00000000ffffff7affffffff",
            INIT_22 => X"fffffff3ffffffffffffff77ffffffff00000060000000000000007e00000000",
            INIT_23 => X"000000220000000000000023000000000000006900000000ffffff9bffffffff",
            INIT_24 => X"fffffffeffffffff000000d80000000000000041000000000000006600000000",
            INIT_25 => X"0000005500000000ffffffbcffffffff00000083000000000000002a00000000",
            INIT_26 => X"000000ab00000000ffffff83ffffffffffffffd4ffffffff0000005c00000000",
            INIT_27 => X"ffffff7bffffffff0000002100000000ffffffedffffffffffffff74ffffffff",
            INIT_28 => X"ffffff6fffffffffffffff43ffffffffffffffc5ffffffffffffff9bffffffff",
            INIT_29 => X"0000006f00000000ffffffc9fffffffffffffef3ffffffff0000001100000000",
            INIT_2A => X"00000036000000000000001b00000000ffffffefffffffff0000003f00000000",
            INIT_2B => X"0000007400000000ffffff9cfffffffffffffff2ffffffff0000001900000000",
            INIT_2C => X"0000000a00000000000000bd000000000000007a00000000ffffffa8ffffffff",
            INIT_2D => X"fffffec8ffffffff000000c500000000ffffff4bffffffffffffffebffffffff",
            INIT_2E => X"ffffff46fffffffffffffff1ffffffffffffffa1ffffffffffffffd2ffffffff",
            INIT_2F => X"ffffffa2ffffffff0000004300000000000000b600000000000000aa00000000",
            INIT_30 => X"fffffffeffffffff0000005200000000ffffffabffffffff0000008100000000",
            INIT_31 => X"ffffff49ffffffff000000ae00000000ffffffa8ffffffff000000bf00000000",
            INIT_32 => X"ffffffe5ffffffff0000004700000000ffffffcbffffffffffffffa4ffffffff",
            INIT_33 => X"0000009500000000ffffffb0ffffffffffffff7effffffff0000009500000000",
            INIT_34 => X"00000045000000000000001900000000000000c600000000000000b300000000",
            INIT_35 => X"0000000d00000000fffffff8ffffffff00000017000000000000010000000000",
            INIT_36 => X"fffffff0fffffffffffffffcfffffffffffffff4ffffffffffffffe4ffffffff",
            INIT_37 => X"ffffffbcffffffffffffff8cfffffffffffffff7ffffffff0000001000000000",
            INIT_38 => X"0000001f00000000ffffffadfffffffffffffffefffffffffffffff8ffffffff",
            INIT_39 => X"0000000000000000fffffff8ffffffffffffffddffffffffffffffb0ffffffff",
            INIT_3A => X"fffffff9ffffffff000000c800000000ffffff80ffffffffffffffd5ffffffff",
            INIT_3B => X"0000002700000000ffffffc5ffffffff0000006100000000ffffff59ffffffff",
            INIT_3C => X"ffffffbbffffffffffffffecffffffff00000074000000000000002700000000",
            INIT_3D => X"00000038000000000000001d000000000000009500000000ffffff32ffffffff",
            INIT_3E => X"00000041000000000000008900000000000000b9000000000000001100000000",
            INIT_3F => X"fffffe01ffffffff0000005300000000ffffff79ffffffff0000000800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffff3bffffffffffffffcdffffffff0000010000000000ffffffebffffffff",
            INIT_41 => X"ffffff2bffffffff00000012000000000000001c000000000000005f00000000",
            INIT_42 => X"ffffffa9ffffffffffffffb2ffffffff00000003000000000000007100000000",
            INIT_43 => X"ffffffa0ffffffff0000008800000000ffffffb1ffffffff0000003900000000",
            INIT_44 => X"ffffffc7ffffffff0000002000000000ffffffd2ffffffff0000001900000000",
            INIT_45 => X"0000008e000000000000000300000000ffffff4effffffff0000001000000000",
            INIT_46 => X"ffffffb3ffffffff0000002e000000000000000a00000000ffffff88ffffffff",
            INIT_47 => X"0000009500000000ffffffa4ffffffff0000001b00000000ffffff83ffffffff",
            INIT_48 => X"0000001b00000000ffffffe5ffffffff0000003900000000ffffff7bffffffff",
            INIT_49 => X"ffffff6fffffffffffffffafffffffffffffffbafffffffffffffef0ffffffff",
            INIT_4A => X"00000013000000000000003f00000000ffffffb5ffffffff0000007700000000",
            INIT_4B => X"0000001b00000000ffffff9fffffffffffffffd5ffffffffffffff94ffffffff",
            INIT_4C => X"ffffff9cffffffffffffffb8ffffffff00000079000000000000001a00000000",
            INIT_4D => X"000000b100000000ffffff21ffffffffffffff4bffffffff0000003100000000",
            INIT_4E => X"ffffff7affffffff000000030000000000000022000000000000003000000000",
            INIT_4F => X"0000004b000000000000003e00000000ffffffa7ffffffff0000010000000000",
            INIT_50 => X"ffffffb5ffffffff0000000d00000000ffffff69ffffffffffffffe8ffffffff",
            INIT_51 => X"ffffffd9ffffffff0000001800000000000000b6000000000000003500000000",
            INIT_52 => X"ffffffffffffffff00000034000000000000007a000000000000001700000000",
            INIT_53 => X"00000000000000000000002300000000fffffff8ffffffffffffffd7ffffffff",
            INIT_54 => X"ffffffa8ffffffff0000006100000000ffffffc2ffffffffffffffd2ffffffff",
            INIT_55 => X"0000000000000000ffffff2effffffff0000008e000000000000003500000000",
            INIT_56 => X"0000000c000000000000008d00000000ffffff75ffffffff000000a900000000",
            INIT_57 => X"0000004000000000ffffffd5ffffffffffffffd0ffffffff0000008500000000",
            INIT_58 => X"000000fe00000000ffffff9affffffffffffffb9fffffffffffffff5ffffffff",
            INIT_59 => X"0000006a000000000000000000000000ffffff9effffffffffffffceffffffff",
            INIT_5A => X"00000097000000000000000f00000000ffffff71ffffffffffffffe4ffffffff",
            INIT_5B => X"ffffff84ffffffff00000046000000000000000b000000000000005b00000000",
            INIT_5C => X"00000084000000000000009e00000000ffffff04ffffffffffffffd1ffffffff",
            INIT_5D => X"ffffffc9ffffffffffffffaaffffffff000000b300000000ffffff61ffffffff",
            INIT_5E => X"ffffff87ffffffff0000009d00000000ffffff7cffffffffffffffbaffffffff",
            INIT_5F => X"ffffffc4ffffffff00000018000000000000004600000000ffffffe6ffffffff",
            INIT_60 => X"0000005600000000ffffffc9ffffffffffffffe6ffffffffffffff8effffffff",
            INIT_61 => X"0000002d000000000000001b00000000ffffff0bffffffffffffff48ffffffff",
            INIT_62 => X"fffffff4ffffffff0000007e00000000ffffffbfffffffff0000003d00000000",
            INIT_63 => X"00000080000000000000002900000000ffffff1dffffffffffffffd5ffffffff",
            INIT_64 => X"fffffff9fffffffffffffff5fffffffffffffed1ffffffffffffff53ffffffff",
            INIT_65 => X"00000047000000000000003300000000ffffffc4ffffffffffffffe9ffffffff",
            INIT_66 => X"ffffffb7ffffffffffffffa7ffffffff000000cb00000000ffffff96ffffffff",
            INIT_67 => X"ffffffadffffffff0000000200000000000000ca00000000000000fa00000000",
            INIT_68 => X"ffffff1dffffffff0000001f00000000ffffff57ffffffff0000002e00000000",
            INIT_69 => X"ffffffdbffffffff0000008900000000ffffffe2ffffffffffffffb9ffffffff",
            INIT_6A => X"00000081000000000000002a00000000ffffffc3ffffffff0000001a00000000",
            INIT_6B => X"ffffffb7ffffffffffffffbfffffffff00000022000000000000004b00000000",
            INIT_6C => X"ffffffd2ffffffffffffff39ffffffffffffff8affffffff0000003000000000",
            INIT_6D => X"fffffff1ffffffff000000b200000000ffffff75ffffffffffffffc0ffffffff",
            INIT_6E => X"fffffff7fffffffffffffea5ffffffff000000cd00000000fffffef9ffffffff",
            INIT_6F => X"0000003800000000ffffff44ffffffffffffffeeffffffffffffff73ffffffff",
            INIT_70 => X"ffffffedffffffff0000005400000000fffffffaffffffff0000008400000000",
            INIT_71 => X"ffffff66ffffffff00000031000000000000009a00000000ffffffe5ffffffff",
            INIT_72 => X"0000003300000000ffffff86ffffffff0000000d000000000000002200000000",
            INIT_73 => X"ffffff4effffffffffffffd0ffffffffffffffc8fffffffffffffe93ffffffff",
            INIT_74 => X"0000002400000000ffffffc6ffffffff0000002700000000ffffffa7ffffffff",
            INIT_75 => X"0000005f00000000ffffff78ffffffff0000004600000000ffffffefffffffff",
            INIT_76 => X"0000000d00000000ffffffadffffffff000000d3000000000000005300000000",
            INIT_77 => X"ffffff20ffffffffffffff26ffffffff0000005b00000000ffffffd4ffffffff",
            INIT_78 => X"0000000e00000000ffffffbbffffffffffffffc3ffffffff0000006300000000",
            INIT_79 => X"fffffffcffffffff00000046000000000000007e00000000ffffffe0ffffffff",
            INIT_7A => X"0000002f0000000000000061000000000000001200000000000000c800000000",
            INIT_7B => X"ffffffdfffffffffffffffa3ffffffff0000005900000000ffffff8affffffff",
            INIT_7C => X"000000bd000000000000000500000000000000b6000000000000002700000000",
            INIT_7D => X"0000000300000000fffffff9fffffffffffffff9ffffffff0000007300000000",
            INIT_7E => X"00000018000000000000001300000000fffffffcffffffff0000000100000000",
            INIT_7F => X"ffffffdcffffffff0000003f00000000fffffff0ffffffff0000000200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE23;


    MEM_IWGHT_LAYER2_INSTANCE24 : if BRAM_NAME = "iwght_layer2_instance24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffd4ffffffff0000001e0000000000000062000000000000007d00000000",
            INIT_01 => X"ffffff25ffffffff0000001b0000000000000004000000000000003200000000",
            INIT_02 => X"0000001a00000000ffffffa9fffffffffffffff9ffffffffffffffb3ffffffff",
            INIT_03 => X"00000094000000000000002300000000ffffff6fffffffff0000003800000000",
            INIT_04 => X"00000007000000000000009a00000000000000cb000000000000002d00000000",
            INIT_05 => X"00000019000000000000000400000000ffffffe1ffffffff0000006600000000",
            INIT_06 => X"fffffff9ffffffff0000000a000000000000003a000000000000001400000000",
            INIT_07 => X"ffffffbcffffffffffffffc6ffffffff00000118000000000000000000000000",
            INIT_08 => X"0000006300000000fffffff9ffffffffffffffc5ffffffff0000002400000000",
            INIT_09 => X"ffffffaafffffffffffffffbffffffffffffffb0ffffffffffffffbbffffffff",
            INIT_0A => X"0000004000000000ffffffebffffffffffffff57ffffffffffffff8cffffffff",
            INIT_0B => X"ffffff82ffffffff0000007b00000000ffffff89ffffffff0000000c00000000",
            INIT_0C => X"ffffff7fffffffff0000000f00000000ffffff71ffffffffffffff2bffffffff",
            INIT_0D => X"000000f9000000000000009300000000ffffffbcffffffffffffff6bffffffff",
            INIT_0E => X"ffffffc1ffffffff0000003100000000ffffff2dffffffffffffff92ffffffff",
            INIT_0F => X"0000003400000000ffffff6bffffffff0000007900000000ffffff96ffffffff",
            INIT_10 => X"ffffffcaffffffff0000006d00000000ffffffb8ffffffff0000005c00000000",
            INIT_11 => X"fffffff8ffffffff00000044000000000000006a00000000000000d500000000",
            INIT_12 => X"fffffff2ffffffffffffffa6fffffffffffffff5ffffffff0000000400000000",
            INIT_13 => X"0000007000000000ffffff96ffffffff00000070000000000000003300000000",
            INIT_14 => X"000000330000000000000049000000000000005b00000000ffffff9effffffff",
            INIT_15 => X"00000071000000000000003600000000ffffff5effffffffffffffa2ffffffff",
            INIT_16 => X"00000061000000000000003d00000000fffffffbffffffffffffff56ffffffff",
            INIT_17 => X"ffffffceffffffff0000006a000000000000001b00000000ffffff67ffffffff",
            INIT_18 => X"0000001600000000fffffff7ffffffffffffff8fffffffffffffffaaffffffff",
            INIT_19 => X"ffffff55ffffffff0000007a00000000000000a800000000ffffffa9ffffffff",
            INIT_1A => X"00000061000000000000008a000000000000010500000000ffffffeaffffffff",
            INIT_1B => X"0000001a00000000ffffffe7ffffffffffffffc0ffffffff0000004500000000",
            INIT_1C => X"0000008a000000000000000e00000000ffffff81ffffffffffffff77ffffffff",
            INIT_1D => X"0000000800000000000000070000000000000038000000000000002100000000",
            INIT_1E => X"000000b100000000ffffffcaffffffff000000ab000000000000002100000000",
            INIT_1F => X"0000001800000000ffffff9affffffff00000000000000000000002e00000000",
            INIT_20 => X"ffffffbeffffffff0000001b00000000ffffffd2ffffffff0000003400000000",
            INIT_21 => X"0000000e00000000ffffff8affffffff0000005900000000ffffffd2ffffffff",
            INIT_22 => X"ffffff44ffffffff00000047000000000000001d00000000ffffff81ffffffff",
            INIT_23 => X"000000b800000000ffffffd2ffffffff000000cb00000000ffffff59ffffffff",
            INIT_24 => X"ffffffecffffffff0000000a00000000ffffffd7ffffffff0000007e00000000",
            INIT_25 => X"ffffffccffffffffffffff75ffffffffffffff94ffffffff0000000600000000",
            INIT_26 => X"ffffff84ffffffffffffffe5ffffffffffffffd9ffffffff0000000a00000000",
            INIT_27 => X"00000023000000000000009e00000000ffffff8bffffffff0000003200000000",
            INIT_28 => X"ffffff91ffffffff0000005e00000000fffffeb4ffffffff0000004500000000",
            INIT_29 => X"ffffffc4ffffffffffffffefffffffff0000003400000000fffffef4ffffffff",
            INIT_2A => X"ffffff5fffffffff0000005100000000ffffffceffffffff0000001d00000000",
            INIT_2B => X"ffffffebffffffffffffffb5ffffffffffffff74fffffffffffffff7ffffffff",
            INIT_2C => X"ffffffadffffffff0000001e000000000000003800000000ffffffe2ffffffff",
            INIT_2D => X"00000023000000000000005000000000ffffffbcffffffff0000000300000000",
            INIT_2E => X"000000b100000000ffffff31ffffffff0000011800000000ffffff91ffffffff",
            INIT_2F => X"0000000600000000ffffffa5ffffffff0000003100000000ffffffd5ffffffff",
            INIT_30 => X"fffffeebffffffffffffffcaffffffffffffffbdffffffffffffff6fffffffff",
            INIT_31 => X"ffffffd3ffffffff0000008900000000ffffffbeffffffffffffff9affffffff",
            INIT_32 => X"ffffffc3ffffffffffffffe9ffffffffffffffd1fffffffffffffd81ffffffff",
            INIT_33 => X"ffffff8effffffffffffff8cffffffff0000005200000000ffffffc3ffffffff",
            INIT_34 => X"0000007500000000ffffff36ffffffff0000004c00000000ffffffccffffffff",
            INIT_35 => X"000000a4000000000000009100000000ffffffe1ffffffff0000008300000000",
            INIT_36 => X"ffffff8affffffff000000b4000000000000002a00000000ffffff0effffffff",
            INIT_37 => X"0000003b000000000000001b000000000000001e000000000000002700000000",
            INIT_38 => X"0000008200000000000000810000000000000029000000000000005700000000",
            INIT_39 => X"0000003400000000ffffffb3ffffffffffffffdeffffffff0000009b00000000",
            INIT_3A => X"0000002800000000ffffff77ffffffff0000002100000000ffffff6affffffff",
            INIT_3B => X"ffffff9fffffffff0000003b000000000000009200000000ffffffceffffffff",
            INIT_3C => X"0000008d00000000fffffffbffffffffffffffb7ffffffff0000008500000000",
            INIT_3D => X"0000007200000000ffffff96ffffffffffffff42fffffffffffffff4ffffffff",
            INIT_3E => X"0000008700000000fffffff4ffffffffffffff37ffffffffffffffb2ffffffff",
            INIT_3F => X"ffffffccffffffffffffffe0ffffffff0000006300000000ffffffafffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffc6ffffffff0000006c00000000ffffffd4ffffffff0000005800000000",
            INIT_41 => X"0000004d0000000000000075000000000000000b00000000ffffff06ffffffff",
            INIT_42 => X"0000000c000000000000002d0000000000000044000000000000007c00000000",
            INIT_43 => X"000000570000000000000061000000000000002700000000ffffffe5ffffffff",
            INIT_44 => X"0000000a00000000ffffffa4ffffffff00000085000000000000005e00000000",
            INIT_45 => X"0000000700000000fffffff4ffffffff0000000800000000ffffff76ffffffff",
            INIT_46 => X"00000011000000000000000a00000000ffffffffffffffff0000000100000000",
            INIT_47 => X"fffffef3ffffffffffffff06fffffffffffffff8fffffffffffffffaffffffff",
            INIT_48 => X"ffffffa2ffffffffffffff72ffffffffffffff08ffffffffffffffcfffffffff",
            INIT_49 => X"0000005d000000000000007a000000000000000e000000000000003700000000",
            INIT_4A => X"0000001000000000ffffff99ffffffff0000005a000000000000001f00000000",
            INIT_4B => X"ffffff47ffffffffffffffe4fffffffffffffee7ffffffff0000009700000000",
            INIT_4C => X"fffffff3ffffffff000000070000000000000049000000000000006a00000000",
            INIT_4D => X"ffffffd0ffffffff0000006300000000ffffffe9ffffffff0000008200000000",
            INIT_4E => X"0000005100000000ffffff6cffffffff000000d200000000ffffff2effffffff",
            INIT_4F => X"fffffff1ffffffff00000025000000000000001100000000fffffffdffffffff",
            INIT_50 => X"0000000900000000ffffff5fffffffffffffffefffffffff0000003100000000",
            INIT_51 => X"ffffffc1ffffffff00000048000000000000008700000000fffffffbffffffff",
            INIT_52 => X"000000a600000000ffffffedffffffff0000003100000000ffffff0affffffff",
            INIT_53 => X"fffffee4ffffffff00000023000000000000007400000000ffffff7bffffffff",
            INIT_54 => X"0000000800000000ffffff88fffffffffffffff4ffffffff000000e000000000",
            INIT_55 => X"ffffffd0ffffffff0000004a000000000000009200000000ffffffecffffffff",
            INIT_56 => X"0000004100000000ffffff7cffffffff0000000d00000000ffffff86ffffffff",
            INIT_57 => X"0000003600000000ffffff8fffffffff0000004400000000fffffff9ffffffff",
            INIT_58 => X"0000009200000000ffffffc5fffffffffffffefaffffffff0000004b00000000",
            INIT_59 => X"0000007e0000000000000050000000000000007d00000000ffffffabffffffff",
            INIT_5A => X"0000001600000000ffffffceffffffffffffffe7ffffffffffffffa7ffffffff",
            INIT_5B => X"0000005900000000000000e80000000000000000000000000000002b00000000",
            INIT_5C => X"ffffffb4ffffffffffffffd2ffffffffffffff4affffffffffffff49ffffffff",
            INIT_5D => X"00000027000000000000002f000000000000002200000000ffffff3affffffff",
            INIT_5E => X"000000b40000000000000096000000000000001800000000ffffffc2ffffffff",
            INIT_5F => X"ffffffd9ffffffff0000005000000000ffffffc9ffffffff0000001d00000000",
            INIT_60 => X"000000bf000000000000003300000000ffffffd6ffffffffffffff38ffffffff",
            INIT_61 => X"00000026000000000000003500000000ffffffc6ffffffffffffff74ffffffff",
            INIT_62 => X"0000006f00000000ffffffdbfffffffffffffff3ffffffff0000001a00000000",
            INIT_63 => X"0000001f00000000fffffff5ffffffffffffffabffffffff0000008600000000",
            INIT_64 => X"fffffebfffffffffffffffb9ffffffff000000aa00000000ffffff89ffffffff",
            INIT_65 => X"ffffff7dffffffffffffffb5ffffffffffffff7affffffffffffff6fffffffff",
            INIT_66 => X"ffffff84ffffffffffffff52ffffffffffffffd1ffffffffffffff56ffffffff",
            INIT_67 => X"0000003e00000000ffffffebffffffffffffffb1ffffffff0000003800000000",
            INIT_68 => X"ffffff99ffffffffffffff44ffffffff00000005000000000000002100000000",
            INIT_69 => X"ffffff55ffffffff0000006b00000000ffffffd0ffffffffffffff99ffffffff",
            INIT_6A => X"ffffffc4ffffffff00000024000000000000006700000000ffffff91ffffffff",
            INIT_6B => X"ffffffc0ffffffff0000007100000000000000dd000000000000004200000000",
            INIT_6C => X"0000004800000000ffffff9dffffffff00000025000000000000006d00000000",
            INIT_6D => X"ffffff41ffffffffffffffdbffffffffffffffb6ffffffffffffffd1ffffffff",
            INIT_6E => X"0000004600000000ffffffe8ffffffff00000079000000000000000700000000",
            INIT_6F => X"fffffffaffffffff000000ac0000000000000011000000000000005600000000",
            INIT_70 => X"0000000200000000ffffffebffffffff00000060000000000000000900000000",
            INIT_71 => X"0000003000000000ffffffc2ffffffff0000002f000000000000003e00000000",
            INIT_72 => X"ffffffddffffffff000000430000000000000075000000000000006700000000",
            INIT_73 => X"0000000d000000000000004800000000ffffffa9ffffffff000000f500000000",
            INIT_74 => X"ffffffe3ffffffff0000004100000000fffffff1ffffffff0000002000000000",
            INIT_75 => X"0000000300000000ffffff9cffffffff000000e0000000000000002400000000",
            INIT_76 => X"0000003400000000ffffff0cffffffffffffff0affffffff0000003900000000",
            INIT_77 => X"ffffffa6ffffffff0000000d00000000fffffff8ffffffffffffff9effffffff",
            INIT_78 => X"0000002c00000000ffffff16ffffffff0000000b00000000ffffff75ffffffff",
            INIT_79 => X"ffffffc6ffffffff00000025000000000000006d000000000000003000000000",
            INIT_7A => X"00000042000000000000005c00000000fffffff7ffffffff0000000b00000000",
            INIT_7B => X"00000034000000000000000f00000000ffffffd9ffffffffffffffa2ffffffff",
            INIT_7C => X"fffffff2ffffffffffffffdbffffffff0000004b00000000ffffffd9ffffffff",
            INIT_7D => X"0000002f00000000fffffff9ffffffffffffffd2ffffffffffffffc3ffffffff",
            INIT_7E => X"ffffffeeffffffffffffffeaffffffffffffff43ffffffff0000006c00000000",
            INIT_7F => X"0000007000000000ffffffeeffffffffffffff33ffffffffffffff3bffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE24;


    MEM_IWGHT_LAYER2_INSTANCE25 : if BRAM_NAME = "iwght_layer2_instance25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffbaffffffffffffffe7fffffffffffffff5ffffffff0000008800000000",
            INIT_01 => X"0000003a00000000fffffff1ffffffffffffffacffffffff000000bd00000000",
            INIT_02 => X"ffffffefffffffff0000000000000000ffffffe9ffffffffffffff93ffffffff",
            INIT_03 => X"000000510000000000000040000000000000002c00000000ffffff65ffffffff",
            INIT_04 => X"00000030000000000000007400000000000000a200000000fffffffdffffffff",
            INIT_05 => X"ffffffa1ffffffff00000035000000000000004900000000fffffea1ffffffff",
            INIT_06 => X"0000002c00000000000000160000000000000006000000000000001b00000000",
            INIT_07 => X"ffffffceffffffff0000004b000000000000000b000000000000001900000000",
            INIT_08 => X"000000c700000000ffffffbbffffffffffffffb4ffffffffffffffd5ffffffff",
            INIT_09 => X"ffffffa3ffffffffffffffbcffffffff0000003500000000ffffff2effffffff",
            INIT_0A => X"fffffff8fffffffffffffff5ffffffffffffffdeffffffff0000003400000000",
            INIT_0B => X"0000002900000000ffffff6affffffff0000009c000000000000000c00000000",
            INIT_0C => X"ffffffa2ffffffff0000007e00000000ffffff67ffffffff0000008600000000",
            INIT_0D => X"000000120000000000000019000000000000000200000000fffffff6ffffffff",
            INIT_0E => X"fffffffcffffffff00000001000000000000000e000000000000000800000000",
            INIT_0F => X"0000000d00000000fffffff8ffffffff0000000100000000fffffff1ffffffff",
            INIT_10 => X"0000001200000000ffffff94ffffffffffffffc6ffffffffffffffd4ffffffff",
            INIT_11 => X"0000009400000000ffffff71ffffffff0000002600000000ffffffdbffffffff",
            INIT_12 => X"ffffffabffffffff0000007d00000000ffffff3effffffffffffffbdffffffff",
            INIT_13 => X"fffffff0fffffffffffffffaffffffff0000001c00000000000000a000000000",
            INIT_14 => X"0000003d00000000ffffffb6ffffffff00000046000000000000004800000000",
            INIT_15 => X"0000008b000000000000006600000000fffffff3ffffffff0000000200000000",
            INIT_16 => X"ffffff76ffffffff000000c900000000fffffe8affffffffffffffa8ffffffff",
            INIT_17 => X"0000000300000000000000d100000000ffffff1bffffffff0000003800000000",
            INIT_18 => X"ffffff8effffffffffffff98ffffffffffffffd6ffffffff000000b300000000",
            INIT_19 => X"0000007200000000ffffff02ffffffffffffffb8ffffffffffffffeaffffffff",
            INIT_1A => X"000000eb00000000ffffffebffffffffffffff7cffffffff0000003400000000",
            INIT_1B => X"ffffffb0ffffffff000000c500000000fffffee9ffffffffffffffe9ffffffff",
            INIT_1C => X"fffffffcffffffffffffffd5ffffffff00000033000000000000004500000000",
            INIT_1D => X"000000cd00000000ffffff39ffffffff0000007c00000000000000e500000000",
            INIT_1E => X"ffffff77ffffffff0000006c00000000ffffff21fffffffffffffffeffffffff",
            INIT_1F => X"ffffffcaffffffff0000001900000000ffffff30ffffffff0000000400000000",
            INIT_20 => X"00000015000000000000007500000000ffffffbcffffffff000000a600000000",
            INIT_21 => X"ffffffe3ffffffffffffffa1ffffffff0000002700000000ffffff5affffffff",
            INIT_22 => X"00000026000000000000008e00000000fffffff4ffffffff0000007100000000",
            INIT_23 => X"0000007a0000000000000053000000000000006900000000ffffffebffffffff",
            INIT_24 => X"ffffff56ffffffffffffffbcffffffffffffff7bffffffffffffffa0ffffffff",
            INIT_25 => X"ffffff8dffffffffffffff87fffffffffffffff8fffffffffffffff0ffffffff",
            INIT_26 => X"0000000800000000000000110000000000000022000000000000010f00000000",
            INIT_27 => X"fffffff9ffffffffffffffb5ffffffffffffff67ffffffff0000007200000000",
            INIT_28 => X"ffffff9bffffffffffffffa8ffffffff0000004200000000ffffff08ffffffff",
            INIT_29 => X"0000002800000000000000a000000000ffffff63fffffffffffffffbffffffff",
            INIT_2A => X"ffffff74ffffffff0000000800000000ffffff77ffffffffffffffd9ffffffff",
            INIT_2B => X"fffffed3ffffffff000000aa000000000000002500000000ffffff82ffffffff",
            INIT_2C => X"ffffff9bffffffff000000150000000000000007000000000000007900000000",
            INIT_2D => X"ffffffe5fffffffffffffff1ffffffff00000026000000000000009c00000000",
            INIT_2E => X"ffffffd8ffffffffffffffe7ffffffffffffffffffffffff0000000300000000",
            INIT_2F => X"00000034000000000000005100000000000000de00000000ffffffd4ffffffff",
            INIT_30 => X"ffffff84ffffffffffffffb5ffffffffffffffabffffffffffffffdbffffffff",
            INIT_31 => X"0000003300000000ffffff44ffffffffffffffc8ffffffffffffffc7ffffffff",
            INIT_32 => X"000000f800000000ffffffbbffffffffffffffc8ffffffff000000d400000000",
            INIT_33 => X"0000005200000000ffffffe6ffffffff0000001a000000000000007e00000000",
            INIT_34 => X"ffffffd5ffffffff0000005e00000000ffffff4effffffff0000000600000000",
            INIT_35 => X"fffffff3ffffffffffffffc8ffffffff00000089000000000000001a00000000",
            INIT_36 => X"0000003300000000ffffffa0ffffffff000000c8000000000000004500000000",
            INIT_37 => X"0000001200000000000000a000000000fffffffbfffffffffffffffeffffffff",
            INIT_38 => X"ffffffd2ffffffffffffff75ffffffff00000008000000000000003600000000",
            INIT_39 => X"0000005b000000000000004b00000000ffffffadffffffff0000003d00000000",
            INIT_3A => X"0000008a00000000ffffffc2ffffffffffffffabffffffff0000001e00000000",
            INIT_3B => X"0000003d00000000ffffffadffffffffffffffeaffffffff0000001700000000",
            INIT_3C => X"fffffffcffffffffffffffeeffffffff0000000b000000000000005a00000000",
            INIT_3D => X"ffffff3fffffffff0000003e000000000000001500000000ffffff5fffffffff",
            INIT_3E => X"ffffffbeffffffff0000000b000000000000007100000000000000ee00000000",
            INIT_3F => X"ffffffc3ffffffffffffffd7ffffffffffffffa5ffffffff0000001700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000bc00000000ffffffbeffffffff0000002200000000ffffffccffffffff",
            INIT_41 => X"ffffffd5ffffffff0000003500000000ffffff8effffffffffffff80ffffffff",
            INIT_42 => X"000000a500000000ffffff82ffffffff0000006900000000ffffffe3ffffffff",
            INIT_43 => X"ffffff8affffffffffffffeaffffffff0000001900000000ffffffd2ffffffff",
            INIT_44 => X"00000048000000000000004b0000000000000092000000000000006000000000",
            INIT_45 => X"ffffff61ffffffffffffff34ffffffffffffffe6ffffffffffffffbeffffffff",
            INIT_46 => X"0000005300000000ffffffadffffffffffffff4fffffffff000000ae00000000",
            INIT_47 => X"0000005c0000000000000046000000000000003d00000000ffffff9effffffff",
            INIT_48 => X"ffffffe4ffffffff0000004f000000000000000500000000ffffffe9ffffffff",
            INIT_49 => X"ffffffeefffffffffffffffcffffffff000000d700000000ffffffddffffffff",
            INIT_4A => X"ffffffc9ffffffffffffffe6ffffffff00000003000000000000002c00000000",
            INIT_4B => X"ffffffccffffffffffffffe0ffffffff0000004200000000ffffffa1ffffffff",
            INIT_4C => X"0000002c00000000ffffff52fffffffffffffff4ffffffff0000001c00000000",
            INIT_4D => X"ffffff9dffffffff0000006c00000000ffffffd2ffffffffffffffe1ffffffff",
            INIT_4E => X"0000001f000000000000007a0000000000000013000000000000000300000000",
            INIT_4F => X"ffffff93ffffffffffffff66ffffffffffffffb8fffffffffffffffbffffffff",
            INIT_50 => X"0000001e000000000000000f00000000ffffff80fffffffffffffff8ffffffff",
            INIT_51 => X"0000006000000000ffffff71ffffffffffffffe4ffffffffffffffdbffffffff",
            INIT_52 => X"fffffff6ffffffff000000570000000000000015000000000000005000000000",
            INIT_53 => X"000000e700000000000000d100000000ffffffc0ffffffffffffffe7ffffffff",
            INIT_54 => X"ffffffd2ffffffff000000dd000000000000001c00000000000000bd00000000",
            INIT_55 => X"fffffffdffffffff0000001b000000000000001300000000ffffffd8ffffffff",
            INIT_56 => X"fffffffcffffffffffffffeeffffffff0000000e00000000fffffff1ffffffff",
            INIT_57 => X"ffffffbafffffffffffffff9ffffffff00000005000000000000000800000000",
            INIT_58 => X"ffffff89ffffffffffffffddffffffff0000005700000000ffffffadffffffff",
            INIT_59 => X"0000002d000000000000008d00000000000000b200000000ffffffa4ffffffff",
            INIT_5A => X"ffffff1cffffffff0000003b000000000000003e00000000ffffffe8ffffffff",
            INIT_5B => X"ffffffb5ffffffff0000001000000000fffffff7ffffffffffffff80ffffffff",
            INIT_5C => X"0000002600000000000000810000000000000046000000000000007800000000",
            INIT_5D => X"ffffff97ffffffffffffffc2ffffffff00000059000000000000006400000000",
            INIT_5E => X"ffffff4affffffff0000003a0000000000000103000000000000003100000000",
            INIT_5F => X"ffffffd4ffffffffffffff00ffffffff000000ec000000000000006f00000000",
            INIT_60 => X"0000008200000000ffffff8dffffffff00000092000000000000007600000000",
            INIT_61 => X"fffffff5ffffffff00000086000000000000008e00000000ffffff7cffffffff",
            INIT_62 => X"0000002b00000000ffffff83ffffffff0000003d000000000000000c00000000",
            INIT_63 => X"ffffff59ffffffffffffff17ffffffff0000006100000000ffffffdcffffffff",
            INIT_64 => X"fffffef2ffffffffffffffd2ffffffffffffff93ffffffffffffffb5ffffffff",
            INIT_65 => X"ffffffaeffffffff000000db00000000ffffffa4ffffffffffffffceffffffff",
            INIT_66 => X"ffffffe6ffffffffffffff88ffffffffffffffceffffffff0000004d00000000",
            INIT_67 => X"000000d300000000000000a100000000ffffff1fffffffff0000003400000000",
            INIT_68 => X"0000001e00000000ffffffd6ffffffff0000001800000000ffffffc7ffffffff",
            INIT_69 => X"0000006600000000ffffff8fffffffffffffff93fffffffffffffff8ffffffff",
            INIT_6A => X"00000001000000000000005900000000000000b8000000000000004b00000000",
            INIT_6B => X"0000003c00000000ffffffe9ffffffffffffff81ffffffff0000006500000000",
            INIT_6C => X"ffffffcbffffffffffffffffffffffffffffffe8ffffffff0000005100000000",
            INIT_6D => X"ffffffc5ffffffff0000003900000000ffffffb8ffffffffffffffb8ffffffff",
            INIT_6E => X"fffffec6ffffffff0000009800000000ffffffb3ffffffff0000009200000000",
            INIT_6F => X"fffffffbffffffffffffffeeffffffffffffffd9ffffffffffffffe7ffffffff",
            INIT_70 => X"0000006f00000000ffffff8dffffffff0000001600000000ffffff5fffffffff",
            INIT_71 => X"fffffff7ffffffffffffff9effffffffffffffe5ffffffff0000001b00000000",
            INIT_72 => X"ffffffa2ffffffffffffffb5ffffffff00000006000000000000004700000000",
            INIT_73 => X"ffffffe5ffffffffffffff10ffffffff0000000900000000ffffff58ffffffff",
            INIT_74 => X"ffffffc8ffffffffffffff11ffffffffffffffe0ffffffff000000fe00000000",
            INIT_75 => X"000000af000000000000000d00000000ffffffadffffffffffffff97ffffffff",
            INIT_76 => X"ffffff9dffffffff0000002800000000ffffffffffffffff0000007200000000",
            INIT_77 => X"ffffff60ffffffff0000005f000000000000002100000000ffffffc8ffffffff",
            INIT_78 => X"ffffffbeffffffffffffff14ffffffff0000007800000000000000b500000000",
            INIT_79 => X"ffffffe0fffffffffffffffaffffffffffffff91ffffffff0000006300000000",
            INIT_7A => X"ffffff9fffffffff0000000400000000ffffff45fffffffffffffe89ffffffff",
            INIT_7B => X"0000002e00000000ffffff52ffffffffffffff45ffffffffffffff61ffffffff",
            INIT_7C => X"ffffff56ffffffff000000ba0000000000000085000000000000000900000000",
            INIT_7D => X"fffffff3ffffffff0000005c00000000ffffffc9fffffffffffffefdffffffff",
            INIT_7E => X"0000008c00000000ffffff97ffffffff0000004300000000000000b800000000",
            INIT_7F => X"fffffff6ffffffff0000003400000000ffffff94ffffffff0000007e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE25;


    MEM_IWGHT_LAYER2_INSTANCE26 : if BRAM_NAME = "iwght_layer2_instance26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004200000000ffffffc9ffffffff0000001e00000000fffffef4ffffffff",
            INIT_01 => X"ffffffefffffffffffffffdafffffffffffffff0ffffffff0000000c00000000",
            INIT_02 => X"ffffffb4fffffffffffffee2fffffffffffffffdffffffff0000002400000000",
            INIT_03 => X"0000003900000000ffffff84fffffffffffffec3ffffffff0000006600000000",
            INIT_04 => X"ffffff79ffffffff00000021000000000000006d00000000ffffff45ffffffff",
            INIT_05 => X"0000002a000000000000001500000000ffffff0cffffffff0000001000000000",
            INIT_06 => X"fffffffdffffffff000000a9000000000000001700000000ffffff07ffffffff",
            INIT_07 => X"00000080000000000000006d000000000000002d00000000ffffff92ffffffff",
            INIT_08 => X"fffffffcffffffffffffffbeffffffff00000027000000000000003000000000",
            INIT_09 => X"000000700000000000000054000000000000001400000000ffffffffffffffff",
            INIT_0A => X"0000009900000000ffffffbdffffffff00000078000000000000002500000000",
            INIT_0B => X"ffffff80ffffffffffffff89ffffffffffffff3affffffff0000007800000000",
            INIT_0C => X"0000002c00000000ffffff8cffffffff0000001e000000000000001500000000",
            INIT_0D => X"0000002f000000000000004100000000ffffffa0fffffffffffffebcffffffff",
            INIT_0E => X"ffffff7cffffffffffffffdfffffffff00000023000000000000007c00000000",
            INIT_0F => X"ffffffafffffffffffffffb1ffffffff0000004200000000ffffff72ffffffff",
            INIT_10 => X"ffffffa2fffffffffffffe9dffffffffffffffbaffffffffffffffb8ffffffff",
            INIT_11 => X"ffffffddffffffffffffff68ffffffffffffff45ffffffffffffff89ffffffff",
            INIT_12 => X"ffffffa0ffffffff0000004200000000ffffff3cffffffffffffff67ffffffff",
            INIT_13 => X"ffffffa1ffffffff000000d9000000000000004600000000ffffff6cffffffff",
            INIT_14 => X"ffffffedffffffff0000005400000000ffffff9dffffffffffffffbeffffffff",
            INIT_15 => X"00000069000000000000000a000000000000006900000000000000bb00000000",
            INIT_16 => X"0000006800000000ffffffe4ffffffff000000f100000000000000d700000000",
            INIT_17 => X"00000015000000000000000000000000ffffff5effffffffffffffefffffffff",
            INIT_18 => X"ffffff91ffffffffffffffdfffffffffffffff98ffffffffffffffdbffffffff",
            INIT_19 => X"0000007f00000000ffffffcdfffffffffffffff8ffffffffffffffdbffffffff",
            INIT_1A => X"0000003700000000ffffff30ffffffffffffff91fffffffffffffff3ffffffff",
            INIT_1B => X"0000005800000000fffffff0ffffffff00000012000000000000006100000000",
            INIT_1C => X"ffffffcdffffffff000000ad00000000ffffff32ffffffff0000005900000000",
            INIT_1D => X"ffffffebffffffff0000001200000000fffffff6ffffffffffffffd5ffffffff",
            INIT_1E => X"fffffff8ffffffff0000000000000000ffffffffffffffff0000000100000000",
            INIT_1F => X"0000000d00000000ffffff61ffffffffffffffefffffffff0000000a00000000",
            INIT_20 => X"00000054000000000000003e00000000ffffffccffffffffffffffbeffffffff",
            INIT_21 => X"00000032000000000000008c00000000000000e3000000000000009f00000000",
            INIT_22 => X"000000b800000000fffffffaffffffff0000004e00000000ffffff91ffffffff",
            INIT_23 => X"0000002f00000000ffffffd7ffffffff0000005d000000000000002500000000",
            INIT_24 => X"000000360000000000000009000000000000001c00000000fffffff4ffffffff",
            INIT_25 => X"fffffff2ffffffffffffff9affffffff0000000000000000ffffffadffffffff",
            INIT_26 => X"ffffff62ffffffff0000008800000000ffffffb7ffffffffffffffb0ffffffff",
            INIT_27 => X"0000001500000000fffffcf0ffffffff000000a100000000ffffff2effffffff",
            INIT_28 => X"0000008e0000000000000012000000000000007200000000000000f100000000",
            INIT_29 => X"0000004100000000ffffffa9ffffffff00000000000000000000000900000000",
            INIT_2A => X"fffffff5ffffffffffffff9dffffffffffffffb6ffffffffffffffebffffffff",
            INIT_2B => X"ffffff68ffffffff00000006000000000000002300000000fffffffeffffffff",
            INIT_2C => X"ffffffe9ffffffff0000008800000000ffffff63ffffffff0000003900000000",
            INIT_2D => X"0000005400000000000000c300000000ffffff50ffffffffffffffb6ffffffff",
            INIT_2E => X"ffffff59ffffffff0000001100000000ffffff9effffffff0000004100000000",
            INIT_2F => X"ffffffe6ffffffff0000001e000000000000003000000000000000a500000000",
            INIT_30 => X"0000008b000000000000001a00000000ffffff9efffffffffffffff4ffffffff",
            INIT_31 => X"00000091000000000000009500000000fffffffaffffffff0000003400000000",
            INIT_32 => X"ffffffeaffffffff00000061000000000000005c00000000ffffff7cffffffff",
            INIT_33 => X"000000ce00000000ffffffc6ffffffff00000025000000000000001700000000",
            INIT_34 => X"ffffffd2ffffffff0000005400000000fffffeefffffffffffffffa8ffffffff",
            INIT_35 => X"00000022000000000000010f000000000000001e00000000ffffffb8ffffffff",
            INIT_36 => X"000000880000000000000024000000000000002900000000000000c600000000",
            INIT_37 => X"ffffffb2ffffffffffffffaeffffffffffffff22fffffffffffffff2ffffffff",
            INIT_38 => X"ffffffcdffffffffffffffeeffffffff00000012000000000000000400000000",
            INIT_39 => X"0000005d000000000000003c00000000ffffffb0ffffffff0000002400000000",
            INIT_3A => X"ffffffe7ffffffff0000008900000000fffffff8ffffffff0000001200000000",
            INIT_3B => X"ffffffcbffffffffffffff6cffffffff0000010500000000ffffffc7ffffffff",
            INIT_3C => X"ffffff8fffffffff0000003300000000ffffffc3ffffffffffffff83ffffffff",
            INIT_3D => X"fffffed0ffffffffffffffdeffffffff0000002b00000000ffffffefffffffff",
            INIT_3E => X"ffffffc1ffffffff0000003d000000000000005f00000000ffffffb0ffffffff",
            INIT_3F => X"fffffefdffffffff0000009100000000ffffffceffffffff0000006200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f300000000000000540000000000000000000000000000005700000000",
            INIT_41 => X"fffffffbffffffffffffffa6ffffffffffffff97ffffffff000000ef00000000",
            INIT_42 => X"ffffffdbffffffff0000001e00000000ffffff27fffffffffffffe98ffffffff",
            INIT_43 => X"ffffffa3ffffffffffffff79ffffffffffffff4fffffffffffffff46ffffffff",
            INIT_44 => X"ffffff69ffffffff0000001100000000ffffffefffffffff000000c200000000",
            INIT_45 => X"00000001000000000000007d00000000ffffffa2ffffffff0000002300000000",
            INIT_46 => X"ffffffaeffffffff00000050000000000000000d00000000ffffffc8ffffffff",
            INIT_47 => X"ffffffaeffffffffffffffd5ffffffff0000001f000000000000001400000000",
            INIT_48 => X"0000005700000000ffffff9bffffffffffffff5cffffffff0000002300000000",
            INIT_49 => X"ffffffbeffffffff0000007900000000ffffff4cffffffffffffff4effffffff",
            INIT_4A => X"ffffffc6ffffffff00000090000000000000000e00000000ffffffa6ffffffff",
            INIT_4B => X"ffffff53ffffffff0000006b000000000000003b00000000000000f700000000",
            INIT_4C => X"000000ce00000000000000ff000000000000003e000000000000003800000000",
            INIT_4D => X"ffffffb1ffffffffffffffe9ffffffffffffff27ffffffffffffff8fffffffff",
            INIT_4E => X"0000002a00000000ffffff4dffffffff000000cd000000000000002e00000000",
            INIT_4F => X"fffffe04ffffffff0000004a00000000ffffff4bffffffff000000a100000000",
            INIT_50 => X"fffffea7ffffffffffffff97ffffffffffffff6fffffffffffffffb4ffffffff",
            INIT_51 => X"0000010200000000000000090000000000000019000000000000001900000000",
            INIT_52 => X"00000023000000000000001d00000000fffffffeffffffff0000011300000000",
            INIT_53 => X"fffffff9ffffffffffffff9cffffffff0000006c000000000000001700000000",
            INIT_54 => X"0000001d0000000000000025000000000000002e000000000000000000000000",
            INIT_55 => X"ffffffc2fffffffffffffff9ffffffffffffff28ffffffffffffff53ffffffff",
            INIT_56 => X"0000006500000000ffffff9effffffffffffffc6ffffffffffffff58ffffffff",
            INIT_57 => X"00000069000000000000000f00000000ffffff0dffffffff0000005600000000",
            INIT_58 => X"ffffffe2ffffffff0000006f00000000fffffd76ffffffff000000a100000000",
            INIT_59 => X"00000050000000000000004e00000000000000a800000000ffffffcbffffffff",
            INIT_5A => X"fffffff3ffffffffffffff7cffffffff0000001e000000000000002a00000000",
            INIT_5B => X"ffffffd1ffffffff0000000f00000000ffffff9affffffff0000001100000000",
            INIT_5C => X"0000000600000000ffffff49ffffffff00000021000000000000009600000000",
            INIT_5D => X"000000df00000000fffffff7ffffffff00000013000000000000003700000000",
            INIT_5E => X"0000006100000000ffffffefffffffffffffffc6ffffffff0000018c00000000",
            INIT_5F => X"ffffffb0ffffffffffffffc0fffffffffffffe74ffffffff0000001e00000000",
            INIT_60 => X"ffffff61ffffffff000000880000000000000045000000000000008600000000",
            INIT_61 => X"0000004c000000000000002000000000ffffffaeffffffff000000eb00000000",
            INIT_62 => X"00000017000000000000003600000000ffffffdcffffffffffffffbdffffffff",
            INIT_63 => X"ffffff87ffffffff0000001200000000fffffffaffffffffffffff95ffffffff",
            INIT_64 => X"ffffff8bfffffffffffffe89ffffffff0000000f00000000000000e900000000",
            INIT_65 => X"fffffff5fffffffffffffff4ffffffff0000000700000000000000ac00000000",
            INIT_66 => X"fffffff7fffffffffffffff8fffffffffffffffbfffffffffffffff9ffffffff",
            INIT_67 => X"00000008000000000000003300000000fffffff8fffffffffffffffdffffffff",
            INIT_68 => X"ffffff59ffffffff00000067000000000000001900000000ffffffbbffffffff",
            INIT_69 => X"ffffffefffffffffffffff80ffffffff00000043000000000000003a00000000",
            INIT_6A => X"0000007800000000fffffecaffffffffffffffbaffffffffffffff08ffffffff",
            INIT_6B => X"00000041000000000000000900000000ffffff6affffffffffffffc8ffffffff",
            INIT_6C => X"ffffff92fffffffffffffe87ffffffffffffffefffffffffffffff60ffffffff",
            INIT_6D => X"ffffff51ffffffff000000a6000000000000007800000000ffffff93ffffffff",
            INIT_6E => X"ffffff87ffffffffffffff44ffffffffffffff8affffffff000000b000000000",
            INIT_6F => X"0000006b000000000000000900000000000000f500000000ffffff53ffffffff",
            INIT_70 => X"0000004b000000000000003d000000000000000700000000ffffff0affffffff",
            INIT_71 => X"0000000a00000000ffffff42fffffffffffffd79fffffffffffffeafffffffff",
            INIT_72 => X"0000001a00000000000000e100000000ffffff4efffffffffffffe29ffffffff",
            INIT_73 => X"ffffffc0ffffffff00000014000000000000001c000000000000004a00000000",
            INIT_74 => X"ffffffb9ffffffff00000036000000000000001600000000ffffff77ffffffff",
            INIT_75 => X"0000007b000000000000003a000000000000003500000000ffffffcfffffffff",
            INIT_76 => X"fffffef8ffffffffffffff68ffffffff000000d7000000000000002100000000",
            INIT_77 => X"0000003a000000000000010f00000000fffffefcffffffff0000001a00000000",
            INIT_78 => X"ffffff6fffffffff0000003c0000000000000034000000000000008100000000",
            INIT_79 => X"ffffffcaffffffffffffffa6ffffffff000000ac000000000000009400000000",
            INIT_7A => X"0000005500000000ffffff2cfffffffffffffed4ffffffffffffffc2ffffffff",
            INIT_7B => X"ffffff47ffffffffffffffe2fffffffffffffdacffffffff0000002d00000000",
            INIT_7C => X"0000008c00000000ffffffcefffffffffffffff5ffffffff0000006200000000",
            INIT_7D => X"ffffff77ffffffff00000070000000000000000d000000000000003b00000000",
            INIT_7E => X"ffffff98ffffffffffffffc3ffffffffffffff90ffffffffffffffb8ffffffff",
            INIT_7F => X"fffffefaffffffff0000003c000000000000009f00000000ffffff39ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE26;


    MEM_IWGHT_LAYER2_INSTANCE27 : if BRAM_NAME = "iwght_layer2_instance27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000008c000000000000003d00000000ffffffaaffffffffffffff3cffffffff",
            INIT_01 => X"ffffff9bffffffff000000be00000000fffffed6ffffffffffffff3affffffff",
            INIT_02 => X"00000033000000000000003d000000000000006a00000000000000d400000000",
            INIT_03 => X"ffffff59ffffffffffffff8dffffffffffffff55ffffffff000000a800000000",
            INIT_04 => X"ffffff3bfffffffffffffed6ffffffffffffffb1ffffffff0000009800000000",
            INIT_05 => X"fffffedbffffffffffffffa9ffffffff0000003600000000fffffeceffffffff",
            INIT_06 => X"0000006e00000000ffffffd5ffffffff0000001700000000000000d100000000",
            INIT_07 => X"ffffffceffffffffffffffcdffffffff0000002f00000000ffffffcfffffffff",
            INIT_08 => X"fffffef3ffffffff000000260000000000000015000000000000004900000000",
            INIT_09 => X"ffffff7cffffffffffffffa4ffffffffffffff87ffffffffffffffb3ffffffff",
            INIT_0A => X"ffffffb2ffffffffffffff9dffffffff000000f100000000ffffffc2ffffffff",
            INIT_0B => X"0000004b0000000000000017000000000000006a000000000000007e00000000",
            INIT_0C => X"0000005e00000000fffffef2ffffffff0000007300000000ffffff47ffffffff",
            INIT_0D => X"ffffff95ffffffff0000002600000000fffffffbffffffff0000002200000000",
            INIT_0E => X"ffffffaeffffffff0000011900000000ffffff59ffffffff0000008900000000",
            INIT_0F => X"fffffff0fffffffffffffffbffffffffffffff7dfffffffffffffe91ffffffff",
            INIT_10 => X"0000005f00000000ffffffb5ffffffffffffff2dffffffff0000005000000000",
            INIT_11 => X"0000004b000000000000000200000000ffffff75ffffffffffffff4effffffff",
            INIT_12 => X"0000005700000000ffffff54ffffffffffffffd4ffffffffffffff83ffffffff",
            INIT_13 => X"ffffffcafffffffffffffffaffffffffffffff2dffffffffffffffebffffffff",
            INIT_14 => X"0000002500000000ffffff0fffffffff0000000900000000ffffffe5ffffffff",
            INIT_15 => X"0000002600000000000000b900000000ffffff2cffffffff000000fc00000000",
            INIT_16 => X"0000004d000000000000009500000000ffffff4fffffffffffffffdaffffffff",
            INIT_17 => X"ffffffa7ffffffffffffffe9ffffffff0000005d00000000000000d100000000",
            INIT_18 => X"ffffff9dffffffffffffffffffffffffffffffa2ffffffff0000001300000000",
            INIT_19 => X"ffffffe6ffffffffffffff42ffffffffffffffebffffffffffffff67ffffffff",
            INIT_1A => X"0000009b00000000000000af00000000ffffff13ffffffff0000001c00000000",
            INIT_1B => X"0000006b00000000ffffffb6ffffffffffffffd8ffffffffffffffc6ffffffff",
            INIT_1C => X"ffffffeeffffffff00000079000000000000002900000000fffffecbffffffff",
            INIT_1D => X"0000001900000000ffffff9fffffffffffffff8effffffffffffffb3ffffffff",
            INIT_1E => X"0000007d00000000ffffffe8fffffffffffffff7ffffffff0000003b00000000",
            INIT_1F => X"000000350000000000000079000000000000000000000000ffffff87ffffffff",
            INIT_20 => X"ffffff95ffffffffffffffebffffffffffffff9bffffffffffffff5bffffffff",
            INIT_21 => X"0000004f00000000ffffffb4ffffffffffffffe8ffffffff0000007a00000000",
            INIT_22 => X"ffffffa5ffffffff000000480000000000000017000000000000000300000000",
            INIT_23 => X"ffffff9cffffffffffffffe3ffffffff0000006d000000000000000000000000",
            INIT_24 => X"0000003700000000000000c100000000ffffffeaffffffff0000000000000000",
            INIT_25 => X"0000005e00000000ffffffedfffffffffffffff4ffffffff0000001a00000000",
            INIT_26 => X"fffffff9ffffffff0000004f00000000ffffffaeffffffffffffff7cffffffff",
            INIT_27 => X"ffffffd3ffffffff0000000400000000ffffffb1ffffffffffffff82ffffffff",
            INIT_28 => X"fffffe0bffffffffffffffdfffffffff0000002800000000fffffffcffffffff",
            INIT_29 => X"ffffffb6ffffffffffffffaaffffffff0000013400000000ffffff90ffffffff",
            INIT_2A => X"0000013700000000ffffff6dffffffffffffffebffffffff0000010700000000",
            INIT_2B => X"ffffffd6ffffffffffffff88ffffffff000000aa00000000fffffff2ffffffff",
            INIT_2C => X"ffffff9dffffffffffffffc7ffffffff0000002e00000000ffffffd6ffffffff",
            INIT_2D => X"0000000300000000000000130000000000000001000000000000009500000000",
            INIT_2E => X"ffffffe7fffffffffffffff2fffffffffffffffdffffffff0000000500000000",
            INIT_2F => X"ffffffd9ffffffffffffffe2ffffffff0000000000000000fffffffaffffffff",
            INIT_30 => X"ffffffb2ffffffff0000013c00000000000000a1000000000000003f00000000",
            INIT_31 => X"ffffffc0fffffffffffffe3effffffff00000017000000000000002600000000",
            INIT_32 => X"00000036000000000000001200000000ffffffc5ffffffff000000b600000000",
            INIT_33 => X"ffffffe6ffffffffffffff6affffffffffffff9fffffffff0000007d00000000",
            INIT_34 => X"ffffff6fffffffff0000003c00000000ffffffa1ffffffffffffff9cffffffff",
            INIT_35 => X"0000004f00000000ffffff76ffffffffffffffcbffffffff0000008b00000000",
            INIT_36 => X"0000002f000000000000007d00000000ffffff97ffffffffffffff00ffffffff",
            INIT_37 => X"fffffedcffffffff0000007f00000000ffffff4bffffffffffffffc8ffffffff",
            INIT_38 => X"00000008000000000000008e00000000ffffff58ffffffffffffff8bffffffff",
            INIT_39 => X"fffffeeeffffffffffffff24ffffffff0000002300000000ffffff59ffffffff",
            INIT_3A => X"00000042000000000000004200000000fffffffcffffffffffffffceffffffff",
            INIT_3B => X"00000020000000000000001c00000000ffffffb3ffffffff000000cd00000000",
            INIT_3C => X"0000006900000000ffffff9cffffffff0000002600000000ffffffd1ffffffff",
            INIT_3D => X"ffffffaeffffffff0000004600000000ffffff72fffffffffffffff5ffffffff",
            INIT_3E => X"ffffffd6ffffffff00000018000000000000009600000000ffffffcfffffffff",
            INIT_3F => X"000000cb00000000ffffffe6ffffffff0000002a00000000ffffffa7ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffa0ffffffffffffffc3ffffffff0000006b00000000ffffff62ffffffff",
            INIT_41 => X"ffffffdfffffffff0000002a00000000ffffff85ffffffff0000005300000000",
            INIT_42 => X"ffffffbdffffffff0000002a00000000000000bf00000000ffffffe4ffffffff",
            INIT_43 => X"ffffffdeffffffff0000005b00000000ffffffd0ffffffffffffffbeffffffff",
            INIT_44 => X"0000004a00000000ffffff91ffffffff0000009c00000000ffffff28ffffffff",
            INIT_45 => X"00000023000000000000009f000000000000001600000000ffffff93ffffffff",
            INIT_46 => X"0000004f00000000ffffffb9ffffffff0000003d00000000ffffffd0ffffffff",
            INIT_47 => X"00000022000000000000006400000000fffffedaffffffff0000007000000000",
            INIT_48 => X"ffffffa7ffffffff0000004500000000000000af000000000000004100000000",
            INIT_49 => X"00000094000000000000003f00000000ffffff92ffffffff0000000b00000000",
            INIT_4A => X"0000001b00000000ffffffb6ffffffffffffffdcffffffff0000004700000000",
            INIT_4B => X"0000004e000000000000002a0000000000000038000000000000008b00000000",
            INIT_4C => X"00000028000000000000002a000000000000002400000000ffffffbaffffffff",
            INIT_4D => X"0000004700000000ffffffb0ffffffffffffff9bffffffff000000d200000000",
            INIT_4E => X"ffffff3cffffffff0000002300000000ffffffe2ffffffffffffff90ffffffff",
            INIT_4F => X"fffffff4ffffffffffffff70ffffffff00000100000000000000000d00000000",
            INIT_50 => X"0000000300000000ffffffcdfffffffffffffebdffffffff0000008700000000",
            INIT_51 => X"ffffffe5ffffffff0000004600000000ffffffb0ffffffffffffff4affffffff",
            INIT_52 => X"0000003500000000ffffff99ffffffff00000088000000000000003d00000000",
            INIT_53 => X"ffffff11ffffffff0000005700000000ffffffd2ffffffff0000005f00000000",
            INIT_54 => X"ffffffecffffffff000000230000000000000027000000000000005300000000",
            INIT_55 => X"ffffffc6ffffffff0000001500000000fffffffbffffffffffffffdeffffffff",
            INIT_56 => X"fffffff7ffffffffffffffcbffffffffffffffc4ffffffff0000000700000000",
            INIT_57 => X"000000530000000000000036000000000000005700000000ffffff4bffffffff",
            INIT_58 => X"000000b300000000000000a80000000000000057000000000000001e00000000",
            INIT_59 => X"0000007600000000ffffffa3ffffffff000000ec000000000000008600000000",
            INIT_5A => X"ffffff9bffffffffffffffe4ffffffffffffffe8ffffffff0000006000000000",
            INIT_5B => X"0000002100000000ffffffafffffffff000000da000000000000002200000000",
            INIT_5C => X"ffffffd7ffffffff0000006600000000ffffff3fffffffff0000001c00000000",
            INIT_5D => X"000000aa000000000000008900000000ffffff45fffffffffffffff4ffffffff",
            INIT_5E => X"fffffeccffffffff0000005400000000ffffff4cffffffff0000001e00000000",
            INIT_5F => X"fffffff4ffffffffffffff5fffffffff0000007b00000000ffffffc2ffffffff",
            INIT_60 => X"ffffff92ffffffffffffff99ffffffff0000009e00000000ffffff86ffffffff",
            INIT_61 => X"0000003600000000ffffffb9ffffffff00000053000000000000006600000000",
            INIT_62 => X"ffffffa7ffffffffffffff63ffffffffffffffcbffffffffffffffb6ffffffff",
            INIT_63 => X"ffffffebffffffff0000004a0000000000000013000000000000004500000000",
            INIT_64 => X"0000001b00000000fffffffeffffffffffffffb7ffffffff0000006700000000",
            INIT_65 => X"0000000500000000ffffff8efffffffffffffff4ffffffff0000007200000000",
            INIT_66 => X"ffffff64fffffffffffffff5ffffffffffffff99ffffffff0000003d00000000",
            INIT_67 => X"00000018000000000000003a0000000000000039000000000000005f00000000",
            INIT_68 => X"0000006200000000fffffefdffffffff00000035000000000000006800000000",
            INIT_69 => X"ffffffc3ffffffff00000004000000000000002400000000ffffffe4ffffffff",
            INIT_6A => X"0000007b00000000ffffffe7ffffffff00000077000000000000000e00000000",
            INIT_6B => X"0000000b000000000000000000000000ffffffdbffffffffffffffd1ffffffff",
            INIT_6C => X"ffffffe2ffffffff0000000300000000fffffff0ffffffffffffffbaffffffff",
            INIT_6D => X"fffffef0ffffffffffffff55fffffffffffffffcffffffff0000005a00000000",
            INIT_6E => X"0000002900000000ffffffa8ffffffff0000002a000000000000002200000000",
            INIT_6F => X"0000006b0000000000000015000000000000001000000000fffffedfffffffff",
            INIT_70 => X"fffffffeffffffff00000064000000000000004600000000ffffffffffffffff",
            INIT_71 => X"0000000a00000000000000c600000000ffffffc4ffffffff0000000200000000",
            INIT_72 => X"0000001e0000000000000006000000000000000b00000000ffffff59ffffffff",
            INIT_73 => X"fffffff2fffffffffffffff9ffffffff0000002000000000ffffffbbffffffff",
            INIT_74 => X"ffffffbbffffffffffffff93ffffffff00000033000000000000008400000000",
            INIT_75 => X"fffffff6fffffffffffffffafffffffffffffffdffffffffffffff9bffffffff",
            INIT_76 => X"fffffff8ffffffff00000002000000000000000d00000000ffffffe9ffffffff",
            INIT_77 => X"0000004500000000ffffffe4fffffffffffffff5ffffffff0000001700000000",
            INIT_78 => X"ffffffcaffffffffffffffb8ffffffffffffff61ffffffff0000008c00000000",
            INIT_79 => X"0000002b0000000000000075000000000000002300000000ffffff90ffffffff",
            INIT_7A => X"ffffff91ffffffff00000039000000000000004800000000fffffee4ffffffff",
            INIT_7B => X"0000001900000000ffffff71ffffffff0000005600000000ffffffedffffffff",
            INIT_7C => X"ffffffc1ffffffff000000b50000000000000065000000000000000100000000",
            INIT_7D => X"fffffffaffffffff0000001e000000000000007c000000000000005200000000",
            INIT_7E => X"000000b2000000000000006700000000ffffff50ffffffff0000007500000000",
            INIT_7F => X"000000840000000000000054000000000000004e00000000fffffef3ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE27;


    MEM_IWGHT_LAYER2_INSTANCE28 : if BRAM_NAME = "iwght_layer2_instance28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffe5ffffffffffffff5cffffffffffffff94ffffffff0000006900000000",
            INIT_01 => X"ffffffc8ffffffff0000008f00000000ffffffb6ffffffffffffffccffffffff",
            INIT_02 => X"ffffff68ffffffff00000044000000000000000b00000000fffffff3ffffffff",
            INIT_03 => X"fffffff6fffffffffffffee9ffffffffffffffd7ffffffffffffffc2ffffffff",
            INIT_04 => X"00000034000000000000006400000000ffffffd9fffffffffffffff6ffffffff",
            INIT_05 => X"ffffffbcffffffff0000006e0000000000000070000000000000003b00000000",
            INIT_06 => X"ffffffd4ffffffffffffffbcffffffffffffffdbffffffff000000e500000000",
            INIT_07 => X"fffffffcffffffff000000170000000000000085000000000000006b00000000",
            INIT_08 => X"0000009d00000000000000b5000000000000002600000000fffffff3ffffffff",
            INIT_09 => X"ffffff64ffffffffffffff8effffffffffffff7ffffffffffffffec9ffffffff",
            INIT_0A => X"fffffecdffffffff0000006400000000fffffec8ffffffff0000009100000000",
            INIT_0B => X"0000003900000000ffffff9cffffffff0000008600000000ffffffedffffffff",
            INIT_0C => X"ffffffb6ffffffff0000001d00000000ffffffdbffffffffffffffd7ffffffff",
            INIT_0D => X"fffffed5ffffffff0000006d00000000ffffffc8fffffffffffffff0ffffffff",
            INIT_0E => X"fffffffefffffffffffffec7ffffffff0000004d000000000000002700000000",
            INIT_0F => X"fffffffcffffffff00000036000000000000006700000000ffffffcdffffffff",
            INIT_10 => X"ffffffffffffffff0000002500000000ffffffdcffffffffffffffc1ffffffff",
            INIT_11 => X"0000003600000000ffffff4fffffffffffffffc6ffffffffffffffc0ffffffff",
            INIT_12 => X"ffffff6bffffffffffffffe1ffffffff0000007200000000ffffffb2ffffffff",
            INIT_13 => X"ffffff9cffffffff000000300000000000000057000000000000003300000000",
            INIT_14 => X"0000003d00000000ffffff85fffffffffffffff2ffffffff0000006b00000000",
            INIT_15 => X"ffffffd1ffffffffffffff13ffffffff0000007100000000000000c400000000",
            INIT_16 => X"ffffff1affffffffffffff00ffffffffffffff74fffffffffffffff1ffffffff",
            INIT_17 => X"ffffffc7ffffffff0000003d00000000ffffff83ffffffff0000000c00000000",
            INIT_18 => X"0000002000000000ffffff92ffffffffffffffdaffffffff0000001100000000",
            INIT_19 => X"00000083000000000000004300000000ffffff99ffffffff0000003d00000000",
            INIT_1A => X"0000003e0000000000000024000000000000002400000000ffffff9effffffff",
            INIT_1B => X"ffffff3bffffffffffffffe5ffffffff0000000000000000ffffff48ffffffff",
            INIT_1C => X"ffffffc5ffffffff0000009900000000ffffffb1ffffffffffffff16ffffffff",
            INIT_1D => X"ffffffd7ffffffffffffff8bffffffffffffff7fffffffff0000008e00000000",
            INIT_1E => X"00000057000000000000001e000000000000002400000000ffffff88ffffffff",
            INIT_1F => X"000000780000000000000049000000000000003a000000000000008e00000000",
            INIT_20 => X"0000002b00000000ffffffdfffffffff0000009d000000000000005300000000",
            INIT_21 => X"ffffffa9ffffffffffffffeaffffffff0000006f000000000000005c00000000",
            INIT_22 => X"00000098000000000000001400000000ffffffacffffffff0000005800000000",
            INIT_23 => X"ffffffbaffffffff0000001300000000ffffffccffffffff0000001f00000000",
            INIT_24 => X"000000b000000000fffffedfffffffff000000d100000000fffffff1ffffffff",
            INIT_25 => X"0000000f00000000ffffffb0ffffffff0000009d000000000000001500000000",
            INIT_26 => X"0000003300000000ffffff8bffffffff0000004c000000000000003300000000",
            INIT_27 => X"fffffeb9ffffffffffffff99fffffffffffffefbffffffff0000001100000000",
            INIT_28 => X"ffffffcdffffffffffffffe7ffffffffffffff87ffffffffffffff91ffffffff",
            INIT_29 => X"0000001800000000ffffffdbffffffff0000004e000000000000003300000000",
            INIT_2A => X"ffffff11ffffffffffffffbcfffffffffffffff6fffffffffffffffeffffffff",
            INIT_2B => X"ffffffadffffffffffffff81ffffffffffffff31ffffffff0000000400000000",
            INIT_2C => X"00000071000000000000006900000000fffffffeffffffff0000001800000000",
            INIT_2D => X"ffffffb1ffffffffffffffa8ffffffff0000009000000000ffffff65ffffffff",
            INIT_2E => X"fffffffaffffffff00000005000000000000006d000000000000003c00000000",
            INIT_2F => X"ffffffa2ffffffffffffff97ffffffff000000d000000000ffffffd2ffffffff",
            INIT_30 => X"00000030000000000000006700000000fffffed7ffffffff0000006300000000",
            INIT_31 => X"ffffffeaffffffff0000008b000000000000004900000000ffffffc8ffffffff",
            INIT_32 => X"ffffffe9ffffffff0000004600000000fffffff7ffffffff0000001a00000000",
            INIT_33 => X"0000000400000000ffffffb0ffffffff00000025000000000000006f00000000",
            INIT_34 => X"0000002d00000000000000250000000000000050000000000000002300000000",
            INIT_35 => X"0000002700000000ffffffaaffffffffffffffd8ffffffffffffffddffffffff",
            INIT_36 => X"00000017000000000000005800000000ffffffa8ffffffffffffff52ffffffff",
            INIT_37 => X"ffffff9afffffffffffffffbffffffffffffff4dfffffffffffffff3ffffffff",
            INIT_38 => X"00000086000000000000003c0000000000000015000000000000002000000000",
            INIT_39 => X"ffffff77ffffffffffffffa9ffffffff00000054000000000000002e00000000",
            INIT_3A => X"0000003d0000000000000074000000000000005400000000ffffffdaffffffff",
            INIT_3B => X"0000000d00000000ffffffefffffffffffffff07ffffffff0000000b00000000",
            INIT_3C => X"fffffff5ffffffff0000002800000000ffffff71ffffffffffffffc9ffffffff",
            INIT_3D => X"fffffff7ffffffff00000006000000000000000200000000fffffeedffffffff",
            INIT_3E => X"fffffffeffffffff0000000c00000000fffffff8ffffffffffffffefffffffff",
            INIT_3F => X"ffffffcfffffffff0000001e0000000000000005000000000000000200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004400000000000000480000000000000058000000000000001700000000",
            INIT_41 => X"0000009e000000000000005100000000ffffffbdffffffffffffff7bffffffff",
            INIT_42 => X"ffffff6dffffffffffffff6dffffffffffffff5dffffffff0000001900000000",
            INIT_43 => X"0000005500000000ffffff4affffffffffffffd6ffffffff0000002900000000",
            INIT_44 => X"ffffff90ffffffff000000860000000000000007000000000000005800000000",
            INIT_45 => X"ffffff31ffffffffffffffb6ffffffff0000005b00000000fffffec7ffffffff",
            INIT_46 => X"000000070000000000000077000000000000007800000000ffffffedffffffff",
            INIT_47 => X"0000007100000000ffffffd5ffffffffffffffebffffffff0000000a00000000",
            INIT_48 => X"ffffff96ffffffff0000003a00000000ffffff5cffffffffffffff2cffffffff",
            INIT_49 => X"0000009a000000000000006e00000000ffffffb2ffffffffffffffd0ffffffff",
            INIT_4A => X"0000001100000000ffffff7cffffffff0000010c00000000ffffffa0ffffffff",
            INIT_4B => X"000000ea00000000ffffff73ffffffffffffff80ffffffff0000006300000000",
            INIT_4C => X"ffffffddffffffffffffff84ffffffffffffffcfffffffffffffffc9ffffffff",
            INIT_4D => X"fffffeefffffffff0000006100000000ffffff86fffffffffffffffaffffffff",
            INIT_4E => X"fffffff6ffffffff000000fe00000000ffffff75ffffffffffffffd6ffffffff",
            INIT_4F => X"0000006200000000ffffff88ffffffff0000000c000000000000002a00000000",
            INIT_50 => X"00000119000000000000005e0000000000000026000000000000000000000000",
            INIT_51 => X"0000005b000000000000002e00000000ffffffd9fffffffffffffeecffffffff",
            INIT_52 => X"0000005200000000000000040000000000000073000000000000001700000000",
            INIT_53 => X"00000050000000000000002200000000ffffffd0ffffffffffffffcaffffffff",
            INIT_54 => X"00000031000000000000003b00000000ffffffa7ffffffff0000003d00000000",
            INIT_55 => X"0000002100000000ffffffc5ffffffff0000001500000000ffffff96ffffffff",
            INIT_56 => X"fffffe4cffffffffffffff0cffffffffffffff9dfffffffffffffe6cffffffff",
            INIT_57 => X"fffffec0ffffffff0000008a00000000fffffeebffffffffffffff43ffffffff",
            INIT_58 => X"ffffff23ffffffffffffffb3ffffffffffffff02ffffffffffffffa4ffffffff",
            INIT_59 => X"00000104000000000000005600000000ffffffe2ffffffff0000007c00000000",
            INIT_5A => X"fffffffaffffffffffffffa4ffffffff0000002a00000000000000c200000000",
            INIT_5B => X"fffffffdfffffffffffffff7ffffffffffffff57ffffffff0000004400000000",
            INIT_5C => X"0000006100000000000000760000000000000004000000000000003400000000",
            INIT_5D => X"ffffffe9ffffffff0000002e000000000000004000000000ffffffd8ffffffff",
            INIT_5E => X"0000000400000000ffffff80ffffffff0000003900000000ffffff94ffffffff",
            INIT_5F => X"000000780000000000000019000000000000003d000000000000002100000000",
            INIT_60 => X"ffffffeeffffffff0000009500000000ffffff4fffffffff0000000f00000000",
            INIT_61 => X"ffffffd9ffffffff0000002300000000ffffff92ffffffffffffff81ffffffff",
            INIT_62 => X"0000004e000000000000002500000000ffffffebffffffff0000000c00000000",
            INIT_63 => X"fffffffdfffffffffffffec8fffffffffffffed8ffffffffffffff6dffffffff",
            INIT_64 => X"0000000800000000ffffff6ffffffffffffffffcffffffffffffff7dffffffff",
            INIT_65 => X"00000020000000000000007200000000ffffffddffffffff0000002100000000",
            INIT_66 => X"0000001000000000ffffff94ffffffff000000d000000000fffffffaffffffff",
            INIT_67 => X"0000001f00000000000000ad00000000fffffed6ffffffffffffffb2ffffffff",
            INIT_68 => X"0000006f00000000ffffff98ffffffffffffffe3ffffffff0000007c00000000",
            INIT_69 => X"ffffffb4ffffffffffffffaaffffffff0000007600000000ffffffc9ffffffff",
            INIT_6A => X"0000007800000000fffffea3fffffffffffffdc4ffffffff000000a100000000",
            INIT_6B => X"00000041000000000000000c000000000000000d000000000000003500000000",
            INIT_6C => X"0000001d0000000000000018000000000000004f000000000000006100000000",
            INIT_6D => X"0000006900000000ffffff76ffffffffffffff32ffffffffffffffd0ffffffff",
            INIT_6E => X"ffffff9effffffffffffffeaffffffff0000007000000000ffffffe6ffffffff",
            INIT_6F => X"ffffffc1ffffffffffffff71ffffffffffffffa5ffffffff000000cb00000000",
            INIT_70 => X"0000002500000000ffffff20ffffffff0000007d000000000000002f00000000",
            INIT_71 => X"000000cc00000000fffffebcffffffffffffff68ffffffffffffff2bffffffff",
            INIT_72 => X"ffffff4dffffffff000000c500000000ffffff9cffffffffffffffefffffffff",
            INIT_73 => X"fffffff1ffffffffffffffc4ffffffffffffffd1ffffffff0000001300000000",
            INIT_74 => X"0000007d00000000ffffffe9ffffffff0000009100000000000000b900000000",
            INIT_75 => X"0000009e00000000fffffef7ffffffff00000041000000000000001900000000",
            INIT_76 => X"ffffffceffffffff0000000b000000000000008d00000000fffffffcffffffff",
            INIT_77 => X"ffffff2fffffffff000000190000000000000078000000000000005a00000000",
            INIT_78 => X"ffffffddffffffffffffffc9ffffffff00000085000000000000001d00000000",
            INIT_79 => X"0000005e000000000000002700000000ffffff66ffffffffffffff79ffffffff",
            INIT_7A => X"ffffffdbffffffffffffffbdffffffff0000007d00000000ffffff42ffffffff",
            INIT_7B => X"ffffffe1ffffffff0000004e0000000000000039000000000000005a00000000",
            INIT_7C => X"ffffff89fffffffffffffef1ffffffffffffff6dffffffff0000005300000000",
            INIT_7D => X"0000007100000000ffffffdfffffffffffffffceffffffffffffffeaffffffff",
            INIT_7E => X"ffffffdcffffffffffffff99ffffffff00000012000000000000007c00000000",
            INIT_7F => X"00000005000000000000004300000000ffffff2fffffffffffffffabffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE28;


    MEM_IWGHT_LAYER2_INSTANCE29 : if BRAM_NAME = "iwght_layer2_instance29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffc4ffffffff000000b300000000ffffff97ffffffffffffff85ffffffff",
            INIT_01 => X"00000026000000000000003c00000000ffffffd5ffffffffffffffdaffffffff",
            INIT_02 => X"ffffffeeffffffffffffffc1ffffffff0000007500000000ffffffb0ffffffff",
            INIT_03 => X"ffffff74ffffffffffffff8affffffffffffffcfffffffffffffffafffffffff",
            INIT_04 => X"0000008d000000000000001d00000000ffffff60ffffffffffffff68ffffffff",
            INIT_05 => X"fffffff3ffffffffffffffeffffffffffffffffdffffffffffffffe7ffffffff",
            INIT_06 => X"fffffff2fffffffffffffff7fffffffffffffff5ffffffff0000000c00000000",
            INIT_07 => X"000000a000000000ffffffddffffffff00000000000000000000000700000000",
            INIT_08 => X"0000003600000000ffffff9affffffff0000008a000000000000007700000000",
            INIT_09 => X"00000015000000000000003300000000ffffff49ffffffffffffff60ffffffff",
            INIT_0A => X"0000007a00000000ffffff55ffffffffffffffa3ffffffff0000006200000000",
            INIT_0B => X"0000005600000000ffffffa5ffffffff0000001000000000ffffffb8ffffffff",
            INIT_0C => X"ffffff63fffffffffffffff1ffffffff00000016000000000000003f00000000",
            INIT_0D => X"ffffff56ffffffff00000023000000000000009300000000ffffff99ffffffff",
            INIT_0E => X"0000000f00000000ffffff47ffffffffffffffa9ffffffffffffffc6ffffffff",
            INIT_0F => X"ffffffe7ffffffff0000007d00000000000000e700000000ffffffbeffffffff",
            INIT_10 => X"0000002700000000ffffff58ffffffff0000007b00000000ffffff79ffffffff",
            INIT_11 => X"0000008d000000000000006e00000000fffffe5effffffffffffffb1ffffffff",
            INIT_12 => X"0000005700000000000000ca000000000000005800000000ffffff6cffffffff",
            INIT_13 => X"0000005a00000000ffffffdcffffffffffffff4dffffffffffffffd3ffffffff",
            INIT_14 => X"ffffffefffffffff0000000800000000ffffffe7ffffffffffffff8fffffffff",
            INIT_15 => X"ffffff34ffffffff0000007900000000ffffff1effffffffffffff81ffffffff",
            INIT_16 => X"ffffffcfffffffff00000039000000000000009d000000000000001300000000",
            INIT_17 => X"ffffff40fffffffffffffd5fffffffffffffff97ffffffff0000001a00000000",
            INIT_18 => X"ffffff6bffffffff0000009700000000ffffffd2ffffffffffffff1effffffff",
            INIT_19 => X"ffffff7bffffffffffffff87ffffffff00000027000000000000006c00000000",
            INIT_1A => X"0000007e00000000000000c600000000ffffff91ffffffff0000014000000000",
            INIT_1B => X"00000088000000000000004e000000000000006200000000fffffffbffffffff",
            INIT_1C => X"00000010000000000000000200000000ffffff9bffffffffffffff45ffffffff",
            INIT_1D => X"ffffffcfffffffff00000083000000000000004100000000ffffff50ffffffff",
            INIT_1E => X"ffffffafffffffffffffffd4ffffffff0000004000000000ffffffc6ffffffff",
            INIT_1F => X"0000004200000000000000ef000000000000002400000000ffffffe9ffffffff",
            INIT_20 => X"0000007300000000ffffffacffffffffffffff5cffffffffffffffc0ffffffff",
            INIT_21 => X"ffffffeeffffffffffffffc6ffffffff0000004800000000ffffffc4ffffffff",
            INIT_22 => X"ffffffeeffffffff0000000400000000fffffff0ffffffff0000006600000000",
            INIT_23 => X"00000082000000000000001100000000ffffffd2ffffffffffffffdfffffffff",
            INIT_24 => X"0000002600000000ffffffa4ffffffff000000aa00000000fffffff5ffffffff",
            INIT_25 => X"0000000a00000000ffffffd6ffffffffffffff93ffffffffffffffb0ffffffff",
            INIT_26 => X"00000048000000000000004e000000000000003900000000ffffff9fffffffff",
            INIT_27 => X"fffffff8ffffffff0000005500000000ffffff90ffffffffffffff9dffffffff",
            INIT_28 => X"ffffffa2ffffffffffffffa0ffffffffffffff7fffffffff000000cd00000000",
            INIT_29 => X"ffffff73ffffffffffffffc8ffffffff00000001000000000000003e00000000",
            INIT_2A => X"000000c200000000fffffff8ffffffff0000002e00000000ffffff86ffffffff",
            INIT_2B => X"ffffff3bffffffff000000130000000000000081000000000000001e00000000",
            INIT_2C => X"ffffffb9ffffffff00000009000000000000005a000000000000009400000000",
            INIT_2D => X"ffffffdaffffffff0000001f00000000ffffffe5ffffffffffffff57ffffffff",
            INIT_2E => X"ffffffa5ffffffffffffffedfffffffffffffff3ffffffffffffffbeffffffff",
            INIT_2F => X"00000089000000000000003c000000000000000f000000000000000200000000",
            INIT_30 => X"0000001800000000000000370000000000000046000000000000005200000000",
            INIT_31 => X"fffffff8ffffffffffffffe7ffffffffffffffd6ffffffff0000001200000000",
            INIT_32 => X"00000095000000000000005c0000000000000053000000000000006b00000000",
            INIT_33 => X"0000007000000000000000b10000000000000017000000000000006e00000000",
            INIT_34 => X"0000009300000000ffffffa2ffffffffffffff11ffffffffffffffd9ffffffff",
            INIT_35 => X"0000003b00000000fffffffaffffffffffffffcbffffffff0000003c00000000",
            INIT_36 => X"0000004800000000ffffffdcfffffffffffffff5ffffffff0000003d00000000",
            INIT_37 => X"0000001c000000000000001200000000ffffff6effffffff0000001b00000000",
            INIT_38 => X"0000002200000000ffffffe0ffffffff0000003a00000000ffffff67ffffffff",
            INIT_39 => X"00000087000000000000004b000000000000007a00000000ffffffe5ffffffff",
            INIT_3A => X"ffffff6cffffffffffffffedffffffffffffff58ffffffff0000000300000000",
            INIT_3B => X"000000190000000000000023000000000000007a00000000ffffff1fffffffff",
            INIT_3C => X"0000003a00000000ffffffabffffffffffffffbbffffffff0000002100000000",
            INIT_3D => X"0000004a000000000000000d000000000000006d00000000ffffff85ffffffff",
            INIT_3E => X"0000000d000000000000003000000000ffffffd0ffffffff0000009d00000000",
            INIT_3F => X"ffffff64ffffffff00000002000000000000005e000000000000008d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffff0effffffffffffffacffffffffffffffa5fffffffffffffff9ffffffff",
            INIT_41 => X"ffffff33ffffffffffffff71ffffffffffffffe6fffffffffffffef8ffffffff",
            INIT_42 => X"ffffffc0ffffffffffffffcaffffffff0000004100000000ffffffe5ffffffff",
            INIT_43 => X"ffffff8effffffffffffffb5ffffffff0000006d000000000000007300000000",
            INIT_44 => X"0000004c00000000ffffffdcffffffffffffffdcffffffffffffff9effffffff",
            INIT_45 => X"fffffe57ffffffff0000000100000000ffffff3cffffffffffffff58ffffffff",
            INIT_46 => X"ffffff9affffffff0000003c00000000fffffefcffffffffffffff5fffffffff",
            INIT_47 => X"ffffff71ffffffffffffff9fffffffff00000000000000000000000700000000",
            INIT_48 => X"0000002400000000fffffffaffffffffffffff4effffffff000000e000000000",
            INIT_49 => X"ffffffc8ffffffff0000003a000000000000002400000000ffffffaeffffffff",
            INIT_4A => X"00000018000000000000008400000000000000a600000000ffffffaaffffffff",
            INIT_4B => X"ffffff2dfffffffffffffff9ffffffff0000001200000000ffffffd6ffffffff",
            INIT_4C => X"fffffed6ffffffffffffff82ffffffffffffff76fffffffffffffedaffffffff",
            INIT_4D => X"0000000c000000000000001d000000000000000f00000000ffffff72ffffffff",
            INIT_4E => X"0000001200000000000000000000000000000008000000000000000d00000000",
            INIT_4F => X"00000002000000000000005f00000000fffffff3fffffffffffffff8ffffffff",
            INIT_50 => X"ffffffe0fffffffffffffff9fffffffffffffffcffffffff0000004c00000000",
            INIT_51 => X"000000f800000000000000760000000000000092000000000000000700000000",
            INIT_52 => X"0000009900000000ffffffd5fffffffffffffffaffffffff0000002700000000",
            INIT_53 => X"ffffffffffffffffffffff81ffffffffffffff91ffffffffffffffaaffffffff",
            INIT_54 => X"ffffff1bffffffffffffff36ffffffffffffffacffffffffffffffacffffffff",
            INIT_55 => X"ffffffe5ffffffffffffff1effffffff0000002b00000000ffffff8cffffffff",
            INIT_56 => X"0000003e00000000ffffff8effffffffffffffdbfffffffffffffffcffffffff",
            INIT_57 => X"ffffff39ffffffffffffff7cffffffff0000000e00000000ffffffaeffffffff",
            INIT_58 => X"ffffffdbffffffffffffff7dffffffffffffffd8ffffffff0000006400000000",
            INIT_59 => X"ffffffe9ffffffff0000005100000000fffffffaffffffffffffffdcffffffff",
            INIT_5A => X"ffffffa7ffffffff00000018000000000000009700000000ffffff45ffffffff",
            INIT_5B => X"ffffff29ffffffffffffff3cffffffff000000be000000000000002f00000000",
            INIT_5C => X"fffffeffffffffffffffff83ffffffff00000021000000000000006d00000000",
            INIT_5D => X"ffffff9dffffffffffffffa1ffffffffffffffaeffffffffffffffdfffffffff",
            INIT_5E => X"0000000100000000000000bc00000000ffffffe2ffffffffffffff7cffffffff",
            INIT_5F => X"ffffff47ffffffff0000003500000000ffffffa4ffffffff0000001100000000",
            INIT_60 => X"0000005700000000ffffffffffffffff0000002f000000000000002f00000000",
            INIT_61 => X"ffffff1dffffffff000000890000000000000092000000000000003700000000",
            INIT_62 => X"0000008a000000000000003d0000000000000020000000000000006200000000",
            INIT_63 => X"0000000600000000ffffffdcffffffff0000004a000000000000007a00000000",
            INIT_64 => X"0000008700000000fffffffaffffffff00000017000000000000000900000000",
            INIT_65 => X"0000000400000000000000ef00000000ffffff7bffffffffffffffafffffffff",
            INIT_66 => X"ffffffedffffffffffffff7affffffffffffffc2ffffffff0000004c00000000",
            INIT_67 => X"0000000a0000000000000194000000000000001800000000ffffffb9ffffffff",
            INIT_68 => X"ffffff9affffffffffffffd0ffffffffffffff4dffffffff0000001300000000",
            INIT_69 => X"0000003c00000000ffffffe6ffffffff00000076000000000000002800000000",
            INIT_6A => X"000000f800000000ffffffccfffffffffffffff8ffffffff0000002f00000000",
            INIT_6B => X"ffffffd0ffffffffffffff3effffffff0000002f00000000ffffffc5ffffffff",
            INIT_6C => X"ffffffecffffffffffffffe6fffffffffffffed8ffffffffffffff5fffffffff",
            INIT_6D => X"0000006400000000ffffffe1ffffffff00000034000000000000007900000000",
            INIT_6E => X"ffffffbfffffffff00000000000000000000007300000000ffffffbfffffffff",
            INIT_6F => X"ffffff62ffffffff0000000a000000000000006600000000ffffffbeffffffff",
            INIT_70 => X"000000b000000000fffffff3ffffffffffffffefffffffffffffffe0ffffffff",
            INIT_71 => X"00000077000000000000001f000000000000005600000000ffffff83ffffffff",
            INIT_72 => X"ffffffd3ffffffff00000023000000000000000a00000000ffffffb6ffffffff",
            INIT_73 => X"0000000100000000ffffffc2ffffffffffffffb7ffffffffffffffbaffffffff",
            INIT_74 => X"0000005600000000fffffff6fffffffffffffecaffffffff0000009a00000000",
            INIT_75 => X"ffffffb5ffffffff0000008f00000000ffffffdefffffffffffffff9ffffffff",
            INIT_76 => X"fffffff9ffffffffffffff7effffffff0000008900000000ffffff93ffffffff",
            INIT_77 => X"0000008f000000000000001e000000000000008c00000000ffffffcfffffffff",
            INIT_78 => X"0000006400000000fffffeeeffffffff0000000100000000ffffffdcffffffff",
            INIT_79 => X"0000006d000000000000003200000000ffffff9affffffff0000006500000000",
            INIT_7A => X"0000008d00000000ffffffe6ffffffffffffff43ffffffff0000008f00000000",
            INIT_7B => X"00000026000000000000002200000000ffffff97ffffffffffffffccffffffff",
            INIT_7C => X"ffffffd2ffffffff000000190000000000000009000000000000002300000000",
            INIT_7D => X"0000004200000000000000c400000000ffffffd3ffffffff0000000f00000000",
            INIT_7E => X"fffffeecffffffffffffff49ffffffffffffff92ffffffff0000001b00000000",
            INIT_7F => X"000000900000000000000066000000000000007a000000000000004a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE29;


    MEM_IWGHT_LAYER2_INSTANCE30 : if BRAM_NAME = "iwght_layer2_instance30" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffff3cffffffffffffff5effffffffffffff97ffffffffffffffb5ffffffff",
            INIT_01 => X"fffffff9ffffffff000000a5000000000000004c00000000fffffe91ffffffff",
            INIT_02 => X"0000002100000000000000c400000000fffffff9ffffffff0000007f00000000",
            INIT_03 => X"ffffff56ffffffff0000002a00000000ffffffe7ffffffff0000007800000000",
            INIT_04 => X"ffffffc6ffffffffffffff4affffffffffffffe2ffffffffffffffb9ffffffff",
            INIT_05 => X"ffffffbeffffffffffffffdbffffffffffffffb8ffffffffffffffefffffffff",
            INIT_06 => X"00000008000000000000006a00000000000000cf00000000ffffff37ffffffff",
            INIT_07 => X"0000001c0000000000000005000000000000001c00000000ffffff6bffffffff",
            INIT_08 => X"ffffff31ffffffffffffffc4ffffffff0000003400000000000000bc00000000",
            INIT_09 => X"0000006800000000ffffffdbffffffff0000007500000000000000a500000000",
            INIT_0A => X"ffffffdeffffffffffffffdfffffffffffffff6dffffffff0000004800000000",
            INIT_0B => X"0000003900000000fffffffbffffffffffffffa9ffffffff0000007700000000",
            INIT_0C => X"ffffffd3fffffffffffffe92ffffffffffffff8effffffff0000002000000000",
            INIT_0D => X"00000000000000000000002b0000000000000026000000000000000200000000",
            INIT_0E => X"ffffffe0ffffffff000000030000000000000039000000000000009700000000",
            INIT_0F => X"0000001300000000ffffffc4ffffffffffffffa2ffffffffffffffaaffffffff",
            INIT_10 => X"0000007700000000ffffffddffffffff00000016000000000000006b00000000",
            INIT_11 => X"ffffff30ffffffffffffff61ffffffff000000bd000000000000007900000000",
            INIT_12 => X"0000008200000000fffffffdffffffffffffff9dffffffffffffff48ffffffff",
            INIT_13 => X"0000003700000000ffffffd6ffffffffffffff73ffffffffffffffebffffffff",
            INIT_14 => X"ffffffadfffffffffffffff5ffffffff00000092000000000000004e00000000",
            INIT_15 => X"ffffffedffffffff0000000b00000000fffffffbffffffffffffff78ffffffff",
            INIT_16 => X"fffffff6fffffffffffffffdffffffff0000001b000000000000001700000000",
            INIT_17 => X"00000044000000000000000000000000fffffffcffffffff0000000e00000000",
            INIT_18 => X"fffffffcffffffff0000004c00000000ffffff9affffffffffffffe8ffffffff",
            INIT_19 => X"ffffffa6ffffffffffffffa7ffffffff0000003f000000000000003700000000",
            INIT_1A => X"ffffff64ffffffff0000007500000000ffffff8affffffff0000007f00000000",
            INIT_1B => X"0000009a000000000000003300000000fffffffafffffffffffffffbffffffff",
            INIT_1C => X"ffffff72ffffffffffffff3dffffffff0000008a000000000000003e00000000",
            INIT_1D => X"000000550000000000000025000000000000003500000000ffffff5dffffffff",
            INIT_1E => X"0000000c0000000000000040000000000000003b00000000ffffffc5ffffffff",
            INIT_1F => X"0000005e00000000fffffe35ffffffff0000000c00000000fffffecdffffffff",
            INIT_20 => X"ffffffe6fffffffffffffff1ffffffff0000003a00000000ffffff1cffffffff",
            INIT_21 => X"000000630000000000000011000000000000006100000000fffffe93ffffffff",
            INIT_22 => X"0000002100000000000000a800000000ffffff36ffffffffffffff6bffffffff",
            INIT_23 => X"ffffff9bffffffff000000530000000000000006000000000000001800000000",
            INIT_24 => X"0000008e00000000ffffff79ffffffffffffff10ffffffffffffffb2ffffffff",
            INIT_25 => X"00000068000000000000002800000000ffffff22ffffffff0000001a00000000",
            INIT_26 => X"00000016000000000000004900000000ffffff8bffffffffffffffcdffffffff",
            INIT_27 => X"ffffff2effffffffffffff4fffffffffffffff62ffffffff0000006500000000",
            INIT_28 => X"ffffffcbffffffff000000010000000000000059000000000000008800000000",
            INIT_29 => X"ffffffebffffffffffffff73fffffffffffffffbffffffff0000000300000000",
            INIT_2A => X"000000be00000000ffffffacffffffffffffff8effffffff0000000000000000",
            INIT_2B => X"0000009600000000ffffffbcffffffff000000d200000000ffffffdfffffffff",
            INIT_2C => X"ffffff49ffffffffffffff3bffffffff00000080000000000000009e00000000",
            INIT_2D => X"ffffffe3ffffffffffffffaaffffffffffffff6fffffffff0000009900000000",
            INIT_2E => X"ffffffc9ffffffff0000002400000000ffffffa9ffffffff0000011900000000",
            INIT_2F => X"ffffff84ffffffff0000002f0000000000000008000000000000004300000000",
            INIT_30 => X"ffffffb9ffffffffffffff9effffffff0000006f000000000000004e00000000",
            INIT_31 => X"ffffffdbffffffffffffffe0ffffffff0000006e000000000000005d00000000",
            INIT_32 => X"0000002700000000000000d800000000ffffff7effffffffffffff91ffffffff",
            INIT_33 => X"ffffffa2ffffffff000000b7000000000000005000000000fffffffbffffffff",
            INIT_34 => X"ffffff30ffffffffffffff1dfffffffffffffe49ffffffffffffffd8ffffffff",
            INIT_35 => X"0000006900000000ffffff1dffffffffffffffceffffffffffffff93ffffffff",
            INIT_36 => X"ffffff87ffffffff0000001c000000000000009600000000ffffffffffffffff",
            INIT_37 => X"0000000e00000000ffffffccffffffffffffff21ffffffff0000003c00000000",
            INIT_38 => X"0000000c000000000000007c00000000ffffff64ffffffff0000006300000000",
            INIT_39 => X"0000009500000000000000b700000000fffffffaffffffff0000008600000000",
            INIT_3A => X"ffffffb9ffffffff0000007c000000000000005400000000ffffff08ffffffff",
            INIT_3B => X"fffffff5ffffffffffffffc3ffffffffffffffa9ffffffffffffffbdffffffff",
            INIT_3C => X"000000d800000000000000f000000000ffffffb9fffffffffffffff8ffffffff",
            INIT_3D => X"fffffefaffffffffffffff94ffffffffffffff64fffffffffffffeebffffffff",
            INIT_3E => X"0000011000000000ffffffd1ffffffff0000001b00000000ffffffa0ffffffff",
            INIT_3F => X"ffffffc5ffffffffffffff9cffffffff00000005000000000000003100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff9ffffffffffffffe6ffffffff00000000000000000000000700000000",
            INIT_41 => X"fffffff9fffffffffffffff6ffffffff0000000000000000fffffffcffffffff",
            INIT_42 => X"ffffffe7fffffffffffffffeffffffffffffffe8ffffffff0000000300000000",
            INIT_43 => X"0000000b00000000ffffffe9ffffffffffffffe5ffffffffffffffe8ffffffff",
            INIT_44 => X"00000000000000000000000900000000ffffffe7ffffffffffffffecffffffff",
            INIT_45 => X"fffffffcffffffff0000000b000000000000000a00000000fffffff0ffffffff",
            INIT_46 => X"0000000b000000000000000400000000ffffffecffffffff0000000400000000",
            INIT_47 => X"ffffffedffffffffffffffeaffffffff00000003000000000000000e00000000",
            INIT_48 => X"0000000a00000000ffffffefffffffff00000003000000000000000a00000000",
            INIT_49 => X"ffffffe1fffffffffffffff7fffffffffffffffaffffffffffffffe7ffffffff",
            INIT_4A => X"00000005000000000000000200000000fffffffcffffffff0000000000000000",
            INIT_4B => X"ffffffddffffffffffffffe8fffffffffffffffcffffffffffffffe9ffffffff",
            INIT_4C => X"fffffffcffffffff0000000500000000ffffffedffffffff0000001600000000",
            INIT_4D => X"fffffff0ffffffffffffffe3ffffffff00000003000000000000000a00000000",
            INIT_4E => X"ffffffe5fffffffffffffffbffffffffffffffedffffffffffffffeeffffffff",
            INIT_4F => X"fffffffbfffffffffffffff5ffffffff0000000200000000ffffffe0ffffffff",
            INIT_50 => X"ffffffe4ffffffffffffffdfffffffffffffffebffffffff0000000700000000",
            INIT_51 => X"fffffff1fffffffffffffff7ffffffff0000000000000000fffffffbffffffff",
            INIT_52 => X"fffffff1ffffffffffffffd9ffffffffffffffffffffffffffffffdeffffffff",
            INIT_53 => X"fffffffcffffffffffffffe0ffffffffffffffe2ffffffffffffffdeffffffff",
            INIT_54 => X"0000000500000000ffffffefffffffff0000000f00000000ffffffecffffffff",
            INIT_55 => X"fffffff3ffffffff00000000000000000000000000000000ffffffeeffffffff",
            INIT_56 => X"fffffff5ffffffff0000000d00000000fffffff8ffffffffffffffebffffffff",
            INIT_57 => X"0000000300000000fffffff4ffffffffffffffedffffffffffffffe8ffffffff",
            INIT_58 => X"fffffffdfffffffffffffff2ffffffff0000000000000000ffffffe0ffffffff",
            INIT_59 => X"000000020000000000000009000000000000000300000000ffffffeeffffffff",
            INIT_5A => X"0000000500000000fffffffefffffffffffffffffffffffffffffff1ffffffff",
            INIT_5B => X"ffffffffffffffff0000000900000000fffffff3ffffffffffffffefffffffff",
            INIT_5C => X"ffffffe6fffffffffffffff7ffffffff0000000500000000fffffff8ffffffff",
            INIT_5D => X"ffffffebfffffffffffffff4ffffffff00000008000000000000000700000000",
            INIT_5E => X"0000000300000000ffffffeeffffffff0000000000000000fffffffbffffffff",
            INIT_5F => X"ffffffedffffffffffffffdfffffffff0000000000000000ffffffecffffffff",
            INIT_60 => X"fffffff9fffffffffffffffeffffffffffffffe9ffffffff0000000100000000",
            INIT_61 => X"ffffffe3ffffffffffffffdeffffffff0000000800000000fffffff7ffffffff",
            INIT_62 => X"fffffffafffffffffffffff0fffffffffffffffcffffffffffffffe8ffffffff",
            INIT_63 => X"0000000800000000fffffff4ffffffff0000000000000000ffffffebffffffff",
            INIT_64 => X"ffffffe9ffffffffffffffeffffffffffffffff7ffffffff0000000000000000",
            INIT_65 => X"fffffffbffffffffffffffe9fffffffffffffff9ffffffff0000000600000000",
            INIT_66 => X"0000000800000000ffffffefffffffff0000001100000000fffffffcffffffff",
            INIT_67 => X"0000000700000000000000060000000000000006000000000000001300000000",
            INIT_68 => X"000000030000000000000008000000000000000500000000ffffffffffffffff",
            INIT_69 => X"fffffff5ffffffffffffffe7ffffffff0000000600000000fffffff1ffffffff",
            INIT_6A => X"fffffffafffffffffffffffbfffffffffffffff3ffffffffffffffefffffffff",
            INIT_6B => X"fffffff2fffffffffffffffbffffffffffffffdffffffffffffffff5ffffffff",
            INIT_6C => X"0000000400000000fffffffcffffffffffffffe8fffffffffffffffcffffffff",
            INIT_6D => X"fffffffffffffffffffffff7fffffffffffffff3ffffffffffffffe3ffffffff",
            INIT_6E => X"00000013000000000000000f000000000000000300000000ffffffefffffffff",
            INIT_6F => X"ffffffeefffffffffffffff4fffffffffffffffeffffffffffffffefffffffff",
            INIT_70 => X"ffffffdbffffffffffffffecfffffffffffffff7ffffffffffffffe1ffffffff",
            INIT_71 => X"ffffffe6fffffffffffffff0fffffffffffffff9ffffffffffffffffffffffff",
            INIT_72 => X"ffffffebffffffffffffffebffffffffffffffeaffffffffffffffe7ffffffff",
            INIT_73 => X"ffffffdbfffffffffffffff8ffffffff0000000d000000000000000b00000000",
            INIT_74 => X"ffffffedffffffff0000001400000000ffffffe0ffffffffffffffe0ffffffff",
            INIT_75 => X"ffffffe9fffffffffffffff1fffffffffffffff2fffffffffffffffbffffffff",
            INIT_76 => X"ffffffe2fffffffffffffffcfffffffffffffffafffffffffffffff1ffffffff",
            INIT_77 => X"fffffff5ffffffffffffffe9ffffffffffffffe4ffffffffffffffe1ffffffff",
            INIT_78 => X"0000000600000000fffffffdfffffffffffffffbffffffffffffffe5ffffffff",
            INIT_79 => X"fffffffdffffffff000000100000000000000007000000000000000300000000",
            INIT_7A => X"ffffffeaffffffffffffffffffffffff0000001000000000fffffff1ffffffff",
            INIT_7B => X"0000000a00000000fffffffeffffffff0000000c00000000fffffffdffffffff",
            INIT_7C => X"ffffffeffffffffffffffffdffffffffffffffebfffffffffffffff5ffffffff",
            INIT_7D => X"0000000200000000fffffffbffffffffffffffffffffffffffffffe4ffffffff",
            INIT_7E => X"fffffffeffffffffffffffffffffffffffffffefffffffffffffffe7ffffffff",
            INIT_7F => X"0000000c00000000fffffffbffffffff0000000000000000ffffffefffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE30;


    MEM_IWGHT_LAYER2_INSTANCE31 : if BRAM_NAME = "iwght_layer2_instance31" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000003000000000000000800000000fffffffaffffffffffffffe3ffffffff",
            INIT_01 => X"fffffff8fffffffffffffffbffffffffffffffeeffffffff0000000500000000",
            INIT_02 => X"0000000500000000fffffffffffffffffffffff2ffffffff0000000200000000",
            INIT_03 => X"fffffff0ffffffff00000006000000000000000300000000fffffff5ffffffff",
            INIT_04 => X"0000000400000000fffffff3ffffffff0000000400000000fffffffcffffffff",
            INIT_05 => X"00000000000000000000000900000000ffffffeefffffffffffffffeffffffff",
            INIT_06 => X"fffffff7ffffffff000000030000000000000009000000000000000000000000",
            INIT_07 => X"0000000300000000ffffffd5fffffffffffffffdffffffffffffffeaffffffff",
            INIT_08 => X"fffffff3ffffffffffffffc4ffffffffffffff8affffffffffffffd0ffffffff",
            INIT_09 => X"ffffff62ffffffffffffffc0ffffffffffffffdefffffffffffffe73ffffffff",
            INIT_0A => X"0000002f00000000ffffffcafffffffffffffeccffffffffffffffc5ffffffff",
            INIT_0B => X"ffffff91ffffffff0000008500000000ffffff9bffffffff0000008d00000000",
            INIT_0C => X"0000005000000000ffffff4effffffff00000029000000000000008500000000",
            INIT_0D => X"ffffffe0ffffffffffffffedffffffff0000001700000000ffffffc3ffffffff",
            INIT_0E => X"ffffff82ffffffff00000056000000000000006500000000ffffff7affffffff",
            INIT_0F => X"ffffffbaffffffff0000002200000000ffffff33fffffffffffffff9ffffffff",
            INIT_10 => X"ffffffc7ffffffff0000000100000000000000b400000000ffffff9effffffff",
            INIT_11 => X"00000007000000000000005400000000ffffff26ffffffffffffff63ffffffff",
            INIT_12 => X"fffffe73ffffffff0000009300000000ffffffc6ffffffff0000009e00000000",
            INIT_13 => X"ffffffa2ffffffffffffffe1ffffffffffffff0efffffffffffffff9ffffffff",
            INIT_14 => X"ffffff53ffffffffffffffecfffffffffffffff6fffffffffffffe34ffffffff",
            INIT_15 => X"000000f800000000ffffff13ffffffffffffff87ffffffff0000006600000000",
            INIT_16 => X"ffffffdbffffffffffffffd7ffffffffffffff92ffffffffffffffedffffffff",
            INIT_17 => X"ffffff29ffffffff0000001800000000ffffffa7ffffffff000000c200000000",
            INIT_18 => X"fffffe03ffffffffffffffd8ffffffffffffffeeffffffff0000001c00000000",
            INIT_19 => X"0000007c00000000ffffff66fffffffffffffee4fffffffffffffef2ffffffff",
            INIT_1A => X"0000001000000000ffffffe2ffffffffffffffeafffffffffffffedbffffffff",
            INIT_1B => X"ffffffe7ffffffffffffffcdffffffffffffffcbfffffffffffffefbffffffff",
            INIT_1C => X"0000001800000000ffffffe1ffffffffffffff79ffffffff0000006700000000",
            INIT_1D => X"000000ae00000000ffffffb5ffffffffffffffc2ffffffff000000ae00000000",
            INIT_1E => X"ffffff85ffffffffffffff8effffffff0000000000000000000000c200000000",
            INIT_1F => X"ffffffadffffffffffffff82ffffffff0000009c000000000000004500000000",
            INIT_20 => X"ffffffb5ffffffffffffff6bffffffffffffff8fffffffff0000005800000000",
            INIT_21 => X"0000001000000000ffffffa2ffffffff0000002f000000000000007a00000000",
            INIT_22 => X"ffffffbbfffffffffffffffcffffffffffffff9bffffffff0000001400000000",
            INIT_23 => X"000000df00000000ffffff55fffffffffffffffcffffffffffffff91ffffffff",
            INIT_24 => X"fffffe91ffffffff0000004300000000fffffff2ffffffff000000c400000000",
            INIT_25 => X"fffffffeffffffff0000000c0000000000000008000000000000001200000000",
            INIT_26 => X"fffffff5fffffffffffffffdffffffff0000000f00000000ffffffefffffffff",
            INIT_27 => X"ffffffadffffffffffffffacffffffff0000000800000000fffffffaffffffff",
            INIT_28 => X"000000520000000000000049000000000000000000000000000000c500000000",
            INIT_29 => X"0000006500000000ffffffd7ffffffffffffffadffffffffffffff8fffffffff",
            INIT_2A => X"ffffffc2ffffffff0000008f00000000ffffffb3ffffffff0000008200000000",
            INIT_2B => X"000000960000000000000035000000000000005e00000000ffffffa3ffffffff",
            INIT_2C => X"0000001f00000000000000000000000000000028000000000000006300000000",
            INIT_2D => X"fffffff1ffffffff0000002500000000ffffffc1fffffffffffffe94ffffffff",
            INIT_2E => X"ffffff3cffffffff00000060000000000000001400000000ffffff25ffffffff",
            INIT_2F => X"0000003b00000000ffffffe5ffffffff000000b9000000000000005f00000000",
            INIT_30 => X"0000003d000000000000002300000000000000f2000000000000002e00000000",
            INIT_31 => X"0000000600000000ffffffecffffffffffffff51ffffffffffffffdaffffffff",
            INIT_32 => X"ffffffa5ffffffff000000de000000000000002f000000000000002800000000",
            INIT_33 => X"0000007400000000ffffff87fffffffffffffffaffffffffffffff9affffffff",
            INIT_34 => X"0000004400000000ffffff8effffffff0000000f000000000000003300000000",
            INIT_35 => X"fffffffeffffffff0000006800000000fffffffcfffffffffffffe86ffffffff",
            INIT_36 => X"0000001a00000000fffffff2ffffffffffffffe4ffffffffffffffa3ffffffff",
            INIT_37 => X"0000006100000000fffffffdffffffff000000a500000000fffffff6ffffffff",
            INIT_38 => X"0000001b00000000ffffffc2ffffffff0000008100000000ffffffb0ffffffff",
            INIT_39 => X"ffffff8dffffffffffffff85ffffffffffffff5cffffffffffffffeaffffffff",
            INIT_3A => X"0000005600000000ffffffefffffffff0000009b00000000ffffffe1ffffffff",
            INIT_3B => X"0000003200000000000000c5000000000000002800000000000000eb00000000",
            INIT_3C => X"ffffffe1ffffffff0000003300000000000000a400000000ffffff51ffffffff",
            INIT_3D => X"0000002700000000ffffffdaffffffff0000004c00000000ffffffeeffffffff",
            INIT_3E => X"000000bc000000000000003a000000000000004300000000ffffffafffffffff",
            INIT_3F => X"0000002e00000000fffffec4ffffffff00000080000000000000004700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000021000000000000006400000000ffffff7dffffffff0000008900000000",
            INIT_41 => X"ffffff9fffffffffffffffe8ffffffff0000003900000000ffffff46ffffffff",
            INIT_42 => X"00000038000000000000008100000000ffffffdbffffffffffffffb9ffffffff",
            INIT_43 => X"ffffff77ffffffffffffffecffffffff00000021000000000000007700000000",
            INIT_44 => X"ffffffdaffffffff0000000f00000000fffffffcffffffff0000005000000000",
            INIT_45 => X"0000004400000000fffffec7ffffffff0000003400000000ffffffaeffffffff",
            INIT_46 => X"fffffff1ffffffffffffffd0ffffffff0000001f00000000ffffff32ffffffff",
            INIT_47 => X"0000004b000000000000001700000000ffffffd0ffffffff000000ce00000000",
            INIT_48 => X"ffffffcbffffffff0000002100000000fffffe35ffffffff000000a200000000",
            INIT_49 => X"fffffffbffffffff0000001e00000000ffffffcaffffffff0000005f00000000",
            INIT_4A => X"fffffef7ffffffff000000d800000000ffffff5bffffffffffffff5bffffffff",
            INIT_4B => X"00000040000000000000002300000000fffffffcffffffffffffffb1ffffffff",
            INIT_4C => X"00000016000000000000013a00000000ffffff07ffffffffffffff25ffffffff",
            INIT_4D => X"0000002c00000000ffffffcaffffffff000000a600000000ffffffdfffffffff",
            INIT_4E => X"ffffff64ffffffff0000009f000000000000007a000000000000007f00000000",
            INIT_4F => X"ffffffe1ffffffffffffffa5ffffffffffffffb8ffffffff0000004d00000000",
            INIT_50 => X"ffffff68fffffffffffffff9ffffffffffffffbfffffffffffffff3bffffffff",
            INIT_51 => X"ffffffe2ffffffff0000003c000000000000004100000000ffffff53ffffffff",
            INIT_52 => X"0000005b000000000000008000000000000000b900000000ffffff8fffffffff",
            INIT_53 => X"ffffffdeffffffff0000001600000000000000b500000000ffffffb3ffffffff",
            INIT_54 => X"0000002500000000ffffff7effffffffffffffbcffffffff0000008000000000",
            INIT_55 => X"ffffff6dffffffffffffffe4ffffffff0000001e000000000000000e00000000",
            INIT_56 => X"fffffe2affffffffffffff9affffffffffffff33ffffffffffffff9effffffff",
            INIT_57 => X"0000004b00000000ffffff48fffffffffffffff6fffffffffffffef6ffffffff",
            INIT_58 => X"ffffff98ffffffffffffffd2ffffffffffffffe9ffffffffffffff57ffffffff",
            INIT_59 => X"ffffffe1ffffffffffffffaaffffffffffffff57ffffffffffffffe9ffffffff",
            INIT_5A => X"0000004700000000ffffffdafffffffffffffe3bfffffffffffffe4effffffff",
            INIT_5B => X"0000007300000000000000a500000000ffffffc8ffffffff0000000000000000",
            INIT_5C => X"00000047000000000000006700000000ffffffbdffffffffffffffc2ffffffff",
            INIT_5D => X"ffffffd7ffffffff0000000a00000000ffffffd5ffffffff0000001300000000",
            INIT_5E => X"00000038000000000000007c00000000fffffff1ffffffff000000af00000000",
            INIT_5F => X"0000002e00000000ffffffb1ffffffff0000006400000000ffffffd5ffffffff",
            INIT_60 => X"ffffffa2ffffffff0000002e00000000ffffffcaffffffff0000005c00000000",
            INIT_61 => X"ffffff94ffffffffffffff19ffffffffffffff80ffffffffffffff7fffffffff",
            INIT_62 => X"0000003f000000000000001800000000ffffffccffffffff0000009800000000",
            INIT_63 => X"ffffffefffffffffffffff79ffffffffffffffa7ffffffff0000004d00000000",
            INIT_64 => X"0000005200000000ffffff8cffffffff00000012000000000000005500000000",
            INIT_65 => X"0000004c000000000000003c00000000ffffff82ffffffff0000002e00000000",
            INIT_66 => X"ffffff52ffffffff00000001000000000000004500000000ffffff47ffffffff",
            INIT_67 => X"ffffffd4ffffffff00000048000000000000004100000000ffffffdcffffffff",
            INIT_68 => X"0000001500000000fffffffaffffffff0000006e00000000ffffffb5ffffffff",
            INIT_69 => X"000000bb00000000ffffff71ffffffffffffff4fffffffff0000001f00000000",
            INIT_6A => X"ffffff13ffffffff0000001400000000ffffff82ffffffff0000001e00000000",
            INIT_6B => X"ffffffeefffffffffffffe67ffffffffffffff64ffffffffffffffdeffffffff",
            INIT_6C => X"00000070000000000000003500000000ffffff2bffffffffffffff2fffffffff",
            INIT_6D => X"fffffff8fffffffffffffffdfffffffffffffff4ffffffff000000cc00000000",
            INIT_6E => X"fffffff5fffffffffffffffafffffffffffffff9ffffffffffffffecffffffff",
            INIT_6F => X"ffffff64ffffffff000000b000000000fffffff7ffffffff0000001500000000",
            INIT_70 => X"0000009000000000ffffff43ffffffffffffffa7ffffffffffffffb1ffffffff",
            INIT_71 => X"0000002800000000ffffff78ffffffff0000004500000000fffffff0ffffffff",
            INIT_72 => X"0000004f00000000ffffffcdffffffffffffff2dfffffffffffffef7ffffffff",
            INIT_73 => X"0000002e00000000fffffeceffffffffffffffd9ffffffffffffffbcffffffff",
            INIT_74 => X"ffffffe1ffffffff0000001c00000000fffffffaffffffff0000002600000000",
            INIT_75 => X"ffffff0bffffffff0000005a00000000ffffffcbffffffff0000005100000000",
            INIT_76 => X"0000000e000000000000003100000000ffffff38ffffffffffffffa8ffffffff",
            INIT_77 => X"ffffffccffffffff000000a700000000000000ab00000000ffffffdeffffffff",
            INIT_78 => X"0000000a00000000ffffffc4fffffffffffffff5ffffffffffffffceffffffff",
            INIT_79 => X"ffffff4effffffff000000c7000000000000000200000000ffffff1cffffffff",
            INIT_7A => X"0000001500000000fffffefbffffffff0000002e000000000000000000000000",
            INIT_7B => X"000000b800000000ffffffa4ffffffffffffffe6ffffffff0000007200000000",
            INIT_7C => X"0000002b0000000000000021000000000000001d000000000000003d00000000",
            INIT_7D => X"ffffffa6ffffffff0000007c00000000ffffff9effffffffffffffeeffffffff",
            INIT_7E => X"ffffff8dffffffff000000fa000000000000003c00000000000000d100000000",
            INIT_7F => X"0000006300000000ffffff8bffffffff00000029000000000000009100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE31;


    MEM_IWGHT_LAYER2_INSTANCE32 : if BRAM_NAME = "iwght_layer2_instance32" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004400000000ffffff68ffffffff0000004f000000000000001400000000",
            INIT_01 => X"000000d800000000ffffff32ffffffffffffff6cffffffff000000e000000000",
            INIT_02 => X"000000c700000000ffffff90ffffffff00000092000000000000007700000000",
            INIT_03 => X"00000031000000000000001200000000000000af000000000000005a00000000",
            INIT_04 => X"ffffff68ffffffff000000dd0000000000000002000000000000004200000000",
            INIT_05 => X"fffffee1fffffffffffffffdffffffff0000000a00000000fffffffcffffffff",
            INIT_06 => X"0000001900000000ffffffecffffffffffffff18ffffffffffffff9effffffff",
            INIT_07 => X"ffffff8fffffffff0000004700000000ffffff60ffffffff0000000e00000000",
            INIT_08 => X"00000035000000000000003b00000000fffffec3ffffffffffffff34ffffffff",
            INIT_09 => X"fffffdeeffffffff000000bb000000000000000d00000000ffffffbdffffffff",
            INIT_0A => X"0000005600000000fffffefdffffffffffffffdaffffffffffffff31ffffffff",
            INIT_0B => X"0000006500000000ffffffadffffffffffffffdcffffffff0000009800000000",
            INIT_0C => X"0000005f000000000000003800000000ffffffbdffffffff000000f100000000",
            INIT_0D => X"00000055000000000000004b00000000fffffef7ffffffff0000003500000000",
            INIT_0E => X"ffffffc6ffffffffffffff59fffffffffffffff9ffffffff0000005a00000000",
            INIT_0F => X"000000ff000000000000002500000000ffffffe9ffffffffffffff9affffffff",
            INIT_10 => X"ffffffdfffffffff000000ba000000000000000300000000ffffffc8ffffffff",
            INIT_11 => X"0000001e0000000000000052000000000000007700000000ffffff9fffffffff",
            INIT_12 => X"0000003100000000000000a800000000ffffffbbffffffffffffffefffffffff",
            INIT_13 => X"000000e500000000fffffff4ffffffff000000cc000000000000007500000000",
            INIT_14 => X"000000c900000000fffffff6ffffffff00000050000000000000005000000000",
            INIT_15 => X"ffffffd3ffffffffffffffe2ffffffff0000009000000000ffffffa3ffffffff",
            INIT_16 => X"ffffffe2ffffffff0000001e00000000ffffffcdffffffff0000003600000000",
            INIT_17 => X"0000002c00000000ffffffafffffffffffffffdfffffffffffffffbeffffffff",
            INIT_18 => X"ffffffbaffffffff00000036000000000000000b000000000000001700000000",
            INIT_19 => X"0000003600000000ffffffedffffffffffffffb1ffffffffffffffb5ffffffff",
            INIT_1A => X"ffffff22ffffffff0000009800000000fffffef3ffffffff0000005800000000",
            INIT_1B => X"0000002d000000000000001500000000000000dd00000000ffffffbcffffffff",
            INIT_1C => X"ffffffa0ffffffff000000010000000000000026000000000000005000000000",
            INIT_1D => X"fffffff7fffffffffffffffefffffffffffffff7ffffffffffffffffffffffff",
            INIT_1E => X"ffffffe9ffffffff0000003e000000000000008700000000fffffee3ffffffff",
            INIT_1F => X"ffffff38ffffffff0000009b000000000000001500000000ffffff25ffffffff",
            INIT_20 => X"000000100000000000000032000000000000007e00000000ffffffdeffffffff",
            INIT_21 => X"0000001900000000ffffff35ffffffffffffffc7ffffffff0000007e00000000",
            INIT_22 => X"ffffff21ffffffff000000e200000000ffffff72ffffffffffffffc3ffffffff",
            INIT_23 => X"ffffffccffffffff000000920000000000000056000000000000000700000000",
            INIT_24 => X"00000014000000000000002600000000ffffffbcffffffffffffff7affffffff",
            INIT_25 => X"000000ca00000000fffffff3ffffffff00000030000000000000000000000000",
            INIT_26 => X"0000002f00000000000000a000000000ffffffd8ffffffff0000001600000000",
            INIT_27 => X"0000001c000000000000001a00000000ffffff91ffffffff0000002900000000",
            INIT_28 => X"00000039000000000000000000000000ffffff98ffffffff000000b900000000",
            INIT_29 => X"ffffff98fffffffffffffeb3ffffffffffffffbfffffffff0000004d00000000",
            INIT_2A => X"ffffff59ffffffff00000062000000000000002800000000ffffff2effffffff",
            INIT_2B => X"0000003100000000fffffeecffffffffffffffd3ffffffff0000002400000000",
            INIT_2C => X"ffffff79ffffffff0000001f000000000000009d000000000000004200000000",
            INIT_2D => X"00000050000000000000002b00000000ffffffc7ffffffff000000b100000000",
            INIT_2E => X"ffffff84ffffffff0000004700000000ffffff4fffffffff000000a700000000",
            INIT_2F => X"000000de00000000ffffffd5ffffffffffffff60ffffffff0000004c00000000",
            INIT_30 => X"ffffffeaffffffff000000ab00000000ffffffe4ffffffffffffff62ffffffff",
            INIT_31 => X"0000000900000000000000a5000000000000009f000000000000004300000000",
            INIT_32 => X"0000002e00000000ffffff70ffffffffffffff3dffffffffffffffbdffffffff",
            INIT_33 => X"ffffff0effffffff000000f300000000fffffff2ffffffffffffffbeffffffff",
            INIT_34 => X"000000b400000000ffffff60ffffffff00000032000000000000000400000000",
            INIT_35 => X"0000000a00000000fffffff8fffffffffffffffdffffffffffffff81ffffffff",
            INIT_36 => X"fffffff7fffffffffffffff4fffffffffffffff3ffffffff0000000800000000",
            INIT_37 => X"ffffffd2ffffffff00000005000000000000001500000000fffffff8ffffffff",
            INIT_38 => X"ffffff74ffffffffffffffa6ffffffff0000007800000000ffffff3dffffffff",
            INIT_39 => X"ffffffe7ffffffff0000000300000000ffffffefffffffff0000013300000000",
            INIT_3A => X"0000005200000000ffffffdaffffffffffffff10ffffffffffffff56ffffffff",
            INIT_3B => X"000000dc000000000000008a000000000000001200000000ffffffa7ffffffff",
            INIT_3C => X"fffffff8ffffffff0000003900000000ffffffe6ffffffffffffffd8ffffffff",
            INIT_3D => X"ffffff87ffffffffffffffcdffffffff0000008f000000000000003c00000000",
            INIT_3E => X"ffffffd2ffffffffffffffffffffffff0000001f000000000000005e00000000",
            INIT_3F => X"00000136000000000000002a00000000ffffffd9ffffffffffffffd5ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ba000000000000006200000000000000ae00000000ffffff89ffffffff",
            INIT_41 => X"ffffff93ffffffffffffff9bffffffffffffffd0ffffffffffffffbcffffffff",
            INIT_42 => X"ffffffe8ffffffffffffffe7ffffffff0000000800000000ffffff72ffffffff",
            INIT_43 => X"0000005e00000000fffffffdffffffff0000004e00000000ffffffcfffffffff",
            INIT_44 => X"0000005800000000000000fa00000000ffffff91ffffffff0000003700000000",
            INIT_45 => X"ffffffefffffffff000000bc00000000ffffffb7ffffffffffffff52ffffffff",
            INIT_46 => X"ffffff67ffffffff00000046000000000000006b000000000000005b00000000",
            INIT_47 => X"0000008c00000000ffffffa7fffffffffffffe57ffffffff0000006700000000",
            INIT_48 => X"0000001000000000ffffffdfffffffff0000000a00000000ffffffd8ffffffff",
            INIT_49 => X"000000380000000000000034000000000000006900000000000000cf00000000",
            INIT_4A => X"00000000000000000000000d00000000ffffffc5ffffffffffffff14ffffffff",
            INIT_4B => X"00000055000000000000007b000000000000003c000000000000007c00000000",
            INIT_4C => X"ffffff52ffffffff0000004000000000ffffffdbffffffffffffffb4ffffffff",
            INIT_4D => X"00000013000000000000008e000000000000003600000000ffffffdcffffffff",
            INIT_4E => X"00000050000000000000003100000000fffffff7ffffffffffffff9cffffffff",
            INIT_4F => X"fffffff8ffffffffffffffa8ffffffff0000008d00000000ffffff5cffffffff",
            INIT_50 => X"fffffffaffffffff0000006d00000000ffffff5ffffffffffffffff8ffffffff",
            INIT_51 => X"ffffffa1ffffffffffffffcfffffffff00000034000000000000002f00000000",
            INIT_52 => X"000000f300000000ffffff44ffffffffffffff3dffffffff000000a600000000",
            INIT_53 => X"ffffffc6ffffffff0000006e00000000ffffff72ffffffff0000006f00000000",
            INIT_54 => X"ffffff5cffffffff0000001a000000000000006f000000000000001c00000000",
            INIT_55 => X"ffffffdcfffffffffffffffdffffffff000000a800000000ffffffe0ffffffff",
            INIT_56 => X"000000c200000000ffffff0bffffffff0000004c000000000000009600000000",
            INIT_57 => X"fffffeb5ffffffff0000005500000000fffffff9ffffffffffffff4affffffff",
            INIT_58 => X"000000e600000000ffffff93ffffffff000000f000000000ffffff35ffffffff",
            INIT_59 => X"fffffff6ffffffff0000007600000000ffffffa6ffffffff0000006200000000",
            INIT_5A => X"fffffef6ffffffffffffff5dffffffffffffffdaffffffffffffffa3ffffffff",
            INIT_5B => X"ffffff94ffffffffffffffc5ffffffff00000000000000000000003600000000",
            INIT_5C => X"ffffff8dffffffff000000c900000000ffffff72ffffffff0000005000000000",
            INIT_5D => X"00000009000000000000001200000000ffffff89ffffffffffffff61ffffffff",
            INIT_5E => X"00000032000000000000002300000000ffffff1dffffffffffffff8dffffffff",
            INIT_5F => X"ffffff87ffffffff0000001a00000000ffffffebffffffffffffff92ffffffff",
            INIT_60 => X"0000008800000000ffffffabffffffff00000024000000000000004600000000",
            INIT_61 => X"ffffffedffffffff0000005300000000ffffffceffffffffffffffd7ffffffff",
            INIT_62 => X"ffffffcfffffffff00000026000000000000001c00000000ffffffe9ffffffff",
            INIT_63 => X"000000e500000000ffffffa3ffffffffffffffe7ffffffff0000002700000000",
            INIT_64 => X"ffffffcfffffffffffffffacffffffffffffff88ffffffff0000007900000000",
            INIT_65 => X"ffffffa9ffffffff0000004600000000000000ff000000000000002900000000",
            INIT_66 => X"ffffff36ffffffff0000007400000000ffffff92ffffffff0000007b00000000",
            INIT_67 => X"ffffff4bfffffffffffffff4ffffffff0000009900000000ffffff74ffffffff",
            INIT_68 => X"000000270000000000000097000000000000000c000000000000001200000000",
            INIT_69 => X"ffffff70fffffffffffffeb7ffffffffffffffccffffffffffffff7affffffff",
            INIT_6A => X"fffffe42ffffffffffffff40ffffffffffffffe0ffffffffffffff8bffffffff",
            INIT_6B => X"fffffff2ffffffffffffff91ffffffff0000001600000000fffffed8ffffffff",
            INIT_6C => X"fffffff3ffffffffffffff71ffffffffffffff7bffffffff0000005900000000",
            INIT_6D => X"0000004100000000ffffffb2ffffffff0000001600000000ffffffb3ffffffff",
            INIT_6E => X"ffffffa6ffffffff0000008400000000ffffffcdffffffff0000006e00000000",
            INIT_6F => X"ffffffa8ffffffffffffffd0ffffffff0000005c000000000000004c00000000",
            INIT_70 => X"0000006f00000000000000220000000000000000000000000000001800000000",
            INIT_71 => X"0000007a000000000000001c0000000000000040000000000000001300000000",
            INIT_72 => X"ffffff6affffffff0000003d00000000ffffff74ffffffff0000007200000000",
            INIT_73 => X"ffffff41ffffffffffffff84ffffffff00000023000000000000004200000000",
            INIT_74 => X"fffffff9ffffffff0000001b00000000000000ab000000000000006000000000",
            INIT_75 => X"ffffff83ffffffffffffffa7ffffffff00000009000000000000008400000000",
            INIT_76 => X"0000000700000000ffffffe9fffffffffffffcfaffffffffffffff8dffffffff",
            INIT_77 => X"ffffffd0ffffffff00000119000000000000002700000000ffffff7affffffff",
            INIT_78 => X"0000004300000000ffffffd6ffffffffffffff06ffffffff0000007700000000",
            INIT_79 => X"ffffff4affffffff00000034000000000000004400000000ffffffceffffffff",
            INIT_7A => X"ffffff6bffffffff0000003e000000000000006600000000ffffff72ffffffff",
            INIT_7B => X"000000e000000000000000bf00000000ffffffb8ffffffffffffff7dffffffff",
            INIT_7C => X"0000003d0000000000000023000000000000009200000000000000a800000000",
            INIT_7D => X"00000013000000000000001600000000fffffff0ffffffffffffff7affffffff",
            INIT_7E => X"fffffffaffffffff00000000000000000000001000000000fffffff0ffffffff",
            INIT_7F => X"0000003b00000000fffffff3ffffffffffffffebffffffffffffffeaffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE32;


    MEM_IWGHT_LAYER2_INSTANCE33 : if BRAM_NAME = "iwght_layer2_instance33" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffeeffffffffffffff96ffffffff0000002800000000ffffffd5ffffffff",
            INIT_01 => X"0000002f000000000000004f0000000000000042000000000000003100000000",
            INIT_02 => X"ffffffe2ffffffff00000023000000000000000000000000ffffff7dffffffff",
            INIT_03 => X"ffffffa0ffffffff0000003e00000000000000ea000000000000002900000000",
            INIT_04 => X"0000007200000000fffffef3ffffffff00000005000000000000000000000000",
            INIT_05 => X"fffffff0ffffffff0000008c000000000000002800000000ffffffddffffffff",
            INIT_06 => X"ffffffdaffffffff0000005200000000fffffff1ffffffff0000007600000000",
            INIT_07 => X"ffffffd4ffffffff000000e0000000000000007600000000ffffffceffffffff",
            INIT_08 => X"ffffff6bffffffffffffff41ffffffff0000003500000000ffffff28ffffffff",
            INIT_09 => X"0000002a00000000fffffff5ffffffffffffffafffffffff0000008600000000",
            INIT_0A => X"ffffff78ffffffff0000000e00000000fffffff5ffffffff0000001f00000000",
            INIT_0B => X"000000f500000000ffffff48ffffffff0000000f00000000ffffff3affffffff",
            INIT_0C => X"ffffff9cffffffff0000008c0000000000000033000000000000008100000000",
            INIT_0D => X"000000470000000000000037000000000000001900000000000000ab00000000",
            INIT_0E => X"000000aa000000000000000000000000ffffffa1ffffffffffffff30ffffffff",
            INIT_0F => X"fffffff3ffffffff0000017400000000ffffff98ffffffff0000000900000000",
            INIT_10 => X"0000013700000000ffffffc7ffffffff00000014000000000000003600000000",
            INIT_11 => X"00000007000000000000000300000000fffffd29ffffffffffffff8fffffffff",
            INIT_12 => X"ffffffd3ffffffff0000001b00000000ffffffbfffffffff0000003800000000",
            INIT_13 => X"ffffffdbffffffffffffff97ffffffffffffff45ffffffff0000003200000000",
            INIT_14 => X"ffffffc8fffffffffffffff0ffffffff0000008e00000000fffffff0ffffffff",
            INIT_15 => X"00000033000000000000005e00000000ffffffbaffffffffffffffc0ffffffff",
            INIT_16 => X"ffffff2bffffffff0000000e00000000000000e100000000ffffff27ffffffff",
            INIT_17 => X"0000002700000000ffffff63fffffffffffffffeffffffff0000009d00000000",
            INIT_18 => X"0000008d0000000000000004000000000000000400000000ffffffafffffffff",
            INIT_19 => X"ffffffc4ffffffffffffffcaffffffff00000029000000000000000900000000",
            INIT_1A => X"ffffffccfffffffffffffff7ffffffffffffffc1ffffffffffffffffffffffff",
            INIT_1B => X"0000003a000000000000003a000000000000008f000000000000005800000000",
            INIT_1C => X"000000b00000000000000082000000000000005200000000ffffffd1ffffffff",
            INIT_1D => X"0000000e000000000000008b0000000000000096000000000000004000000000",
            INIT_1E => X"ffffffc1fffffffffffffffdffffffffffffff8effffffff0000005b00000000",
            INIT_1F => X"0000005300000000ffffffa0ffffffff0000009f00000000ffffff82ffffffff",
            INIT_20 => X"ffffffdafffffffffffffe8cffffffffffffff19fffffffffffffd34ffffffff",
            INIT_21 => X"0000002800000000ffffff82ffffffff0000007700000000fffffdd1ffffffff",
            INIT_22 => X"0000004a000000000000003400000000ffffff56ffffffff0000000a00000000",
            INIT_23 => X"ffffff7dffffffff00000000000000000000005400000000fffffff2ffffffff",
            INIT_24 => X"ffffffd0ffffffff0000002500000000ffffff0cffffffffffffff54ffffffff",
            INIT_25 => X"ffffff90ffffffff00000004000000000000010700000000fffffff1ffffffff",
            INIT_26 => X"ffffff90ffffffff00000024000000000000009a00000000ffffff79ffffffff",
            INIT_27 => X"0000002c00000000ffffff74ffffffff0000003700000000ffffffcdffffffff",
            INIT_28 => X"fffffebdffffffffffffffe0ffffffffffffff5efffffffffffffe39ffffffff",
            INIT_29 => X"ffffffccfffffffffffffeb6ffffffffffffff82fffffffffffffefcffffffff",
            INIT_2A => X"0000008300000000ffffffd2ffffffff0000009700000000ffffff96ffffffff",
            INIT_2B => X"0000003c00000000ffffffceffffffffffffffd7ffffffff000001a900000000",
            INIT_2C => X"0000001e000000000000001c0000000000000000000000000000001f00000000",
            INIT_2D => X"0000002d0000000000000078000000000000007700000000ffffff90ffffffff",
            INIT_2E => X"0000001000000000fffffff9ffffffff00000095000000000000003900000000",
            INIT_2F => X"00000022000000000000003300000000ffffff31ffffffffffffff3cffffffff",
            INIT_30 => X"ffffffb0ffffffff000000a9000000000000003d00000000000000b200000000",
            INIT_31 => X"fffffe8bffffffffffffff52fffffffffffffe0afffffffffffffe94ffffffff",
            INIT_32 => X"fffffebeffffffffffffff2fffffffffffffff59fffffffffffffd32ffffffff",
            INIT_33 => X"ffffffc7ffffffff00000013000000000000002400000000ffffff2effffffff",
            INIT_34 => X"fffffee4ffffffff00000059000000000000002a000000000000003b00000000",
            INIT_35 => X"ffffff94ffffffff000000a300000000fffffe82fffffffffffffff2ffffffff",
            INIT_36 => X"00000016000000000000008100000000000000ce000000000000001500000000",
            INIT_37 => X"ffffff9dffffffff000000e100000000fffffefeffffffffffffffb1ffffffff",
            INIT_38 => X"000000970000000000000048000000000000003700000000ffffff30ffffffff",
            INIT_39 => X"00000054000000000000003f000000000000008b000000000000007600000000",
            INIT_3A => X"0000010400000000ffffff99ffffffff0000008a000000000000003d00000000",
            INIT_3B => X"ffffff98ffffffff0000004500000000fffffe9dffffffffffffff43ffffffff",
            INIT_3C => X"000000850000000000000079000000000000001400000000ffffff7cffffffff",
            INIT_3D => X"00000077000000000000000c00000000ffffff43ffffffff0000001a00000000",
            INIT_3E => X"0000001e000000000000001a000000000000004500000000fffffff6ffffffff",
            INIT_3F => X"0000009700000000ffffffabffffffff0000002000000000ffffffb2ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000005000000000000004600000000ffffff8cffffffff0000008800000000",
            INIT_41 => X"000000320000000000000023000000000000001100000000ffffff1cffffffff",
            INIT_42 => X"0000004600000000ffffffa1ffffffff0000007000000000ffffff95ffffffff",
            INIT_43 => X"ffffff53fffffffffffffeeeffffffffffffffc2ffffffffffffffd0ffffffff",
            INIT_44 => X"ffffff3dffffffff0000002f00000000ffffffc5ffffffff0000001500000000",
            INIT_45 => X"fffffff5ffffffffffffffedffffffff0000000300000000ffffffaeffffffff",
            INIT_46 => X"0000000a00000000fffffffeffffffff00000005000000000000000f00000000",
            INIT_47 => X"ffffff51fffffffffffffed9ffffffff0000001100000000ffffffebffffffff",
            INIT_48 => X"ffffffaefffffffffffffda1fffffffffffffed8ffffffffffffff32ffffffff",
            INIT_49 => X"ffffff2fffffffff0000004f00000000ffffff4cfffffffffffffec8ffffffff",
            INIT_4A => X"00000058000000000000002600000000ffffff42ffffffffffffff51ffffffff",
            INIT_4B => X"ffffffdbffffffff0000008d00000000000000f8000000000000001400000000",
            INIT_4C => X"0000008300000000ffffffd5ffffffffffffffc1ffffffff000000ef00000000",
            INIT_4D => X"0000002800000000000000c80000000000000009000000000000003d00000000",
            INIT_4E => X"ffffff69ffffffff000000ff00000000ffffffe5fffffffffffffdd6ffffffff",
            INIT_4F => X"0000001a000000000000000e00000000ffffff10ffffffff0000006a00000000",
            INIT_50 => X"ffffffd4ffffffffffffffa6fffffffffffffe31ffffffffffffffcbffffffff",
            INIT_51 => X"0000006c00000000ffffff79ffffffffffffffc0ffffffff0000002f00000000",
            INIT_52 => X"ffffff40fffffffffffffff9ffffffff00000000000000000000001600000000",
            INIT_53 => X"000000c2000000000000008400000000ffffffc4ffffffff000000a500000000",
            INIT_54 => X"ffffffdbffffffff00000038000000000000006b000000000000002d00000000",
            INIT_55 => X"ffffff6effffffff00000029000000000000008f000000000000004400000000",
            INIT_56 => X"fffffe79fffffffffffffff0ffffffffffffff0dffffffff0000005e00000000",
            INIT_57 => X"ffffff5dffffffff0000006f000000000000008f000000000000008800000000",
            INIT_58 => X"ffffffcaffffffffffffff71ffffffffffffffcbffffffffffffffedffffffff",
            INIT_59 => X"ffffffa7ffffffff0000001d0000000000000076000000000000003f00000000",
            INIT_5A => X"ffffffdeffffffff0000005000000000ffffffd8ffffffff0000000b00000000",
            INIT_5B => X"ffffff77ffffffff0000007a00000000fffffff6fffffffffffffecaffffffff",
            INIT_5C => X"0000004000000000ffffff2efffffffffffffff5ffffffff0000005e00000000",
            INIT_5D => X"000000d1000000000000004500000000fffffe39ffffffff0000000200000000",
            INIT_5E => X"ffffffbeffffffff00000048000000000000002d00000000ffffff85ffffffff",
            INIT_5F => X"000000000000000000000069000000000000003600000000ffffff89ffffffff",
            INIT_60 => X"0000001b00000000ffffffb7ffffffffffffff7bffffffff0000006a00000000",
            INIT_61 => X"ffffffacffffffffffffff8affffffff0000004900000000fffffecbffffffff",
            INIT_62 => X"000000f600000000ffffff83ffffffff00000062000000000000006300000000",
            INIT_63 => X"fffffff3ffffffff0000002400000000fffffffcffffffff0000002500000000",
            INIT_64 => X"000000a600000000ffffff9fffffffff0000000200000000ffffff82ffffffff",
            INIT_65 => X"ffffffcbffffffff0000006a0000000000000058000000000000000000000000",
            INIT_66 => X"00000027000000000000006400000000ffffff12ffffffff0000001500000000",
            INIT_67 => X"0000006000000000ffffffd2ffffffffffffff0fffffffff000000e900000000",
            INIT_68 => X"00000038000000000000007a00000000ffffffaaffffffffffffff62ffffffff",
            INIT_69 => X"0000004500000000ffffffc4ffffffff00000030000000000000000000000000",
            INIT_6A => X"ffffffdbffffffffffffff66ffffffffffffff54ffffffff0000009000000000",
            INIT_6B => X"ffffffd3ffffffffffffff8dfffffffffffffefdfffffffffffffff2ffffffff",
            INIT_6C => X"0000002000000000ffffffe0ffffffffffffff82ffffffff0000008a00000000",
            INIT_6D => X"000000df00000000ffffff7dffffffff0000005f00000000fffffeffffffffff",
            INIT_6E => X"ffffff27ffffffff0000000e00000000ffffff93ffffffff0000009100000000",
            INIT_6F => X"000000b400000000ffffffcdffffffffffffff42ffffffffffffff84ffffffff",
            INIT_70 => X"000000140000000000000043000000000000000f00000000ffffffc0ffffffff",
            INIT_71 => X"0000004700000000000000c600000000000000a200000000000000e000000000",
            INIT_72 => X"0000002c000000000000000000000000ffffff9dffffffff0000007d00000000",
            INIT_73 => X"0000006e000000000000004900000000ffffffa3ffffffff0000001100000000",
            INIT_74 => X"00000004000000000000006f0000000000000148000000000000006400000000",
            INIT_75 => X"000000a700000000ffffffc8ffffffff000000cd00000000ffffffd3ffffffff",
            INIT_76 => X"ffffff53ffffffffffffffeafffffffffffffff3ffffffffffffff5dffffffff",
            INIT_77 => X"0000001400000000fffffe8affffffffffffff6bffffffffffffffd1ffffffff",
            INIT_78 => X"ffffff9affffffffffffff63ffffffff0000001600000000ffffff98ffffffff",
            INIT_79 => X"ffffffdfffffffffffffffdeffffffff00000048000000000000002c00000000",
            INIT_7A => X"0000003f00000000000000300000000000000005000000000000005f00000000",
            INIT_7B => X"ffffffbeffffffff00000028000000000000002d000000000000000000000000",
            INIT_7C => X"ffffff90ffffffff00000051000000000000003e000000000000000d00000000",
            INIT_7D => X"000000b200000000000000ae00000000ffffffb4ffffffffffffffabffffffff",
            INIT_7E => X"0000002900000000ffffffd7ffffffff0000001100000000ffffff53ffffffff",
            INIT_7F => X"000000b800000000000000f800000000ffffffc6fffffffffffffef0ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE33;


    MEM_IWGHT_LAYER2_INSTANCE34 : if BRAM_NAME = "iwght_layer2_instance34" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffa7ffffffffffffff62ffffffffffffffc7ffffffff000000a000000000",
            INIT_01 => X"ffffff58ffffffffffffffeefffffffffffffef0fffffffffffffe1dffffffff",
            INIT_02 => X"0000001900000000ffffffa4ffffffffffffff5dffffffff0000009700000000",
            INIT_03 => X"ffffff88ffffffff000000ca00000000ffffff2effffffffffffffc2ffffffff",
            INIT_04 => X"0000003a00000000fffffefbffffffffffffffadfffffffffffffe5dffffffff",
            INIT_05 => X"ffffffb3ffffffff0000007800000000000000a600000000ffffffe9ffffffff",
            INIT_06 => X"0000001c00000000ffffffe4ffffffffffffff79ffffffffffffffe0ffffffff",
            INIT_07 => X"ffffff72ffffffffffffff56ffffffffffffff18ffffffff0000009e00000000",
            INIT_08 => X"ffffff98ffffffffffffffb7ffffffffffffffe3ffffffff0000000600000000",
            INIT_09 => X"0000001500000000fffffff6ffffffff0000008b000000000000007800000000",
            INIT_0A => X"000000660000000000000084000000000000006200000000ffffffb0ffffffff",
            INIT_0B => X"ffffffe4ffffffff000000540000000000000042000000000000006400000000",
            INIT_0C => X"fffffffeffffffffffffff9affffffff00000031000000000000008000000000",
            INIT_0D => X"00000000000000000000000500000000ffffffebffffffff0000006a00000000",
            INIT_0E => X"fffffff7fffffffffffffffaffffffff0000000700000000fffffff3ffffffff",
            INIT_0F => X"0000000000000000ffffff95ffffffff0000000d000000000000000d00000000",
            INIT_10 => X"00000093000000000000006c000000000000004300000000ffffffffffffffff",
            INIT_11 => X"000000c100000000ffffffd5ffffffff00000021000000000000007a00000000",
            INIT_12 => X"ffffffdbffffffffffffffe4ffffffffffffffe5ffffffff0000005400000000",
            INIT_13 => X"fffffef1fffffffffffffef2ffffffff0000004900000000ffffff75ffffffff",
            INIT_14 => X"ffffff80ffffffff0000003800000000ffffffd3ffffffff0000000c00000000",
            INIT_15 => X"0000003d000000000000001300000000ffffffd6ffffffffffffffcfffffffff",
            INIT_16 => X"0000004a000000000000007b00000000ffffffd8ffffffff0000000000000000",
            INIT_17 => X"ffffffd0ffffffff0000002000000000000000ad00000000fffffffbffffffff",
            INIT_18 => X"0000001900000000fffffff4ffffffffffffff99ffffffffffffffd3ffffffff",
            INIT_19 => X"0000008e000000000000009700000000fffffeccffffffff0000006200000000",
            INIT_1A => X"0000004b00000000ffffffdfffffffffffffffc2ffffffffffffff3fffffffff",
            INIT_1B => X"0000001e00000000ffffffb4ffffffff0000009900000000ffffffd9ffffffff",
            INIT_1C => X"0000008500000000ffffffcbffffffff0000009600000000fffffed2ffffffff",
            INIT_1D => X"000000050000000000000010000000000000008500000000ffffff7dffffffff",
            INIT_1E => X"fffffffaffffffff00000064000000000000005b00000000ffffffd9ffffffff",
            INIT_1F => X"fffffff7ffffffff0000009400000000ffffffc9ffffffffffffffb4ffffffff",
            INIT_20 => X"0000003800000000ffffff6fffffffffffffff6bffffffff0000007b00000000",
            INIT_21 => X"fffffffdffffffffffffffe0ffffffffffffffacfffffffffffffedbffffffff",
            INIT_22 => X"0000007d00000000ffffffa9ffffffffffffffcbffffffff0000018800000000",
            INIT_23 => X"ffffffe0ffffffff00000054000000000000004900000000ffffff15ffffffff",
            INIT_24 => X"0000007d000000000000005f000000000000001d00000000ffffffc6ffffffff",
            INIT_25 => X"ffffff0effffffffffffffb2ffffffff0000000b00000000ffffffdbffffffff",
            INIT_26 => X"0000006100000000ffffff56ffffffffffffff6dffffffffffffffbcffffffff",
            INIT_27 => X"0000008e0000000000000058000000000000001b000000000000008b00000000",
            INIT_28 => X"00000008000000000000003800000000000000c3000000000000005100000000",
            INIT_29 => X"ffffff51ffffffff00000006000000000000005e00000000ffffff7bffffffff",
            INIT_2A => X"ffffff30ffffffffffffff8dffffffff000000cc00000000ffffffd0ffffffff",
            INIT_2B => X"00000004000000000000004c000000000000003d00000000fffffff3ffffffff",
            INIT_2C => X"0000003400000000ffffffcdffffffffffffff8cffffffffffffffc2ffffffff",
            INIT_2D => X"ffffff65ffffffff0000004e00000000ffffff6dffffffffffffffe3ffffffff",
            INIT_2E => X"ffffff84ffffffffffffffd2ffffffffffffff93ffffffffffffffb5ffffffff",
            INIT_2F => X"00000020000000000000001900000000fffffefaffffffff000000a900000000",
            INIT_30 => X"ffffffa6ffffffff0000007a00000000ffffff91ffffffff0000007000000000",
            INIT_31 => X"ffffffe1ffffffffffffffa5ffffffffffffffc8ffffffff0000006300000000",
            INIT_32 => X"00000035000000000000000d000000000000000500000000ffffffd2ffffffff",
            INIT_33 => X"0000004f00000000ffffff0dfffffffffffffeecffffffffffffff9dffffffff",
            INIT_34 => X"ffffff8affffffff0000006600000000fffffec1ffffffff0000001400000000",
            INIT_35 => X"ffffffcdffffffff0000009a00000000ffffffe1ffffffff0000001b00000000",
            INIT_36 => X"ffffff59ffffffffffffffadffffffffffffff99ffffffffffffffdaffffffff",
            INIT_37 => X"0000000f00000000000000a400000000ffffffa8ffffffff0000000e00000000",
            INIT_38 => X"ffffffbeffffffff0000003400000000ffffffe3ffffffff0000003800000000",
            INIT_39 => X"fffffffdffffffffffffffdbffffffff0000000e00000000ffffffcbffffffff",
            INIT_3A => X"0000004c00000000ffffffdcfffffffffffffff9ffffffffffffff48ffffffff",
            INIT_3B => X"ffffffe5ffffffff0000010b00000000ffffffefffffffff0000008f00000000",
            INIT_3C => X"0000000400000000ffffff5dffffffff000000c1000000000000005c00000000",
            INIT_3D => X"0000005c00000000ffffff8bffffffffffffffabffffffff000000eb00000000",
            INIT_3E => X"00000008000000000000018600000000ffffff48ffffffffffffffa4ffffffff",
            INIT_3F => X"ffffffd8ffffffff0000003b00000000ffffff97ffffffffffffff84ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffcfffffffff0000004400000000ffffff4cffffffffffffffa7ffffffff",
            INIT_41 => X"000000070000000000000000000000000000003a000000000000008900000000",
            INIT_42 => X"ffffff4cffffffffffffffd8ffffffff0000007e00000000fffffffeffffffff",
            INIT_43 => X"ffffff33ffffffff0000009f000000000000006900000000ffffff5affffffff",
            INIT_44 => X"0000000600000000ffffffdaffffffff0000003d00000000ffffffb0ffffffff",
            INIT_45 => X"ffffff84ffffffff000000420000000000000086000000000000000600000000",
            INIT_46 => X"fffffff4ffffffffffffff51ffffffff00000047000000000000002500000000",
            INIT_47 => X"ffffffb8ffffffff0000003700000000ffffffeaffffffffffffff59ffffffff",
            INIT_48 => X"fffffef7ffffffffffffffdfffffffffffffff28ffffffffffffff7effffffff",
            INIT_49 => X"fffffff8ffffffffffffff6cffffffff0000003900000000ffffffadffffffff",
            INIT_4A => X"ffffffaeffffffffffffffebffffffff0000000900000000ffffffe1ffffffff",
            INIT_4B => X"fffffffaffffffff0000001f00000000ffffff1affffffff0000001900000000",
            INIT_4C => X"ffffffc5ffffffffffffffb2ffffffff0000002b00000000ffffffddffffffff",
            INIT_4D => X"0000001e00000000ffffffebffffffffffffff33ffffffff0000001700000000",
            INIT_4E => X"ffffffc0ffffffff0000003900000000ffffffb0ffffffffffffffeeffffffff",
            INIT_4F => X"fffffff7ffffffff0000002e0000000000000067000000000000007500000000",
            INIT_50 => X"ffffffc2ffffffff0000005c0000000000000082000000000000010e00000000",
            INIT_51 => X"ffffffccffffffffffffff8cffffffff00000013000000000000000b00000000",
            INIT_52 => X"ffffffbaffffffff00000041000000000000009400000000ffffff74ffffffff",
            INIT_53 => X"0000008b000000000000007500000000000000aa000000000000001000000000",
            INIT_54 => X"00000069000000000000002c00000000fffffff8ffffffff0000000800000000",
            INIT_55 => X"fffffffdffffffff0000000a0000000000000007000000000000006400000000",
            INIT_56 => X"0000000300000000fffffffefffffffffffffff5fffffffffffffff3ffffffff",
            INIT_57 => X"00000004000000000000001f00000000fffffffdffffffff0000000500000000",
            INIT_58 => X"0000000700000000ffffffd3fffffffffffffff7ffffffffffffffdaffffffff",
            INIT_59 => X"fffffffafffffffffffffefdffffffffffffff30ffffffffffffffe0ffffffff",
            INIT_5A => X"fffffef5ffffffffffffff9effffffffffffffb6ffffffff0000001800000000",
            INIT_5B => X"ffffff43ffffffff0000017c000000000000002300000000fffffffbffffffff",
            INIT_5C => X"0000006100000000ffffffd5ffffffffffffffdaffffffff0000002500000000",
            INIT_5D => X"0000008a00000000fffffff1ffffffffffffff12ffffffffffffffc0ffffffff",
            INIT_5E => X"00000057000000000000003500000000fffffe7fffffffff000000b200000000",
            INIT_5F => X"ffffff2fffffffff0000009100000000000000b600000000ffffffa5ffffffff",
            INIT_60 => X"ffffffb6ffffffffffffffb8ffffffff0000008200000000000000e000000000",
            INIT_61 => X"fffffed1ffffffff00000047000000000000002c000000000000010400000000",
            INIT_62 => X"ffffffc0ffffffffffffff54ffffffffffffffa0ffffffff0000006f00000000",
            INIT_63 => X"ffffff81ffffffff0000000300000000fffffff3fffffffffffffe81ffffffff",
            INIT_64 => X"0000004700000000ffffffe2ffffffff0000006d00000000000000c600000000",
            INIT_65 => X"0000002a00000000ffffffc1fffffffffffffff1ffffffffffffffbcffffffff",
            INIT_66 => X"ffffff8cffffffff0000003c00000000ffffffc1ffffffffffffff41ffffffff",
            INIT_67 => X"ffffffc4ffffffffffffffdfffffffffffffff82ffffffff0000003500000000",
            INIT_68 => X"000000ec000000000000004a00000000fffffff7ffffffff0000018200000000",
            INIT_69 => X"ffffffa7ffffffffffffffd6ffffffffffffff2fffffffff0000000300000000",
            INIT_6A => X"0000011400000000ffffffb6ffffffffffffff4bffffffff0000004f00000000",
            INIT_6B => X"ffffffacffffffffffffff88ffffffffffffff9bffffffffffffffafffffffff",
            INIT_6C => X"0000006600000000fffffffaffffffff0000000700000000ffffff19ffffffff",
            INIT_6D => X"ffffffc5ffffffff0000010a000000000000002c000000000000002a00000000",
            INIT_6E => X"0000000e000000000000002a00000000fffffff6ffffffff0000003400000000",
            INIT_6F => X"0000005a000000000000001b00000000ffffff25fffffffffffffffdffffffff",
            INIT_70 => X"000000130000000000000018000000000000008500000000ffffffb8ffffffff",
            INIT_71 => X"ffffffb8fffffffffffffff1ffffffff000000ba000000000000005100000000",
            INIT_72 => X"ffffff69ffffffffffffffd5ffffffffffffff6bffffffff0000007200000000",
            INIT_73 => X"ffffff9fffffffff000000d70000000000000078000000000000009d00000000",
            INIT_74 => X"fffffeccffffffffffffff5cfffffffffffffe9affffffff0000001200000000",
            INIT_75 => X"ffffffb0fffffffffffffff1ffffffffffffffadffffffffffffff0effffffff",
            INIT_76 => X"ffffffa7ffffffff0000005d000000000000006b00000000fffffea9ffffffff",
            INIT_77 => X"fffffed0ffffffff000000680000000000000008000000000000001200000000",
            INIT_78 => X"ffffff9bffffffff0000009e000000000000008a00000000fffffff8ffffffff",
            INIT_79 => X"ffffffb0ffffffffffffff8ffffffffffffffffbffffffffffffff3effffffff",
            INIT_7A => X"ffffff80ffffffffffffff7fffffffff0000002b00000000000000ad00000000",
            INIT_7B => X"ffffff34ffffffff0000002300000000000000c900000000ffffffd1ffffffff",
            INIT_7C => X"ffffff65ffffffff000000a5000000000000008000000000fffffef7ffffffff",
            INIT_7D => X"ffffff73ffffffffffffffe2ffffffff000000a1000000000000002000000000",
            INIT_7E => X"ffffffdaffffffff0000003900000000ffffffbfffffffffffffff80ffffffff",
            INIT_7F => X"0000000f000000000000000e000000000000006000000000ffffff62ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE34;


    MEM_IWGHT_LAYER2_INSTANCE35 : if BRAM_NAME = "iwght_layer2_instance35" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004500000000ffffffccffffffff00000085000000000000007100000000",
            INIT_01 => X"000000e100000000ffffffd7ffffffff00000022000000000000001e00000000",
            INIT_02 => X"ffffffd1ffffffff0000004b00000000ffffffebffffffff0000004200000000",
            INIT_03 => X"ffffff7effffffff000000a700000000ffffffb9ffffffffffffffe1ffffffff",
            INIT_04 => X"0000002500000000000000060000000000000010000000000000004600000000",
            INIT_05 => X"00000064000000000000003a00000000ffffff5bfffffffffffffffdffffffff",
            INIT_06 => X"ffffff98fffffffffffffff8ffffffffffffffeeffffffffffffff42ffffffff",
            INIT_07 => X"00000059000000000000004400000000ffffff2bffffffff0000001800000000",
            INIT_08 => X"ffffff60ffffffff0000006800000000ffffff59ffffffffffffffe1ffffffff",
            INIT_09 => X"ffffffffffffffff0000000700000000ffffffedffffffff0000003300000000",
            INIT_0A => X"ffffffd5ffffffff0000002f00000000ffffff45ffffffff0000001d00000000",
            INIT_0B => X"0000002900000000000000090000000000000000000000000000007900000000",
            INIT_0C => X"ffffff61ffffffffffffffedffffffffffffff7fffffffff0000005300000000",
            INIT_0D => X"ffffffa8fffffffffffffffdffffffffffffff32ffffffffffffff8effffffff",
            INIT_0E => X"ffffffc1ffffffff00000062000000000000007d00000000ffffffc7ffffffff",
            INIT_0F => X"ffffffd7ffffffff0000001400000000ffffffa5ffffffff0000004c00000000",
            INIT_10 => X"ffffffbbffffffff00000057000000000000007f00000000ffffff97ffffffff",
            INIT_11 => X"0000004700000000ffffffcaffffffffffffffd1ffffffff0000001000000000",
            INIT_12 => X"ffffffbfffffffff00000038000000000000002c000000000000006300000000",
            INIT_13 => X"0000000b00000000ffffff7cfffffffffffffff9ffffffff0000008500000000",
            INIT_14 => X"ffffffedffffffff000000520000000000000022000000000000001400000000",
            INIT_15 => X"0000008a000000000000001300000000000000d3000000000000000000000000",
            INIT_16 => X"00000045000000000000002800000000ffffffb9ffffffff0000004700000000",
            INIT_17 => X"ffffff66ffffffff0000002900000000ffffffc9ffffffff0000000d00000000",
            INIT_18 => X"ffffffe1ffffffffffffff6effffffff0000004100000000ffffffc5ffffffff",
            INIT_19 => X"ffffffe0ffffffffffffffdeffffffff00000018000000000000006700000000",
            INIT_1A => X"0000006b000000000000004c000000000000001700000000000000db00000000",
            INIT_1B => X"ffffffd1ffffffff00000070000000000000002e00000000fffffffaffffffff",
            INIT_1C => X"fffffe65ffffffffffffffb0fffffffffffffeffffffffffffffffeaffffffff",
            INIT_1D => X"00000003000000000000000f00000000fffffff5ffffffffffffff2effffffff",
            INIT_1E => X"0000000c0000000000000003000000000000001600000000ffffffe7ffffffff",
            INIT_1F => X"0000000400000000ffffff89ffffffff0000001200000000fffffff4ffffffff",
            INIT_20 => X"000000490000000000000038000000000000005700000000ffffffa0ffffffff",
            INIT_21 => X"ffffffd2ffffffff000000d00000000000000072000000000000007e00000000",
            INIT_22 => X"ffffffd8ffffffffffffff81ffffffffffffff6affffffffffffffcbffffffff",
            INIT_23 => X"00000003000000000000009700000000ffffffcaffffffff0000000a00000000",
            INIT_24 => X"ffffff4bffffffffffffffcfffffffffffffff90ffffffffffffffd7ffffffff",
            INIT_25 => X"ffffffacffffffff0000000b00000000ffffff42ffffffffffffffb0ffffffff",
            INIT_26 => X"0000007100000000fffffff0ffffffff0000000e00000000ffffffc3ffffffff",
            INIT_27 => X"0000003c00000000fffffff2ffffffffffffff76ffffffff0000002800000000",
            INIT_28 => X"0000000e000000000000001800000000ffffffd0ffffffffffffff7fffffffff",
            INIT_29 => X"ffffffc0ffffffff0000003d00000000ffffffe6ffffffffffffff80ffffffff",
            INIT_2A => X"0000001d000000000000002d00000000000000f700000000fffffec1ffffffff",
            INIT_2B => X"0000006200000000ffffff54ffffffff0000009a00000000ffffff5fffffffff",
            INIT_2C => X"ffffffdeffffffff0000008700000000ffffffebffffffff0000000200000000",
            INIT_2D => X"ffffffafffffffff0000000200000000ffffffcbfffffffffffffff5ffffffff",
            INIT_2E => X"0000000000000000ffffff76ffffffff00000046000000000000009b00000000",
            INIT_2F => X"0000009900000000ffffffefffffffff0000000f000000000000004900000000",
            INIT_30 => X"ffffffb3ffffffff0000000600000000ffffffc5fffffffffffffef5ffffffff",
            INIT_31 => X"ffffffcaffffffffffffffb7ffffffff0000000200000000ffffffdfffffffff",
            INIT_32 => X"0000009600000000ffffffe3ffffffffffffffd3ffffffffffffffe6ffffffff",
            INIT_33 => X"0000001e00000000ffffffc7ffffffff00000006000000000000006500000000",
            INIT_34 => X"0000001b000000000000001600000000ffffffc4ffffffffffffffdfffffffff",
            INIT_35 => X"0000007d00000000fffffffeffffffff00000034000000000000003000000000",
            INIT_36 => X"0000002d000000000000000300000000ffffff9ffffffffffffffffdffffffff",
            INIT_37 => X"ffffff68ffffffffffffff6fffffffff0000000300000000ffffff5effffffff",
            INIT_38 => X"ffffffacffffffffffffff87ffffffff0000007000000000ffffff98ffffffff",
            INIT_39 => X"fffffe6effffffffffffffa2ffffffffffffffa0ffffffffffffffbcffffffff",
            INIT_3A => X"fffffe86fffffffffffffffefffffffffffffed1ffffffff0000000d00000000",
            INIT_3B => X"ffffffbbffffffff0000000200000000ffffffdcffffffff0000004700000000",
            INIT_3C => X"ffffffbaffffffffffffff8effffffff00000016000000000000001c00000000",
            INIT_3D => X"0000005d000000000000005100000000ffffffe3fffffffffffffff7ffffffff",
            INIT_3E => X"0000006a000000000000002d000000000000006a00000000ffffff7dffffffff",
            INIT_3F => X"ffffffd7ffffffff000000c900000000ffffffefffffffffffffffd1ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000030000000000000006f00000000ffffff9dffffffff0000004500000000",
            INIT_41 => X"ffffff54ffffffff0000005800000000ffffffc0ffffffff0000006c00000000",
            INIT_42 => X"0000000e00000000000000d00000000000000002000000000000003400000000",
            INIT_43 => X"ffffffeeffffffffffffff0affffffff0000001e00000000ffffffebffffffff",
            INIT_44 => X"fffffff0ffffffff0000003d00000000ffffffcaffffffff0000004500000000",
            INIT_45 => X"ffffffe3ffffffff00000007000000000000001400000000ffffffceffffffff",
            INIT_46 => X"ffffffc5ffffffff000000d900000000ffffffb7ffffffff0000009d00000000",
            INIT_47 => X"ffffff81ffffffffffffffccffffffff0000005700000000ffffff49ffffffff",
            INIT_48 => X"0000002c00000000fffffff5ffffffff00000075000000000000002e00000000",
            INIT_49 => X"00000038000000000000008300000000ffffff37ffffffff0000004400000000",
            INIT_4A => X"0000005f00000000fffffff9ffffffff0000002e000000000000003200000000",
            INIT_4B => X"00000010000000000000003a000000000000002000000000ffffff6bffffffff",
            INIT_4C => X"0000000d00000000ffffff93ffffffffffffffb3ffffffffffffff99ffffffff",
            INIT_4D => X"0000002a000000000000002400000000ffffffd7ffffffffffffffa1ffffffff",
            INIT_4E => X"0000003400000000ffffffc6ffffffff0000007a000000000000007800000000",
            INIT_4F => X"0000000c0000000000000006000000000000009600000000ffffffd0ffffffff",
            INIT_50 => X"ffffffaaffffffff0000002a00000000ffffff55ffffffffffffffa3ffffffff",
            INIT_51 => X"0000005100000000000000490000000000000003000000000000001200000000",
            INIT_52 => X"000000900000000000000002000000000000002f000000000000005400000000",
            INIT_53 => X"0000007700000000ffffffd4ffffffff0000008500000000ffffff63ffffffff",
            INIT_54 => X"0000000700000000ffffff7effffffffffffffaeffffffffffffffd6ffffffff",
            INIT_55 => X"ffffff97ffffffff00000032000000000000002400000000ffffffc9ffffffff",
            INIT_56 => X"0000013500000000ffffffd5ffffffff0000001200000000000000f500000000",
            INIT_57 => X"0000000b000000000000000500000000ffffffb6ffffffffffffffb6ffffffff",
            INIT_58 => X"ffffffcfffffffff00000005000000000000000300000000ffffffbcffffffff",
            INIT_59 => X"ffffffe9ffffffffffffff8dffffffff00000000000000000000000800000000",
            INIT_5A => X"00000016000000000000002a00000000ffffffe2ffffffff0000006e00000000",
            INIT_5B => X"fffffff1ffffffffffffffa4ffffffff0000003f00000000ffffff5fffffffff",
            INIT_5C => X"00000020000000000000007000000000000000fc000000000000001100000000",
            INIT_5D => X"0000002300000000000000a0000000000000009100000000fffffffeffffffff",
            INIT_5E => X"0000003300000000ffffff5cffffffffffffffb2ffffffffffffff9fffffffff",
            INIT_5F => X"ffffffdfffffffff0000002d0000000000000054000000000000003200000000",
            INIT_60 => X"00000018000000000000008600000000ffffffaeffffffff0000006400000000",
            INIT_61 => X"fffffff4ffffffff0000000e0000000000000008000000000000002e00000000",
            INIT_62 => X"0000002a00000000ffffff83ffffffff00000037000000000000002c00000000",
            INIT_63 => X"0000000100000000000000e700000000000000d8000000000000005100000000",
            INIT_64 => X"0000002600000000fffffffaffffffffffffffc5ffffffff0000003b00000000",
            INIT_65 => X"0000000b0000000000000000000000000000000d00000000ffffff99ffffffff",
            INIT_66 => X"0000001c00000000fffffff8fffffffffffffff9ffffffff0000001600000000",
            INIT_67 => X"00000046000000000000002d00000000fffffffefffffffffffffffeffffffff",
            INIT_68 => X"ffffffdeffffffff000000470000000000000042000000000000000300000000",
            INIT_69 => X"ffffff56ffffffff000000200000000000000040000000000000008d00000000",
            INIT_6A => X"ffffff76ffffffffffffffdcffffffff0000002d00000000ffffff2effffffff",
            INIT_6B => X"000000be000000000000001d00000000ffffff8ffffffffffffffff7ffffffff",
            INIT_6C => X"0000001500000000ffffff99ffffffffffffffc7fffffffffffffffdffffffff",
            INIT_6D => X"0000001a000000000000001d000000000000008c000000000000001600000000",
            INIT_6E => X"000000bc00000000ffffffa8ffffffff0000007d00000000ffffffb5ffffffff",
            INIT_6F => X"ffffff8bffffffff00000001000000000000008900000000ffffffeeffffffff",
            INIT_70 => X"000000da0000000000000053000000000000009b000000000000005400000000",
            INIT_71 => X"ffffff9dffffffff000000060000000000000047000000000000001500000000",
            INIT_72 => X"0000006e00000000ffffffd8ffffffff0000005200000000ffffffbcffffffff",
            INIT_73 => X"ffffffe9ffffffffffffff4effffffff0000008700000000000000b700000000",
            INIT_74 => X"0000007600000000ffffff70fffffffffffffe9affffffff0000008c00000000",
            INIT_75 => X"ffffffaaffffffffffffffcfffffffffffffff27ffffffffffffff7cffffffff",
            INIT_76 => X"ffffff24ffffffff0000008f00000000ffffffe3fffffffffffffedeffffffff",
            INIT_77 => X"00000046000000000000000100000000fffffff9ffffffffffffffcbffffffff",
            INIT_78 => X"ffffffcdffffffff0000002e00000000ffffffe6ffffffffffffffcbffffffff",
            INIT_79 => X"ffffff71ffffffffffffffb6ffffffff0000003d000000000000000300000000",
            INIT_7A => X"000000dd000000000000007e00000000ffffffccffffffffffffff82ffffffff",
            INIT_7B => X"ffffffdfffffffff00000030000000000000000000000000ffffffb2ffffffff",
            INIT_7C => X"ffffffb3ffffffff00000032000000000000001e00000000fffffffeffffffff",
            INIT_7D => X"fffffff9ffffffffffffffbdffffffff0000006900000000ffffff77ffffffff",
            INIT_7E => X"00000002000000000000001900000000ffffffd8ffffffff0000007b00000000",
            INIT_7F => X"0000000f0000000000000059000000000000004a000000000000004c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE35;


    MEM_IWGHT_LAYER2_INSTANCE36 : if BRAM_NAME = "iwght_layer2_instance36" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffebffffffffffffffedfffffffffffffff9ffffffff0000003a00000000",
            INIT_01 => X"000000160000000000000070000000000000006b00000000ffffffcdffffffff",
            INIT_02 => X"000000970000000000000003000000000000005d000000000000000000000000",
            INIT_03 => X"0000008300000000ffffff6dffffffffffffffb4ffffffffffffff3effffffff",
            INIT_04 => X"00000016000000000000005000000000ffffffb2ffffffff0000000300000000",
            INIT_05 => X"000000ae00000000000000350000000000000013000000000000000b00000000",
            INIT_06 => X"00000028000000000000001200000000ffffff8cffffffff0000004c00000000",
            INIT_07 => X"00000018000000000000004200000000ffffffe3ffffffff0000001800000000",
            INIT_08 => X"0000006400000000ffffff99fffffffffffffff6ffffffff0000000c00000000",
            INIT_09 => X"ffffff8bffffffff0000004f0000000000000007000000000000001400000000",
            INIT_0A => X"ffffff84ffffffff0000003f000000000000005c00000000ffffff78ffffffff",
            INIT_0B => X"00000053000000000000004b00000000ffffffe9ffffffffffffffccffffffff",
            INIT_0C => X"00000027000000000000001a0000000000000030000000000000003e00000000",
            INIT_0D => X"ffffff4efffffffffffffff7ffffffff0000002d00000000ffffff50ffffffff",
            INIT_0E => X"00000097000000000000000600000000fffffff3ffffffffffffffc5ffffffff",
            INIT_0F => X"ffffffe0ffffffffffffffaaffffffff0000003e00000000ffffffadffffffff",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE36;


    MEM_IWGHT_LAYER3_INSTANCE0 : if BRAM_NAME = "iwght_layer3_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000d03500000000fffe9044fffffffffffe8cefffffffffffffa5f9ffffffff",
            INIT_01 => X"0000025400000000000055e400000000fffffde2ffffffff0001bca900000000",
            INIT_02 => X"fffffff0ffffffff000000060000000000000a5b00000000ffffa58dffffffff",
            INIT_03 => X"ffffff61ffffffffffffff27ffffffff0000005a00000000000000f000000000",
            INIT_04 => X"fffffff9ffffffffffffffb1ffffffff0000001a00000000ffffffeaffffffff",
            INIT_05 => X"0000006f00000000ffffff11ffffffffffffff0bffffffffffffffe8ffffffff",
            INIT_06 => X"0000006d000000000000002300000000ffffffe3ffffffff0000000000000000",
            INIT_07 => X"00000002000000000000005000000000ffffffcbffffffff0000006f00000000",
            INIT_08 => X"00000040000000000000002700000000fffffedbffffffff0000000200000000",
            INIT_09 => X"0000002100000000ffffffd9ffffffffffffffb7ffffffffffffffbbffffffff",
            INIT_0A => X"ffffffaeffffffffffffffe1ffffffffffffff90ffffffffffffff44ffffffff",
            INIT_0B => X"ffffffa3ffffffffffffffedfffffffffffffff5ffffffff0000005400000000",
            INIT_0C => X"0000003a000000000000000800000000ffffff98ffffffff0000001f00000000",
            INIT_0D => X"ffffff92ffffffffffffff5cffffffffffffffdbfffffffffffffffbffffffff",
            INIT_0E => X"ffffff51ffffffff0000001800000000ffffffffffffffff0000009800000000",
            INIT_0F => X"0000003300000000ffffff7affffffff000000ae00000000ffffff1effffffff",
            INIT_10 => X"ffffffdeffffffff00000024000000000000002d00000000ffffffe6ffffffff",
            INIT_11 => X"ffffff93ffffffffffffffe1ffffffff0000001f00000000ffffffcfffffffff",
            INIT_12 => X"0000003200000000ffffffecffffffffffffffddffffffff0000000900000000",
            INIT_13 => X"0000001000000000ffffff37ffffffff0000003800000000ffffffd5ffffffff",
            INIT_14 => X"00000033000000000000001200000000ffffffecffffffff0000001700000000",
            INIT_15 => X"0000008700000000ffffffa4ffffffffffffffd2ffffffff0000005400000000",
            INIT_16 => X"0000001f00000000000000cc00000000ffffffacffffffffffffffe4ffffffff",
            INIT_17 => X"0000001200000000ffffffffffffffff0000002a000000000000002d00000000",
            INIT_18 => X"00000010000000000000003f000000000000007a00000000ffffffbdffffffff",
            INIT_19 => X"0000009700000000ffffffc6ffffffffffffff93ffffffff0000004100000000",
            INIT_1A => X"fffffff1ffffffff00000073000000000000005300000000fffffff9ffffffff",
            INIT_1B => X"fffffff1fffffffffffffffafffffffffffffffcffffffff0000000200000000",
            INIT_1C => X"ffffffd1fffffffffffffffdffffffff0000002c00000000ffffff90ffffffff",
            INIT_1D => X"ffffffdeffffffffffffffcffffffffffffffff9ffffffffffffffe7ffffffff",
            INIT_1E => X"ffffffeeffffffff0000004100000000ffffffa9fffffffffffffff4ffffffff",
            INIT_1F => X"ffffffe0ffffffffffffffd5ffffffff0000001f000000000000001f00000000",
            INIT_20 => X"ffffffd8ffffffffffffff7fffffffff0000000800000000ffffffefffffffff",
            INIT_21 => X"ffffff8cffffffff0000003e00000000ffffffabfffffffffffffffaffffffff",
            INIT_22 => X"0000003900000000fffffff5ffffffff0000000f00000000ffffff3fffffffff",
            INIT_23 => X"ffffffecffffffff00000113000000000000003400000000000000c200000000",
            INIT_24 => X"ffffffd7ffffffff0000005400000000ffffffd7ffffffffffffffe6ffffffff",
            INIT_25 => X"0000002e000000000000002000000000ffffffe9ffffffffffffff6fffffffff",
            INIT_26 => X"000000160000000000000027000000000000002f00000000ffffffe9ffffffff",
            INIT_27 => X"0000001600000000ffffffabffffffff00000078000000000000003100000000",
            INIT_28 => X"ffffffcaffffffffffffff84ffffffffffffff68ffffffff0000001b00000000",
            INIT_29 => X"fffffff7ffffffff0000000200000000ffffff98ffffffffffffffe0ffffffff",
            INIT_2A => X"000000a6000000000000003b000000000000008c000000000000004800000000",
            INIT_2B => X"ffffffd1fffffffffffffffbffffffff0000000f000000000000005200000000",
            INIT_2C => X"ffffffb6fffffffffffffff2ffffffffffffffd0fffffffffffffff0ffffffff",
            INIT_2D => X"ffffffadffffffff00000003000000000000002400000000ffffff9bffffffff",
            INIT_2E => X"ffffff51ffffffffffffffecfffffffffffffe36ffffffff0000000200000000",
            INIT_2F => X"ffffffa1ffffffffffffff68ffffffff0000004000000000ffffffcdffffffff",
            INIT_30 => X"ffffffcbffffffffffffffeeffffffffffffff97ffffffff0000000900000000",
            INIT_31 => X"ffffff9effffffffffffff6fffffffff0000002c000000000000003a00000000",
            INIT_32 => X"ffffff8cffffffff0000000200000000ffffffecffffffffffffff35ffffffff",
            INIT_33 => X"ffffffbbffffffffffffffceffffffff0000000f000000000000000b00000000",
            INIT_34 => X"ffffffc0ffffffffffffffc6ffffffff0000006800000000fffffffcffffffff",
            INIT_35 => X"fffffeceffffffffffffffc5ffffffffffffffabfffffffffffffeaaffffffff",
            INIT_36 => X"000000120000000000000044000000000000000f000000000000001600000000",
            INIT_37 => X"0000001700000000ffffffdaffffffff00000011000000000000005d00000000",
            INIT_38 => X"ffffffccffffffff00000004000000000000000c00000000ffffffafffffffff",
            INIT_39 => X"ffffff5affffffffffffff45ffffffff00000005000000000000003800000000",
            INIT_3A => X"ffffffbdffffffff0000005200000000ffffff9bffffffff0000000d00000000",
            INIT_3B => X"00000002000000000000004f00000000ffffffeafffffffffffffff0ffffffff",
            INIT_3C => X"00000005000000000000004200000000ffffff6cffffffffffffffb4ffffffff",
            INIT_3D => X"ffffffc7ffffffff00000020000000000000002300000000ffffffdcffffffff",
            INIT_3E => X"0000006900000000ffffffe2ffffffff0000007b00000000fffffffdffffffff",
            INIT_3F => X"ffffff89ffffffff00000011000000000000002d000000000000001200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001100000000000000350000000000000082000000000000000300000000",
            INIT_41 => X"0000004d000000000000005700000000fffffed9ffffffffffffffb5ffffffff",
            INIT_42 => X"ffffff74fffffffffffffff9ffffffff0000005000000000ffffff9bffffffff",
            INIT_43 => X"0000002400000000000000c100000000ffffffbdffffffffffffff52ffffffff",
            INIT_44 => X"0000003a0000000000000023000000000000004f00000000ffffffe8ffffffff",
            INIT_45 => X"ffffff37ffffffffffffffc2ffffffff0000000a00000000fffffec2ffffffff",
            INIT_46 => X"ffffffa9ffffffff0000005000000000ffffffc5fffffffffffffffcffffffff",
            INIT_47 => X"00000010000000000000009f0000000000000023000000000000008f00000000",
            INIT_48 => X"ffffffd8ffffffff00000043000000000000009c00000000ffffff64ffffffff",
            INIT_49 => X"fffffff3ffffffffffffff3fffffffff0000004c00000000ffffff61ffffffff",
            INIT_4A => X"00000014000000000000004d00000000ffffffe9ffffffffffffffaaffffffff",
            INIT_4B => X"ffffffffffffffff0000004b00000000fffffffdffffffffffffffceffffffff",
            INIT_4C => X"0000005700000000ffffffb4ffffffffffffffd3ffffffffffffff0bffffffff",
            INIT_4D => X"ffffff7bffffffff00000065000000000000008e00000000fffffffeffffffff",
            INIT_4E => X"ffffff90ffffffff0000001f000000000000007f00000000fffffff4ffffffff",
            INIT_4F => X"ffffffdbfffffffffffffff4ffffffffffffffdfffffffffffffffc4ffffffff",
            INIT_50 => X"ffffffeeffffffff0000009300000000ffffff72fffffffffffffff2ffffffff",
            INIT_51 => X"0000004d000000000000004700000000ffffff94fffffffffffffffcffffffff",
            INIT_52 => X"ffffff80fffffffffffffffeffffffffffffffe4ffffffff0000000b00000000",
            INIT_53 => X"ffffffbdffffffff000000450000000000000015000000000000004f00000000",
            INIT_54 => X"ffffffbcffffffff000000e400000000ffffffb7ffffffff0000000c00000000",
            INIT_55 => X"ffffffcdffffffff0000002900000000ffffffdaffffffffffffff63ffffffff",
            INIT_56 => X"ffffff89ffffffff00000024000000000000008a000000000000000300000000",
            INIT_57 => X"0000000400000000ffffffbffffffffffffffffaffffffff0000000500000000",
            INIT_58 => X"ffffff2fffffffffffffffa7fffffffffffffe40ffffffffffffffe3ffffffff",
            INIT_59 => X"0000000700000000ffffff14ffffffffffffff99ffffffffffffffa2ffffffff",
            INIT_5A => X"ffffffc3ffffffffffffffc9ffffffff0000004c00000000fffffff6ffffffff",
            INIT_5B => X"0000003100000000ffffff95fffffffffffffffffffffffffffffffbffffffff",
            INIT_5C => X"ffffff64ffffffff0000002a00000000ffffff81ffffffffffffff4affffffff",
            INIT_5D => X"ffffff77ffffffffffffffdbffffffff0000006f00000000ffffff93ffffffff",
            INIT_5E => X"fffffff3fffffffffffffffaffffffffffffff13ffffffffffffffaeffffffff",
            INIT_5F => X"ffffffdaffffffffffffffc7ffffffff0000000e000000000000009200000000",
            INIT_60 => X"ffffff80ffffffff0000003900000000ffffff36fffffffffffffffaffffffff",
            INIT_61 => X"fffffff1fffffffffffffffdffffffffffffff8fffffffff0000007100000000",
            INIT_62 => X"000000190000000000000008000000000000003700000000ffffff47ffffffff",
            INIT_63 => X"ffffff92ffffffff0000003e00000000ffffff90ffffffffffffff9cffffffff",
            INIT_64 => X"fffffffbffffffff0000002600000000fffffff5ffffffff0000001200000000",
            INIT_65 => X"fffffff3ffffffff0000002100000000ffffffdfffffffffffffff55ffffffff",
            INIT_66 => X"ffffffffffffffff0000004d00000000ffffffd0ffffffff0000000700000000",
            INIT_67 => X"0000000a000000000000001400000000ffffffaaffffffff000000c900000000",
            INIT_68 => X"0000002d00000000ffffff6cffffffffffffffc7ffffffffffffffc0ffffffff",
            INIT_69 => X"fffffffaffffffff0000000e00000000ffffff72ffffffff0000002900000000",
            INIT_6A => X"0000006600000000000000fd00000000ffffff18ffffffffffffffc3ffffffff",
            INIT_6B => X"00000003000000000000002800000000fffffffafffffffffffffffbffffffff",
            INIT_6C => X"00000014000000000000004900000000ffffff16ffffffff0000000500000000",
            INIT_6D => X"ffffff93ffffffffffffffa5ffffffff0000003500000000ffffff90ffffffff",
            INIT_6E => X"fffffffbffffffffffffff86ffffffff00000070000000000000004300000000",
            INIT_6F => X"ffffffb5ffffffff0000003000000000ffffff65ffffffff0000004700000000",
            INIT_70 => X"0000007e00000000ffffffa8ffffffff00000097000000000000000900000000",
            INIT_71 => X"ffffff95ffffffff0000000500000000ffffff80ffffffffffffffb1ffffffff",
            INIT_72 => X"0000002400000000fffffff9ffffffff0000001d00000000ffffff86ffffffff",
            INIT_73 => X"ffffffb8ffffffff0000009300000000ffffffa4ffffffff0000002b00000000",
            INIT_74 => X"ffffffc3ffffffff00000038000000000000001b000000000000001400000000",
            INIT_75 => X"ffffffd4ffffffffffffffc8ffffffffffffffebffffffffffffff9dffffffff",
            INIT_76 => X"0000002b00000000ffffffccffffffff0000001500000000ffffffebffffffff",
            INIT_77 => X"00000006000000000000000900000000ffffffa8ffffffff000000ac00000000",
            INIT_78 => X"0000001b00000000ffffffa4ffffffff0000003100000000ffffffe1ffffffff",
            INIT_79 => X"0000000b00000000ffffff2cfffffffffffffffaffffffffffffffe9ffffffff",
            INIT_7A => X"0000000c00000000000000f1000000000000003200000000ffffff55ffffffff",
            INIT_7B => X"fffffff4ffffffff00000033000000000000000700000000ffffffbdffffffff",
            INIT_7C => X"ffffffd5ffffffff0000001e000000000000002a00000000ffffff7cffffffff",
            INIT_7D => X"0000001400000000ffffffd9ffffffffffffffd0ffffffff0000004700000000",
            INIT_7E => X"0000003200000000ffffffcdffffffffffffff0effffffff0000002200000000",
            INIT_7F => X"0000002b000000000000002d000000000000000600000000ffffffa9ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE0;


    MEM_IWGHT_LAYER3_INSTANCE1 : if BRAM_NAME = "iwght_layer3_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004a00000000ffffffa6ffffffffffffffddffffffffffffffe0ffffffff",
            INIT_01 => X"ffffff69ffffffffffffffc6ffffffffffffff1fffffffff0000007600000000",
            INIT_02 => X"ffffffd7fffffffffffffff4ffffffffffffffe1ffffffffffffffdfffffffff",
            INIT_03 => X"ffffffc6ffffffff00000097000000000000003d000000000000000c00000000",
            INIT_04 => X"ffffff7cffffffff000000300000000000000090000000000000001200000000",
            INIT_05 => X"00000036000000000000005c00000000fffffff3ffffffffffffffc5ffffffff",
            INIT_06 => X"0000002700000000ffffffb6fffffffffffffff2ffffffff0000000900000000",
            INIT_07 => X"fffffff6ffffffffffffffd9ffffffffffffffe1ffffffff0000007900000000",
            INIT_08 => X"ffffffefffffffff0000000300000000ffffffacffffffffffffffe2ffffffff",
            INIT_09 => X"ffffffd8ffffffffffffffe0ffffffffffffffc1ffffffffffffff43ffffffff",
            INIT_0A => X"ffffffcdffffffff00000049000000000000003a000000000000006800000000",
            INIT_0B => X"0000001000000000ffffff64ffffffffffffffefffffffffffffffdfffffffff",
            INIT_0C => X"ffffff94ffffffff0000000d00000000fffffef4ffffffff000000a700000000",
            INIT_0D => X"ffffff62ffffffffffffff9cffffffff0000005700000000ffffffbeffffffff",
            INIT_0E => X"ffffff82ffffffffffffffc7ffffffff0000004a00000000ffffff5dffffffff",
            INIT_0F => X"ffffffebffffffff0000005e00000000ffffff95ffffffffffffff26ffffffff",
            INIT_10 => X"ffffff62ffffffff0000001f00000000fffffff6ffffffff0000000600000000",
            INIT_11 => X"0000000d00000000000000c000000000ffffff9fffffffff000000b200000000",
            INIT_12 => X"ffffffc4fffffffffffffff6ffffffff00000011000000000000003f00000000",
            INIT_13 => X"00000013000000000000008200000000ffffff8bffffffffffffff3dffffffff",
            INIT_14 => X"ffffffcbffffffffffffff92ffffffff0000001000000000ffffffebffffffff",
            INIT_15 => X"0000008800000000ffffffffffffffff0000005e00000000fffffff0ffffffff",
            INIT_16 => X"ffffffa6ffffffff0000002500000000ffffffbdfffffffffffffff4ffffffff",
            INIT_17 => X"ffffffefffffffff0000005a00000000fffffffaffffffff0000004600000000",
            INIT_18 => X"00000023000000000000001800000000ffffff90fffffffffffffff8ffffffff",
            INIT_19 => X"0000005700000000ffffffdeffffffff0000000f00000000ffffff8dffffffff",
            INIT_1A => X"fffffffbffffffffffffffe0ffffffff0000007800000000000000b600000000",
            INIT_1B => X"00000000000000000000005e00000000fffffffdffffffffffffffcbffffffff",
            INIT_1C => X"ffffffd9ffffffffffffff9effffffffffffffc8ffffffffffffffbbffffffff",
            INIT_1D => X"ffffff9afffffffffffffff4ffffffffffffffe2ffffffff0000002e00000000",
            INIT_1E => X"fffffffbffffffffffffffeefffffffffffffee6ffffffff0000002200000000",
            INIT_1F => X"ffffffefffffffffffffffd8ffffffffffffff90ffffffff0000001c00000000",
            INIT_20 => X"0000000b00000000fffffff4ffffffffffffff83ffffffff0000001500000000",
            INIT_21 => X"0000007b00000000ffffff7effffffffffffff7cffffffffffffff8cffffffff",
            INIT_22 => X"0000005200000000ffffffeeffffffffffffff94ffffffff0000002c00000000",
            INIT_23 => X"0000003c00000000ffffff09ffffffffffffffccffffffff0000008400000000",
            INIT_24 => X"ffffffc8ffffffffffffffeeffffffff0000005d000000000000001100000000",
            INIT_25 => X"0000002000000000ffffff82ffffffffffffff32ffffffffffffff28ffffffff",
            INIT_26 => X"ffffffa3fffffffffffffff1ffffffff00000038000000000000000d00000000",
            INIT_27 => X"ffffffe6ffffffff0000008200000000ffffff3cfffffffffffffffeffffffff",
            INIT_28 => X"0000001600000000ffffff81ffffffffffffffacffffffffffffffb0ffffffff",
            INIT_29 => X"0000003500000000ffffff86ffffffff0000000400000000ffffffd6ffffffff",
            INIT_2A => X"0000006000000000ffffff4ffffffffffffffff6fffffffffffffff6ffffffff",
            INIT_2B => X"ffffffdfffffffffffffffd9fffffffffffffff6ffffffff0000000a00000000",
            INIT_2C => X"ffffffb0ffffffffffffffd5ffffffffffffff67ffffffffffffff9cffffffff",
            INIT_2D => X"000000740000000000000057000000000000003400000000ffffffa9ffffffff",
            INIT_2E => X"00000028000000000000001000000000ffffffcafffffffffffffff4ffffffff",
            INIT_2F => X"ffffff86ffffffffffffffebffffffffffffff55ffffffff0000005b00000000",
            INIT_30 => X"0000007200000000ffffffeeffffffff0000000800000000ffffffe7ffffffff",
            INIT_31 => X"0000003f00000000000000720000000000000018000000000000003800000000",
            INIT_32 => X"00000041000000000000001800000000fffffff4fffffffffffffffaffffffff",
            INIT_33 => X"00000051000000000000007d000000000000002a000000000000014e00000000",
            INIT_34 => X"0000000800000000ffffffb5ffffffff0000005700000000ffffffe5ffffffff",
            INIT_35 => X"ffffffbfffffffffffffffc0ffffffff0000003e00000000ffffffacffffffff",
            INIT_36 => X"00000068000000000000000a00000000fffffff9ffffffff0000001300000000",
            INIT_37 => X"fffffff4ffffffff0000001c000000000000000e00000000ffffffe2ffffffff",
            INIT_38 => X"00000046000000000000001500000000ffffffa9fffffffffffffffdffffffff",
            INIT_39 => X"000000a600000000ffffff23ffffffff0000008b00000000ffffff68ffffffff",
            INIT_3A => X"ffffff60ffffffff0000006b0000000000000035000000000000002300000000",
            INIT_3B => X"0000001b00000000ffffffc4ffffffffffffffefffffffffffffff92ffffffff",
            INIT_3C => X"ffffffe6ffffffffffffffe9ffffffff00000000000000000000008d00000000",
            INIT_3D => X"0000003800000000ffffffcaffffffffffffffadffffffff0000000700000000",
            INIT_3E => X"ffffffebffffffffffffff4affffffffffffff3fffffffffffffffffffffffff",
            INIT_3F => X"fffffff8fffffffffffffff6ffffffffffffffa2ffffffff0000002000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008300000000ffffffb7ffffffff00000031000000000000001900000000",
            INIT_41 => X"ffffffbfffffffff0000002200000000fffffed2fffffffffffffffbffffffff",
            INIT_42 => X"00000000000000000000000000000000fffffffbffffffffffffffddffffffff",
            INIT_43 => X"0000000100000000ffffff77ffffffff00000031000000000000007300000000",
            INIT_44 => X"0000003000000000ffffff7fffffffff0000004000000000ffffffddffffffff",
            INIT_45 => X"0000009200000000ffffffc7ffffffffffffffe0ffffffffffffff50ffffffff",
            INIT_46 => X"ffffff48ffffffffffffffc7ffffffff0000002800000000ffffffedffffffff",
            INIT_47 => X"ffffffecffffffff0000005f00000000ffffffebffffffffffffffe5ffffffff",
            INIT_48 => X"fffffffaffffffff00000037000000000000003c00000000ffffffe8ffffffff",
            INIT_49 => X"ffffff77ffffffffffffffd0ffffffff0000003a00000000fffffff7ffffffff",
            INIT_4A => X"0000002300000000ffffff68ffffffffffffffd2fffffffffffffed1ffffffff",
            INIT_4B => X"0000004f00000000ffffff51fffffffffffffff6ffffffffffffff1effffffff",
            INIT_4C => X"ffffffaeffffffffffffffdbffffffff0000006f00000000000000b500000000",
            INIT_4D => X"ffffffd0ffffffffffffff13ffffffff00000008000000000000001a00000000",
            INIT_4E => X"ffffffb4fffffffffffffff8ffffffffffffffd0ffffffffffffffb0ffffffff",
            INIT_4F => X"00000050000000000000005c00000000ffffffc9ffffffff0000001300000000",
            INIT_50 => X"ffffffeaffffffff00000056000000000000002200000000fffffff8ffffffff",
            INIT_51 => X"ffffff64ffffffff0000002d00000000fffffea5fffffffffffffffdffffffff",
            INIT_52 => X"ffffff5bffffffffffffffe6ffffffffffffffdcffffffffffffffd1ffffffff",
            INIT_53 => X"0000003600000000fffffefbffffffff00000063000000000000001a00000000",
            INIT_54 => X"0000001100000000fffffff0ffffffff0000003a00000000ffffffefffffffff",
            INIT_55 => X"0000004c00000000ffffff5effffffffffffff8fffffffff0000008a00000000",
            INIT_56 => X"fffffedcffffffff000000ca00000000ffffffd4ffffffff0000000c00000000",
            INIT_57 => X"0000000900000000ffffffdbffffffff00000065000000000000005800000000",
            INIT_58 => X"ffffffe5ffffffffffffffdfffffffffffffffa2ffffffff0000006000000000",
            INIT_59 => X"ffffff3cfffffffffffffee6ffffffff0000000700000000ffffffb6ffffffff",
            INIT_5A => X"fffffff6ffffffffffffff2dfffffffffffffe61ffffffffffffffdcffffffff",
            INIT_5B => X"ffffffc0ffffffffffffff6fffffffff0000001700000000ffffffdfffffffff",
            INIT_5C => X"ffffff54ffffffff00000043000000000000000a00000000ffffffbfffffffff",
            INIT_5D => X"ffffffd2ffffffffffffff3cffffffff00000006000000000000003600000000",
            INIT_5E => X"fffffff2ffffffff00000020000000000000001e00000000ffffff78ffffffff",
            INIT_5F => X"0000009700000000fffffffbffffffffffffffe7ffffffffffffffd4ffffffff",
            INIT_60 => X"000000100000000000000042000000000000006800000000ffffffffffffffff",
            INIT_61 => X"00000010000000000000006500000000fffffff8ffffffff000000e000000000",
            INIT_62 => X"ffffff93ffffffffffffffecffffffff0000000000000000ffffff9dffffffff",
            INIT_63 => X"0000004000000000ffffff2bffffffff0000003400000000fffffe96ffffffff",
            INIT_64 => X"0000006100000000fffffff4ffffffff0000002700000000fffffff8ffffffff",
            INIT_65 => X"0000000900000000fffffff4ffffffff0000000000000000ffffff62ffffffff",
            INIT_66 => X"ffffff93ffffffff00000031000000000000002500000000fffffffbffffffff",
            INIT_67 => X"ffffffe9ffffffffffffffe6ffffffffffffff42ffffffffffffffd7ffffffff",
            INIT_68 => X"0000000d000000000000006b000000000000006900000000ffffffffffffffff",
            INIT_69 => X"ffffff88ffffffffffffff96ffffffff0000002e00000000ffffff92ffffffff",
            INIT_6A => X"0000008100000000ffffff82fffffffffffffed7ffffffff0000000d00000000",
            INIT_6B => X"0000001b00000000ffffffd9ffffffff0000000b00000000ffffffe4ffffffff",
            INIT_6C => X"ffffffecffffffffffffffaaffffffff000000c0000000000000009c00000000",
            INIT_6D => X"0000003100000000ffffffdcffffffffffffffc4ffffffffffffff44ffffffff",
            INIT_6E => X"ffffff66fffffffffffffe8dffffffffffffffd2ffffffffffffff6dffffffff",
            INIT_6F => X"0000007500000000ffffffa8ffffffffffffffd9ffffffff0000001600000000",
            INIT_70 => X"0000004800000000fffffff1fffffffffffffd7effffffff0000000300000000",
            INIT_71 => X"ffffff25ffffffffffffffedffffffff00000019000000000000001200000000",
            INIT_72 => X"fffffef8ffffffffffffffedffffffffffffffa9ffffffffffffff21ffffffff",
            INIT_73 => X"0000003500000000ffffffe7ffffffff0000001d00000000ffffffafffffffff",
            INIT_74 => X"0000009800000000ffffffa5ffffffff0000006d00000000fffffff3ffffffff",
            INIT_75 => X"0000006900000000ffffff36ffffffffffffffe2fffffffffffffef2ffffffff",
            INIT_76 => X"0000000000000000ffffff9effffffff0000000500000000ffffffecffffffff",
            INIT_77 => X"ffffffeeffffffff0000005200000000ffffff1cffffffff0000000d00000000",
            INIT_78 => X"ffffffbfffffffffffffffa5ffffffff0000008e00000000ffffff6fffffffff",
            INIT_79 => X"ffffff47ffffffffffffffc7ffffffff000000b800000000fffffffbffffffff",
            INIT_7A => X"ffffff40ffffffffffffff7effffffffffffff55ffffffff0000006400000000",
            INIT_7B => X"0000002a00000000ffffff06fffffffffffffff3ffffffff0000005000000000",
            INIT_7C => X"0000005a00000000ffffff83ffffffffffffffedffffffffffffff39ffffffff",
            INIT_7D => X"ffffffd9ffffffffffffff9fffffffffffffffffffffffffffffff16ffffffff",
            INIT_7E => X"00000040000000000000009f00000000ffffffd2ffffffff000000de00000000",
            INIT_7F => X"000000000000000000000056000000000000003100000000ffffff55ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE1;


    MEM_IWGHT_LAYER3_INSTANCE2 : if BRAM_NAME = "iwght_layer3_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffffdffffffff00000092000000000000000a000000000000000a00000000",
            INIT_01 => X"0000000c00000000000000c600000000ffffff8cffffffffffffff41ffffffff",
            INIT_02 => X"ffffffb7ffffffff0000000800000000ffffffe2ffffffffffffffdcffffffff",
            INIT_03 => X"0000002b00000000fffffe1bffffffff0000001900000000ffffffc8ffffffff",
            INIT_04 => X"0000003f000000000000006a00000000ffffffdbffffffff0000001600000000",
            INIT_05 => X"0000009300000000ffffffc4ffffffff0000003b00000000fffffe37ffffffff",
            INIT_06 => X"00000031000000000000007100000000ffffffaafffffffffffffffaffffffff",
            INIT_07 => X"fffffff4ffffffff000000b700000000ffffff34ffffffffffffff99ffffffff",
            INIT_08 => X"00000049000000000000006f00000000ffffff88ffffffffffffffe2ffffffff",
            INIT_09 => X"0000001c000000000000002b000000000000009300000000fffffffcffffffff",
            INIT_0A => X"0000000000000000fffffff6ffffffff0000001500000000ffffff98ffffffff",
            INIT_0B => X"0000000000000000ffffff6afffffffffffffff2ffffffff0000004100000000",
            INIT_0C => X"ffffffe6ffffffff0000000000000000ffffff9dffffffff0000000100000000",
            INIT_0D => X"ffffff8dffffffffffffffc0ffffffff0000005000000000ffffff3cffffffff",
            INIT_0E => X"ffffff8affffffff000000860000000000000068000000000000000700000000",
            INIT_0F => X"0000005100000000ffffffadffffffff00000006000000000000009500000000",
            INIT_10 => X"ffffffecffffffff0000007800000000ffffff89ffffffff0000000000000000",
            INIT_11 => X"ffffffa2ffffffff0000004a000000000000001e00000000ffffffe1ffffffff",
            INIT_12 => X"ffffff1affffffffffffffecffffffff0000003c00000000ffffff7effffffff",
            INIT_13 => X"00000006000000000000006d00000000ffffff7dffffffffffffff25ffffffff",
            INIT_14 => X"000000db000000000000006500000000ffffffedffffffff0000000400000000",
            INIT_15 => X"00000053000000000000004e000000000000000800000000fffffdf9ffffffff",
            INIT_16 => X"ffffff55ffffffff0000003d000000000000003800000000ffffffe7ffffffff",
            INIT_17 => X"00000010000000000000007700000000ffffff7effffffffffffffddffffffff",
            INIT_18 => X"ffffffe9ffffffff00000013000000000000000700000000fffffff4ffffffff",
            INIT_19 => X"0000003300000000ffffff9fffffffff0000002f00000000ffffffdfffffffff",
            INIT_1A => X"0000003c00000000ffffffafffffffffffffffb1ffffffffffffff75ffffffff",
            INIT_1B => X"00000000000000000000003c0000000000000003000000000000009b00000000",
            INIT_1C => X"ffffff77ffffffffffffff62ffffffffffffffedfffffffffffffecaffffffff",
            INIT_1D => X"ffffffceffffffffffffffedffffffffffffff98ffffffffffffff38ffffffff",
            INIT_1E => X"000000450000000000000002000000000000003c00000000ffffff2bffffffff",
            INIT_1F => X"0000001f00000000ffffffbeffffffff00000041000000000000005000000000",
            INIT_20 => X"ffffffe7ffffffff0000006900000000fffffeceffffffff0000000700000000",
            INIT_21 => X"0000000300000000ffffff62ffffffff0000001500000000ffffff95ffffffff",
            INIT_22 => X"0000004c000000000000001800000000ffffffdbffffffffffffff68ffffffff",
            INIT_23 => X"0000001800000000ffffffabffffffffffffffe3fffffffffffffea8ffffffff",
            INIT_24 => X"ffffffd1ffffffff0000001200000000ffffffdefffffffffffffffaffffffff",
            INIT_25 => X"ffffff32ffffffff00000004000000000000003300000000fffffff2ffffffff",
            INIT_26 => X"ffffffbaffffffffffffffe6ffffffff00000041000000000000001b00000000",
            INIT_27 => X"0000000300000000ffffffcaffffffff0000003400000000ffffffd0ffffffff",
            INIT_28 => X"ffffffceffffffffffffffd1ffffffff0000001200000000ffffffbfffffffff",
            INIT_29 => X"0000001f000000000000004a00000000fffffff5ffffffff0000000700000000",
            INIT_2A => X"ffffffebffffffff0000008c00000000ffffffdfffffffffffffff85ffffffff",
            INIT_2B => X"fffffff4ffffffffffffff72ffffffff0000001400000000ffffffb1ffffffff",
            INIT_2C => X"0000000500000000ffffffddffffffffffffffa3ffffffff0000001400000000",
            INIT_2D => X"fffffff1fffffffffffffffbffffffffffffffe1ffffffffffffffe7ffffffff",
            INIT_2E => X"0000001e00000000fffffff2ffffffff0000010500000000ffffffd8ffffffff",
            INIT_2F => X"ffffffb7ffffffff0000001e00000000ffffffd7ffffffff0000000200000000",
            INIT_30 => X"ffffffc8ffffffffffffffbdffffffffffffffeeffffffffffffffe8ffffffff",
            INIT_31 => X"0000001000000000ffffffc0ffffffffffffffbcffffffffffffffdcffffffff",
            INIT_32 => X"ffffff79ffffffff00000003000000000000002000000000ffffffadffffffff",
            INIT_33 => X"ffffffd7ffffffffffffff5dfffffffffffffff5ffffffffffffff84ffffffff",
            INIT_34 => X"ffffffdcffffffffffffffefffffffff0000001d000000000000000000000000",
            INIT_35 => X"ffffff97ffffffff0000001e000000000000005400000000ffffffd7ffffffff",
            INIT_36 => X"0000003100000000fffffff9ffffffffffffffa5ffffffffffffffeaffffffff",
            INIT_37 => X"0000000e00000000ffffffb3ffffffff00000054000000000000001700000000",
            INIT_38 => X"ffffffc4ffffffff0000006a00000000ffffffe0ffffffff0000003200000000",
            INIT_39 => X"0000005c000000000000002700000000ffffffe8ffffffff0000006000000000",
            INIT_3A => X"00000005000000000000005600000000ffffffe7ffffffffffffff9dffffffff",
            INIT_3B => X"0000000e00000000ffffffe9ffffffff0000000c00000000ffffffe8ffffffff",
            INIT_3C => X"00000022000000000000000400000000ffffffb0ffffffffffffff98ffffffff",
            INIT_3D => X"0000001400000000ffffffffffffffff00000008000000000000003700000000",
            INIT_3E => X"ffffffa0ffffffffffffffd1ffffffffffffffbdfffffffffffffffaffffffff",
            INIT_3F => X"ffffffe1ffffffffffffffb2fffffffffffffff9ffffffffffffffd3ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003100000000ffffff96ffffffffffffff91ffffffff0000000200000000",
            INIT_41 => X"0000006b00000000ffffffa8ffffffffffffff8bffffffffffffffd2ffffffff",
            INIT_42 => X"ffffffdeffffffffffffffeaffffffffffffffb9ffffffffffffffebffffffff",
            INIT_43 => X"ffffff85ffffffffffffff66ffffffffffffffbcffffffffffffffbbffffffff",
            INIT_44 => X"ffffffd2ffffffffffffffd0ffffffff00000078000000000000001300000000",
            INIT_45 => X"0000000f00000000ffffff71ffffffff0000000400000000ffffff9bffffffff",
            INIT_46 => X"0000000d00000000ffffffe8fffffffffffffffbfffffffffffffff6ffffffff",
            INIT_47 => X"ffffffecffffffff0000003e00000000ffffffa9ffffffff0000002500000000",
            INIT_48 => X"0000001100000000ffffff8fffffffffffffff79ffffffffffffff7effffffff",
            INIT_49 => X"0000008a000000000000000c00000000ffffffd7fffffffffffffff5ffffffff",
            INIT_4A => X"fffffffcffffffff0000005f00000000ffffffe0ffffffffffffff8cffffffff",
            INIT_4B => X"ffffffb9fffffffffffffff2fffffffffffffffaffffffff0000002700000000",
            INIT_4C => X"ffffffecffffffff0000003200000000ffffffadffffffff0000003400000000",
            INIT_4D => X"0000004b000000000000000700000000ffffff9fffffffff0000006200000000",
            INIT_4E => X"ffffffd7ffffffff00000010000000000000004300000000ffffffd3ffffffff",
            INIT_4F => X"ffffffdeffffffffffffffdfffffffffffffffbcffffffff0000004e00000000",
            INIT_50 => X"0000000500000000fffffffeffffffff0000001b00000000ffffffdeffffffff",
            INIT_51 => X"0000002700000000fffffff9ffffffffffffff97ffffffff0000002c00000000",
            INIT_52 => X"00000045000000000000000000000000ffffff95ffffffff0000001600000000",
            INIT_53 => X"fffffff3fffffffffffffea6ffffffff0000006d00000000ffffffcfffffffff",
            INIT_54 => X"ffffff9effffffff0000006900000000ffffff51ffffffffffffffecffffffff",
            INIT_55 => X"ffffffcbffffffff00000000000000000000004f00000000ffffff56ffffffff",
            INIT_56 => X"0000000d00000000000000bd00000000ffffffb8ffffffff0000001200000000",
            INIT_57 => X"0000000200000000ffffffa5ffffffff0000000b00000000ffffffe6ffffffff",
            INIT_58 => X"fffffff8fffffffffffffff0ffffffffffffff4fffffffffffffffcdffffffff",
            INIT_59 => X"0000003c000000000000001400000000ffffffecffffffff0000003100000000",
            INIT_5A => X"0000000600000000000000440000000000000046000000000000000100000000",
            INIT_5B => X"fffffff5ffffffff0000000200000000ffffffe9ffffffffffffffe8ffffffff",
            INIT_5C => X"0000002200000000ffffff72ffffffffffffffecffffffff0000000000000000",
            INIT_5D => X"ffffffe5fffffffffffffffbffffffffffffffe0fffffffffffffff5ffffffff",
            INIT_5E => X"fffffffdffffffffffffffe0ffffffffffffffc3ffffffff0000004d00000000",
            INIT_5F => X"ffffffc1ffffffff0000000c00000000fffffff5ffffffffffffffecffffffff",
            INIT_60 => X"0000001b000000000000002b000000000000006800000000ffffffecffffffff",
            INIT_61 => X"0000000700000000ffffffc8ffffffffffffff72ffffffffffffffedffffffff",
            INIT_62 => X"ffffff45ffffffffffffffe8ffffffff0000001900000000ffffffceffffffff",
            INIT_63 => X"ffffffb3ffffffffffffff70ffffffff0000006600000000ffffffdaffffffff",
            INIT_64 => X"ffffff9bffffffff0000002a00000000ffffffc0ffffffffffffffffffffffff",
            INIT_65 => X"fffffffbffffffff0000000f00000000ffffffe0ffffffffffffff86ffffffff",
            INIT_66 => X"ffffffc8ffffffffffffff7cffffffff0000002d000000000000000500000000",
            INIT_67 => X"fffffffdffffffffffffffe4ffffffffffffffaafffffffffffffff6ffffffff",
            INIT_68 => X"0000004400000000fffffff0ffffffff0000002f00000000ffffffeaffffffff",
            INIT_69 => X"ffffffecffffffff0000001a00000000fffffff6ffffffff0000004300000000",
            INIT_6A => X"00000053000000000000004d00000000ffffffd2ffffffffffffffb2ffffffff",
            INIT_6B => X"ffffffcfffffffffffffffffffffffffffffffe5fffffffffffffff8ffffffff",
            INIT_6C => X"0000002800000000ffffffb3ffffffffffffffc7ffffffff0000003000000000",
            INIT_6D => X"0000007f0000000000000029000000000000004a000000000000001e00000000",
            INIT_6E => X"0000003c00000000ffffffcaffffffffffffff95fffffffffffffff1ffffffff",
            INIT_6F => X"0000003b00000000ffffffcbffffffff00000000000000000000000400000000",
            INIT_70 => X"0000002e00000000ffffff5cffffffffffffffa0fffffffffffffff2ffffffff",
            INIT_71 => X"ffffffbfffffffffffffff68ffffffff0000002600000000ffffff7dffffffff",
            INIT_72 => X"0000000000000000ffffffebffffffffffffffb3ffffffffffffff7cffffffff",
            INIT_73 => X"ffffff64ffffffffffffffdeffffffff0000002d00000000000000c600000000",
            INIT_74 => X"ffffffd9ffffffff0000003a0000000000000017000000000000000d00000000",
            INIT_75 => X"ffffffc5ffffffff0000003200000000ffffffc6ffffffffffffff6dffffffff",
            INIT_76 => X"0000003a00000000ffffffdeffffffffffffffdbffffffff0000001000000000",
            INIT_77 => X"00000019000000000000001b0000000000000005000000000000000700000000",
            INIT_78 => X"0000004100000000ffffffdaffffffffffffff67ffffffffffffff45ffffffff",
            INIT_79 => X"ffffffccffffffff0000000f0000000000000001000000000000000d00000000",
            INIT_7A => X"0000004600000000000000500000000000000040000000000000007200000000",
            INIT_7B => X"ffffffe8ffffffffffffffdcffffffff0000000b000000000000003400000000",
            INIT_7C => X"ffffffeaffffffff0000005e00000000ffffff49ffffffff0000006800000000",
            INIT_7D => X"00000019000000000000003b00000000ffffffdbffffffff0000003500000000",
            INIT_7E => X"ffffffdcffffffff00000000000000000000000000000000ffffffe0ffffffff",
            INIT_7F => X"ffffffacffffffffffffffe5ffffffffffffffe7ffffffffffffffb9ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE2;


    MEM_IWGHT_LAYER3_INSTANCE3 : if BRAM_NAME = "iwght_layer3_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001c00000000ffffff9dffffffffffffff65ffffffff0000000400000000",
            INIT_01 => X"fffffff9ffffffffffffffe4ffffffffffffff95ffffffff0000005b00000000",
            INIT_02 => X"ffffffdfffffffff0000000a00000000ffffffb7ffffffff0000003600000000",
            INIT_03 => X"ffffff6dfffffffffffffe56ffffffff0000003500000000ffffff59ffffffff",
            INIT_04 => X"ffffffbaffffffff0000003f00000000ffffffdfffffffff0000001100000000",
            INIT_05 => X"ffffffb1ffffffff0000000b000000000000000e00000000fffffffdffffffff",
            INIT_06 => X"0000001f0000000000000081000000000000002f000000000000000600000000",
            INIT_07 => X"fffffffbffffffffffffff4fffffffffffffffefffffffff0000005400000000",
            INIT_08 => X"fffffff3ffffffff0000000e00000000ffffff55ffffffffffffffa8ffffffff",
            INIT_09 => X"00000010000000000000006f00000000ffffffa9ffffffffffffffc9ffffffff",
            INIT_0A => X"0000004e000000000000003d000000000000000b00000000ffffff3cffffffff",
            INIT_0B => X"ffffffa3ffffffff000000a1000000000000001200000000ffffffe1ffffffff",
            INIT_0C => X"0000000a00000000000000a7000000000000005800000000fffffea2ffffffff",
            INIT_0D => X"ffffffb1ffffffff000000070000000000000008000000000000001600000000",
            INIT_0E => X"0000000f00000000ffffff85fffffffffffffee9ffffffff0000001400000000",
            INIT_0F => X"0000003500000000fffffffaffffffffffffff87ffffffff0000002e00000000",
            INIT_10 => X"0000004c00000000ffffff6dffffffff0000000d000000000000001100000000",
            INIT_11 => X"0000001a00000000ffffff7cffffffffffffffcaffffffff0000003d00000000",
            INIT_12 => X"ffffff7bffffffff0000000a00000000fffffffaffffffff0000003d00000000",
            INIT_13 => X"ffffff91ffffffff0000002700000000ffffffcdffffffff0000003900000000",
            INIT_14 => X"ffffffb2ffffffff00000002000000000000005f00000000ffffffe6ffffffff",
            INIT_15 => X"000000850000000000000016000000000000000000000000000000ae00000000",
            INIT_16 => X"0000000d00000000ffffffc7ffffffff0000001400000000ffffffe8ffffffff",
            INIT_17 => X"fffffff9ffffffffffffff7fffffffff0000001e00000000fffffffdffffffff",
            INIT_18 => X"0000001a00000000ffffffcefffffffffffffff4ffffffffffffff9effffffff",
            INIT_19 => X"ffffffceffffffff0000001500000000ffffff73ffffffffffffffffffffffff",
            INIT_1A => X"ffffffcdffffffff0000000e00000000ffffffb0ffffffffffffff83ffffffff",
            INIT_1B => X"ffffffabffffffff0000001a000000000000001800000000ffffffe0ffffffff",
            INIT_1C => X"ffffff82ffffffff0000001600000000fffffff9fffffffffffffefaffffffff",
            INIT_1D => X"ffffffd1ffffffff0000004a0000000000000005000000000000000000000000",
            INIT_1E => X"fffffff3ffffffffffffffccffffffffffffffadffffffff0000005300000000",
            INIT_1F => X"0000004300000000ffffffd4ffffffffffffffaeffffffff0000000300000000",
            INIT_20 => X"0000003f00000000ffffffa9fffffffffffffffdffffffff0000001300000000",
            INIT_21 => X"ffffffe4ffffffffffffffa8ffffffffffffff5dffffffff0000001800000000",
            INIT_22 => X"0000002200000000ffffffecffffffffffffffc2ffffffff0000000700000000",
            INIT_23 => X"ffffff99ffffffff000000a1000000000000004c00000000000000d300000000",
            INIT_24 => X"ffffffbbfffffffffffffffcffffffff00000035000000000000000900000000",
            INIT_25 => X"ffffff39ffffffff0000000c000000000000001c000000000000001600000000",
            INIT_26 => X"ffffffebffffffffffffffaaffffffffffffffa9ffffffff0000001000000000",
            INIT_27 => X"0000000600000000ffffffcbffffffff0000000e000000000000001e00000000",
            INIT_28 => X"ffffffedffffffffffffffd2ffffffffffffff7dffffffffffffffaaffffffff",
            INIT_29 => X"ffffffe1ffffffff000000240000000000000000000000000000001b00000000",
            INIT_2A => X"0000001a00000000000000a500000000ffffffa7ffffffffffffffb1ffffffff",
            INIT_2B => X"0000005a00000000ffffffdcffffffff0000000500000000ffffffacffffffff",
            INIT_2C => X"00000001000000000000005100000000ffffffe1ffffffffffffff0cffffffff",
            INIT_2D => X"ffffffbcffffffff0000002a0000000000000049000000000000004600000000",
            INIT_2E => X"ffffff7bffffffffffffffbdfffffffffffffecdffffffff0000003c00000000",
            INIT_2F => X"ffffffdcffffffffffffffdcffffffffffffff8fffffffffffffffb9ffffffff",
            INIT_30 => X"0000004100000000ffffffeeffffffff0000000400000000fffffffdffffffff",
            INIT_31 => X"0000000d000000000000000200000000ffffff1dffffffff0000001500000000",
            INIT_32 => X"fffffff0fffffffffffffff6ffffffffffffff83ffffffff0000003f00000000",
            INIT_33 => X"ffffffc8fffffffffffffefcffffffffffffffe4ffffffffffffff3fffffffff",
            INIT_34 => X"ffffffc5ffffffffffffffeaffffffffffffffe5ffffffffffffffffffffffff",
            INIT_35 => X"ffffff9effffffff0000002f00000000ffffffb1ffffffffffffffecffffffff",
            INIT_36 => X"0000003700000000ffffffe5fffffffffffffffaffffffff0000000e00000000",
            INIT_37 => X"fffffff8ffffffffffffffc7ffffffffffffffb5ffffffff0000000000000000",
            INIT_38 => X"0000005300000000ffffffbfffffffffffffffecffffffffffffffe0ffffffff",
            INIT_39 => X"fffffffaffffffffffffffe3ffffffff00000007000000000000005400000000",
            INIT_3A => X"fffffff4ffffffff0000004600000000ffffffb5ffffffffffffff8bffffffff",
            INIT_3B => X"ffffffd1ffffffff0000000b00000000fffffff2ffffffffffffffa7ffffffff",
            INIT_3C => X"0000004000000000ffffffbdffffffffffffffe7ffffffffffffffddffffffff",
            INIT_3D => X"0000001e000000000000000f00000000ffffffb0ffffffff0000002400000000",
            INIT_3E => X"0000000e00000000ffffffeaffffffffffffff6ffffffffffffffffaffffffff",
            INIT_3F => X"ffffffb3ffffffffffffffe8ffffffff0000005600000000ffffffebffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffd9ffffffff0000005800000000fffffff3ffffffff0000000400000000",
            INIT_41 => X"ffffffeaffffffffffffffdffffffffffffffff6ffffffffffffffcbffffffff",
            INIT_42 => X"ffffffceffffffffffffffe9ffffffff0000003b00000000ffffffecffffffff",
            INIT_43 => X"ffffffc3ffffffffffffff70ffffffffffffffaaffffffffffffffa6ffffffff",
            INIT_44 => X"00000001000000000000000700000000ffffffecffffffff0000000000000000",
            INIT_45 => X"ffffffe7ffffffffffffffe0ffffffff00000053000000000000000800000000",
            INIT_46 => X"fffffff1fffffffffffffff3fffffffffffffffbfffffffffffffffbffffffff",
            INIT_47 => X"ffffffe6ffffffffffffffc3ffffffffffffffdbffffffffffffffeeffffffff",
            INIT_48 => X"0000002000000000ffffff86ffffffff0000002b00000000ffffffe9ffffffff",
            INIT_49 => X"fffffff7ffffffff000000400000000000000014000000000000001600000000",
            INIT_4A => X"ffffffafffffffff0000001e00000000fffffff5ffffffffffffff76ffffffff",
            INIT_4B => X"ffffffbdffffffffffffffe6ffffffffffffffedffffffffffffffdaffffffff",
            INIT_4C => X"0000002100000000ffffff5fffffffff00000005000000000000005a00000000",
            INIT_4D => X"0000002d000000000000000f00000000ffffffe9ffffffff0000000e00000000",
            INIT_4E => X"000000000000000000000039000000000000000400000000ffffffb1ffffffff",
            INIT_4F => X"ffffffe4ffffffff00000032000000000000002600000000ffffffb1ffffffff",
            INIT_50 => X"ffffffc5ffffffffffffffddffffffff0000003500000000fffffffcffffffff",
            INIT_51 => X"ffffffcfffffffffffffffb8ffffffffffffffafffffffff0000006600000000",
            INIT_52 => X"fffffff0ffffffff00000008000000000000000d000000000000001d00000000",
            INIT_53 => X"ffffffd2ffffffffffffffabffffffffffffffbaffffffffffffff2cffffffff",
            INIT_54 => X"ffffff94ffffffff0000001700000000fffffff4ffffffffffffffeeffffffff",
            INIT_55 => X"0000002e0000000000000001000000000000000000000000ffffff8bffffffff",
            INIT_56 => X"ffffffdeffffffffffffffe4ffffffff0000004200000000fffffff5ffffffff",
            INIT_57 => X"ffffffe1ffffffff000000310000000000000022000000000000001500000000",
            INIT_58 => X"0000001b00000000ffffffcdffffffffffffffd4ffffffffffffffceffffffff",
            INIT_59 => X"ffffffd8ffffffff00000025000000000000000a00000000fffffffeffffffff",
            INIT_5A => X"ffffffceffffffffffffff82fffffffffffffff7ffffffffffffff91ffffffff",
            INIT_5B => X"ffffffd6ffffffffffffffb9ffffffffffffffe9ffffffff0000001400000000",
            INIT_5C => X"0000000d00000000ffffffd1ffffffffffffffd1ffffffffffffff6fffffffff",
            INIT_5D => X"00000000000000000000000e00000000ffffffd1ffffffff0000002f00000000",
            INIT_5E => X"ffffffffffffffffffffffd9ffffffffffffff66ffffffff0000001000000000",
            INIT_5F => X"ffffff87ffffffff0000000d00000000ffffffdfffffffff0000005200000000",
            INIT_60 => X"ffffffdcffffffffffffffe4ffffffff0000001c00000000ffffffe5ffffffff",
            INIT_61 => X"0000001900000000ffffff8cffffffff0000001400000000ffffff93ffffffff",
            INIT_62 => X"ffffffdeffffffff00000004000000000000003e000000000000000600000000",
            INIT_63 => X"0000004b000000000000009400000000fffffffaffffffff0000002d00000000",
            INIT_64 => X"0000001800000000ffffffe7ffffffffffffffb7fffffffffffffff4ffffffff",
            INIT_65 => X"ffffff70fffffffffffffff7ffffffff00000045000000000000004000000000",
            INIT_66 => X"0000000600000000ffffff93fffffffffffffff2ffffffff0000000e00000000",
            INIT_67 => X"0000000e00000000000000160000000000000015000000000000005200000000",
            INIT_68 => X"0000002400000000ffffffbaffffffffffffffe1ffffffffffffffb1ffffffff",
            INIT_69 => X"0000002b000000000000001100000000ffffffbaffffffffffffffd8ffffffff",
            INIT_6A => X"ffffffe2ffffffff00000050000000000000007400000000ffffffd4ffffffff",
            INIT_6B => X"fffffff1ffffffffffffffaaffffffff0000000100000000ffffffeaffffffff",
            INIT_6C => X"ffffffdfffffffff0000001d00000000ffffffb7fffffffffffffeb2ffffffff",
            INIT_6D => X"0000003400000000fffffff2ffffffffffffff8affffffff0000002500000000",
            INIT_6E => X"ffffffadffffffffffffffbaffffffffffffffd1ffffffffffffffcdffffffff",
            INIT_6F => X"ffffffd8ffffffffffffff3affffffff0000001000000000ffffffc4ffffffff",
            INIT_70 => X"ffffff85ffffffffffffff9effffffff0000003300000000fffffff6ffffffff",
            INIT_71 => X"0000002500000000ffffffebffffffff0000003100000000ffffff7affffffff",
            INIT_72 => X"ffffffdbffffffff0000000e00000000ffffffc4ffffffff0000001400000000",
            INIT_73 => X"0000000400000000ffffff94ffffffffffffff9affffffff0000003900000000",
            INIT_74 => X"ffffff98ffffffff00000008000000000000002b000000000000000300000000",
            INIT_75 => X"0000000f00000000000000200000000000000058000000000000007a00000000",
            INIT_76 => X"ffffffdeffffffffffffff80ffffffffffffffd0ffffffff0000000000000000",
            INIT_77 => X"fffffff3ffffffffffffffafffffffff0000003a00000000ffffffd0ffffffff",
            INIT_78 => X"fffffff5ffffffffffffff70fffffffffffffffeffffffffffffffa9ffffffff",
            INIT_79 => X"00000000000000000000004200000000ffffffc1ffffffffffffffeeffffffff",
            INIT_7A => X"ffffff97ffffffffffffffe9fffffffffffffffbffffffff0000000000000000",
            INIT_7B => X"0000003f000000000000002800000000ffffffecffffffffffffff8affffffff",
            INIT_7C => X"ffffffeaffffffff00000006000000000000001000000000fffffff6ffffffff",
            INIT_7D => X"00000026000000000000000700000000ffffff8fffffffff0000001800000000",
            INIT_7E => X"0000000100000000ffffff51ffffffffffffff86ffffffff0000003d00000000",
            INIT_7F => X"ffffffa3ffffffffffffffe1ffffffffffffffddffffffff0000002e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE3;


    MEM_IWGHT_LAYER3_INSTANCE4 : if BRAM_NAME = "iwght_layer3_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffadffffffffffffff13ffffffff0000003b00000000ffffffeaffffffff",
            INIT_01 => X"00000022000000000000002f00000000ffffffaeffffffffffffffa8ffffffff",
            INIT_02 => X"00000000000000000000000f0000000000000036000000000000001100000000",
            INIT_03 => X"ffffffd9ffffffffffffffb2ffffffffffffffbbffffffffffffffe8ffffffff",
            INIT_04 => X"ffffffcaffffffff00000000000000000000001a000000000000000100000000",
            INIT_05 => X"0000000b0000000000000000000000000000001e000000000000001a00000000",
            INIT_06 => X"ffffffeeffffffffffffff9affffffffffffffcfffffffff0000001500000000",
            INIT_07 => X"0000001400000000ffffffeeffffffff0000002500000000ffffffe4ffffffff",
            INIT_08 => X"0000000200000000ffffffb7ffffffff0000007200000000ffffffa8ffffffff",
            INIT_09 => X"ffffffc9ffffffff0000005300000000ffffffd6ffffffffffffffdfffffffff",
            INIT_0A => X"ffffffdaffffffffffffffd1ffffffffffffff9bffffffffffffffa2ffffffff",
            INIT_0B => X"00000005000000000000003700000000ffffffeeffffffffffffffe5ffffffff",
            INIT_0C => X"0000002e000000000000000000000000fffffffeffffffffffffffd3ffffffff",
            INIT_0D => X"0000003300000000ffffffd5ffffffffffffff5ffffffffffffffffcffffffff",
            INIT_0E => X"0000001f000000000000005b00000000ffffff99ffffffff0000001200000000",
            INIT_0F => X"ffffffabffffffffffffffe7fffffffffffffff6ffffffffffffffeeffffffff",
            INIT_10 => X"ffffffd3ffffffffffffffeeffffffff00000070000000000000000100000000",
            INIT_11 => X"0000000500000000fffffff5ffffffffffffff67ffffffffffffffe3ffffffff",
            INIT_12 => X"ffffffc9ffffffff00000016000000000000002500000000fffffffbffffffff",
            INIT_13 => X"0000002800000000000000750000000000000010000000000000007a00000000",
            INIT_14 => X"ffffffdeffffffff0000002000000000ffffffadffffffff0000001700000000",
            INIT_15 => X"ffffff95fffffffffffffffffffffffffffffff7ffffffff0000000f00000000",
            INIT_16 => X"0000005d0000000000000004000000000000000200000000fffffff9ffffffff",
            INIT_17 => X"0000001400000000ffffffd8ffffffff0000001300000000ffffff95ffffffff",
            INIT_18 => X"0000000500000000000000590000000000000018000000000000000500000000",
            INIT_19 => X"0000003400000000ffffffb0ffffffffffffff8bffffffff0000003800000000",
            INIT_1A => X"fffffff7ffffffff00000007000000000000000a00000000ffffff93ffffffff",
            INIT_1B => X"0000003a000000000000001100000000fffffff4ffffffff0000001300000000",
            INIT_1C => X"ffffffdaffffffffffffffb5ffffffffffffffddffffffffffffffc7ffffffff",
            INIT_1D => X"0000003d000000000000001000000000ffffffb3ffffffff0000005900000000",
            INIT_1E => X"00000002000000000000004b00000000ffffffb4ffffffffffffff9dffffffff",
            INIT_1F => X"fffffffcffffffffffffffa0ffffffffffffffd6ffffffff0000000000000000",
            INIT_20 => X"ffffffe6ffffffffffffffd2ffffffffffffffd9fffffffffffffff6ffffffff",
            INIT_21 => X"0000000000000000ffffff67ffffffff00000029000000000000003000000000",
            INIT_22 => X"00000051000000000000001900000000ffffffa7ffffffff0000000100000000",
            INIT_23 => X"fffffffaffffffffffffff99ffffffffffffff96ffffffffffffff8dffffffff",
            INIT_24 => X"ffffffd0ffffffffffffffd5fffffffffffffffbffffffff0000001e00000000",
            INIT_25 => X"ffffff88ffffffff0000001a00000000ffffffedffffffff0000006600000000",
            INIT_26 => X"0000000d000000000000002500000000ffffffcaffffffff0000001500000000",
            INIT_27 => X"fffffff4fffffffffffffff6ffffffff0000003b00000000ffffff84ffffffff",
            INIT_28 => X"0000000b000000000000000f00000000fffffff6ffffffffffffff9fffffffff",
            INIT_29 => X"fffffff1ffffffff0000001700000000ffffffbdffffffffffffffbbffffffff",
            INIT_2A => X"ffffffc8ffffffffffffff78ffffffffffffffeeffffffff0000002600000000",
            INIT_2B => X"fffffffeffffffffffffffa4ffffffff0000000000000000ffffffe4ffffffff",
            INIT_2C => X"0000004600000000ffffffe5fffffffffffffff1ffffffffffffff77ffffffff",
            INIT_2D => X"fffffffeffffffffffffffcaffffffff00000000000000000000000200000000",
            INIT_2E => X"fffffffcffffffffffffffe2ffffffff0000002400000000ffffffbdffffffff",
            INIT_2F => X"ffffffacffffffffffffffe4fffffffffffffff4ffffffff0000000000000000",
            INIT_30 => X"0000004200000000ffffffd8ffffffffffffffe1fffffffffffffffeffffffff",
            INIT_31 => X"0000005d000000000000000900000000ffffffebffffffff0000000b00000000",
            INIT_32 => X"0000004700000000fffffffcfffffffffffffff0ffffffff0000001300000000",
            INIT_33 => X"ffffffc5ffffffffffffff57ffffffffffffffeeffffffff0000000100000000",
            INIT_34 => X"ffffffb7ffffffffffffffdfffffffffffffffe9fffffffffffffff5ffffffff",
            INIT_35 => X"00000040000000000000004400000000ffffffcaffffffff0000000300000000",
            INIT_36 => X"ffffffefffffffffffffffe9ffffffff0000003100000000fffffff2ffffffff",
            INIT_37 => X"fffffffdffffffffffffffebffffffff0000005300000000ffffffd0ffffffff",
            INIT_38 => X"ffffffdeffffffffffffffebffffffff0000001b00000000ffffffe5ffffffff",
            INIT_39 => X"ffffffc4ffffffff0000003500000000ffffffeeffffffff0000000b00000000",
            INIT_3A => X"ffffffe7ffffffffffffffbeffffffff00000042000000000000005b00000000",
            INIT_3B => X"ffffffd6fffffffffffffff3ffffffff0000000600000000ffffffc2ffffffff",
            INIT_3C => X"00000036000000000000001e00000000ffffffd8ffffffffffffffe8ffffffff",
            INIT_3D => X"0000002300000000ffffffdaffffffff00000022000000000000001700000000",
            INIT_3E => X"0000002100000000ffffffe0ffffffffffffffd0ffffffff0000001700000000",
            INIT_3F => X"ffffff8affffffffffffffa2ffffffffffffff86ffffffffffffffeaffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffe5fffffffffffffffaffffffff0000000500000000ffffffdaffffffff",
            INIT_41 => X"fffffff7ffffffffffffffeaffffffffffffff1dfffffffffffffff2ffffffff",
            INIT_42 => X"ffffffb9fffffffffffffff4fffffffffffffff0ffffffffffffffc6ffffffff",
            INIT_43 => X"ffffffb2ffffffffffffffd7ffffffff0000000f000000000000000500000000",
            INIT_44 => X"0000004200000000ffffffa2ffffffffffffffc0fffffffffffffffeffffffff",
            INIT_45 => X"000000260000000000000039000000000000003500000000ffffffe6ffffffff",
            INIT_46 => X"0000002d000000000000005500000000fffffff8fffffffffffffff7ffffffff",
            INIT_47 => X"0000000400000000ffffffd4ffffffffffffffe7ffffffffffffff97ffffffff",
            INIT_48 => X"ffffffddffffffffffffff94ffffffff0000004f00000000ffffffe6ffffffff",
            INIT_49 => X"00000024000000000000005300000000ffffffd3ffffffffffffff89ffffffff",
            INIT_4A => X"ffffff81fffffffffffffef4ffffffffffffff83ffffffff0000003700000000",
            INIT_4B => X"00000004000000000000002900000000fffffffeffffffff0000003a00000000",
            INIT_4C => X"ffffffafffffffffffffffe4ffffffff00000007000000000000000000000000",
            INIT_4D => X"0000003000000000ffffffa2ffffffffffffffdfffffffffffffffdeffffffff",
            INIT_4E => X"0000000700000000ffffffdaffffffffffffff9effffffffffffffb9ffffffff",
            INIT_4F => X"00000020000000000000003f00000000ffffffeeffffffffffffff94ffffffff",
            INIT_50 => X"ffffffe2ffffffffffffffa1ffffffff0000005a000000000000001100000000",
            INIT_51 => X"ffffff95ffffffff0000006400000000ffffff6bffffffff0000008200000000",
            INIT_52 => X"00000003000000000000001200000000ffffffb5ffffffffffffffe7ffffffff",
            INIT_53 => X"ffffff7dffffffff0000004000000000ffffffaafffffffffffffea2ffffffff",
            INIT_54 => X"0000000000000000fffffff3ffffffffffffffe8ffffffff0000000700000000",
            INIT_55 => X"ffffffcdffffffff00000019000000000000007600000000ffffffbcffffffff",
            INIT_56 => X"ffffffdcffffffffffffffddffffffffffffff2affffffff0000001500000000",
            INIT_57 => X"ffffffeaffffffffffffffd3ffffffffffffffefffffffffffffff72ffffffff",
            INIT_58 => X"0000002f00000000ffffff7cffffffffffffffd2ffffffffffffffb4ffffffff",
            INIT_59 => X"00000020000000000000002b00000000ffffffb8ffffffffffffff84ffffffff",
            INIT_5A => X"0000007700000000ffffff0dffffffffffffffe2ffffffff0000003300000000",
            INIT_5B => X"ffffffe9ffffffff00000042000000000000000a000000000000003400000000",
            INIT_5C => X"00000021000000000000001b000000000000005c000000000000001d00000000",
            INIT_5D => X"ffffffc2ffffffffffffff8cffffffffffffffccffffffffffffffa4ffffffff",
            INIT_5E => X"ffffff5effffffffffffffd6fffffffffffffefdffffffff0000001900000000",
            INIT_5F => X"ffffffefffffffff0000001a0000000000000085000000000000002200000000",
            INIT_60 => X"ffffff8bffffffff000000550000000000000082000000000000001200000000",
            INIT_61 => X"ffffffb6ffffffffffffffeeffffffff0000003400000000ffffffd1ffffffff",
            INIT_62 => X"ffffffd6ffffffffffffffffffffffffffffffa1ffffffffffffffecffffffff",
            INIT_63 => X"ffffffc6fffffffffffffff7ffffffffffffffb9ffffffffffffffd2ffffffff",
            INIT_64 => X"ffffff9dffffffff0000003200000000ffffffafffffffff0000000500000000",
            INIT_65 => X"ffffff84fffffffffffffffbfffffffffffffffdffffffff0000002b00000000",
            INIT_66 => X"ffffffd6ffffffffffffffb3ffffffffffffff97fffffffffffffffcffffffff",
            INIT_67 => X"fffffff2ffffffff00000014000000000000003f00000000ffffffdeffffffff",
            INIT_68 => X"ffffffe0ffffffffffffffbbffffffff00000064000000000000002c00000000",
            INIT_69 => X"0000001d000000000000005800000000ffffffaaffffffffffffffbeffffffff",
            INIT_6A => X"0000003500000000ffffff8cffffffffffffffedffffffff0000004d00000000",
            INIT_6B => X"0000005c00000000ffffffbaffffffffffffffe6ffffffff0000004800000000",
            INIT_6C => X"ffffff78ffffffffffffffdbffffffff0000000400000000ffffff87ffffffff",
            INIT_6D => X"ffffff68fffffffffffffffcffffffff0000002200000000ffffff86ffffffff",
            INIT_6E => X"ffffffa8fffffffffffffff7ffffffffffffff89ffffffffffffffccffffffff",
            INIT_6F => X"0000001d0000000000000000000000000000003c000000000000002800000000",
            INIT_70 => X"ffffffbaffffffffffffff8bffffffffffffffebffffffffffffffeeffffffff",
            INIT_71 => X"0000000a000000000000005900000000ffffff6ffffffffffffffff8ffffffff",
            INIT_72 => X"0000002e00000000ffffffffffffffff00000014000000000000004a00000000",
            INIT_73 => X"ffffffdfffffffffffffffacffffffffffffff8ffffffffffffffff0ffffffff",
            INIT_74 => X"00000029000000000000003100000000ffffffc4fffffffffffffffaffffffff",
            INIT_75 => X"ffffff8cffffffffffffffe5ffffffffffffffe5ffffffffffffff6dffffffff",
            INIT_76 => X"0000002700000000fffffff5ffffffffffffffe3ffffffff0000000600000000",
            INIT_77 => X"ffffffedffffffffffffffd5ffffffff0000002800000000ffffffacffffffff",
            INIT_78 => X"fffffff2ffffffff00000051000000000000000900000000000000a100000000",
            INIT_79 => X"00000044000000000000000300000000ffffffb1ffffffffffffff84ffffffff",
            INIT_7A => X"ffffffaeffffffff0000001e00000000fffffffaffffffff000000a300000000",
            INIT_7B => X"0000001b000000000000001900000000fffffffbffffffff0000002900000000",
            INIT_7C => X"0000002e0000000000000064000000000000003f000000000000007000000000",
            INIT_7D => X"0000004d000000000000002a000000000000004300000000ffffffc0ffffffff",
            INIT_7E => X"0000001f00000000ffffffc0ffffffffffffff1dffffffffffffffb0ffffffff",
            INIT_7F => X"00000037000000000000000700000000ffffff9effffffffffffffb4ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE4;


    MEM_IWGHT_LAYER3_INSTANCE5 : if BRAM_NAME = "iwght_layer3_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003800000000ffffff7effffffff00000019000000000000000200000000",
            INIT_01 => X"ffffff38ffffffffffffffdfffffffff00000011000000000000001e00000000",
            INIT_02 => X"fffffffcfffffffffffffffdffffffff0000004000000000ffffffdeffffffff",
            INIT_03 => X"ffffff96ffffffffffffff2bffffffffffffffaaffffffff0000000800000000",
            INIT_04 => X"ffffffffffffffffffffffe2ffffffffffffff99fffffffffffffff1ffffffff",
            INIT_05 => X"0000002c00000000ffffffa5ffffffff0000003400000000ffffffdcffffffff",
            INIT_06 => X"0000003200000000ffffff2fffffffffffffff97ffffffff0000001200000000",
            INIT_07 => X"0000000d00000000ffffffd5ffffffffffffffe0ffffffffffffff3fffffffff",
            INIT_08 => X"ffffffadffffffff0000000e00000000ffffff7affffffff000000ab00000000",
            INIT_09 => X"ffffffd2ffffffff0000002000000000ffffff45ffffffff0000004300000000",
            INIT_0A => X"ffffffe7ffffffff0000000000000000ffffffc6ffffffffffffffddffffffff",
            INIT_0B => X"fffffff9ffffffff000000160000000000000016000000000000003b00000000",
            INIT_0C => X"0000000b0000000000000004000000000000003f00000000ffffff99ffffffff",
            INIT_0D => X"00000028000000000000004b00000000ffffff85ffffffffffffffc4ffffffff",
            INIT_0E => X"0000002800000000ffffffe6ffffffffffffff0affffffffffffff94ffffffff",
            INIT_0F => X"0000003f00000000ffffffb0ffffffff0000006800000000ffffffd6ffffffff",
            INIT_10 => X"ffffff74ffffffffffffffc4ffffffffffffffe1fffffffffffffffaffffffff",
            INIT_11 => X"ffffff6cffffffffffffff7dffffffffffffffafffffffffffffffcbffffffff",
            INIT_12 => X"fffffff4fffffffffffffff3ffffffff00000027000000000000003500000000",
            INIT_13 => X"ffffffb3ffffffff0000000e00000000ffffffd1ffffffff0000003e00000000",
            INIT_14 => X"0000001600000000ffffffbdffffffffffffffe1ffffffffffffffebffffffff",
            INIT_15 => X"ffffffcbffffffffffffff8affffffff0000000d00000000ffffffe1ffffffff",
            INIT_16 => X"0000005600000000ffffffe5ffffffffffffff65ffffffff0000000d00000000",
            INIT_17 => X"0000000600000000ffffffe3ffffffff0000001900000000ffffff92ffffffff",
            INIT_18 => X"00000037000000000000000600000000ffffffdbffffffff000000ae00000000",
            INIT_19 => X"ffffffc7ffffffff0000005000000000ffffffceffffffff0000003e00000000",
            INIT_1A => X"0000001100000000ffffffc9ffffffff0000000900000000ffffffb9ffffffff",
            INIT_1B => X"0000003900000000ffffffd2ffffffff00000017000000000000003a00000000",
            INIT_1C => X"fffffff6ffffffff00000038000000000000003c00000000ffffffcfffffffff",
            INIT_1D => X"0000000c000000000000005300000000ffffffdaffffffff0000000200000000",
            INIT_1E => X"0000000f00000000ffffffe2ffffffff0000003600000000fffffff2ffffffff",
            INIT_1F => X"0000004300000000ffffffeeffffffff0000008a00000000ffffffc5ffffffff",
            INIT_20 => X"fffffff3fffffffffffffffcffffffffffffffc8ffffffff0000000500000000",
            INIT_21 => X"ffffffaeffffffffffffff87fffffffffffffee9ffffffff0000004c00000000",
            INIT_22 => X"ffffffeaffffffff000000160000000000000024000000000000006400000000",
            INIT_23 => X"ffffffaeffffffffffffff2effffffffffffff92fffffffffffffffeffffffff",
            INIT_24 => X"ffffffc6ffffffffffffff4effffffffffffff47ffffffff0000000100000000",
            INIT_25 => X"0000001200000000000000080000000000000004000000000000003a00000000",
            INIT_26 => X"ffffff9bffffffffffffffeeffffffffffffffc3fffffffffffffff9ffffffff",
            INIT_27 => X"0000001600000000ffffffd4ffffffff0000003100000000ffffffd5ffffffff",
            INIT_28 => X"fffffff5ffffffff000000640000000000000017000000000000007c00000000",
            INIT_29 => X"0000002c000000000000000d00000000ffffffb0ffffffffffffff88ffffffff",
            INIT_2A => X"ffffffecfffffffffffffff0ffffffff0000001000000000ffffff70ffffffff",
            INIT_2B => X"ffffffd3ffffffff00000069000000000000001200000000fffffff9ffffffff",
            INIT_2C => X"ffffffddffffffff00000001000000000000003b000000000000003800000000",
            INIT_2D => X"ffffffbaffffffff0000001a000000000000003c00000000ffffffcaffffffff",
            INIT_2E => X"ffffffa6ffffffffffffffa0ffffffff000000af000000000000002600000000",
            INIT_2F => X"00000023000000000000002700000000ffffff5cffffffff0000001d00000000",
            INIT_30 => X"ffffff37fffffffffffffff0ffffffffffffff5cffffffffffffffeeffffffff",
            INIT_31 => X"ffffffa2ffffffff0000004d00000000ffffffe3fffffffffffffffeffffffff",
            INIT_32 => X"0000006600000000fffffffaffffffff00000030000000000000004200000000",
            INIT_33 => X"ffffffcdffffffffffffffb4ffffffffffffffaaffffffffffffffadffffffff",
            INIT_34 => X"ffffffc0ffffffffffffff8affffffffffffff76ffffffffffffffe6ffffffff",
            INIT_35 => X"ffffff3fffffffffffffffa5ffffffffffffffe9ffffffff000000bd00000000",
            INIT_36 => X"0000002600000000ffffffc4ffffffffffffffd7fffffffffffffff1ffffffff",
            INIT_37 => X"ffffffeefffffffffffffffdffffffff0000000d00000000ffffff71ffffffff",
            INIT_38 => X"0000001b000000000000000d00000000ffffffd0ffffffffffffffb6ffffffff",
            INIT_39 => X"00000001000000000000000e00000000ffffff4fffffffff0000000b00000000",
            INIT_3A => X"ffffffb0ffffffffffffff9cffffffffffffffd2ffffffffffffff37ffffffff",
            INIT_3B => X"ffffff75ffffffffffffffd4ffffffff00000004000000000000001800000000",
            INIT_3C => X"ffffffbbffffffffffffffb3ffffffff0000006200000000ffffff5affffffff",
            INIT_3D => X"ffffffa5ffffffff0000001800000000ffffffafffffffff0000002300000000",
            INIT_3E => X"ffffffcdffffffffffffffe7ffffffffffffffc2ffffffff0000001000000000",
            INIT_3F => X"0000005b0000000000000004000000000000002200000000ffffffb3ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffff5affffffffffffff8bffffffffffffffe2ffffffff0000000100000000",
            INIT_41 => X"ffffffdcffffffffffffff91ffffffffffffff67ffffffffffffffe5ffffffff",
            INIT_42 => X"00000025000000000000000b0000000000000024000000000000002a00000000",
            INIT_43 => X"fffffff3ffffffffffffffa0ffffffffffffffbbffffffffffffffd9ffffffff",
            INIT_44 => X"0000003a00000000ffffff33ffffffff00000007000000000000000100000000",
            INIT_45 => X"0000003800000000ffffffdfffffffffffffffe4ffffffff0000009c00000000",
            INIT_46 => X"0000001600000000ffffffc0ffffffffffffff58fffffffffffffff7ffffffff",
            INIT_47 => X"0000001800000000ffffffeeffffffffffffffd2ffffffffffffff9effffffff",
            INIT_48 => X"0000005300000000ffffffd5ffffffffffffffd0ffffffff0000009a00000000",
            INIT_49 => X"00000028000000000000002b00000000ffffffa2ffffffff0000000700000000",
            INIT_4A => X"ffffffb0ffffffff00000070000000000000001d00000000fffffe62ffffffff",
            INIT_4B => X"00000031000000000000001000000000fffffff5ffffffffffffffd6ffffffff",
            INIT_4C => X"ffffffbaffffffff00000058000000000000002200000000ffffffc0ffffffff",
            INIT_4D => X"0000002000000000ffffffc1ffffffffffffffc8ffffffff0000001400000000",
            INIT_4E => X"ffffffedffffffffffffff69ffffffff0000001b000000000000000000000000",
            INIT_4F => X"00000011000000000000002500000000ffffffc6ffffffffffffffe0ffffffff",
            INIT_50 => X"ffffffdeffffffffffffff5fffffffff00000026000000000000000200000000",
            INIT_51 => X"ffffffd3ffffffffffffffe7fffffffffffffea7ffffffff0000001800000000",
            INIT_52 => X"ffffffbafffffffffffffff0fffffffffffffff0ffffffff0000002a00000000",
            INIT_53 => X"0000003900000000ffffff8fffffffffffffffb2ffffffffffffff82ffffffff",
            INIT_54 => X"ffffffb1ffffffffffffffefffffffffffffffc0ffffffff0000000f00000000",
            INIT_55 => X"0000000a000000000000004100000000ffffffd4ffffffffffffffc5ffffffff",
            INIT_56 => X"ffffffccffffffffffffffa7ffffffff0000006800000000fffffffbffffffff",
            INIT_57 => X"0000000400000000fffffff7ffffffff0000000800000000ffffffe8ffffffff",
            INIT_58 => X"fffffff6ffffffffffffffdfffffffffffffffc7ffffffffffffffd2ffffffff",
            INIT_59 => X"0000001300000000ffffffceffffffffffffffe0ffffffff0000001a00000000",
            INIT_5A => X"ffffffefffffffffffffffffffffffffffffff99ffffffff0000001c00000000",
            INIT_5B => X"ffffffc1ffffffffffffff92ffffffffffffffffffffffffffffffdbffffffff",
            INIT_5C => X"0000004b000000000000004500000000ffffffe8ffffffffffffffc0ffffffff",
            INIT_5D => X"00000052000000000000001d0000000000000001000000000000002b00000000",
            INIT_5E => X"fffffffcffffffffffffff54ffffffffffffffdeffffffffffffffa4ffffffff",
            INIT_5F => X"ffffffe1fffffffffffffffbffffffff0000002d00000000ffffffbcffffffff",
            INIT_60 => X"ffffffdffffffffffffffff8ffffffffffffffafffffffffffffffe8ffffffff",
            INIT_61 => X"00000004000000000000006500000000ffffff9effffffff0000005800000000",
            INIT_62 => X"0000003300000000ffffffecffffffff0000004900000000fffffffaffffffff",
            INIT_63 => X"0000004500000000fffffeb1ffffffffffffff9effffffffffffff9effffffff",
            INIT_64 => X"ffffffd3ffffffffffffffb8ffffffffffffff9effffffff0000000300000000",
            INIT_65 => X"ffffffe3ffffffff00000023000000000000003400000000ffffffc8ffffffff",
            INIT_66 => X"ffffffe2fffffffffffffff7ffffffff0000000300000000fffffffbffffffff",
            INIT_67 => X"fffffffaffffffff00000015000000000000002700000000ffffff8fffffffff",
            INIT_68 => X"0000000e00000000ffffff94ffffffffffffffb4fffffffffffffffaffffffff",
            INIT_69 => X"fffffff0fffffffffffffffcffffffff0000000d000000000000003d00000000",
            INIT_6A => X"ffffff90ffffffff0000002100000000ffffffb9ffffffffffffffa0ffffffff",
            INIT_6B => X"ffffff9effffffff0000001800000000fffffff8ffffffffffffffa9ffffffff",
            INIT_6C => X"0000001a00000000ffffff9bffffffffffffffe1ffffffffffffff4dffffffff",
            INIT_6D => X"000000710000000000000064000000000000005f000000000000003a00000000",
            INIT_6E => X"ffffffc1ffffffffffffffc0ffffffff0000002f00000000ffffffdfffffffff",
            INIT_6F => X"0000001f0000000000000014000000000000000900000000ffffff9fffffffff",
            INIT_70 => X"ffffffdcffffffff0000002a000000000000000400000000ffffffe4ffffffff",
            INIT_71 => X"ffffffc8fffffffffffffff3ffffffffffffffb0ffffffffffffffe0ffffffff",
            INIT_72 => X"ffffff93ffffffffffffffe9ffffffffffffffe8ffffffff0000002100000000",
            INIT_73 => X"0000001c00000000ffffff16ffffffffffffffbcffffffffffffff54ffffffff",
            INIT_74 => X"fffffff4ffffffffffffffcdfffffffffffffffeffffffffffffffeeffffffff",
            INIT_75 => X"ffffffc1ffffffffffffff87ffffffffffffffd8ffffffff0000004700000000",
            INIT_76 => X"0000001b00000000ffffff7dfffffffffffffffaffffffff0000000200000000",
            INIT_77 => X"fffffff6ffffffff0000004200000000fffffff2ffffffffffffffdaffffffff",
            INIT_78 => X"0000002d00000000000000100000000000000023000000000000001d00000000",
            INIT_79 => X"ffffffc9fffffffffffffff8fffffffffffffff2ffffffffffffffeaffffffff",
            INIT_7A => X"ffffffa0ffffffffffffffc3ffffffff00000005000000000000003500000000",
            INIT_7B => X"ffffffa1ffffffff0000002e00000000ffffffeeffffffffffffffc3ffffffff",
            INIT_7C => X"0000005000000000fffffff3ffffffffffffffc2ffffffffffffff89ffffffff",
            INIT_7D => X"0000003500000000fffffffbffffffff00000043000000000000002100000000",
            INIT_7E => X"ffffffe3ffffffffffffff9effffffff0000002e000000000000001500000000",
            INIT_7F => X"00000049000000000000000d00000000ffffffddffffffffffffff8cffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE5;


    MEM_IWGHT_LAYER3_INSTANCE6 : if BRAM_NAME = "iwght_layer3_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001200000000ffffff9bffffffffffffffffffffffff0000000500000000",
            INIT_01 => X"0000000b00000000fffffff8ffffffff000000ba00000000ffffffe1ffffffff",
            INIT_02 => X"ffffffffffffffff000000100000000000000037000000000000002700000000",
            INIT_03 => X"00000040000000000000001e00000000ffffffd3ffffffffffffff79ffffffff",
            INIT_04 => X"ffffff9bffffffffffffffe2ffffffffffffff7affffffff0000001200000000",
            INIT_05 => X"ffffff8effffffff0000002d0000000000000018000000000000000700000000",
            INIT_06 => X"ffffffffffffffffffffff77ffffffff0000001d00000000fffffff3ffffffff",
            INIT_07 => X"fffffffcffffffff0000002b00000000ffffffebffffffff0000001800000000",
            INIT_08 => X"ffffffddffffffffffffffb4ffffffffffffffe5ffffffff0000004100000000",
            INIT_09 => X"00000072000000000000002300000000ffffffc7ffffffff0000003500000000",
            INIT_0A => X"ffffffbeffffffff0000002d00000000fffffff1ffffffff0000002f00000000",
            INIT_0B => X"ffffffa9ffffffffffffffc9ffffffff00000000000000000000000000000000",
            INIT_0C => X"ffffffd9ffffffffffffffc7ffffffff0000000600000000ffffff58ffffffff",
            INIT_0D => X"fffffffbffffffff0000003500000000ffffffcbffffffff0000001300000000",
            INIT_0E => X"ffffffc6ffffffffffffffb8ffffffff0000006800000000fffffff3ffffffff",
            INIT_0F => X"fffffff1ffffffffffffffb4ffffffff0000001700000000ffffffc5ffffffff",
            INIT_10 => X"ffffff62ffffffffffffff75ffffffffffffffa9ffffffffffffffdaffffffff",
            INIT_11 => X"0000004a00000000ffffff9effffffff0000005800000000ffffff84ffffffff",
            INIT_12 => X"0000006100000000fffffff2ffffffff0000001900000000ffffffccffffffff",
            INIT_13 => X"0000006700000000ffffff77ffffffffffffff80ffffffffffffff58ffffffff",
            INIT_14 => X"ffffffaffffffffffffffff9ffffffffffffff90fffffffffffffff7ffffffff",
            INIT_15 => X"ffffffccffffffff0000001a000000000000007c00000000ffffffb4ffffffff",
            INIT_16 => X"ffffffcfffffffff0000000800000000fffffff6ffffffff0000001200000000",
            INIT_17 => X"00000005000000000000003e00000000ffffffe4ffffffffffffffbeffffffff",
            INIT_18 => X"ffffffc1ffffffffffffffc4ffffffffffffffeaffffffff0000004000000000",
            INIT_19 => X"00000004000000000000000100000000ffffffb8ffffffff0000005b00000000",
            INIT_1A => X"ffffff7bfffffffffffffff3fffffffffffffff1ffffffffffffffd3ffffffff",
            INIT_1B => X"ffffff8bffffffff0000001d000000000000000300000000ffffffc1ffffffff",
            INIT_1C => X"ffffffdbffffffffffffff45fffffffffffffffdffffffff0000008d00000000",
            INIT_1D => X"ffffffe2ffffffff0000003800000000ffffffc4ffffffff0000003000000000",
            INIT_1E => X"0000000800000000ffffff8cffffffff0000003600000000ffffffe4ffffffff",
            INIT_1F => X"fffffff9ffffffffffffffafffffffff0000000000000000ffffffffffffffff",
            INIT_20 => X"ffffffbfffffffffffffffc9ffffffff00000028000000000000000300000000",
            INIT_21 => X"0000002800000000ffffffcbfffffffffffffdebffffffffffffff82ffffffff",
            INIT_22 => X"0000003b00000000ffffffefffffffff00000039000000000000002100000000",
            INIT_23 => X"0000001200000000ffffff93ffffffffffffff9dffffffffffffffc7ffffffff",
            INIT_24 => X"ffffff90ffffffff0000002300000000ffffffd7ffffffff0000000500000000",
            INIT_25 => X"ffffffe4fffffffffffffffafffffffffffffff4ffffffff0000006f00000000",
            INIT_26 => X"ffffffebffffffffffffff94ffffffffffffffd7fffffffffffffffbffffffff",
            INIT_27 => X"00000009000000000000002b000000000000000200000000ffffffbcffffffff",
            INIT_28 => X"0000001300000000ffffffbcffffffffffffffe3ffffffffffffffc2ffffffff",
            INIT_29 => X"ffffff9dffffffff0000003c00000000fffffff1ffffffff0000005100000000",
            INIT_2A => X"ffffff8ffffffffffffffff6ffffffffffffffeafffffffffffffff3ffffffff",
            INIT_2B => X"ffffffceffffffff0000000800000000ffffffe6ffffffffffffffe4ffffffff",
            INIT_2C => X"0000002500000000ffffffb8ffffffff0000000400000000ffffff6effffffff",
            INIT_2D => X"fffffffcffffffffffffffd1fffffffffffffff6ffffffff0000001d00000000",
            INIT_2E => X"00000005000000000000002500000000ffffffe5ffffffff0000000000000000",
            INIT_2F => X"0000000200000000ffffffe0ffffffffffffff87ffffffffffffff57ffffffff",
            INIT_30 => X"fffffffdffffffffffffffbdffffffff0000006300000000ffffffd5ffffffff",
            INIT_31 => X"0000000e00000000ffffffa8ffffffffffffff9effffffffffffffa2ffffffff",
            INIT_32 => X"000000380000000000000017000000000000003e000000000000001800000000",
            INIT_33 => X"0000003300000000ffffffb6ffffffffffffffe1ffffffffffffffdaffffffff",
            INIT_34 => X"ffffffabffffffff0000003a00000000ffffffe0ffffffff0000000600000000",
            INIT_35 => X"00000022000000000000003700000000fffffffcffffffffffffffc7ffffffff",
            INIT_36 => X"0000000700000000ffffffb1ffffffff0000000d000000000000000800000000",
            INIT_37 => X"0000001900000000ffffffb6ffffffff0000003500000000ffffffe5ffffffff",
            INIT_38 => X"0000002c00000000ffffffd4ffffffffffffffe4ffffffff0000003400000000",
            INIT_39 => X"0000003700000000fffffff5ffffffffffffff7dffffffff0000000000000000",
            INIT_3A => X"fffffff9ffffffffffffffcfffffffff0000005700000000ffffffcfffffffff",
            INIT_3B => X"ffffffdaffffffff0000000700000000ffffffe8ffffffff0000000600000000",
            INIT_3C => X"ffffff7dffffffffffffffd3fffffffffffffff1ffffffff0000005c00000000",
            INIT_3D => X"00000011000000000000001100000000ffffffecffffffff0000005d00000000",
            INIT_3E => X"00000030000000000000001a00000000ffffffd1ffffffffffffffb7ffffffff",
            INIT_3F => X"0000001a00000000ffffffd8ffffffffffffffe0ffffffffffffffb0ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffafffffffffffffff76ffffffffffffffc5fffffffffffffff8ffffffff",
            INIT_41 => X"0000006500000000ffffff82ffffffff00000021000000000000006000000000",
            INIT_42 => X"ffffffc6fffffffffffffff2ffffffffffffffccffffffffffffffabffffffff",
            INIT_43 => X"0000005b00000000ffffffd4ffffffffffffffa1ffffffffffffff60ffffffff",
            INIT_44 => X"ffffff91ffffffffffffffe2ffffffffffffffc1ffffffff0000000800000000",
            INIT_45 => X"ffffffeeffffffff0000000000000000ffffffeefffffffffffffee7ffffffff",
            INIT_46 => X"ffffffe1fffffffffffffff2ffffffffffffffd3fffffffffffffff7ffffffff",
            INIT_47 => X"0000001300000000000000050000000000000013000000000000002f00000000",
            INIT_48 => X"ffffffe3ffffffff0000003e0000000000000000000000000000002600000000",
            INIT_49 => X"0000000800000000ffffffa6ffffffffffffff73ffffffff0000000400000000",
            INIT_4A => X"ffffff8cffffffffffffff94ffffffff0000002900000000fffffff2ffffffff",
            INIT_4B => X"fffffff2ffffffffffffffc7ffffffff00000001000000000000000300000000",
            INIT_4C => X"0000000600000000ffffff4fffffffffffffffefffffffff000000d500000000",
            INIT_4D => X"0000001b00000000ffffffecffffffffffffffabffffffff0000001100000000",
            INIT_4E => X"0000000b0000000000000025000000000000002d00000000ffffffcfffffffff",
            INIT_4F => X"ffffffe1ffffffffffffffeffffffffffffffff6ffffffffffffffc9ffffffff",
            INIT_50 => X"00000043000000000000003e00000000ffffffe9ffffffffffffffecffffffff",
            INIT_51 => X"fffffff1ffffffff0000003200000000ffffffa9ffffffffffffffb2ffffffff",
            INIT_52 => X"0000007600000000ffffffefffffffff0000000000000000ffffffe6ffffffff",
            INIT_53 => X"ffffffd0fffffffffffffed0ffffffff0000000000000000ffffff51ffffffff",
            INIT_54 => X"ffffffaaffffffffffffff9fffffffffffffffe8fffffffffffffff6ffffffff",
            INIT_55 => X"ffffff9affffffff0000000500000000fffffff5ffffffffffffff76ffffffff",
            INIT_56 => X"0000001200000000ffffffa9ffffffff0000000c00000000fffffff1ffffffff",
            INIT_57 => X"fffffff6ffffffffffffffb7ffffffff0000004100000000ffffff75ffffffff",
            INIT_58 => X"0000000900000000ffffffecffffffff0000001900000000fffffff5ffffffff",
            INIT_59 => X"ffffffc1ffffffff0000002d00000000ffffffb2ffffffff0000003f00000000",
            INIT_5A => X"0000000800000000fffffff2ffffffff0000005e000000000000000c00000000",
            INIT_5B => X"ffffffb0ffffffff0000000a00000000ffffffe7ffffffffffffffcfffffffff",
            INIT_5C => X"0000003a00000000ffffffeaffffffff0000000e00000000ffffffbdffffffff",
            INIT_5D => X"0000004600000000fffffffdffffffffffffffd2ffffffff0000003600000000",
            INIT_5E => X"0000001e000000000000000600000000fffffffbfffffffffffffff6ffffffff",
            INIT_5F => X"ffffff5effffffffffffffe9ffffffffffffff6fffffffffffffffbdffffffff",
            INIT_60 => X"0000004c00000000ffffffbcffffffff00000027000000000000000000000000",
            INIT_61 => X"ffffff7bffffffff0000002d00000000fffffff5ffffffffffffffcaffffffff",
            INIT_62 => X"ffffffbbffffffff00000011000000000000000900000000ffffffd1ffffffff",
            INIT_63 => X"0000000000000000ffffff57ffffffff00000054000000000000000000000000",
            INIT_64 => X"ffffff92ffffffff0000001300000000fffffeccffffffff0000000900000000",
            INIT_65 => X"ffffff6bffffffff0000002e000000000000001d000000000000004100000000",
            INIT_66 => X"ffffffdaffffffffffffff39ffffffffffffffb5ffffffff0000000700000000",
            INIT_67 => X"fffffffeffffffffffffff9effffffff00000035000000000000001d00000000",
            INIT_68 => X"fffffff6ffffffff0000005600000000ffffff5affffffffffffffb1ffffffff",
            INIT_69 => X"ffffffd1ffffffffffffffdbffffffffffffffe5ffffffff000000b000000000",
            INIT_6A => X"0000005400000000ffffff94ffffffff0000002a00000000000000a100000000",
            INIT_6B => X"0000000d000000000000000d000000000000000100000000ffffff0dffffffff",
            INIT_6C => X"0000000e00000000ffffffefffffffffffffff0fffffffffffffff86ffffffff",
            INIT_6D => X"0000000a000000000000002e00000000ffffffccffffffffffffffc9ffffffff",
            INIT_6E => X"ffffff68ffffffffffffffccffffffffffffff7affffffffffffffbeffffffff",
            INIT_6F => X"ffffffd2ffffffffffffffe1ffffffffffffff9fffffffff0000004600000000",
            INIT_70 => X"ffffff9effffffff0000001600000000ffffff3fffffffff0000000f00000000",
            INIT_71 => X"ffffff18fffffffffffffef0ffffffffffffffefffffffff000000c300000000",
            INIT_72 => X"ffffffdeffffffff0000000e00000000ffffff82ffffffff0000006100000000",
            INIT_73 => X"ffffff72ffffffff0000008900000000000000f9000000000000007600000000",
            INIT_74 => X"ffffffc7ffffffffffffffeaffffffffffffff79ffffffffffffffedffffffff",
            INIT_75 => X"ffffffbffffffffffffffff5fffffffffffffff1ffffffffffffffabffffffff",
            INIT_76 => X"ffffffa0ffffffffffffffaaffffffffffffffe7fffffffffffffff0ffffffff",
            INIT_77 => X"0000000000000000ffffff8bffffffff0000001d000000000000007000000000",
            INIT_78 => X"0000003900000000000000f000000000ffffff64ffffffffffffff9effffffff",
            INIT_79 => X"ffffff84ffffffff00000013000000000000000400000000ffffff58ffffffff",
            INIT_7A => X"0000001b00000000ffffff87ffffffff0000002f000000000000000300000000",
            INIT_7B => X"0000005500000000ffffffe9fffffffffffffff8ffffffffffffffbeffffffff",
            INIT_7C => X"ffffff97ffffffff0000008f000000000000006800000000000000a800000000",
            INIT_7D => X"ffffff91ffffffffffffff10ffffffff0000003400000000fffffff3ffffffff",
            INIT_7E => X"0000000100000000ffffff44fffffffffffffec0fffffffffffffff7ffffffff",
            INIT_7F => X"fffffff9ffffffff0000008100000000ffffff8fffffffff0000002c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE6;


    MEM_IWGHT_LAYER3_INSTANCE7 : if BRAM_NAME = "iwght_layer3_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffff02ffffffffffffff89ffffffffffffffacffffffff0000001b00000000",
            INIT_01 => X"ffffffc1ffffffff0000002600000000ffffffc8ffffffffffffffffffffffff",
            INIT_02 => X"ffffffefffffffff0000001400000000ffffffd2ffffffffffffffd3ffffffff",
            INIT_03 => X"0000001800000000fffffffbffffffff0000003100000000ffffff16ffffffff",
            INIT_04 => X"fffffffbffffffffffffffd9fffffffffffffff4ffffffff0000000e00000000",
            INIT_05 => X"0000006900000000fffffff8ffffffff0000003b00000000fffffff6ffffffff",
            INIT_06 => X"00000002000000000000001d00000000fffffff3ffffffffffffffeaffffffff",
            INIT_07 => X"ffffffecffffffffffffff8affffffffffffffa0ffffffffffffff3affffffff",
            INIT_08 => X"0000004c000000000000002c000000000000007400000000ffffffafffffffff",
            INIT_09 => X"fffffffaffffffff0000004e00000000fffffff2ffffffff0000001400000000",
            INIT_0A => X"00000035000000000000000f00000000ffffff1dffffffffffffffaaffffffff",
            INIT_0B => X"00000039000000000000005900000000fffffff5ffffffffffffff84ffffffff",
            INIT_0C => X"00000096000000000000000e00000000ffffffecffffffff0000007200000000",
            INIT_0D => X"0000001100000000ffffff86ffffffffffffffd3ffffffff0000004b00000000",
            INIT_0E => X"0000003f00000000ffffffa2fffffffffffffeeeffffffff0000001400000000",
            INIT_0F => X"ffffffa9ffffffff00000064000000000000002500000000ffffffc6ffffffff",
            INIT_10 => X"ffffffe9ffffffffffffffe4ffffffffffffffb5ffffffff0000000900000000",
            INIT_11 => X"0000001100000000fffffef5ffffffffffffff63ffffffffffffff5effffffff",
            INIT_12 => X"ffffffd2ffffffff0000001400000000ffffff62ffffffff0000004000000000",
            INIT_13 => X"0000001100000000ffffff4dffffffff0000001f00000000ffffff76ffffffff",
            INIT_14 => X"0000004200000000ffffffdfffffffff00000068000000000000000300000000",
            INIT_15 => X"ffffffbbffffffffffffffd3ffffffff00000020000000000000005600000000",
            INIT_16 => X"fffffff9ffffffffffffff6fffffffffffffffb6ffffffff0000001200000000",
            INIT_17 => X"0000001800000000ffffffeaffffffff0000004c000000000000005700000000",
            INIT_18 => X"ffffffb2fffffffffffffff7ffffffffffffffe6ffffffffffffff7dffffffff",
            INIT_19 => X"fffffffcffffffff0000000b00000000fffffff0ffffffff0000007300000000",
            INIT_1A => X"fffffffdffffffffffffff21ffffffffffffffcbffffffff0000001300000000",
            INIT_1B => X"ffffff93ffffffff00000051000000000000000300000000ffffff94ffffffff",
            INIT_1C => X"000000a200000000ffffffd4ffffffffffffff65ffffffff0000003700000000",
            INIT_1D => X"0000006800000000fffffffaffffffffffffff93ffffffffffffffcbffffffff",
            INIT_1E => X"fffffff6ffffffff0000005200000000ffffff51ffffffff0000001f00000000",
            INIT_1F => X"fffffff4ffffffff0000001600000000ffffffa7ffffffffffffffbaffffffff",
            INIT_20 => X"0000002900000000ffffffedffffffffffffff7cffffffff0000000600000000",
            INIT_21 => X"0000003100000000ffffff72ffffffffffffff83ffffffffffffffeeffffffff",
            INIT_22 => X"00000001000000000000000200000000ffffff9affffffff0000003300000000",
            INIT_23 => X"fffffff7ffffffff000000b6000000000000008300000000fffffeffffffffff",
            INIT_24 => X"0000002f00000000ffffff7affffffffffffff83fffffffffffffff2ffffffff",
            INIT_25 => X"0000006300000000ffffff96ffffffffffffffc9ffffffffffffffdcffffffff",
            INIT_26 => X"000000a100000000fffffef6ffffffff00000000000000000000000000000000",
            INIT_27 => X"0000001a00000000ffffffa7ffffffff0000004b00000000ffffffdfffffffff",
            INIT_28 => X"0000007500000000ffffff80ffffffffffffffdaffffffffffffff30ffffffff",
            INIT_29 => X"0000003600000000000000c000000000ffffffd2ffffffffffffff9dffffffff",
            INIT_2A => X"0000006800000000ffffff5effffffff000000d4000000000000004500000000",
            INIT_2B => X"ffffffc2ffffffffffffffc9ffffffff0000001600000000ffffff37ffffffff",
            INIT_2C => X"0000009000000000000000ae00000000ffffff49ffffffff0000002f00000000",
            INIT_2D => X"0000000a00000000ffffff67ffffffffffffffb1ffffffff0000007200000000",
            INIT_2E => X"0000001600000000ffffff30fffffffffffffdebfffffffffffffff0ffffffff",
            INIT_2F => X"fffffefaffffffff00000017000000000000001400000000ffffffd7ffffffff",
            INIT_30 => X"ffffffd9ffffffffffffffb9ffffffffffffffd8ffffffff0000000200000000",
            INIT_31 => X"ffffffd6ffffffffffffff43ffffffffffffffd5ffffffffffffffffffffffff",
            INIT_32 => X"ffffff9bfffffffffffffff6ffffffffffffff7fffffffff0000002f00000000",
            INIT_33 => X"ffffffedffffffffffffff77ffffffff0000003700000000ffffff98ffffffff",
            INIT_34 => X"ffffffbfffffffffffffffd6ffffffffffffffd2ffffffffffffffe9ffffffff",
            INIT_35 => X"ffffff65fffffffffffffff5ffffffff0000003e00000000fffffe14ffffffff",
            INIT_36 => X"fffffff7ffffffff00000030000000000000001d000000000000001300000000",
            INIT_37 => X"0000000600000000ffffffadffffffff00000002000000000000000900000000",
            INIT_38 => X"0000002d000000000000006000000000ffffff95ffffffffffffff12ffffffff",
            INIT_39 => X"00000039000000000000005b00000000fffffffbffffffff0000001e00000000",
            INIT_3A => X"0000001b00000000ffffffa9ffffffffffffffcbffffffffffffff34ffffffff",
            INIT_3B => X"ffffff26ffffffff00000043000000000000001700000000ffffff8bffffffff",
            INIT_3C => X"0000005b00000000ffffffb2ffffffffffffff50ffffffff0000006600000000",
            INIT_3D => X"00000010000000000000004f00000000ffffffbfffffffff0000007500000000",
            INIT_3E => X"0000002a00000000ffffff87ffffffffffffffd9fffffffffffffff2ffffffff",
            INIT_3F => X"ffffffc0ffffffff00000077000000000000003f000000000000000b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003700000000ffffffa6ffffffffffffff83fffffffffffffffbffffffff",
            INIT_41 => X"0000000f00000000ffffffabffffffff00000036000000000000006800000000",
            INIT_42 => X"0000005b00000000ffffffedffffffffffffff9cffffffff0000004500000000",
            INIT_43 => X"0000002e0000000000000033000000000000004d00000000ffffffdcffffffff",
            INIT_44 => X"ffffffb8ffffffffffffff8effffffffffffff90ffffffffffffffe6ffffffff",
            INIT_45 => X"ffffffd6ffffffff0000002300000000ffffffeaffffffffffffffb4ffffffff",
            INIT_46 => X"ffffffe5ffffffffffffffe9ffffffffffffff7bffffffff0000001300000000",
            INIT_47 => X"ffffffefffffffffffffffe9ffffffff0000002900000000ffffff3dffffffff",
            INIT_48 => X"ffffff70fffffffffffffff6fffffffffffffff5ffffffffffffff19ffffffff",
            INIT_49 => X"00000030000000000000004500000000ffffffc2ffffffffffffffe7ffffffff",
            INIT_4A => X"ffffffe9ffffffffffffffbdffffffff00000020000000000000007600000000",
            INIT_4B => X"ffffff48ffffffff00000016000000000000000a00000000ffffff55ffffffff",
            INIT_4C => X"0000000f00000000ffffffb1ffffffff0000000e00000000ffffffb3ffffffff",
            INIT_4D => X"00000033000000000000000200000000fffffec7ffffffffffffffe9ffffffff",
            INIT_4E => X"0000001c000000000000000000000000ffffffbaffffffffffffff4effffffff",
            INIT_4F => X"ffffffa1ffffffffffffffbdffffffff00000013000000000000002500000000",
            INIT_50 => X"0000002c0000000000000064000000000000003000000000ffffffebffffffff",
            INIT_51 => X"ffffffe2ffffffffffffffd7ffffffff00000041000000000000003900000000",
            INIT_52 => X"ffffffe3ffffffff0000000b0000000000000013000000000000002700000000",
            INIT_53 => X"fffffff2ffffffff0000004800000000ffffffb2ffffffffffffff91ffffffff",
            INIT_54 => X"ffffffdcfffffffffffffffcffffffffffffff8effffffff0000000900000000",
            INIT_55 => X"ffffff8affffffff0000004f000000000000002800000000ffffffd3ffffffff",
            INIT_56 => X"fffffff1ffffffffffffff80ffffffff0000000a000000000000000000000000",
            INIT_57 => X"0000000f00000000ffffffddfffffffffffffffcffffffffffffffe7ffffffff",
            INIT_58 => X"ffffff6cfffffffffffffff3ffffffff0000001000000000ffffffb1ffffffff",
            INIT_59 => X"00000011000000000000002e00000000ffffff8effffffff0000000400000000",
            INIT_5A => X"ffffffa7ffffffff0000005c000000000000004a00000000ffffffbaffffffff",
            INIT_5B => X"ffffffd1ffffffff0000002500000000ffffffeaffffffffffffffb6ffffffff",
            INIT_5C => X"0000000700000000ffffffb4ffffffffffffffa5ffffffffffffff5bffffffff",
            INIT_5D => X"00000024000000000000003100000000ffffffd3ffffffff0000001d00000000",
            INIT_5E => X"0000003e00000000ffffffd2ffffffff0000008e00000000fffffedcffffffff",
            INIT_5F => X"fffffec6ffffffff0000001b000000000000006800000000fffffff3ffffffff",
            INIT_60 => X"00000017000000000000001e000000000000003b00000000fffffff7ffffffff",
            INIT_61 => X"0000003200000000fffffff2ffffffffffffffb4ffffffff0000007b00000000",
            INIT_62 => X"fffffffafffffffffffffffeffffffffffffffe0ffffffff0000002e00000000",
            INIT_63 => X"0000004d00000000ffffff8effffffff0000003700000000fffffeb1ffffffff",
            INIT_64 => X"ffffff30ffffffffffffffebffffffffffffff3bffffffff0000001300000000",
            INIT_65 => X"ffffff3ffffffffffffffff0ffffffff0000000f00000000fffffffcffffffff",
            INIT_66 => X"ffffffebffffffffffffff9afffffffffffffff4ffffffffffffffebffffffff",
            INIT_67 => X"fffffff9ffffffff00000001000000000000003b00000000ffffffd0ffffffff",
            INIT_68 => X"fffffff9ffffffff0000001000000000fffffff4ffffffff0000000600000000",
            INIT_69 => X"ffffffb7ffffffff0000005700000000ffffffd8ffffffffffffffe7ffffffff",
            INIT_6A => X"ffffffeeffffffffffffff29ffffffffffffff6affffffffffffffc1ffffffff",
            INIT_6B => X"ffffffdfffffffff00000027000000000000000900000000ffffff4affffffff",
            INIT_6C => X"ffffffabffffffffffffffcaffffffffffffff9affffffff0000000e00000000",
            INIT_6D => X"ffffffb1ffffffff0000005f00000000ffffff95ffffffffffffffdcffffffff",
            INIT_6E => X"0000001a00000000ffffff83ffffffffffffffaaffffffffffffffb8ffffffff",
            INIT_6F => X"ffffffd6ffffffffffffffa4ffffffff00000065000000000000007400000000",
            INIT_70 => X"ffffffc3ffffffffffffffddffffffffffffff48ffffffff0000000200000000",
            INIT_71 => X"ffffffb1fffffffffffffffdffffffffffffff7fffffffff0000005d00000000",
            INIT_72 => X"0000000f00000000ffffffecfffffffffffffff8ffffffff0000008000000000",
            INIT_73 => X"00000009000000000000002700000000ffffff89ffffffff0000002300000000",
            INIT_74 => X"ffffffecffffffff00000029000000000000000a00000000fffffffeffffffff",
            INIT_75 => X"ffffffc3fffffffffffffff9fffffffffffffff6ffffffffffffff80ffffffff",
            INIT_76 => X"0000000300000000ffffffdfffffffffffffffb9fffffffffffffff8ffffffff",
            INIT_77 => X"0000000b00000000ffffffabffffffff0000000500000000ffffff9dffffffff",
            INIT_78 => X"ffffff7bffffffff0000003d0000000000000089000000000000000e00000000",
            INIT_79 => X"ffffffaeffffffffffffffefffffffff0000007e00000000ffffffc8ffffffff",
            INIT_7A => X"0000001c0000000000000050000000000000002600000000fffffde5ffffffff",
            INIT_7B => X"00000031000000000000001200000000fffffff1ffffffffffffffdaffffffff",
            INIT_7C => X"0000001c00000000000000180000000000000085000000000000000400000000",
            INIT_7D => X"ffffffc9ffffffffffffffd6ffffffff00000052000000000000003200000000",
            INIT_7E => X"000000760000000000000000000000000000007400000000ffffffa2ffffffff",
            INIT_7F => X"0000004d00000000ffffffabffffffffffffff42ffffffff0000003c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE7;


    MEM_IWGHT_LAYER3_INSTANCE8 : if BRAM_NAME = "iwght_layer3_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff3ffffffffffffffbaffffffff0000003f000000000000000200000000",
            INIT_01 => X"ffffffe6ffffffffffffffedffffffffffffff8effffffffffffffc7ffffffff",
            INIT_02 => X"ffffff6bffffffffffffffedffffffff0000003100000000ffffff6dffffffff",
            INIT_03 => X"0000002a00000000000000cb0000000000000006000000000000000100000000",
            INIT_04 => X"fffffff6ffffffff0000000800000000ffffffa5ffffffffffffffeaffffffff",
            INIT_05 => X"ffffff8effffffff0000003f00000000ffffff9fffffffff0000000800000000",
            INIT_06 => X"ffffffe1fffffffffffffff5ffffffffffffffedffffffff0000000400000000",
            INIT_07 => X"ffffffe5fffffffffffffff8ffffffff0000005000000000ffffffc8ffffffff",
            INIT_08 => X"ffffffa9ffffffffffffff44ffffffff0000006b000000000000004900000000",
            INIT_09 => X"ffffff5efffffffffffffff0ffffffff0000001400000000fffffffaffffffff",
            INIT_0A => X"ffffffc6ffffffff0000008100000000ffffffc6ffffffff0000000f00000000",
            INIT_0B => X"0000004f00000000ffffffddffffffff00000009000000000000002000000000",
            INIT_0C => X"ffffffe8ffffffffffffff99ffffffffffffffccffffffffffffff99ffffffff",
            INIT_0D => X"ffffff8affffffff0000004d00000000fffffee2fffffffffffffff3ffffffff",
            INIT_0E => X"000000480000000000000007000000000000007a00000000ffffff80ffffffff",
            INIT_0F => X"fffffffaffffffffffffff91ffffffff0000000900000000ffffff6dffffffff",
            INIT_10 => X"ffffffb5ffffffffffffff88fffffffffffffff2fffffffffffffff8ffffffff",
            INIT_11 => X"ffffff63ffffffffffffffc3ffffffff0000000c00000000ffffffa2ffffffff",
            INIT_12 => X"ffffff79ffffffff00000005000000000000008700000000ffffffe9ffffffff",
            INIT_13 => X"0000003d0000000000000044000000000000000f00000000ffffffb9ffffffff",
            INIT_14 => X"0000004d000000000000001200000000ffffffebfffffffffffffff5ffffffff",
            INIT_15 => X"ffffffe8ffffffff0000003d00000000ffffffd5ffffffff0000000d00000000",
            INIT_16 => X"ffffff5cffffffffffffffabffffffffffffff94ffffffffffffffeaffffffff",
            INIT_17 => X"0000000b00000000ffffffd6ffffffffffffffaaffffffff0000004200000000",
            INIT_18 => X"ffffff73ffffffff000000020000000000000043000000000000005500000000",
            INIT_19 => X"ffffffaaffffffffffffffffffffffffffffffe7ffffffff0000000f00000000",
            INIT_1A => X"ffffff73ffffffff0000001d00000000fffffff2ffffffffffffffb9ffffffff",
            INIT_1B => X"ffffffe5ffffffffffffff6cffffffff00000001000000000000001c00000000",
            INIT_1C => X"000000330000000000000017000000000000002900000000ffffffd6ffffffff",
            INIT_1D => X"fffffff2ffffffffffffffc1ffffffffffffffe2ffffffffffffffebffffffff",
            INIT_1E => X"000000500000000000000049000000000000009f00000000ffffffa9ffffffff",
            INIT_1F => X"0000004000000000ffffffadffffffff0000002600000000ffffff4bffffffff",
            INIT_20 => X"ffffff8bffffffff0000002e000000000000000600000000fffffffbffffffff",
            INIT_21 => X"ffffffd3ffffffffffffff74ffffffffffffff25ffffffffffffffb5ffffffff",
            INIT_22 => X"ffffffc9ffffffff0000000b000000000000003e00000000ffffffffffffffff",
            INIT_23 => X"ffffffe1ffffffffffffffb6ffffffffffffff31ffffffffffffffafffffffff",
            INIT_24 => X"00000022000000000000000700000000fffffeffffffffffffffffdeffffffff",
            INIT_25 => X"000000a700000000ffffffcdffffffff0000001c000000000000008c00000000",
            INIT_26 => X"0000001f000000000000000600000000ffffffa2fffffffffffffff8ffffffff",
            INIT_27 => X"fffffffcffffffffffffff90ffffffff0000003200000000ffffffb0ffffffff",
            INIT_28 => X"000000b5000000000000006a000000000000000d000000000000007300000000",
            INIT_29 => X"ffffffd1ffffffff0000005000000000ffffff86ffffffff0000001c00000000",
            INIT_2A => X"0000001200000000fffffe2efffffffffffffffdffffffffffffffa0ffffffff",
            INIT_2B => X"ffffffbeffffffff00000006000000000000000a000000000000001300000000",
            INIT_2C => X"ffffffeeffffffff0000000e0000000000000033000000000000003200000000",
            INIT_2D => X"ffffffb8ffffffff0000003d0000000000000000000000000000003a00000000",
            INIT_2E => X"000000570000000000000021000000000000006800000000ffffffa2ffffffff",
            INIT_2F => X"00000078000000000000003500000000ffffffb9ffffffff0000003a00000000",
            INIT_30 => X"ffffffc3ffffffffffffff20ffffffffffffff0ffffffffffffffff8ffffffff",
            INIT_31 => X"ffffff66ffffffff0000002b000000000000004900000000ffffffe3ffffffff",
            INIT_32 => X"000001120000000000000002000000000000001e000000000000002000000000",
            INIT_33 => X"ffffffd2ffffffffffffff66ffffffffffffffa2ffffffff0000009400000000",
            INIT_34 => X"0000003f00000000ffffff4bffffffffffffffc4ffffffffffffffebffffffff",
            INIT_35 => X"ffffff4fffffffff0000001000000000ffffff80ffffffffffffffdbffffffff",
            INIT_36 => X"0000003a00000000ffffff77fffffffffffffff0ffffffff0000001600000000",
            INIT_37 => X"00000012000000000000005500000000fffffff7ffffffffffffff88ffffffff",
            INIT_38 => X"ffffffffffffffff0000007200000000ffffff83ffffffff0000009100000000",
            INIT_39 => X"ffffffd8ffffffffffffff40ffffffffffffff81fffffffffffffff3ffffffff",
            INIT_3A => X"fffffff4ffffffff0000003300000000ffffff97ffffffffffffff27ffffffff",
            INIT_3B => X"ffffffb2ffffffffffffffa6ffffffffffffffebffffffff0000005b00000000",
            INIT_3C => X"ffffff65ffffffffffffff52ffffffff0000006100000000ffffffc6ffffffff",
            INIT_3D => X"0000000300000000ffffffabffffffffffffffd1ffffffffffffffa2ffffffff",
            INIT_3E => X"ffffffebffffffff0000003700000000ffffffffffffffff0000000000000000",
            INIT_3F => X"0000001d000000000000007c00000000ffffffbfffffffff0000000d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffff5fffffffffffffffd4ffffffff0000004100000000ffffffefffffffff",
            INIT_41 => X"ffffff4afffffffffffffff0fffffffffffffe7dffffffffffffff3dffffffff",
            INIT_42 => X"0000002800000000ffffffe6ffffffff00000050000000000000001100000000",
            INIT_43 => X"0000006600000000fffffefdffffffffffffffe5ffffffff0000002100000000",
            INIT_44 => X"0000001600000000ffffff73ffffffffffffff85ffffffff0000001600000000",
            INIT_45 => X"fffffff1fffffffffffffffcffffffff0000001c000000000000009200000000",
            INIT_46 => X"ffffffedffffffffffffff9effffffffffffff84ffffffff0000001800000000",
            INIT_47 => X"ffffffefffffffff0000000700000000ffffff95ffffffffffffff38ffffffff",
            INIT_48 => X"ffffffe2ffffffffffffffecffffffffffffffd1ffffffff0000004500000000",
            INIT_49 => X"0000002b00000000ffffff4dffffffffffffffd5ffffffff0000000600000000",
            INIT_4A => X"ffffff9effffffff0000007d00000000fffffff5ffffffff0000002300000000",
            INIT_4B => X"ffffffbcffffffff0000001a0000000000000004000000000000007100000000",
            INIT_4C => X"ffffff68ffffffff0000001c000000000000005900000000ffffff72ffffffff",
            INIT_4D => X"0000003c00000000ffffffefffffffff0000001500000000ffffffebffffffff",
            INIT_4E => X"fffffffeffffffff0000008d000000000000002300000000ffffffcbffffffff",
            INIT_4F => X"0000003c000000000000001d00000000ffffff87ffffffffffffffb9ffffffff",
            INIT_50 => X"ffffffdcffffffffffffffcfffffffff000000b600000000fffffff9ffffffff",
            INIT_51 => X"ffffffdfffffffff0000000300000000fffffef5ffffffffffffff9bffffffff",
            INIT_52 => X"0000007d00000000ffffffe9ffffffffffffffceffffffff0000004400000000",
            INIT_53 => X"ffffffd8ffffffffffffff46fffffffffffffea7ffffffffffffffbdffffffff",
            INIT_54 => X"0000001500000000ffffffa1ffffffff0000003100000000fffffff2ffffffff",
            INIT_55 => X"ffffff87ffffffff00000035000000000000006b00000000ffffff7effffffff",
            INIT_56 => X"0000000b000000000000005b00000000ffffffdaffffffff0000001100000000",
            INIT_57 => X"000000030000000000000015000000000000006300000000ffffffc7ffffffff",
            INIT_58 => X"0000009d000000000000008500000000ffffffb8ffffffff0000003800000000",
            INIT_59 => X"ffffff84ffffffffffffffc0ffffffffffffff84ffffffffffffffa9ffffffff",
            INIT_5A => X"0000001300000000ffffff6fffffffff0000000600000000ffffff69ffffffff",
            INIT_5B => X"ffffffddfffffffffffffff2ffffffff00000014000000000000004f00000000",
            INIT_5C => X"00000019000000000000003b00000000fffffff8fffffffffffffef9ffffffff",
            INIT_5D => X"ffffffc5ffffffff0000006f000000000000007f00000000ffffffbeffffffff",
            INIT_5E => X"ffffffb4ffffffff0000003f00000000000000d9000000000000007800000000",
            INIT_5F => X"00000041000000000000008400000000ffffffb9ffffffff0000001200000000",
            INIT_60 => X"ffffffdcffffffffffffff9bffffffffffffffd2fffffffffffffff4ffffffff",
            INIT_61 => X"ffffff69ffffffffffffffc0ffffffffffffffe2fffffffffffffff1ffffffff",
            INIT_62 => X"ffffff6cffffffff0000000d0000000000000005000000000000005e00000000",
            INIT_63 => X"ffffff8effffffff0000004900000000ffffff5dffffffff0000003000000000",
            INIT_64 => X"000000a000000000ffffff93ffffffff0000000f000000000000000000000000",
            INIT_65 => X"ffffff30ffffffffffffffbaffffffff0000000d00000000fffffff1ffffffff",
            INIT_66 => X"ffffffe9ffffffffffffff63ffffffffffffffe7ffffffffffffffedffffffff",
            INIT_67 => X"0000000300000000ffffff8bffffffffffffffcdffffffff0000002900000000",
            INIT_68 => X"0000002e000000000000000b000000000000000f00000000ffffffe2ffffffff",
            INIT_69 => X"00000034000000000000001d00000000ffffff7effffffffffffffbeffffffff",
            INIT_6A => X"ffffffe4ffffffffffffff3affffffff0000002900000000ffffffeaffffffff",
            INIT_6B => X"ffffff5cffffffff00000021000000000000001100000000ffffffffffffffff",
            INIT_6C => X"fffffff1ffffffff0000000b000000000000003c000000000000006900000000",
            INIT_6D => X"ffffffdbfffffffffffffff7ffffffffffffff5fffffffffffffffd4ffffffff",
            INIT_6E => X"0000001700000000fffffff2ffffffffffffffeaffffffff0000000c00000000",
            INIT_6F => X"fffffff2ffffffff0000009500000000ffffff22fffffffffffffef7ffffffff",
            INIT_70 => X"000000240000000000000038000000000000006000000000ffffffe3ffffffff",
            INIT_71 => X"ffffff74fffffffffffffff6ffffffff0000000f00000000ffffff47ffffffff",
            INIT_72 => X"ffffffaafffffffffffffffffffffffffffffffaffffffff0000008300000000",
            INIT_73 => X"0000005600000000ffffff4affffffffffffff82ffffffff0000001300000000",
            INIT_74 => X"ffffffddffffffffffffffc4ffffffff0000000f000000000000000a00000000",
            INIT_75 => X"0000004f00000000ffffffb0ffffffff0000001900000000ffffff9cffffffff",
            INIT_76 => X"0000006300000000ffffffc3ffffffffffffffa2ffffffffffffffedffffffff",
            INIT_77 => X"0000000600000000ffffffe5ffffffffffffff9dffffffffffffff99ffffffff",
            INIT_78 => X"000000450000000000000053000000000000000e00000000fffffff8ffffffff",
            INIT_79 => X"0000003700000000ffffffa7ffffffffffffff83ffffffffffffffffffffffff",
            INIT_7A => X"ffffff59ffffffff0000003f000000000000005100000000ffffff01ffffffff",
            INIT_7B => X"ffffffd2ffffffff0000005a000000000000000300000000ffffffe1ffffffff",
            INIT_7C => X"ffffffd5ffffffff000000970000000000000008000000000000002000000000",
            INIT_7D => X"0000004f000000000000000700000000ffffffa3ffffffff0000002a00000000",
            INIT_7E => X"ffffffa5ffffffff0000006900000000ffffffd7ffffffffffffffeeffffffff",
            INIT_7F => X"ffffffffffffffff0000005200000000ffffffc8ffffffffffffff71ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE8;


    MEM_IWGHT_LAYER3_INSTANCE9 : if BRAM_NAME = "iwght_layer3_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffa8ffffffffffffff39ffffffff0000006800000000ffffffe0ffffffff",
            INIT_01 => X"fffffff2ffffffffffffffe8ffffffffffffffd6ffffffffffffffb7ffffffff",
            INIT_02 => X"0000009700000000000000030000000000000025000000000000000a00000000",
            INIT_03 => X"fffffff7ffffffff0000012100000000ffffffe7ffffffff000000f500000000",
            INIT_04 => X"ffffffefffffffff00000061000000000000003f00000000ffffffdeffffffff",
            INIT_05 => X"ffffffc3ffffffffffffff8fffffffff0000008900000000ffffff97ffffffff",
            INIT_06 => X"ffffffc1ffffffff0000001500000000fffffed5fffffffffffffff9ffffffff",
            INIT_07 => X"fffffffaffffffffffffffcaffffffff0000002e000000000000000900000000",
            INIT_08 => X"fffffff5ffffffffffffff9bffffffffffffffe4ffffffff0000002000000000",
            INIT_09 => X"ffffffe4ffffffffffffff41ffffffffffffffacffffffff0000000400000000",
            INIT_0A => X"0000002800000000fffffff8ffffffff0000008000000000fffffff2ffffffff",
            INIT_0B => X"0000007900000000ffffffd7ffffffff00000003000000000000007b00000000",
            INIT_0C => X"ffffff36ffffffffffffffa0ffffffff0000002000000000ffffff3fffffffff",
            INIT_0D => X"ffffff6bffffffffffffff66ffffffff0000000900000000ffffffb5ffffffff",
            INIT_0E => X"ffffffbeffffffff0000002b00000000fffffeaaffffffff0000005700000000",
            INIT_0F => X"000000bb00000000000000dd00000000ffffffb5ffffffff0000000800000000",
            INIT_10 => X"0000003f00000000ffffffd8ffffffff00000000000000000000000300000000",
            INIT_11 => X"ffffff9effffffffffffffc8ffffffff000000c3000000000000003400000000",
            INIT_12 => X"fffffff6ffffffff0000000800000000ffffff63ffffffffffffff90ffffffff",
            INIT_13 => X"0000001c000000000000005f00000000ffffffa7fffffffffffffff1ffffffff",
            INIT_14 => X"ffffffd2ffffffff0000004900000000fffffff8ffffffff0000000900000000",
            INIT_15 => X"ffffffb4ffffffff0000002600000000ffffff54ffffffffffffffbfffffffff",
            INIT_16 => X"0000002900000000ffffff70ffffffff0000003200000000fffffff6ffffffff",
            INIT_17 => X"0000001300000000ffffffc8ffffffffffffffb8ffffffff0000001b00000000",
            INIT_18 => X"ffffffa4ffffffff00000019000000000000001800000000fffffff1ffffffff",
            INIT_19 => X"ffffffd6ffffffffffffff79fffffffffffffff2ffffffffffffff73ffffffff",
            INIT_1A => X"ffffffb3ffffffffffffffcdffffffff0000006d00000000fffffea5ffffffff",
            INIT_1B => X"000000090000000000000000000000000000000f00000000ffffffdaffffffff",
            INIT_1C => X"ffffff83ffffffff0000004100000000ffffffd8ffffffff0000003a00000000",
            INIT_1D => X"ffffffb3ffffffffffffffeeffffffff0000001900000000ffffff98ffffffff",
            INIT_1E => X"000000d4000000000000003900000000ffffff7bffffffff0000008f00000000",
            INIT_1F => X"ffffffa7ffffffffffffffa5ffffffffffffffecffffffff0000000b00000000",
            INIT_20 => X"ffffff9effffffffffffff22ffffffffffffffddffffffffffffffe6ffffffff",
            INIT_21 => X"ffffffd7ffffffffffffffadffffffffffffff7afffffffffffffffcffffffff",
            INIT_22 => X"0000006800000000fffffff1fffffffffffffff2ffffffff0000002200000000",
            INIT_23 => X"fffffff3ffffffffffffff40ffffffffffffffddffffffff0000003300000000",
            INIT_24 => X"ffffffccffffffffffffffafffffffffffffff55ffffffff0000000400000000",
            INIT_25 => X"ffffff36ffffffff0000007b00000000ffffffb4ffffffffffffffe3ffffffff",
            INIT_26 => X"ffffffb1ffffffff0000001d00000000ffffffebffffffff0000001200000000",
            INIT_27 => X"ffffffecffffffffffffffd8ffffffffffffffdcffffffff0000001100000000",
            INIT_28 => X"ffffff94ffffffff0000003700000000ffffff7fffffffffffffffe6ffffffff",
            INIT_29 => X"ffffffc8ffffffffffffff8affffffffffffff96ffffffffffffffdcffffffff",
            INIT_2A => X"ffffffb3ffffffffffffffc5ffffffffffffffffffffffffffffff69ffffffff",
            INIT_2B => X"0000001400000000fffffff6ffffffff0000000200000000ffffff73ffffffff",
            INIT_2C => X"fffffebbfffffffffffffff1ffffffff0000006d00000000ffffffb8ffffffff",
            INIT_2D => X"ffffffd0ffffffff00000075000000000000000b00000000ffffff8fffffffff",
            INIT_2E => X"ffffffbaffffffff00000050000000000000003d000000000000009b00000000",
            INIT_2F => X"0000005800000000ffffffc9ffffffff0000004200000000ffffffb3ffffffff",
            INIT_30 => X"fffffff5ffffffffffffffdfffffffffffffffc7fffffffffffffff4ffffffff",
            INIT_31 => X"ffffff43ffffffff0000004f00000000000000dc000000000000004f00000000",
            INIT_32 => X"00000019000000000000001700000000ffffffeaffffffffffffff9bffffffff",
            INIT_33 => X"ffffffa2fffffffffffffee4ffffffff0000004800000000ffffff88ffffffff",
            INIT_34 => X"ffffffc7ffffffff00000019000000000000000d00000000fffffffcffffffff",
            INIT_35 => X"ffffffa2ffffffffffffffbfffffffffffffff98ffffffffffffffecffffffff",
            INIT_36 => X"fffffffcffffffffffffffcaffffffffffffffadffffffff0000000100000000",
            INIT_37 => X"fffffffcffffffffffffffd2ffffffffffffff9cffffffffffffff3bffffffff",
            INIT_38 => X"ffffffaafffffffffffffff2ffffffff0000003f00000000ffffffe0ffffffff",
            INIT_39 => X"ffffffdbfffffffffffffee3fffffffffffffff4fffffffffffffeecffffffff",
            INIT_3A => X"00000060000000000000000400000000fffffff2ffffffff0000002b00000000",
            INIT_3B => X"0000001d0000000000000075000000000000001600000000000000af00000000",
            INIT_3C => X"ffffff78ffffffffffffff94ffffffffffffffbfffffffff0000000e00000000",
            INIT_3D => X"ffffffb6ffffffffffffff6cffffffff0000006f00000000ffffffd9ffffffff",
            INIT_3E => X"ffffff9cffffffff0000001200000000ffffff4affffffff0000002000000000",
            INIT_3F => X"fffffffeffffffffffffffc5ffffffff0000006d000000000000003e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff7ffffffffffffff67ffffffffffffff87ffffffff0000001100000000",
            INIT_41 => X"fffffffafffffffffffffff6ffffffff0000004f000000000000005e00000000",
            INIT_42 => X"ffffffa3ffffffff0000000600000000ffffffedffffffff0000004b00000000",
            INIT_43 => X"0000001a000000000000018c000000000000002700000000ffffff59ffffffff",
            INIT_44 => X"ffffffddffffffff00000007000000000000006c00000000fffffffcffffffff",
            INIT_45 => X"ffffffa7ffffffff0000005700000000ffffff60ffffffff0000001f00000000",
            INIT_46 => X"000000260000000000000050000000000000009000000000ffffffedffffffff",
            INIT_47 => X"fffffff9ffffffffffffffb4ffffffffffffffe1ffffffff0000001a00000000",
            INIT_48 => X"0000001400000000ffffffdcffffffff0000007e00000000ffffff6effffffff",
            INIT_49 => X"0000000500000000fffffef4ffffffff0000006200000000ffffffb1ffffffff",
            INIT_4A => X"fffffffdffffffffffffffb5ffffffffffffffd2ffffffffffffffdcffffffff",
            INIT_4B => X"000000e900000000ffffffb8ffffffffffffffe9ffffffff0000004000000000",
            INIT_4C => X"ffffffd8ffffffff0000005d00000000ffffff9dfffffffffffffff9ffffffff",
            INIT_4D => X"0000001200000000ffffffbfffffffffffffffd0ffffffffffffffd8ffffffff",
            INIT_4E => X"0000002300000000ffffffe3ffffffff0000000900000000000000dd00000000",
            INIT_4F => X"ffffff5effffffff0000000a0000000000000000000000000000000800000000",
            INIT_50 => X"0000003800000000ffffffe8ffffffffffffff60ffffffffffffffedffffffff",
            INIT_51 => X"000000c100000000fffffff8ffffffff0000009b00000000ffffffcfffffffff",
            INIT_52 => X"0000002b00000000fffffff9ffffffffffffffebffffffff0000005900000000",
            INIT_53 => X"ffffffc1ffffffff000000bd000000000000001f00000000fffffe73ffffffff",
            INIT_54 => X"ffffff96ffffffffffffff81ffffffffffffffdbffffffff0000000900000000",
            INIT_55 => X"ffffff8dffffffff0000004000000000ffffffd5ffffffff0000009300000000",
            INIT_56 => X"0000000a00000000ffffffe7ffffffff0000002f00000000fffffffdffffffff",
            INIT_57 => X"0000000f00000000ffffffcaffffffffffffffe7ffffffff0000004100000000",
            INIT_58 => X"ffffffd4ffffffffffffffefffffffff00000084000000000000001200000000",
            INIT_59 => X"ffffffa7ffffffffffffffb2fffffffffffffff6ffffffffffffffbeffffffff",
            INIT_5A => X"00000058000000000000000200000000ffffffd5ffffffffffffffdaffffffff",
            INIT_5B => X"0000004c000000000000002000000000ffffffebffffffffffffffb8ffffffff",
            INIT_5C => X"0000000500000000ffffff9effffffff00000055000000000000005e00000000",
            INIT_5D => X"ffffff57ffffffffffffff42ffffffff00000035000000000000001800000000",
            INIT_5E => X"00000055000000000000000b00000000fffffff5ffffffff000000da00000000",
            INIT_5F => X"fffffff0ffffffff00000000000000000000004000000000ffffffeaffffffff",
            INIT_60 => X"ffffffdfffffffff0000000c00000000ffffffe1ffffffff0000000c00000000",
            INIT_61 => X"000000410000000000000019000000000000005a00000000ffffff9fffffffff",
            INIT_62 => X"ffffffd3fffffffffffffff0ffffffff0000002b00000000fffffff2ffffffff",
            INIT_63 => X"ffffff68ffffffff0000010d0000000000000029000000000000001e00000000",
            INIT_64 => X"ffffff44ffffffff00000032000000000000004d000000000000000000000000",
            INIT_65 => X"ffffff5cfffffffffffffef0fffffffffffffec8ffffffff0000004900000000",
            INIT_66 => X"0000002200000000ffffff57ffffffffffffffe7fffffffffffffff7ffffffff",
            INIT_67 => X"0000001700000000ffffffd5ffffffffffffff89ffffffffffffffcdffffffff",
            INIT_68 => X"000000520000000000000021000000000000001200000000ffffffd8ffffffff",
            INIT_69 => X"ffffff57fffffffffffffed2ffffffffffffffa8ffffffffffffff93ffffffff",
            INIT_6A => X"ffffff4ffffffffffffffee2ffffffffffffffa1ffffffff0000002f00000000",
            INIT_6B => X"0000002800000000ffffff7dffffffff0000000200000000ffffffedffffffff",
            INIT_6C => X"0000001400000000ffffff78fffffffffffffee1ffffffff000000bb00000000",
            INIT_6D => X"0000007100000000ffffffa3ffffffffffffffe4ffffffff0000008b00000000",
            INIT_6E => X"ffffff9effffffffffffffa4fffffffffffffed5ffffffffffffffc3ffffffff",
            INIT_6F => X"ffffff63ffffffffffffff3cffffffff00000099000000000000002300000000",
            INIT_70 => X"000000260000000000000027000000000000002200000000ffffffe5ffffffff",
            INIT_71 => X"000000e1000000000000000400000000ffffffe6ffffffff0000001f00000000",
            INIT_72 => X"ffffffbbfffffffffffffff2ffffffff0000000500000000ffffff5cffffffff",
            INIT_73 => X"ffffffbeffffffffffffff0dffffffff0000010500000000ffffff3fffffffff",
            INIT_74 => X"ffffffaeffffffff00000015000000000000003f000000000000000600000000",
            INIT_75 => X"0000000e00000000ffffffd1ffffffffffffffd6fffffffffffffff6ffffffff",
            INIT_76 => X"ffffff3dffffffff00000051000000000000003c00000000fffffff3ffffffff",
            INIT_77 => X"0000000e00000000ffffff1fffffffffffffff7affffffff0000000e00000000",
            INIT_78 => X"ffffff57ffffffff0000000400000000ffffffefffffffff0000001000000000",
            INIT_79 => X"ffffff65ffffffffffffff96fffffffffffffffeffffffffffffffb9ffffffff",
            INIT_7A => X"0000008c000000000000000600000000ffffff71ffffffff0000008f00000000",
            INIT_7B => X"000000aa000000000000006b000000000000000300000000ffffffd6ffffffff",
            INIT_7C => X"0000007300000000000000c700000000ffffff90ffffffffffffff2cffffffff",
            INIT_7D => X"ffffff8dffffffffffffff66ffffffff00000045000000000000002500000000",
            INIT_7E => X"0000002600000000ffffff5bfffffffffffffd8effffffff0000009800000000",
            INIT_7F => X"ffffff55ffffffff000000110000000000000074000000000000009f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE9;


    MEM_IWGHT_LAYER3_INSTANCE10 : if BRAM_NAME = "iwght_layer3_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffffffffffff0000007a0000000000000046000000000000000d00000000",
            INIT_01 => X"0000015d00000000ffffffafffffffff000000ed00000000ffffffe2ffffffff",
            INIT_02 => X"ffffffa5ffffffff0000001400000000ffffff9affffffffffffff55ffffffff",
            INIT_03 => X"ffffff3bffffffff0000007800000000ffffff45ffffffffffffffbbffffffff",
            INIT_04 => X"ffffff12ffffffffffffffb3ffffffff0000001900000000ffffffe7ffffffff",
            INIT_05 => X"ffffff85ffffffffffffff89ffffffffffffffd1ffffffff0000003100000000",
            INIT_06 => X"ffffff62ffffffff00000013000000000000007100000000fffffff8ffffffff",
            INIT_07 => X"0000000500000000ffffff1fffffffffffffffe8ffffffff0000000b00000000",
            INIT_08 => X"ffffffdeffffffffffffffbdffffffffffffffe6ffffffffffffff46ffffffff",
            INIT_09 => X"0000002100000000ffffffc2ffffffffffffffc1ffffffff0000002800000000",
            INIT_0A => X"0000005d00000000fffffefcffffffffffffff92ffffffff000000c000000000",
            INIT_0B => X"ffffffe2ffffffffffffff94ffffffff00000006000000000000009400000000",
            INIT_0C => X"0000008900000000ffffff6affffffff0000004d00000000000000aa00000000",
            INIT_0D => X"ffffffbcffffffffffffffacffffffff0000005100000000fffffff8ffffffff",
            INIT_0E => X"00000072000000000000000500000000ffffff09ffffffffffffff88ffffffff",
            INIT_0F => X"0000008300000000ffffffc8ffffffff00000097000000000000002d00000000",
            INIT_10 => X"00000014000000000000009d00000000ffffffd9ffffffff0000000700000000",
            INIT_11 => X"000000e200000000ffffffa5ffffffff000000ab00000000ffffffe4ffffffff",
            INIT_12 => X"ffffff7efffffffffffffff6ffffffff0000002f00000000ffffffa2ffffffff",
            INIT_13 => X"00000007000000000000007000000000ffffffb4ffffffff0000003100000000",
            INIT_14 => X"0000004e000000000000006b000000000000007100000000ffffffeeffffffff",
            INIT_15 => X"ffffffc9fffffffffffffff8ffffffffffffff68ffffffffffffffa0ffffffff",
            INIT_16 => X"ffffffbfffffffffffffffd1ffffffffffffffdeffffffff0000000400000000",
            INIT_17 => X"00000008000000000000000000000000fffffff0ffffffffffffffe3ffffffff",
            INIT_18 => X"00000040000000000000003700000000ffffffd5ffffffff0000001100000000",
            INIT_19 => X"ffffffe8ffffffffffffff8affffffffffffffbcffffffffffffffe8ffffffff",
            INIT_1A => X"ffffffedfffffffffffffff5ffffffff0000008600000000ffffff9cffffffff",
            INIT_1B => X"ffffffe8fffffffffffffff8fffffffffffffffbffffffff0000004f00000000",
            INIT_1C => X"ffffffbcffffffff0000007b000000000000002b000000000000007400000000",
            INIT_1D => X"00000049000000000000003c000000000000004c00000000ffffffcdffffffff",
            INIT_1E => X"ffffffbfffffffff0000006400000000ffffffe0ffffffff0000001000000000",
            INIT_1F => X"ffffff7affffffffffffff87ffffffffffffffdcffffffff0000002800000000",
            INIT_20 => X"0000006500000000ffffff54ffffffff0000003100000000ffffffe8ffffffff",
            INIT_21 => X"0000004d000000000000002300000000fffffee0ffffffffffffffc5ffffffff",
            INIT_22 => X"fffffff8fffffffffffffff4ffffffff0000000f000000000000004100000000",
            INIT_23 => X"0000000600000000ffffff4fffffffffffffffbdffffffff0000000500000000",
            INIT_24 => X"00000033000000000000002c000000000000002b00000000ffffffebffffffff",
            INIT_25 => X"0000000f00000000ffffffc4ffffffffffffffb4ffffffffffffffe9ffffffff",
            INIT_26 => X"0000003600000000ffffff9cffffffff000000a600000000fffffff9ffffffff",
            INIT_27 => X"00000016000000000000002000000000ffffff46fffffffffffffff5ffffffff",
            INIT_28 => X"ffffffa8fffffffffffffff7ffffffffffffff3bfffffffffffffff2ffffffff",
            INIT_29 => X"ffffff91ffffffffffffff45ffffffff0000002c000000000000000f00000000",
            INIT_2A => X"ffffffecffffffffffffffb4ffffffffffffff9affffffff0000000000000000",
            INIT_2B => X"0000002000000000ffffffd9fffffffffffffffaffffffff0000003600000000",
            INIT_2C => X"00000004000000000000002900000000ffffff6bffffffffffffffe8ffffffff",
            INIT_2D => X"0000000e00000000ffffff96ffffffff00000045000000000000003900000000",
            INIT_2E => X"ffffffeeffffffff0000002300000000ffffffc3ffffffffffffffaaffffffff",
            INIT_2F => X"0000004600000000ffffffa6ffffffffffffff91ffffffff0000002f00000000",
            INIT_30 => X"000000de000000000000003700000000ffffffc5ffffffff0000000f00000000",
            INIT_31 => X"0000007800000000fffffff5ffffffffffffffe6fffffffffffffffeffffffff",
            INIT_32 => X"ffffffcbfffffffffffffffeffffffff00000003000000000000008600000000",
            INIT_33 => X"ffffffaeffffffffffffffcdffffffffffffffc8ffffffffffffff8cffffffff",
            INIT_34 => X"0000005200000000ffffffd6ffffffffffffffdfffffffffffffffeeffffffff",
            INIT_35 => X"ffffffb9ffffffff0000004700000000fffffffcffffffffffffff8bffffffff",
            INIT_36 => X"0000006d000000000000002900000000ffffffddffffffffffffffffffffffff",
            INIT_37 => X"fffffff9ffffffffffffffbcffffffffffffffcbffffffffffffffeeffffffff",
            INIT_38 => X"fffffffaffffffff000000a300000000ffffff06ffffffffffffffa5ffffffff",
            INIT_39 => X"ffffff47ffffffffffffff53ffffffff0000004f000000000000008000000000",
            INIT_3A => X"ffffffaaffffffffffffffb8ffffffffffffffedffffffffffffff32ffffffff",
            INIT_3B => X"ffffffeeffffffff000000490000000000000000000000000000001400000000",
            INIT_3C => X"ffffffbefffffffffffffff0ffffffffffffffdeffffffff0000004100000000",
            INIT_3D => X"ffffffc5ffffffff0000002d000000000000001300000000ffffffffffffffff",
            INIT_3E => X"00000036000000000000001d000000000000002f000000000000000e00000000",
            INIT_3F => X"ffffffdbffffffff0000004c00000000ffffffabffffffffffffffabffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004a000000000000003b000000000000005000000000fffffff1ffffffff",
            INIT_41 => X"ffffff71ffffffff0000008f00000000ffffffbaffffffffffffffd8ffffffff",
            INIT_42 => X"ffffffbaffffffffffffffe9ffffffff0000000500000000ffffff39ffffffff",
            INIT_43 => X"ffffffd4ffffffffffffff9bffffffffffffff82ffffffffffffffbaffffffff",
            INIT_44 => X"00000015000000000000003f000000000000002300000000fffffff3ffffffff",
            INIT_45 => X"000000a6000000000000004a00000000ffffff2affffffffffffffd7ffffffff",
            INIT_46 => X"ffffff87ffffffffffffffb8ffffffff0000009400000000fffffff6ffffffff",
            INIT_47 => X"fffffff1ffffffff0000005a00000000ffffff47ffffffffffffffd7ffffffff",
            INIT_48 => X"ffffffe9ffffffffffffff77ffffffffffffff5cffffffff0000000800000000",
            INIT_49 => X"ffffff24ffffffffffffffafffffffff0000006a00000000ffffffa5ffffffff",
            INIT_4A => X"ffffffaafffffffffffffff9ffffffffffffff67ffffffffffffff8fffffffff",
            INIT_4B => X"ffffffcbfffffffffffffff2ffffffff00000017000000000000002600000000",
            INIT_4C => X"ffffff48fffffffffffffffbffffffffffffffb3ffffffff0000004700000000",
            INIT_4D => X"ffffffe0fffffffffffffff6ffffffffffffffdcffffffffffffff8effffffff",
            INIT_4E => X"ffffffd2ffffffff0000003000000000fffffe44ffffffff0000003a00000000",
            INIT_4F => X"ffffffaeffffffff0000000900000000fffffffdffffffff0000004400000000",
            INIT_50 => X"0000007d000000000000004f00000000ffffffa0ffffffff0000000b00000000",
            INIT_51 => X"ffffffa8ffffffff0000000800000000ffffff42ffffffff0000006100000000",
            INIT_52 => X"0000006300000000ffffffeeffffffffffffffb8ffffffff0000000000000000",
            INIT_53 => X"ffffffc6ffffffff0000001f00000000ffffff8dffffffffffffffe6ffffffff",
            INIT_54 => X"ffffffe7ffffffff0000007500000000ffffff98fffffffffffffff2ffffffff",
            INIT_55 => X"ffffff6effffffffffffff98ffffffffffffff85ffffffffffffffe7ffffffff",
            INIT_56 => X"0000000100000000ffffffe5ffffffffffffffc6ffffffffffffffe4ffffffff",
            INIT_57 => X"ffffffeaffffffffffffff9cffffffffffffff3cffffffff0000002400000000",
            INIT_58 => X"00000014000000000000003200000000ffffff15ffffffff0000001400000000",
            INIT_59 => X"0000009e00000000ffffff89ffffffff000000a7000000000000002200000000",
            INIT_5A => X"ffffffc0ffffffffffffff80ffffffff00000052000000000000001700000000",
            INIT_5B => X"ffffff79ffffffffffffffccffffffff00000006000000000000002800000000",
            INIT_5C => X"ffffffd8ffffffffffffffbeffffffffffffff68ffffffff0000004200000000",
            INIT_5D => X"ffffffcaffffffffffffffddffffffff0000003e00000000ffffff1effffffff",
            INIT_5E => X"ffffff67ffffffff000000af000000000000003d00000000ffffff9fffffffff",
            INIT_5F => X"000000110000000000000033000000000000000f00000000ffffffd8ffffffff",
            INIT_60 => X"000000950000000000000060000000000000003f000000000000000600000000",
            INIT_61 => X"0000002200000000000000410000000000000062000000000000007b00000000",
            INIT_62 => X"0000002700000000ffffffefffffffffffffff9dfffffffffffffff9ffffffff",
            INIT_63 => X"0000001f000000000000001d00000000ffffffc3ffffffffffffff43ffffffff",
            INIT_64 => X"0000005b00000000ffffffc4ffffffffffffffbcffffffff0000001500000000",
            INIT_65 => X"0000003400000000ffffffaefffffffffffffffdffffffffffffffc7ffffffff",
            INIT_66 => X"0000003c00000000fffffff2ffffffffffffffedfffffffffffffffbffffffff",
            INIT_67 => X"ffffffe7ffffffff0000002600000000ffffffd1ffffffff0000005200000000",
            INIT_68 => X"ffffff6affffffff0000005c000000000000008a000000000000002f00000000",
            INIT_69 => X"000000e600000000ffffffa1ffffffff0000005800000000ffffff84ffffffff",
            INIT_6A => X"ffffff54ffffffffffffffc8ffffffff0000003e00000000fffffed9ffffffff",
            INIT_6B => X"ffffff81ffffffffffffffa6ffffffff0000001700000000ffffffc8ffffffff",
            INIT_6C => X"ffffffb8ffffffffffffff65ffffffffffffff8bffffffffffffffd1ffffffff",
            INIT_6D => X"fffffffdffffffff0000002700000000ffffffefffffffffffffff16ffffffff",
            INIT_6E => X"ffffff7cffffffff0000000d00000000ffffff70ffffffff0000004e00000000",
            INIT_6F => X"ffffffe3ffffffff0000005100000000ffffffbdffffffff0000002e00000000",
            INIT_70 => X"0000000000000000000000370000000000000107000000000000000300000000",
            INIT_71 => X"0000001b0000000000000033000000000000007a00000000ffffff98ffffffff",
            INIT_72 => X"ffffffa4ffffffff00000016000000000000000f00000000ffffff9fffffffff",
            INIT_73 => X"0000007e00000000fffffef2ffffffffffffffdeffffffffffffff1bffffffff",
            INIT_74 => X"0000002b00000000ffffffe4ffffffffffffffe4fffffffffffffff6ffffffff",
            INIT_75 => X"0000000a00000000ffffffafffffffff00000026000000000000002b00000000",
            INIT_76 => X"ffffff36ffffffff0000001c0000000000000029000000000000000700000000",
            INIT_77 => X"fffffff7ffffffff0000005700000000ffffff50ffffffffffffffafffffffff",
            INIT_78 => X"ffffff6dffffffffffffff73ffffffff0000000b000000000000001c00000000",
            INIT_79 => X"ffffffafffffffffffffffb4ffffffff000000e5000000000000005200000000",
            INIT_7A => X"ffffff7affffffffffffffeaffffffffffffff92ffffffff0000001400000000",
            INIT_7B => X"ffffffe9ffffffffffffffa7ffffffffffffffe8ffffffffffffffceffffffff",
            INIT_7C => X"0000000000000000ffffff98ffffffff00000066000000000000005a00000000",
            INIT_7D => X"ffffffb7fffffffffffffffeffffffffffffffecfffffffffffffee6ffffffff",
            INIT_7E => X"ffffffc5ffffffffffffffc9fffffffffffffeffffffffff0000000a00000000",
            INIT_7F => X"ffffffefffffffff0000005c000000000000006200000000ffffffbeffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE10;


    MEM_IWGHT_LAYER3_INSTANCE11 : if BRAM_NAME = "iwght_layer3_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffef4ffffffffffffffecffffffffffffff79fffffffffffffff4ffffffff",
            INIT_01 => X"ffffffc0ffffffff0000003500000000ffffff90ffffffffffffff7fffffffff",
            INIT_02 => X"0000008200000000fffffff2ffffffff0000001d000000000000000a00000000",
            INIT_03 => X"0000003900000000fffffed7ffffffff00000034000000000000001300000000",
            INIT_04 => X"0000002000000000fffffffeffffffffffffff9affffffff0000001100000000",
            INIT_05 => X"ffffffabffffffffffffffeaffffffffffffffebffffffffffffff94ffffffff",
            INIT_06 => X"ffffff7fffffffffffffffe9ffffffff00000037000000000000001000000000",
            INIT_07 => X"0000000b000000000000007300000000fffffffeffffffff0000003a00000000",
            INIT_08 => X"ffffff59ffffffffffffff9fffffffff00000010000000000000003500000000",
            INIT_09 => X"fffffff8ffffffff0000003e00000000000000d6000000000000002100000000",
            INIT_0A => X"00000066000000000000000e00000000ffffff77fffffffffffffff6ffffffff",
            INIT_0B => X"ffffffc3ffffffffffffffdaffffffff0000000400000000ffffffb7ffffffff",
            INIT_0C => X"00000011000000000000005c00000000ffffffc9ffffffff0000006000000000",
            INIT_0D => X"0000005000000000ffffffb6ffffffff0000001e00000000ffffff42ffffffff",
            INIT_0E => X"ffffffe0ffffffffffffffbfffffffffffffff62ffffffff0000000800000000",
            INIT_0F => X"ffffffe6ffffffffffffff92ffffffffffffffebffffffff0000004500000000",
            INIT_10 => X"ffffff17ffffffffffffff90ffffffffffffff34ffffffff0000000100000000",
            INIT_11 => X"ffffff52ffffffff0000000900000000ffffff7effffffffffffffc6ffffffff",
            INIT_12 => X"ffffffb5ffffffff0000000f00000000fffffffcffffffffffffffc1ffffffff",
            INIT_13 => X"0000004300000000ffffff56ffffffff0000000b00000000ffffff95ffffffff",
            INIT_14 => X"00000085000000000000008900000000ffffff53ffffffff0000000900000000",
            INIT_15 => X"0000002300000000ffffff86ffffffff00000006000000000000006400000000",
            INIT_16 => X"ffffffbdffffffff0000004100000000fffffff6ffffffff0000001000000000",
            INIT_17 => X"ffffffe8ffffffff0000007900000000ffffff79ffffffff0000003e00000000",
            INIT_18 => X"ffffff8effffffffffffff89ffffffff00000008000000000000000800000000",
            INIT_19 => X"fffffff5ffffffffffffffccffffffff0000009f00000000ffffffbdffffffff",
            INIT_1A => X"ffffffe2ffffffffffffff33ffffffffffffff1bffffffffffffff9effffffff",
            INIT_1B => X"0000000800000000ffffff89ffffffffffffffefffffffff0000002f00000000",
            INIT_1C => X"0000003100000000ffffff2cffffffff0000002a00000000ffffff89ffffffff",
            INIT_1D => X"ffffffc7ffffffff00000000000000000000000d00000000ffffff67ffffffff",
            INIT_1E => X"fffffff2ffffffff0000001700000000ffffff83ffffffffffffffeaffffffff",
            INIT_1F => X"0000007900000000000000310000000000000029000000000000008300000000",
            INIT_20 => X"0000004400000000ffffffa1ffffffffffffffa8ffffffffffffffe4ffffffff",
            INIT_21 => X"fffffff2ffffffffffffffebffffffff0000004b00000000ffffff20ffffffff",
            INIT_22 => X"fffffffbffffffffffffffa5ffffffff",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE11;


    MEM_IFMAP_LAYER0_INSTANCE0 : if BRAM_NAME = "ifmap_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a600000000000000a5000000000000009f000000000000009e00000000",
            INIT_01 => X"0000009f00000000000000a2000000000000009c00000000000000a000000000",
            INIT_02 => X"000000a000000000000000a1000000000000009f000000000000009e00000000",
            INIT_03 => X"000000aa00000000000000a900000000000000a600000000000000a100000000",
            INIT_04 => X"000000a000000000000000a000000000000000a200000000000000a700000000",
            INIT_05 => X"0000009400000000000000960000000000000095000000000000009c00000000",
            INIT_06 => X"0000008d000000000000008c000000000000008f000000000000009500000000",
            INIT_07 => X"00000074000000000000007e0000000000000089000000000000008f00000000",
            INIT_08 => X"000000a6000000000000009f0000000000000097000000000000009800000000",
            INIT_09 => X"000000a200000000000000a400000000000000a000000000000000a200000000",
            INIT_0A => X"0000009f000000000000009b000000000000009c00000000000000a300000000",
            INIT_0B => X"000000ab00000000000000ab00000000000000aa00000000000000a300000000",
            INIT_0C => X"00000097000000000000009a00000000000000a000000000000000a900000000",
            INIT_0D => X"0000008d000000000000008c000000000000008b000000000000009100000000",
            INIT_0E => X"0000008e00000000000000910000000000000093000000000000009500000000",
            INIT_0F => X"00000077000000000000007d0000000000000088000000000000008f00000000",
            INIT_10 => X"000000a7000000000000009e0000000000000097000000000000009700000000",
            INIT_11 => X"000000a500000000000000a500000000000000a300000000000000a000000000",
            INIT_12 => X"0000009d000000000000009e00000000000000a200000000000000a300000000",
            INIT_13 => X"000000a900000000000000a700000000000000a600000000000000a100000000",
            INIT_14 => X"000000790000000000000091000000000000009f00000000000000aa00000000",
            INIT_15 => X"0000007200000000000000650000000000000062000000000000006e00000000",
            INIT_16 => X"0000008c000000000000008f0000000000000086000000000000007800000000",
            INIT_17 => X"000000780000000000000082000000000000008b000000000000008e00000000",
            INIT_18 => X"000000ae00000000000000a0000000000000009b000000000000009b00000000",
            INIT_19 => X"000000a900000000000000a900000000000000a700000000000000a700000000",
            INIT_1A => X"000000bf00000000000000a700000000000000a500000000000000a500000000",
            INIT_1B => X"000000a400000000000000a2000000000000009d00000000000000b100000000",
            INIT_1C => X"0000006700000000000000680000000000000095000000000000009e00000000",
            INIT_1D => X"0000004a0000000000000050000000000000005c000000000000006200000000",
            INIT_1E => X"0000008400000000000000710000000000000053000000000000005600000000",
            INIT_1F => X"0000007f0000000000000088000000000000008c000000000000008c00000000",
            INIT_20 => X"000000aa00000000000000a1000000000000009c000000000000009b00000000",
            INIT_21 => X"000000a600000000000000a900000000000000a300000000000000a900000000",
            INIT_22 => X"000000f600000000000000ad00000000000000a400000000000000a400000000",
            INIT_23 => X"0000008e0000000000000092000000000000009700000000000000c300000000",
            INIT_24 => X"000000710000000000000055000000000000004e000000000000006f00000000",
            INIT_25 => X"0000005d0000000000000061000000000000006a000000000000007000000000",
            INIT_26 => X"0000006900000000000000550000000000000054000000000000004a00000000",
            INIT_27 => X"000000810000000000000085000000000000008a000000000000008000000000",
            INIT_28 => X"0000009300000000000000820000000000000085000000000000009400000000",
            INIT_29 => X"000000a700000000000000a700000000000000a500000000000000a100000000",
            INIT_2A => X"000000b400000000000000a300000000000000a500000000000000a300000000",
            INIT_2B => X"0000004200000000000000610000000000000080000000000000009d00000000",
            INIT_2C => X"0000007600000000000000590000000000000042000000000000004500000000",
            INIT_2D => X"0000005e00000000000000720000000000000077000000000000007a00000000",
            INIT_2E => X"00000043000000000000003a000000000000005b000000000000006300000000",
            INIT_2F => X"00000086000000000000008a000000000000008c000000000000006c00000000",
            INIT_30 => X"00000058000000000000002f000000000000006d000000000000007f00000000",
            INIT_31 => X"000000aa00000000000000a800000000000000aa000000000000009900000000",
            INIT_32 => X"0000009300000000000000a400000000000000a600000000000000a900000000",
            INIT_33 => X"000000440000000000000064000000000000007f000000000000008100000000",
            INIT_34 => X"0000008400000000000000530000000000000048000000000000004e00000000",
            INIT_35 => X"0000006b0000000000000069000000000000007c000000000000009200000000",
            INIT_36 => X"0000002e000000000000003f0000000000000055000000000000007300000000",
            INIT_37 => X"00000086000000000000008d0000000000000084000000000000004f00000000",
            INIT_38 => X"00000046000000000000002a0000000000000063000000000000008300000000",
            INIT_39 => X"000000a800000000000000a500000000000000a7000000000000008f00000000",
            INIT_3A => X"00000078000000000000008c00000000000000a100000000000000ab00000000",
            INIT_3B => X"0000005800000000000000740000000000000090000000000000008200000000",
            INIT_3C => X"0000007c000000000000004d0000000000000055000000000000005b00000000",
            INIT_3D => X"0000006a0000000000000066000000000000008800000000000000a300000000",
            INIT_3E => X"0000003100000000000000360000000000000055000000000000006400000000",
            INIT_3F => X"00000088000000000000008a000000000000006b000000000000003900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007c0000000000000036000000000000006700000000000000aa00000000",
            INIT_41 => X"000000a600000000000000a300000000000000a1000000000000009900000000",
            INIT_42 => X"0000007d000000000000007100000000000000ae00000000000000a500000000",
            INIT_43 => X"000000560000000000000079000000000000009c000000000000009d00000000",
            INIT_44 => X"0000005100000000000000500000000000000054000000000000005200000000",
            INIT_45 => X"0000005700000000000000710000000000000092000000000000008a00000000",
            INIT_46 => X"0000003800000000000000470000000000000056000000000000005300000000",
            INIT_47 => X"000000890000000000000085000000000000004a000000000000002800000000",
            INIT_48 => X"0000009a000000000000005e000000000000008600000000000000b400000000",
            INIT_49 => X"00000099000000000000009c000000000000009e00000000000000ae00000000",
            INIT_4A => X"0000009c00000000000000cf00000000000000ed00000000000000cf00000000",
            INIT_4B => X"0000005d000000000000007d000000000000009400000000000000ae00000000",
            INIT_4C => X"0000004c000000000000003b000000000000004a000000000000005600000000",
            INIT_4D => X"0000006a0000000000000085000000000000008f000000000000008900000000",
            INIT_4E => X"0000004b00000000000000540000000000000057000000000000005600000000",
            INIT_4F => X"00000084000000000000005f0000000000000028000000000000003200000000",
            INIT_50 => X"000000a5000000000000008e000000000000006c00000000000000b700000000",
            INIT_51 => X"0000007a000000000000009f000000000000009b00000000000000b100000000",
            INIT_52 => X"000000a400000000000000dc00000000000000ed00000000000000d500000000",
            INIT_53 => X"00000078000000000000007d000000000000009c00000000000000b700000000",
            INIT_54 => X"0000005b000000000000002d0000000000000050000000000000004e00000000",
            INIT_55 => X"0000006b000000000000009b000000000000009d00000000000000af00000000",
            INIT_56 => X"0000004e00000000000000580000000000000067000000000000005700000000",
            INIT_57 => X"00000068000000000000003b0000000000000029000000000000003b00000000",
            INIT_58 => X"000000aa0000000000000087000000000000006400000000000000bc00000000",
            INIT_59 => X"0000008600000000000000ad00000000000000a600000000000000bb00000000",
            INIT_5A => X"000000aa00000000000000c700000000000000c2000000000000007500000000",
            INIT_5B => X"00000075000000000000008600000000000000bd00000000000000b900000000",
            INIT_5C => X"0000007d00000000000000260000000000000054000000000000006600000000",
            INIT_5D => X"0000005d000000000000009200000000000000a000000000000000d200000000",
            INIT_5E => X"000000550000000000000068000000000000005e000000000000005300000000",
            INIT_5F => X"0000004c000000000000003e0000000000000037000000000000004900000000",
            INIT_60 => X"000000af000000000000007f000000000000005a00000000000000bd00000000",
            INIT_61 => X"0000009f00000000000000b200000000000000a600000000000000ae00000000",
            INIT_62 => X"0000008900000000000000a800000000000000a8000000000000006100000000",
            INIT_63 => X"0000007b00000000000000a000000000000000d800000000000000ba00000000",
            INIT_64 => X"0000009600000000000000320000000000000073000000000000007800000000",
            INIT_65 => X"0000005b000000000000007b000000000000009b00000000000000c200000000",
            INIT_66 => X"00000056000000000000005f0000000000000054000000000000005400000000",
            INIT_67 => X"00000049000000000000004f0000000000000049000000000000005400000000",
            INIT_68 => X"000000b90000000000000098000000000000005d00000000000000bd00000000",
            INIT_69 => X"000000a700000000000000ad0000000000000088000000000000007700000000",
            INIT_6A => X"000000a700000000000000910000000000000093000000000000006700000000",
            INIT_6B => X"0000008d00000000000000b400000000000000e200000000000000bd00000000",
            INIT_6C => X"0000009a00000000000000470000000000000075000000000000007e00000000",
            INIT_6D => X"000000570000000000000072000000000000009500000000000000ba00000000",
            INIT_6E => X"0000006300000000000000500000000000000048000000000000005000000000",
            INIT_6F => X"0000005e0000000000000061000000000000005a000000000000006400000000",
            INIT_70 => X"000000ba00000000000000a8000000000000006c00000000000000c200000000",
            INIT_71 => X"000000a7000000000000009c0000000000000063000000000000006900000000",
            INIT_72 => X"000000c6000000000000008a0000000000000073000000000000006400000000",
            INIT_73 => X"0000009a000000000000009100000000000000ac00000000000000be00000000",
            INIT_74 => X"0000009800000000000000470000000000000067000000000000009200000000",
            INIT_75 => X"0000006e0000000000000082000000000000008900000000000000b300000000",
            INIT_76 => X"0000006d000000000000005f000000000000005b000000000000005500000000",
            INIT_77 => X"0000007500000000000000610000000000000064000000000000007300000000",
            INIT_78 => X"000000b800000000000000ac000000000000008400000000000000c500000000",
            INIT_79 => X"0000009b000000000000008c000000000000004e000000000000008200000000",
            INIT_7A => X"000000e6000000000000008f0000000000000082000000000000007300000000",
            INIT_7B => X"000000830000000000000087000000000000009100000000000000f200000000",
            INIT_7C => X"00000090000000000000005f000000000000006c000000000000007900000000",
            INIT_7D => X"000000570000000000000070000000000000009800000000000000a800000000",
            INIT_7E => X"0000007000000000000000690000000000000057000000000000004700000000",
            INIT_7F => X"0000008800000000000000790000000000000067000000000000007800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE0;


    MEM_IFMAP_LAYER0_INSTANCE1 : if BRAM_NAME = "ifmap_layer0_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bf00000000000000a8000000000000009200000000000000cb00000000",
            INIT_01 => X"0000008a000000000000007e000000000000004e00000000000000a800000000",
            INIT_02 => X"000000ad000000000000009a0000000000000060000000000000008a00000000",
            INIT_03 => X"000000710000000000000071000000000000008c00000000000000a200000000",
            INIT_04 => X"000000ab00000000000000700000000000000069000000000000006500000000",
            INIT_05 => X"0000006d00000000000000870000000000000094000000000000009c00000000",
            INIT_06 => X"00000065000000000000005e000000000000004f000000000000004e00000000",
            INIT_07 => X"000000900000000000000097000000000000007d000000000000006b00000000",
            INIT_08 => X"000000b700000000000000a400000000000000a300000000000000d600000000",
            INIT_09 => X"0000009c0000000000000060000000000000005e00000000000000b000000000",
            INIT_0A => X"000000760000000000000081000000000000006a000000000000009400000000",
            INIT_0B => X"0000007300000000000000660000000000000074000000000000007200000000",
            INIT_0C => X"0000007600000000000000900000000000000065000000000000005600000000",
            INIT_0D => X"0000004b00000000000000850000000000000080000000000000004400000000",
            INIT_0E => X"000000660000000000000047000000000000003a000000000000003c00000000",
            INIT_0F => X"0000008c0000000000000096000000000000008f000000000000007400000000",
            INIT_10 => X"000000ad00000000000000a700000000000000b200000000000000d400000000",
            INIT_11 => X"0000008d0000000000000056000000000000007c00000000000000b000000000",
            INIT_12 => X"0000004d00000000000000680000000000000087000000000000009900000000",
            INIT_13 => X"000000930000000000000081000000000000007c000000000000008600000000",
            INIT_14 => X"000000840000000000000096000000000000005c000000000000005500000000",
            INIT_15 => X"00000040000000000000004b000000000000006b000000000000007500000000",
            INIT_16 => X"0000008500000000000000560000000000000041000000000000002c00000000",
            INIT_17 => X"00000097000000000000009a00000000000000a0000000000000009b00000000",
            INIT_18 => X"000000ae00000000000000ab00000000000000bb00000000000000c700000000",
            INIT_19 => X"000000770000000000000056000000000000009000000000000000b100000000",
            INIT_1A => X"0000004600000000000000900000000000000089000000000000007a00000000",
            INIT_1B => X"000000b80000000000000091000000000000006c000000000000008100000000",
            INIT_1C => X"0000008900000000000000830000000000000049000000000000007400000000",
            INIT_1D => X"0000003400000000000000330000000000000059000000000000008600000000",
            INIT_1E => X"000000a30000000000000079000000000000005a000000000000002f00000000",
            INIT_1F => X"00000095000000000000009e00000000000000a400000000000000ab00000000",
            INIT_20 => X"000000b100000000000000b300000000000000c300000000000000a500000000",
            INIT_21 => X"000000830000000000000063000000000000009800000000000000b500000000",
            INIT_22 => X"00000050000000000000005d000000000000006700000000000000ab00000000",
            INIT_23 => X"000000bf00000000000000b2000000000000007a000000000000005d00000000",
            INIT_24 => X"0000005700000000000000590000000000000064000000000000009600000000",
            INIT_25 => X"000000180000000000000026000000000000002e000000000000003c00000000",
            INIT_26 => X"00000090000000000000006c000000000000003c000000000000002e00000000",
            INIT_27 => X"00000078000000000000007f0000000000000080000000000000009000000000",
            INIT_28 => X"000000b200000000000000b100000000000000c3000000000000007500000000",
            INIT_29 => X"000000960000000000000053000000000000008a00000000000000b500000000",
            INIT_2A => X"00000086000000000000008500000000000000db00000000000000f500000000",
            INIT_2B => X"000000c200000000000000be00000000000000b0000000000000009500000000",
            INIT_2C => X"0000003d000000000000006e000000000000007d00000000000000a800000000",
            INIT_2D => X"0000003a00000000000000310000000000000022000000000000002300000000",
            INIT_2E => X"000000480000000000000045000000000000003a000000000000003d00000000",
            INIT_2F => X"00000037000000000000003b0000000000000045000000000000004e00000000",
            INIT_30 => X"000000b000000000000000ae00000000000000af000000000000004f00000000",
            INIT_31 => X"000000d3000000000000006d000000000000008c00000000000000b100000000",
            INIT_32 => X"0000007c00000000000000d000000000000000fc00000000000000fd00000000",
            INIT_33 => X"0000007a0000000000000074000000000000007c000000000000007200000000",
            INIT_34 => X"0000003c00000000000000440000000000000044000000000000006800000000",
            INIT_35 => X"0000003800000000000000330000000000000032000000000000003400000000",
            INIT_36 => X"00000033000000000000002b0000000000000033000000000000003800000000",
            INIT_37 => X"0000002a000000000000002b0000000000000030000000000000003b00000000",
            INIT_38 => X"000000a800000000000000900000000000000060000000000000002900000000",
            INIT_39 => X"000000f600000000000000a500000000000000a500000000000000b200000000",
            INIT_3A => X"0000003c000000000000006e00000000000000e300000000000000fd00000000",
            INIT_3B => X"0000003000000000000000310000000000000031000000000000003500000000",
            INIT_3C => X"0000002a000000000000002e000000000000002a000000000000002d00000000",
            INIT_3D => X"0000002b000000000000002e000000000000002e000000000000002600000000",
            INIT_3E => X"00000032000000000000002e000000000000002e000000000000002a00000000",
            INIT_3F => X"0000002d00000000000000330000000000000035000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000083000000000000003b000000000000001d000000000000001d00000000",
            INIT_41 => X"000000fe00000000000000c2000000000000008400000000000000a600000000",
            INIT_42 => X"00000032000000000000003d000000000000008d00000000000000f100000000",
            INIT_43 => X"0000003200000000000000310000000000000033000000000000003200000000",
            INIT_44 => X"000000220000000000000027000000000000002a000000000000002f00000000",
            INIT_45 => X"0000002a00000000000000260000000000000027000000000000002300000000",
            INIT_46 => X"0000003b000000000000003e0000000000000038000000000000002d00000000",
            INIT_47 => X"00000033000000000000002e0000000000000032000000000000003800000000",
            INIT_48 => X"000000490000000000000022000000000000001e000000000000003000000000",
            INIT_49 => X"0000010000000000000000d70000000000000080000000000000008000000000",
            INIT_4A => X"000000320000000000000036000000000000004200000000000000bb00000000",
            INIT_4B => X"0000002d000000000000002e0000000000000034000000000000003400000000",
            INIT_4C => X"0000002700000000000000240000000000000029000000000000002b00000000",
            INIT_4D => X"0000002e000000000000002b0000000000000028000000000000002800000000",
            INIT_4E => X"0000003b0000000000000040000000000000003e000000000000003b00000000",
            INIT_4F => X"0000005300000000000000460000000000000032000000000000003600000000",
            INIT_50 => X"00000029000000000000001f0000000000000023000000000000003400000000",
            INIT_51 => X"000000f000000000000000e00000000000000080000000000000004200000000",
            INIT_52 => X"000000380000000000000031000000000000003a000000000000007c00000000",
            INIT_53 => X"0000002f000000000000002c000000000000002c000000000000003600000000",
            INIT_54 => X"0000002c000000000000002b000000000000002b000000000000002e00000000",
            INIT_55 => X"0000003a0000000000000036000000000000002d000000000000002c00000000",
            INIT_56 => X"00000024000000000000002b000000000000002e000000000000003600000000",
            INIT_57 => X"0000004c00000000000000550000000000000049000000000000003300000000",
            INIT_58 => X"00000023000000000000001d0000000000000023000000000000003200000000",
            INIT_59 => X"000000d300000000000000ca000000000000004e000000000000002c00000000",
            INIT_5A => X"0000003000000000000000360000000000000041000000000000006100000000",
            INIT_5B => X"0000002d00000000000000280000000000000030000000000000003a00000000",
            INIT_5C => X"0000002e000000000000002f0000000000000030000000000000002f00000000",
            INIT_5D => X"0000003000000000000000270000000000000027000000000000003300000000",
            INIT_5E => X"00000028000000000000001c0000000000000027000000000000002f00000000",
            INIT_5F => X"00000033000000000000002e0000000000000043000000000000004300000000",
            INIT_60 => X"0000002100000000000000200000000000000023000000000000003200000000",
            INIT_61 => X"000000aa0000000000000068000000000000002e000000000000002900000000",
            INIT_62 => X"0000003500000000000000340000000000000036000000000000004000000000",
            INIT_63 => X"0000002d0000000000000036000000000000003a000000000000003d00000000",
            INIT_64 => X"00000031000000000000002e0000000000000029000000000000002a00000000",
            INIT_65 => X"000000270000000000000028000000000000002a000000000000002e00000000",
            INIT_66 => X"0000003f000000000000002c0000000000000028000000000000002500000000",
            INIT_67 => X"00000033000000000000000f000000000000001f000000000000002f00000000",
            INIT_68 => X"00000026000000000000001f000000000000002a000000000000004400000000",
            INIT_69 => X"00000047000000000000002a000000000000002b000000000000002500000000",
            INIT_6A => X"00000026000000000000001b000000000000001f000000000000003100000000",
            INIT_6B => X"00000035000000000000003a0000000000000038000000000000003100000000",
            INIT_6C => X"000000350000000000000039000000000000003c000000000000003800000000",
            INIT_6D => X"000000210000000000000027000000000000002d000000000000003200000000",
            INIT_6E => X"00000049000000000000004f000000000000003e000000000000002a00000000",
            INIT_6F => X"00000028000000000000000d0000000000000026000000000000003800000000",
            INIT_70 => X"0000002b00000000000000230000000000000031000000000000003d00000000",
            INIT_71 => X"00000028000000000000002c000000000000002a000000000000002700000000",
            INIT_72 => X"0000001e0000000000000017000000000000001b000000000000002a00000000",
            INIT_73 => X"0000002f0000000000000024000000000000001d000000000000001b00000000",
            INIT_74 => X"0000004b0000000000000042000000000000003e000000000000003800000000",
            INIT_75 => X"0000002b000000000000002b0000000000000031000000000000004500000000",
            INIT_76 => X"0000005d000000000000006d0000000000000055000000000000003c00000000",
            INIT_77 => X"00000014000000000000001d000000000000001a000000000000003c00000000",
            INIT_78 => X"0000002b000000000000002d0000000000000038000000000000003600000000",
            INIT_79 => X"0000002600000000000000280000000000000028000000000000002800000000",
            INIT_7A => X"0000001d0000000000000016000000000000001a000000000000002400000000",
            INIT_7B => X"000000120000000000000013000000000000001d000000000000001900000000",
            INIT_7C => X"0000004a000000000000003d000000000000002f000000000000002000000000",
            INIT_7D => X"0000002d00000000000000340000000000000035000000000000004200000000",
            INIT_7E => X"0000005900000000000000690000000000000059000000000000004300000000",
            INIT_7F => X"0000001500000000000000220000000000000018000000000000003000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE1;


    MEM_IFMAP_LAYER0_INSTANCE2 : if BRAM_NAME = "ifmap_layer0_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000760000000000000074000000000000006f000000000000007000000000",
            INIT_01 => X"000000710000000000000073000000000000006d000000000000007000000000",
            INIT_02 => X"0000006f00000000000000740000000000000071000000000000006f00000000",
            INIT_03 => X"0000007700000000000000750000000000000075000000000000006f00000000",
            INIT_04 => X"00000070000000000000006f0000000000000071000000000000007500000000",
            INIT_05 => X"0000006a000000000000006b000000000000006b000000000000006d00000000",
            INIT_06 => X"0000006100000000000000620000000000000065000000000000006b00000000",
            INIT_07 => X"00000055000000000000005b000000000000005f000000000000006100000000",
            INIT_08 => X"000000740000000000000072000000000000006e000000000000007000000000",
            INIT_09 => X"0000007200000000000000750000000000000071000000000000007000000000",
            INIT_0A => X"0000006e000000000000006f000000000000006e000000000000007400000000",
            INIT_0B => X"0000007300000000000000750000000000000077000000000000007100000000",
            INIT_0C => X"000000730000000000000070000000000000006f000000000000007300000000",
            INIT_0D => X"0000006400000000000000660000000000000068000000000000006e00000000",
            INIT_0E => X"0000006100000000000000660000000000000066000000000000006900000000",
            INIT_0F => X"00000058000000000000005b000000000000005f000000000000006200000000",
            INIT_10 => X"0000006f000000000000006f000000000000006d000000000000006e00000000",
            INIT_11 => X"0000007500000000000000750000000000000073000000000000006a00000000",
            INIT_12 => X"0000006d00000000000000720000000000000073000000000000007300000000",
            INIT_13 => X"0000007100000000000000720000000000000073000000000000006f00000000",
            INIT_14 => X"00000060000000000000006f0000000000000072000000000000007400000000",
            INIT_15 => X"00000055000000000000004d000000000000004e000000000000005a00000000",
            INIT_16 => X"0000006300000000000000670000000000000060000000000000005600000000",
            INIT_17 => X"00000059000000000000005f0000000000000062000000000000006300000000",
            INIT_18 => X"00000070000000000000006d000000000000006e000000000000006b00000000",
            INIT_19 => X"0000007700000000000000780000000000000075000000000000006e00000000",
            INIT_1A => X"00000092000000000000007b0000000000000075000000000000007300000000",
            INIT_1B => X"000000720000000000000073000000000000006f000000000000008200000000",
            INIT_1C => X"000000570000000000000050000000000000006f000000000000007000000000",
            INIT_1D => X"0000003f000000000000004b000000000000005a000000000000005a00000000",
            INIT_1E => X"000000620000000000000055000000000000003e000000000000004600000000",
            INIT_1F => X"0000005e00000000000000630000000000000065000000000000006600000000",
            INIT_20 => X"0000007200000000000000730000000000000072000000000000006b00000000",
            INIT_21 => X"0000007400000000000000780000000000000071000000000000007200000000",
            INIT_22 => X"000000d600000000000000800000000000000074000000000000007100000000",
            INIT_23 => X"0000006c000000000000006f0000000000000072000000000000009c00000000",
            INIT_24 => X"0000006700000000000000450000000000000035000000000000005000000000",
            INIT_25 => X"0000005e00000000000000660000000000000072000000000000006e00000000",
            INIT_26 => X"000000530000000000000049000000000000004e000000000000004800000000",
            INIT_27 => X"0000005d000000000000005e0000000000000065000000000000006000000000",
            INIT_28 => X"0000007000000000000000640000000000000068000000000000006d00000000",
            INIT_29 => X"0000007300000000000000740000000000000071000000000000007300000000",
            INIT_2A => X"0000008a00000000000000760000000000000074000000000000006f00000000",
            INIT_2B => X"00000032000000000000004b0000000000000066000000000000007a00000000",
            INIT_2C => X"0000007100000000000000530000000000000038000000000000003a00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007900000000",
            INIT_2E => X"0000003a000000000000003a000000000000005b000000000000006400000000",
            INIT_2F => X"0000005f00000000000000620000000000000069000000000000005400000000",
            INIT_30 => X"0000004a0000000000000025000000000000005f000000000000006400000000",
            INIT_31 => X"0000007600000000000000730000000000000076000000000000007500000000",
            INIT_32 => X"0000006b00000000000000780000000000000074000000000000007500000000",
            INIT_33 => X"000000430000000000000057000000000000006c000000000000006200000000",
            INIT_34 => X"000000820000000000000054000000000000004b000000000000005300000000",
            INIT_35 => X"0000006600000000000000630000000000000076000000000000008e00000000",
            INIT_36 => X"0000002f00000000000000470000000000000053000000000000006f00000000",
            INIT_37 => X"0000005d00000000000000630000000000000062000000000000003d00000000",
            INIT_38 => X"00000040000000000000002b0000000000000060000000000000007300000000",
            INIT_39 => X"0000007400000000000000720000000000000075000000000000006f00000000",
            INIT_3A => X"0000005e000000000000006d0000000000000071000000000000007700000000",
            INIT_3B => X"00000057000000000000006a0000000000000083000000000000006e00000000",
            INIT_3C => X"00000076000000000000004d0000000000000058000000000000005f00000000",
            INIT_3D => X"00000062000000000000005d000000000000007c000000000000009900000000",
            INIT_3E => X"00000035000000000000003c0000000000000051000000000000005d00000000",
            INIT_3F => X"0000006100000000000000670000000000000053000000000000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000079000000000000003a000000000000006900000000000000a100000000",
            INIT_41 => X"0000007a00000000000000750000000000000071000000000000007c00000000",
            INIT_42 => X"0000006900000000000000590000000000000087000000000000007900000000",
            INIT_43 => X"00000050000000000000006f000000000000008f000000000000008d00000000",
            INIT_44 => X"00000047000000000000004e0000000000000055000000000000005100000000",
            INIT_45 => X"0000004f00000000000000670000000000000087000000000000007d00000000",
            INIT_46 => X"0000003900000000000000490000000000000052000000000000004d00000000",
            INIT_47 => X"00000067000000000000006a000000000000003b000000000000002300000000",
            INIT_48 => X"0000009a0000000000000064000000000000008b00000000000000b000000000",
            INIT_49 => X"0000007600000000000000740000000000000074000000000000009500000000",
            INIT_4A => X"0000008300000000000000b400000000000000d600000000000000b400000000",
            INIT_4B => X"00000055000000000000006e0000000000000083000000000000009900000000",
            INIT_4C => X"000000440000000000000039000000000000004a000000000000005400000000",
            INIT_4D => X"00000062000000000000007c0000000000000085000000000000007d00000000",
            INIT_4E => X"0000004c00000000000000550000000000000055000000000000005100000000",
            INIT_4F => X"00000067000000000000004b000000000000001e000000000000003100000000",
            INIT_50 => X"000000a90000000000000097000000000000007400000000000000b700000000",
            INIT_51 => X"0000005900000000000000760000000000000070000000000000009c00000000",
            INIT_52 => X"0000008700000000000000bf00000000000000e000000000000000c500000000",
            INIT_53 => X"0000006f000000000000006c0000000000000089000000000000009f00000000",
            INIT_54 => X"00000055000000000000002c0000000000000050000000000000004c00000000",
            INIT_55 => X"000000640000000000000093000000000000009300000000000000a500000000",
            INIT_56 => X"0000004f00000000000000580000000000000066000000000000005300000000",
            INIT_57 => X"00000051000000000000002e0000000000000024000000000000003b00000000",
            INIT_58 => X"000000af0000000000000090000000000000006c00000000000000bf00000000",
            INIT_59 => X"0000005d000000000000007b000000000000007800000000000000a700000000",
            INIT_5A => X"0000008e00000000000000ab00000000000000b6000000000000005f00000000",
            INIT_5B => X"0000006b000000000000007700000000000000ab00000000000000a100000000",
            INIT_5C => X"0000007900000000000000260000000000000054000000000000006200000000",
            INIT_5D => X"00000059000000000000008b000000000000009800000000000000c900000000",
            INIT_5E => X"000000570000000000000068000000000000005d000000000000005000000000",
            INIT_5F => X"0000003800000000000000370000000000000035000000000000004b00000000",
            INIT_60 => X"000000b40000000000000086000000000000006000000000000000c200000000",
            INIT_61 => X"0000006d000000000000007b000000000000007b000000000000009c00000000",
            INIT_62 => X"000000720000000000000090000000000000009a000000000000004400000000",
            INIT_63 => X"00000071000000000000009500000000000000ca00000000000000a600000000",
            INIT_64 => X"0000009300000000000000320000000000000072000000000000007200000000",
            INIT_65 => X"000000580000000000000076000000000000009500000000000000bb00000000",
            INIT_66 => X"00000057000000000000005f0000000000000054000000000000005300000000",
            INIT_67 => X"00000037000000000000004a0000000000000049000000000000005700000000",
            INIT_68 => X"000000bc000000000000009a000000000000005f00000000000000c000000000",
            INIT_69 => X"00000074000000000000007c000000000000006a000000000000006e00000000",
            INIT_6A => X"00000095000000000000007d0000000000000084000000000000004800000000",
            INIT_6B => X"0000008300000000000000ac00000000000000d800000000000000ae00000000",
            INIT_6C => X"0000009800000000000000470000000000000072000000000000007500000000",
            INIT_6D => X"00000055000000000000006e000000000000009000000000000000b500000000",
            INIT_6E => X"0000006400000000000000500000000000000049000000000000005000000000",
            INIT_6F => X"0000004900000000000000590000000000000058000000000000006500000000",
            INIT_70 => X"000000ba00000000000000a7000000000000006b00000000000000c400000000",
            INIT_71 => X"0000007a00000000000000770000000000000059000000000000006d00000000",
            INIT_72 => X"000000b9000000000000007b000000000000006a000000000000004a00000000",
            INIT_73 => X"0000008f000000000000008c00000000000000a500000000000000b400000000",
            INIT_74 => X"0000009800000000000000470000000000000064000000000000008800000000",
            INIT_75 => X"0000006d0000000000000080000000000000008500000000000000af00000000",
            INIT_76 => X"0000006e0000000000000060000000000000005d000000000000005600000000",
            INIT_77 => X"0000005f00000000000000550000000000000060000000000000007400000000",
            INIT_78 => X"000000b200000000000000a7000000000000008100000000000000c500000000",
            INIT_79 => X"0000007d00000000000000780000000000000053000000000000008900000000",
            INIT_7A => X"000000dd00000000000000830000000000000078000000000000005e00000000",
            INIT_7B => X"000000790000000000000082000000000000008a00000000000000ec00000000",
            INIT_7C => X"0000008600000000000000580000000000000068000000000000007000000000",
            INIT_7D => X"00000055000000000000006c0000000000000093000000000000009f00000000",
            INIT_7E => X"0000006d00000000000000680000000000000058000000000000004800000000",
            INIT_7F => X"0000006800000000000000600000000000000056000000000000006e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE2;


    MEM_IFMAP_LAYER0_INSTANCE3 : if BRAM_NAME = "ifmap_layer0_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b600000000000000a4000000000000009200000000000000cb00000000",
            INIT_01 => X"0000007e000000000000007d000000000000005600000000000000aa00000000",
            INIT_02 => X"000000a3000000000000008f0000000000000050000000000000007900000000",
            INIT_03 => X"0000006a000000000000006a0000000000000084000000000000009800000000",
            INIT_04 => X"0000008f000000000000005a0000000000000065000000000000006500000000",
            INIT_05 => X"000000690000000000000082000000000000008d000000000000008a00000000",
            INIT_06 => X"0000005b000000000000005d000000000000004f000000000000004c00000000",
            INIT_07 => X"00000068000000000000006c0000000000000058000000000000005300000000",
            INIT_08 => X"000000b800000000000000a700000000000000a600000000000000d700000000",
            INIT_09 => X"000000950000000000000060000000000000006600000000000000b600000000",
            INIT_0A => X"000000690000000000000074000000000000005d000000000000008900000000",
            INIT_0B => X"0000006e000000000000005b0000000000000069000000000000006600000000",
            INIT_0C => X"0000006000000000000000800000000000000067000000000000005b00000000",
            INIT_0D => X"00000045000000000000007e0000000000000078000000000000003800000000",
            INIT_0E => X"0000005d00000000000000460000000000000038000000000000003800000000",
            INIT_0F => X"0000006e00000000000000740000000000000070000000000000005e00000000",
            INIT_10 => X"000000b500000000000000af00000000000000b800000000000000d300000000",
            INIT_11 => X"0000008b0000000000000058000000000000008300000000000000b800000000",
            INIT_12 => X"00000040000000000000005a0000000000000080000000000000009400000000",
            INIT_13 => X"0000008f0000000000000075000000000000006f000000000000007900000000",
            INIT_14 => X"00000075000000000000008b0000000000000060000000000000005c00000000",
            INIT_15 => X"0000003b00000000000000440000000000000063000000000000006d00000000",
            INIT_16 => X"000000690000000000000045000000000000003e000000000000002900000000",
            INIT_17 => X"0000006f00000000000000730000000000000078000000000000007700000000",
            INIT_18 => X"000000b300000000000000b000000000000000bd00000000000000c000000000",
            INIT_19 => X"00000079000000000000005a000000000000009500000000000000b600000000",
            INIT_1A => X"0000003b00000000000000860000000000000088000000000000007c00000000",
            INIT_1B => X"000000b000000000000000860000000000000061000000000000007600000000",
            INIT_1C => X"0000007c0000000000000077000000000000004b000000000000007600000000",
            INIT_1D => X"0000003300000000000000310000000000000056000000000000008100000000",
            INIT_1E => X"00000076000000000000005b000000000000005a000000000000003100000000",
            INIT_1F => X"0000006b000000000000006f0000000000000071000000000000007900000000",
            INIT_20 => X"000000ad00000000000000b200000000000000c1000000000000009c00000000",
            INIT_21 => X"000000870000000000000067000000000000009d00000000000000b500000000",
            INIT_22 => X"0000004d000000000000005a000000000000006900000000000000af00000000",
            INIT_23 => X"000000b600000000000000ad0000000000000076000000000000005a00000000",
            INIT_24 => X"0000004d000000000000004e0000000000000064000000000000009400000000",
            INIT_25 => X"00000021000000000000002e0000000000000034000000000000003d00000000",
            INIT_26 => X"0000007d00000000000000640000000000000047000000000000003900000000",
            INIT_27 => X"000000690000000000000071000000000000006d000000000000007b00000000",
            INIT_28 => X"000000a900000000000000b200000000000000c8000000000000007800000000",
            INIT_29 => X"000000990000000000000057000000000000009000000000000000b300000000",
            INIT_2A => X"0000008d000000000000008c00000000000000de00000000000000f700000000",
            INIT_2B => X"000000c000000000000000c400000000000000b6000000000000009c00000000",
            INIT_2C => X"0000003e000000000000006d000000000000008500000000000000ac00000000",
            INIT_2D => X"0000005100000000000000460000000000000036000000000000003100000000",
            INIT_2E => X"0000006500000000000000630000000000000054000000000000005500000000",
            INIT_2F => X"0000005a000000000000005c0000000000000060000000000000006800000000",
            INIT_30 => X"000000ac00000000000000b700000000000000c5000000000000006900000000",
            INIT_31 => X"000000d30000000000000070000000000000009200000000000000b100000000",
            INIT_32 => X"0000008f00000000000000e000000000000000fd00000000000000fc00000000",
            INIT_33 => X"000000850000000000000085000000000000008d000000000000008400000000",
            INIT_34 => X"000000520000000000000057000000000000005d000000000000007c00000000",
            INIT_35 => X"0000005d00000000000000550000000000000054000000000000005400000000",
            INIT_36 => X"000000680000000000000060000000000000005b000000000000005e00000000",
            INIT_37 => X"0000005f00000000000000610000000000000061000000000000006c00000000",
            INIT_38 => X"000000ae00000000000000a80000000000000089000000000000005900000000",
            INIT_39 => X"000000f500000000000000a600000000000000aa00000000000000b600000000",
            INIT_3A => X"00000058000000000000008800000000000000e700000000000000fb00000000",
            INIT_3B => X"00000048000000000000004b000000000000004c000000000000005000000000",
            INIT_3C => X"0000005200000000000000510000000000000051000000000000004f00000000",
            INIT_3D => X"000000570000000000000059000000000000005a000000000000005600000000",
            INIT_3E => X"00000060000000000000005e000000000000005d000000000000005900000000",
            INIT_3F => X"0000005a000000000000005f000000000000005e000000000000006000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009900000000000000660000000000000057000000000000005b00000000",
            INIT_41 => X"000000fa00000000000000bd000000000000008800000000000000b300000000",
            INIT_42 => X"00000054000000000000005e000000000000009f00000000000000f500000000",
            INIT_43 => X"0000005400000000000000530000000000000055000000000000005400000000",
            INIT_44 => X"0000004f00000000000000520000000000000054000000000000005600000000",
            INIT_45 => X"0000005900000000000000550000000000000056000000000000005300000000",
            INIT_46 => X"0000006500000000000000670000000000000067000000000000005c00000000",
            INIT_47 => X"00000067000000000000005e0000000000000063000000000000006600000000",
            INIT_48 => X"0000006a0000000000000055000000000000005e000000000000006f00000000",
            INIT_49 => X"000000fd00000000000000d50000000000000088000000000000009400000000",
            INIT_4A => X"00000058000000000000005b000000000000005d00000000000000c600000000",
            INIT_4B => X"000000520000000000000053000000000000005a000000000000005a00000000",
            INIT_4C => X"0000005300000000000000500000000000000051000000000000005200000000",
            INIT_4D => X"0000005f000000000000005c0000000000000059000000000000005600000000",
            INIT_4E => X"0000006c000000000000006d000000000000006e000000000000006c00000000",
            INIT_4F => X"00000089000000000000007b0000000000000069000000000000006c00000000",
            INIT_50 => X"0000005300000000000000560000000000000063000000000000007200000000",
            INIT_51 => X"000000f500000000000000e50000000000000091000000000000005f00000000",
            INIT_52 => X"0000005e0000000000000057000000000000005c000000000000008f00000000",
            INIT_53 => X"0000005300000000000000520000000000000052000000000000005c00000000",
            INIT_54 => X"0000005800000000000000560000000000000053000000000000005400000000",
            INIT_55 => X"0000006e000000000000006a0000000000000061000000000000005a00000000",
            INIT_56 => X"0000005b000000000000005f0000000000000061000000000000006900000000",
            INIT_57 => X"0000007d000000000000008a0000000000000082000000000000006c00000000",
            INIT_58 => X"0000005600000000000000590000000000000062000000000000006e00000000",
            INIT_59 => X"000000e400000000000000db000000000000006a000000000000005300000000",
            INIT_5A => X"00000057000000000000005e0000000000000068000000000000007e00000000",
            INIT_5B => X"0000005200000000000000500000000000000057000000000000006100000000",
            INIT_5C => X"0000005900000000000000590000000000000057000000000000005400000000",
            INIT_5D => X"00000066000000000000005d000000000000005c000000000000006100000000",
            INIT_5E => X"000000650000000000000055000000000000005d000000000000006500000000",
            INIT_5F => X"000000600000000000000062000000000000007e000000000000008100000000",
            INIT_60 => X"00000058000000000000005c0000000000000061000000000000006c00000000",
            INIT_61 => X"000000c500000000000000850000000000000054000000000000005800000000",
            INIT_62 => X"0000005f000000000000005e0000000000000061000000000000006400000000",
            INIT_63 => X"0000005300000000000000600000000000000064000000000000006700000000",
            INIT_64 => X"0000005c00000000000000580000000000000050000000000000004f00000000",
            INIT_65 => X"0000005c000000000000005d000000000000005f000000000000005c00000000",
            INIT_66 => X"0000007d0000000000000066000000000000005d000000000000005a00000000",
            INIT_67 => X"0000005d000000000000003c000000000000005a000000000000006e00000000",
            INIT_68 => X"0000005b00000000000000580000000000000064000000000000007c00000000",
            INIT_69 => X"0000006b000000000000004f0000000000000059000000000000005700000000",
            INIT_6A => X"000000520000000000000047000000000000004d000000000000005900000000",
            INIT_6B => X"0000005c00000000000000660000000000000064000000000000005d00000000",
            INIT_6C => X"0000006100000000000000630000000000000063000000000000005e00000000",
            INIT_6D => X"000000530000000000000058000000000000005e000000000000005f00000000",
            INIT_6E => X"0000008300000000000000840000000000000070000000000000005b00000000",
            INIT_6F => X"0000005500000000000000400000000000000061000000000000007400000000",
            INIT_70 => X"0000005b00000000000000550000000000000066000000000000007400000000",
            INIT_71 => X"000000510000000000000058000000000000005c000000000000005a00000000",
            INIT_72 => X"0000004a00000000000000430000000000000048000000000000005500000000",
            INIT_73 => X"0000005600000000000000500000000000000049000000000000004700000000",
            INIT_74 => X"00000077000000000000006d0000000000000065000000000000005f00000000",
            INIT_75 => X"000000580000000000000058000000000000005f000000000000007100000000",
            INIT_76 => X"00000091000000000000009c0000000000000082000000000000006900000000",
            INIT_77 => X"0000004000000000000000520000000000000052000000000000007300000000",
            INIT_78 => X"0000005600000000000000590000000000000069000000000000006b00000000",
            INIT_79 => X"000000510000000000000057000000000000005c000000000000005900000000",
            INIT_7A => X"0000004900000000000000420000000000000045000000000000004f00000000",
            INIT_7B => X"0000003a000000000000003f0000000000000049000000000000004500000000",
            INIT_7C => X"0000007700000000000000680000000000000057000000000000004600000000",
            INIT_7D => X"00000057000000000000005f0000000000000060000000000000006f00000000",
            INIT_7E => X"0000008700000000000000920000000000000083000000000000006d00000000",
            INIT_7F => X"000000430000000000000054000000000000004d000000000000006300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE3;


    MEM_IFMAP_LAYER0_INSTANCE4 : if BRAM_NAME = "ifmap_layer0_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000350000000000000033000000000000002f000000000000003100000000",
            INIT_01 => X"0000002d000000000000002f0000000000000029000000000000002e00000000",
            INIT_02 => X"0000003400000000000000290000000000000029000000000000002c00000000",
            INIT_03 => X"0000002c000000000000002d0000000000000029000000000000003100000000",
            INIT_04 => X"0000002b00000000000000270000000000000026000000000000002800000000",
            INIT_05 => X"0000002b000000000000002d000000000000002d000000000000002c00000000",
            INIT_06 => X"00000029000000000000002b0000000000000027000000000000002c00000000",
            INIT_07 => X"0000002100000000000000240000000000000024000000000000002600000000",
            INIT_08 => X"00000038000000000000002d0000000000000028000000000000003300000000",
            INIT_09 => X"0000002d000000000000002f000000000000002b000000000000003100000000",
            INIT_0A => X"0000003600000000000000290000000000000026000000000000002e00000000",
            INIT_0B => X"0000002100000000000000280000000000000029000000000000003400000000",
            INIT_0C => X"0000003200000000000000290000000000000021000000000000001e00000000",
            INIT_0D => X"0000003000000000000000340000000000000037000000000000003500000000",
            INIT_0E => X"00000026000000000000002d000000000000002e000000000000003200000000",
            INIT_0F => X"000000220000000000000020000000000000001f000000000000002200000000",
            INIT_10 => X"0000003000000000000000240000000000000021000000000000002f00000000",
            INIT_11 => X"0000002d000000000000002d000000000000002c000000000000002a00000000",
            INIT_12 => X"000000390000000000000030000000000000002b000000000000002b00000000",
            INIT_13 => X"0000002300000000000000250000000000000026000000000000003300000000",
            INIT_14 => X"000000310000000000000036000000000000002f000000000000002700000000",
            INIT_15 => X"00000032000000000000002f0000000000000032000000000000003400000000",
            INIT_16 => X"0000002700000000000000330000000000000037000000000000003000000000",
            INIT_17 => X"0000002100000000000000220000000000000022000000000000002300000000",
            INIT_18 => X"0000002c000000000000001f0000000000000020000000000000002800000000",
            INIT_19 => X"000000300000000000000030000000000000002e000000000000002b00000000",
            INIT_1A => X"0000005f0000000000000039000000000000002d000000000000002c00000000",
            INIT_1B => X"00000036000000000000002f0000000000000029000000000000004b00000000",
            INIT_1C => X"00000041000000000000002f0000000000000043000000000000003a00000000",
            INIT_1D => X"0000003200000000000000420000000000000054000000000000004c00000000",
            INIT_1E => X"0000002e000000000000002d0000000000000027000000000000003400000000",
            INIT_1F => X"0000002400000000000000270000000000000027000000000000002b00000000",
            INIT_20 => X"0000002f00000000000000310000000000000030000000000000002900000000",
            INIT_21 => X"0000002c000000000000002f0000000000000028000000000000002b00000000",
            INIT_22 => X"000000a4000000000000003b000000000000002a000000000000002900000000",
            INIT_23 => X"00000047000000000000003c0000000000000038000000000000006b00000000",
            INIT_24 => X"000000620000000000000038000000000000001f000000000000003200000000",
            INIT_25 => X"0000005d00000000000000690000000000000076000000000000006f00000000",
            INIT_26 => X"0000002d000000000000002f0000000000000046000000000000004300000000",
            INIT_27 => X"000000240000000000000024000000000000002e000000000000003000000000",
            INIT_28 => X"0000003500000000000000390000000000000040000000000000003600000000",
            INIT_29 => X"0000002900000000000000290000000000000027000000000000002c00000000",
            INIT_2A => X"00000055000000000000002a0000000000000027000000000000002500000000",
            INIT_2B => X"0000001f000000000000002b000000000000003a000000000000004e00000000",
            INIT_2C => X"0000006e000000000000004c000000000000002d000000000000002b00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007800000000",
            INIT_2E => X"00000025000000000000002f0000000000000056000000000000006100000000",
            INIT_2F => X"00000028000000000000002c000000000000003a000000000000003100000000",
            INIT_30 => X"0000001c00000000000000110000000000000050000000000000003900000000",
            INIT_31 => X"0000002b0000000000000028000000000000002b000000000000003000000000",
            INIT_32 => X"0000003400000000000000270000000000000025000000000000002a00000000",
            INIT_33 => X"000000390000000000000046000000000000004b000000000000003b00000000",
            INIT_34 => X"00000079000000000000004a0000000000000040000000000000004800000000",
            INIT_35 => X"0000005e000000000000005a000000000000006c000000000000008400000000",
            INIT_36 => X"000000270000000000000045000000000000004d000000000000006700000000",
            INIT_37 => X"000000270000000000000030000000000000003a000000000000002400000000",
            INIT_38 => X"000000290000000000000026000000000000005c000000000000005a00000000",
            INIT_39 => X"000000270000000000000024000000000000002a000000000000003800000000",
            INIT_3A => X"0000003100000000000000330000000000000033000000000000003100000000",
            INIT_3B => X"0000004f000000000000005d000000000000006b000000000000004d00000000",
            INIT_3C => X"0000006b00000000000000450000000000000052000000000000005800000000",
            INIT_3D => X"0000005800000000000000510000000000000070000000000000008c00000000",
            INIT_3E => X"00000031000000000000003a000000000000004a000000000000005400000000",
            INIT_3F => X"0000002700000000000000330000000000000032000000000000002000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000071000000000000003b0000000000000069000000000000009000000000",
            INIT_41 => X"000000320000000000000029000000000000002b000000000000005200000000",
            INIT_42 => X"0000004e000000000000003b000000000000005f000000000000004200000000",
            INIT_43 => X"0000004a00000000000000650000000000000080000000000000007900000000",
            INIT_44 => X"0000003d00000000000000490000000000000052000000000000004d00000000",
            INIT_45 => X"00000046000000000000005d000000000000007b000000000000007000000000",
            INIT_46 => X"000000350000000000000043000000000000004c000000000000004500000000",
            INIT_47 => X"0000002d000000000000003b0000000000000023000000000000001b00000000",
            INIT_48 => X"000000950000000000000069000000000000008f00000000000000a300000000",
            INIT_49 => X"0000003c000000000000002f0000000000000033000000000000007000000000",
            INIT_4A => X"0000007700000000000000a600000000000000c6000000000000009200000000",
            INIT_4B => X"0000004f000000000000006b000000000000007d000000000000009100000000",
            INIT_4C => X"0000003a00000000000000350000000000000047000000000000004f00000000",
            INIT_4D => X"000000590000000000000072000000000000007a000000000000007000000000",
            INIT_4E => X"00000047000000000000004e000000000000004e000000000000004a00000000",
            INIT_4F => X"00000039000000000000002c000000000000000f000000000000002b00000000",
            INIT_50 => X"000000a8000000000000009e000000000000007a00000000000000af00000000",
            INIT_51 => X"0000002f00000000000000330000000000000032000000000000007a00000000",
            INIT_52 => X"0000008300000000000000bc00000000000000e200000000000000b300000000",
            INIT_53 => X"0000006800000000000000680000000000000084000000000000009b00000000",
            INIT_54 => X"0000004d0000000000000028000000000000004d000000000000004500000000",
            INIT_55 => X"0000005c000000000000008a0000000000000089000000000000009a00000000",
            INIT_56 => X"00000049000000000000004f0000000000000060000000000000004d00000000",
            INIT_57 => X"0000002e000000000000001f0000000000000021000000000000003b00000000",
            INIT_58 => X"000000b20000000000000099000000000000007400000000000000bd00000000",
            INIT_59 => X"0000002c0000000000000037000000000000003b000000000000008800000000",
            INIT_5A => X"0000008500000000000000a400000000000000bc000000000000005000000000",
            INIT_5B => X"0000005f000000000000006a000000000000009f000000000000009700000000",
            INIT_5C => X"000000710000000000000022000000000000004f000000000000005900000000",
            INIT_5D => X"000000520000000000000082000000000000008e00000000000000c000000000",
            INIT_5E => X"00000051000000000000005e0000000000000058000000000000004b00000000",
            INIT_5F => X"0000001a00000000000000300000000000000037000000000000004e00000000",
            INIT_60 => X"000000b90000000000000090000000000000006900000000000000c200000000",
            INIT_61 => X"0000002f00000000000000350000000000000044000000000000008500000000",
            INIT_62 => X"0000005e000000000000007e0000000000000098000000000000002c00000000",
            INIT_63 => X"00000062000000000000008100000000000000b7000000000000009400000000",
            INIT_64 => X"0000008c000000000000002f000000000000006d000000000000006900000000",
            INIT_65 => X"00000053000000000000006f000000000000008c00000000000000b200000000",
            INIT_66 => X"0000005100000000000000550000000000000050000000000000004f00000000",
            INIT_67 => X"0000001800000000000000400000000000000049000000000000005900000000",
            INIT_68 => X"000000c000000000000000a3000000000000006700000000000000c100000000",
            INIT_69 => X"00000032000000000000003a0000000000000042000000000000006200000000",
            INIT_6A => X"0000007f00000000000000670000000000000078000000000000002700000000",
            INIT_6B => X"00000075000000000000009d00000000000000c8000000000000009b00000000",
            INIT_6C => X"000000930000000000000044000000000000006d000000000000006b00000000",
            INIT_6D => X"000000500000000000000068000000000000008800000000000000ae00000000",
            INIT_6E => X"0000005e00000000000000480000000000000046000000000000004c00000000",
            INIT_6F => X"0000002200000000000000450000000000000051000000000000006300000000",
            INIT_70 => X"000000bc00000000000000ac000000000000007000000000000000c400000000",
            INIT_71 => X"00000037000000000000003e0000000000000043000000000000006d00000000",
            INIT_72 => X"000000a900000000000000670000000000000058000000000000002200000000",
            INIT_73 => X"00000086000000000000008c000000000000009f00000000000000a900000000",
            INIT_74 => X"000000950000000000000046000000000000005f000000000000007d00000000",
            INIT_75 => X"00000069000000000000007a000000000000007f00000000000000aa00000000",
            INIT_76 => X"00000068000000000000005a000000000000005b000000000000005300000000",
            INIT_77 => X"0000002f00000000000000350000000000000050000000000000006f00000000",
            INIT_78 => X"000000b500000000000000ae000000000000008800000000000000c500000000",
            INIT_79 => X"0000004d0000000000000058000000000000004d000000000000008e00000000",
            INIT_7A => X"000000d30000000000000074000000000000005d000000000000003400000000",
            INIT_7B => X"000000700000000000000082000000000000008900000000000000e600000000",
            INIT_7C => X"00000076000000000000004b000000000000005f000000000000006500000000",
            INIT_7D => X"000000500000000000000065000000000000008a000000000000009200000000",
            INIT_7E => X"0000006300000000000000630000000000000057000000000000004400000000",
            INIT_7F => X"0000003000000000000000300000000000000036000000000000005d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE4;


    MEM_IFMAP_LAYER0_INSTANCE5 : if BRAM_NAME = "ifmap_layer0_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bc00000000000000b200000000000000a000000000000000cc00000000",
            INIT_01 => X"00000071000000000000007e000000000000005a00000000000000ac00000000",
            INIT_02 => X"0000009b00000000000000850000000000000025000000000000005200000000",
            INIT_03 => X"0000005a00000000000000580000000000000075000000000000008d00000000",
            INIT_04 => X"00000068000000000000003a0000000000000057000000000000005c00000000",
            INIT_05 => X"000000610000000000000076000000000000007e000000000000006d00000000",
            INIT_06 => X"00000052000000000000005e000000000000004d000000000000004800000000",
            INIT_07 => X"0000002e0000000000000037000000000000002d000000000000003700000000",
            INIT_08 => X"000000c200000000000000b800000000000000b400000000000000d700000000",
            INIT_09 => X"000000910000000000000066000000000000006900000000000000ba00000000",
            INIT_0A => X"0000005f0000000000000069000000000000003d000000000000006f00000000",
            INIT_0B => X"0000006200000000000000490000000000000059000000000000005900000000",
            INIT_0C => X"000000400000000000000066000000000000005f000000000000005800000000",
            INIT_0D => X"0000003d00000000000000730000000000000069000000000000002000000000",
            INIT_0E => X"0000004e00000000000000410000000000000035000000000000003300000000",
            INIT_0F => X"0000003600000000000000400000000000000044000000000000004000000000",
            INIT_10 => X"000000c100000000000000bd00000000000000c000000000000000cd00000000",
            INIT_11 => X"0000008f0000000000000060000000000000008500000000000000bc00000000",
            INIT_12 => X"000000370000000000000050000000000000006f000000000000008d00000000",
            INIT_13 => X"0000008500000000000000640000000000000060000000000000006c00000000",
            INIT_14 => X"0000005d0000000000000078000000000000005d000000000000005d00000000",
            INIT_15 => X"00000034000000000000003a0000000000000056000000000000005c00000000",
            INIT_16 => X"0000003b0000000000000028000000000000003c000000000000002700000000",
            INIT_17 => X"0000002e000000000000002d0000000000000036000000000000003e00000000",
            INIT_18 => X"000000b900000000000000b500000000000000bb00000000000000b400000000",
            INIT_19 => X"000000840000000000000063000000000000009800000000000000b800000000",
            INIT_1A => X"00000033000000000000007e0000000000000087000000000000008200000000",
            INIT_1B => X"000000a8000000000000007b0000000000000056000000000000006c00000000",
            INIT_1C => X"0000006900000000000000670000000000000049000000000000007600000000",
            INIT_1D => X"00000032000000000000002c000000000000004e000000000000007600000000",
            INIT_1E => X"00000044000000000000003c000000000000005d000000000000003400000000",
            INIT_1F => X"0000002e00000000000000320000000000000034000000000000004000000000",
            INIT_20 => X"000000ac00000000000000af00000000000000bb000000000000009200000000",
            INIT_21 => X"00000092000000000000006f00000000000000a000000000000000b400000000",
            INIT_22 => X"000000490000000000000057000000000000006f00000000000000b900000000",
            INIT_23 => X"000000b100000000000000ad0000000000000074000000000000005600000000",
            INIT_24 => X"0000003f00000000000000420000000000000065000000000000009400000000",
            INIT_25 => X"0000002900000000000000330000000000000036000000000000003900000000",
            INIT_26 => X"00000052000000000000004b0000000000000053000000000000004500000000",
            INIT_27 => X"0000003f0000000000000045000000000000003d000000000000004c00000000",
            INIT_28 => X"000000a800000000000000b000000000000000c8000000000000007c00000000",
            INIT_29 => X"0000009f000000000000005b000000000000009300000000000000b300000000",
            INIT_2A => X"00000093000000000000009000000000000000e100000000000000fa00000000",
            INIT_2B => X"000000c500000000000000d000000000000000c000000000000000a400000000",
            INIT_2C => X"0000003e000000000000006d000000000000008f00000000000000b500000000",
            INIT_2D => X"0000006600000000000000570000000000000044000000000000003a00000000",
            INIT_2E => X"00000077000000000000007a000000000000006f000000000000006e00000000",
            INIT_2F => X"0000007300000000000000700000000000000070000000000000007800000000",
            INIT_30 => X"000000b100000000000000c000000000000000d5000000000000008500000000",
            INIT_31 => X"000000d10000000000000071000000000000009600000000000000b600000000",
            INIT_32 => X"0000009d00000000000000e800000000000000fc00000000000000f700000000",
            INIT_33 => X"00000098000000000000009c00000000000000a2000000000000009500000000",
            INIT_34 => X"0000006500000000000000680000000000000077000000000000009400000000",
            INIT_35 => X"0000007d0000000000000073000000000000006e000000000000006f00000000",
            INIT_36 => X"0000008d00000000000000870000000000000082000000000000008300000000",
            INIT_37 => X"0000008400000000000000890000000000000084000000000000008e00000000",
            INIT_38 => X"000000bc00000000000000bc00000000000000a8000000000000008700000000",
            INIT_39 => X"000000ed00000000000000a400000000000000ae00000000000000c000000000",
            INIT_3A => X"0000006f000000000000009900000000000000e400000000000000f100000000",
            INIT_3B => X"00000065000000000000006b0000000000000069000000000000006900000000",
            INIT_3C => X"0000007400000000000000710000000000000078000000000000007300000000",
            INIT_3D => X"00000080000000000000007e000000000000007d000000000000007d00000000",
            INIT_3E => X"000000890000000000000089000000000000008b000000000000008400000000",
            INIT_3F => X"00000085000000000000008b0000000000000086000000000000008700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b000000000000000860000000000000082000000000000008d00000000",
            INIT_41 => X"000000f200000000000000b5000000000000008900000000000000bf00000000",
            INIT_42 => X"00000076000000000000007f00000000000000af00000000000000f500000000",
            INIT_43 => X"0000007400000000000000780000000000000079000000000000007700000000",
            INIT_44 => X"0000007100000000000000730000000000000075000000000000007500000000",
            INIT_45 => X"00000082000000000000007d000000000000007d000000000000007800000000",
            INIT_46 => X"0000008e000000000000008e0000000000000091000000000000008600000000",
            INIT_47 => X"00000095000000000000008c0000000000000090000000000000009200000000",
            INIT_48 => X"00000088000000000000007c000000000000008c00000000000000a200000000",
            INIT_49 => X"000000f900000000000000d1000000000000008f00000000000000a700000000",
            INIT_4A => X"0000007d0000000000000080000000000000007600000000000000cd00000000",
            INIT_4B => X"000000730000000000000079000000000000007f000000000000007f00000000",
            INIT_4C => X"0000007500000000000000710000000000000070000000000000007100000000",
            INIT_4D => X"0000008a00000000000000860000000000000083000000000000007b00000000",
            INIT_4E => X"0000009500000000000000930000000000000098000000000000009600000000",
            INIT_4F => X"000000b600000000000000a70000000000000098000000000000009a00000000",
            INIT_50 => X"0000007a0000000000000082000000000000009300000000000000a500000000",
            INIT_51 => X"000000f700000000000000ea00000000000000a4000000000000007e00000000",
            INIT_52 => X"00000083000000000000007b0000000000000072000000000000009900000000",
            INIT_53 => X"0000007700000000000000770000000000000077000000000000008100000000",
            INIT_54 => X"0000007f000000000000007b0000000000000077000000000000007700000000",
            INIT_55 => X"0000009a0000000000000096000000000000008d000000000000008300000000",
            INIT_56 => X"0000008a000000000000008c000000000000008d000000000000009600000000",
            INIT_57 => X"000000a900000000000000b600000000000000b2000000000000009e00000000",
            INIT_58 => X"00000085000000000000008a000000000000009500000000000000a200000000",
            INIT_59 => X"000000ea00000000000000e9000000000000008a000000000000007e00000000",
            INIT_5A => X"0000007c0000000000000081000000000000007e000000000000008c00000000",
            INIT_5B => X"000000770000000000000074000000000000007b000000000000008500000000",
            INIT_5C => X"000000840000000000000082000000000000007e000000000000007a00000000",
            INIT_5D => X"00000094000000000000008b000000000000008a000000000000008c00000000",
            INIT_5E => X"000000990000000000000085000000000000008b000000000000009300000000",
            INIT_5F => X"0000008b000000000000008e00000000000000b000000000000000b600000000",
            INIT_60 => X"0000008d000000000000008f000000000000009300000000000000a100000000",
            INIT_61 => X"000000d3000000000000009f000000000000007d000000000000008a00000000",
            INIT_62 => X"0000008200000000000000800000000000000079000000000000007700000000",
            INIT_63 => X"0000007800000000000000830000000000000087000000000000008b00000000",
            INIT_64 => X"0000008700000000000000820000000000000078000000000000007600000000",
            INIT_65 => X"00000088000000000000008a000000000000008b000000000000008800000000",
            INIT_66 => X"000000b20000000000000097000000000000008a000000000000008700000000",
            INIT_67 => X"000000880000000000000067000000000000008c00000000000000a400000000",
            INIT_68 => X"000000920000000000000089000000000000009400000000000000b100000000",
            INIT_69 => X"0000008500000000000000710000000000000084000000000000008b00000000",
            INIT_6A => X"0000007500000000000000690000000000000069000000000000007200000000",
            INIT_6B => X"0000008000000000000000890000000000000087000000000000008000000000",
            INIT_6C => X"0000008a000000000000008b0000000000000089000000000000008300000000",
            INIT_6D => X"0000007d00000000000000830000000000000088000000000000008900000000",
            INIT_6E => X"000000b500000000000000b3000000000000009a000000000000008500000000",
            INIT_6F => X"0000007f000000000000006c000000000000009200000000000000a800000000",
            INIT_70 => X"0000008f0000000000000084000000000000009400000000000000a800000000",
            INIT_71 => X"00000070000000000000007d0000000000000086000000000000008b00000000",
            INIT_72 => X"0000006d00000000000000660000000000000068000000000000007300000000",
            INIT_73 => X"000000780000000000000073000000000000006c000000000000006a00000000",
            INIT_74 => X"0000009c00000000000000900000000000000087000000000000008000000000",
            INIT_75 => X"0000007f000000000000007f0000000000000086000000000000009800000000",
            INIT_76 => X"000000be00000000000000c500000000000000aa000000000000009000000000",
            INIT_77 => X"0000006b000000000000007e000000000000008200000000000000a400000000",
            INIT_78 => X"000000860000000000000084000000000000009500000000000000a000000000",
            INIT_79 => X"00000073000000000000007b0000000000000084000000000000008600000000",
            INIT_7A => X"0000006c00000000000000650000000000000069000000000000007200000000",
            INIT_7B => X"000000590000000000000062000000000000006c000000000000006800000000",
            INIT_7C => X"0000009800000000000000890000000000000076000000000000006400000000",
            INIT_7D => X"0000007b00000000000000820000000000000083000000000000009100000000",
            INIT_7E => X"000000af00000000000000b600000000000000a7000000000000009100000000",
            INIT_7F => X"0000006e0000000000000081000000000000007c000000000000009100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE5;


    MEM_IFMAP_LAYER1_INSTANCE0 : if BRAM_NAME = "ifmap_layer1_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000021000000000000001f000000000000002f000000000000001800000000",
            INIT_01 => X"0000002c00000000000000240000000000000028000000000000001900000000",
            INIT_02 => X"0000001900000000000000080000000000000000000000000000001b00000000",
            INIT_03 => X"0000001c0000000000000027000000000000002a000000000000002800000000",
            INIT_04 => X"000000190000000000000021000000000000001d000000000000003b00000000",
            INIT_05 => X"0000001300000000000000100000000000000013000000000000001b00000000",
            INIT_06 => X"0000000b00000000000000080000000000000000000000000000000f00000000",
            INIT_07 => X"000000000000000000000000000000000000001b000000000000001000000000",
            INIT_08 => X"000000220000000000000014000000000000002b000000000000002100000000",
            INIT_09 => X"000000000000000000000009000000000000002c000000000000003400000000",
            INIT_0A => X"0000000000000000000000030000000000000012000000000000000700000000",
            INIT_0B => X"0000001b00000000000000000000000000000030000000000000002000000000",
            INIT_0C => X"0000000c000000000000000f0000000000000012000000000000001d00000000",
            INIT_0D => X"0000003200000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000100000000000000030000000000000000e00000000",
            INIT_0F => X"0000000000000000000000120000000000000000000000000000002000000000",
            INIT_10 => X"0000002a00000000000000370000000000000000000000000000000000000000",
            INIT_11 => X"0000001c000000000000001b0000000000000000000000000000001d00000000",
            INIT_12 => X"0000000000000000000000000000000000000021000000000000000e00000000",
            INIT_13 => X"0000002f000000000000000f0000000000000032000000000000000000000000",
            INIT_14 => X"00000034000000000000002b0000000000000041000000000000003000000000",
            INIT_15 => X"0000000000000000000000350000000000000005000000000000000000000000",
            INIT_16 => X"00000002000000000000000b0000000000000015000000000000001200000000",
            INIT_17 => X"000000000000000000000000000000000000005c000000000000001900000000",
            INIT_18 => X"0000000000000000000000380000000000000019000000000000000000000000",
            INIT_19 => X"0000000400000000000000080000000000000025000000000000002f00000000",
            INIT_1A => X"0000000000000000000000320000000000000000000000000000000f00000000",
            INIT_1B => X"0000001900000000000000000000000000000000000000000000002000000000",
            INIT_1C => X"000000260000000000000000000000000000003b000000000000001400000000",
            INIT_1D => X"0000003d00000000000000040000000000000000000000000000003700000000",
            INIT_1E => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_1F => X"0000000f00000000000000420000000000000028000000000000000000000000",
            INIT_20 => X"0000004200000000000000110000000000000019000000000000000000000000",
            INIT_21 => X"0000000c00000000000000020000000000000027000000000000001900000000",
            INIT_22 => X"0000000c0000000000000000000000000000003b000000000000000000000000",
            INIT_23 => X"0000000000000000000000190000000000000006000000000000000000000000",
            INIT_24 => X"00000000000000000000001e0000000000000023000000000000000300000000",
            INIT_25 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_26 => X"0000000000000000000000020000000000000000000000000000004000000000",
            INIT_27 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"00000008000000000000002b0000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_3F => X"0000001e00000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000100000000000000000000000000000000000000000000001300000000",
            INIT_41 => X"00000000000000000000000a000000000000000e00000000000000b700000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000022000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000023000000000000000000000000",
            INIT_4A => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000008700000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"000000000000000000000000000000000000001500000000000000a700000000",
            INIT_4D => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000004e00000000000000000000000000000000000000000000000b00000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"000000480000000000000000000000000000005a000000000000005f00000000",
            INIT_55 => X"0000002300000000000000000000000000000002000000000000000300000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_57 => X"0000000000000000000000990000000000000000000000000000000000000000",
            INIT_58 => X"0000003e00000000000000240000000000000000000000000000000000000000",
            INIT_59 => X"000000000000000000000000000000000000003a000000000000006d00000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"000000000000000000000047000000000000003f000000000000000c00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000860000000000000000000000000000000000000000",
            INIT_62 => X"0000007500000000000000bf0000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000050000000000000006300000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000740000000000000000000000000000000000000000",
            INIT_66 => X"000000000000000000000000000000000000005c000000000000002e00000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000005f00000000000000590000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000590000000000000000000000000000000000000000",
            INIT_6D => X"0000001a000000000000006e000000000000000d000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000013000000000000002100000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"00000020000000000000002e0000000000000000000000000000000000000000",
            INIT_71 => X"0000002700000000000000250000000000000023000000000000003600000000",
            INIT_72 => X"0000000d0000000000000025000000000000002d000000000000002800000000",
            INIT_73 => X"0000001700000000000000240000000000000028000000000000001100000000",
            INIT_74 => X"0000003a00000000000000240000000000000028000000000000001300000000",
            INIT_75 => X"0000000000000000000000000000000000000042000000000000001c00000000",
            INIT_76 => X"0000000000000000000000150000000000000001000000000000000000000000",
            INIT_77 => X"0000000c0000000000000025000000000000000d000000000000000000000000",
            INIT_78 => X"00000022000000000000002b0000000000000063000000000000000000000000",
            INIT_79 => X"000000000000000000000000000000000000000b000000000000003b00000000",
            INIT_7A => X"000000000000000000000000000000000000003d000000000000002100000000",
            INIT_7B => X"00000000000000000000001b0000000000000021000000000000000000000000",
            INIT_7C => X"0000000000000000000000360000000000000004000000000000006200000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000004800000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000009700000000",
            INIT_7F => X"000000000000000000000000000000000000006f000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE0;


    MEM_IFMAP_LAYER1_INSTANCE1 : if BRAM_NAME = "ifmap_layer1_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001e000000000000000000000000000000f0000000000000000000000000",
            INIT_01 => X"000000e800000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000005100000000",
            INIT_04 => X"0000000000000000000000540000000000000044000000000000007000000000",
            INIT_05 => X"00000000000000000000012e0000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_07 => X"0000000000000000000000060000000000000000000000000000002b00000000",
            INIT_08 => X"0000000000000000000000000000000000000063000000000000005b00000000",
            INIT_09 => X"00000000000000000000000000000000000000bd000000000000000000000000",
            INIT_0A => X"0000001100000000000000000000000000000002000000000000000000000000",
            INIT_0B => X"0000008000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_0D => X"0000002800000000000000000000000000000000000000000000008700000000",
            INIT_0E => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_0F => X"0000003800000000000000070000000000000000000000000000000000000000",
            INIT_10 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_11 => X"0000001e000000000000002f0000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_13 => X"0000006d000000000000006a0000000000000000000000000000003d00000000",
            INIT_14 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_15 => X"00000004000000000000002d000000000000001a000000000000000000000000",
            INIT_16 => X"000000fb00000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"00000000000000000000003f0000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000002000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"00000000000000000000005d0000000000000000000000000000002a00000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000003f00000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"000000000000000000000000000000000000000000000000000000d800000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"000000fa00000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000100000000000000000000000000000000000000000000000700000000",
            INIT_29 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000700000000000000040000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000060000000000000001000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000003700000000000000000000000000000000000000000000000500000000",
            INIT_2F => X"0000000000000000000000560000000000000053000000000000001c00000000",
            INIT_30 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000003500000000000000500000000000000005000000000000000500000000",
            INIT_32 => X"000000000000000000000000000000000000002500000000000000a700000000",
            INIT_33 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_34 => X"00000008000000000000000c0000000000000052000000000000000f00000000",
            INIT_35 => X"000000000000000000000000000000000000003e000000000000000300000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000120000000000000000000000000000000800000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000023000000000000004100000000",
            INIT_3B => X"000000000000000000000000000000000000002a000000000000000000000000",
            INIT_3C => X"00000000000000000000004b0000000000000001000000000000000000000000",
            INIT_3D => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_3F => X"0000003900000000000000000000000000000015000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_41 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000020000000000000032000000000000002300000000",
            INIT_43 => X"0000001000000000000000190000000000000006000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000004a00000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"00000000000000000000001d0000000000000071000000000000006300000000",
            INIT_49 => X"000000310000000000000003000000000000003b000000000000008200000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_4B => X"0000000000000000000000000000000000000055000000000000000000000000",
            INIT_4C => X"0000000000000000000000170000000000000000000000000000003400000000",
            INIT_4D => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_4E => X"0000001f00000000000000050000000000000009000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_50 => X"00000034000000000000001d0000000000000000000000000000000000000000",
            INIT_51 => X"0000003300000000000000320000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_53 => X"000000aa00000000000000b1000000000000009c000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000003600000000",
            INIT_55 => X"0000000000000000000000000000000000000009000000000000000700000000",
            INIT_56 => X"0000006200000000000000000000000000000017000000000000002e00000000",
            INIT_57 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_5A => X"0000000200000000000000000000000000000000000000000000000b00000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_5D => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"000000000000000000000007000000000000001e000000000000009c00000000",
            INIT_5F => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000330000000000000023000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"000000a000000000000000060000000000000011000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"00000000000000000000004a0000000000000000000000000000000000000000",
            INIT_69 => X"0000007800000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"000000000000000000000000000000000000000a000000000000000900000000",
            INIT_6B => X"0000000000000000000000500000000000000000000000000000000c00000000",
            INIT_6C => X"0000000000000000000000000000000000000080000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000001900000000000000000000000000000002000000000000001400000000",
            INIT_6F => X"000000000000000000000000000000000000000d000000000000002600000000",
            INIT_70 => X"00000000000000000000001d0000000000000000000000000000004f00000000",
            INIT_71 => X"0000000000000000000000320000000000000015000000000000000000000000",
            INIT_72 => X"0000003400000000000000000000000000000000000000000000002a00000000",
            INIT_73 => X"0000004300000000000000000000000000000019000000000000000000000000",
            INIT_74 => X"0000000000000000000000190000000000000000000000000000000000000000",
            INIT_75 => X"0000002c000000000000000a0000000000000000000000000000000000000000",
            INIT_76 => X"00000000000000000000003d0000000000000062000000000000000000000000",
            INIT_77 => X"0000004b00000000000000000000000000000000000000000000000f00000000",
            INIT_78 => X"0000000000000000000000000000000000000039000000000000000000000000",
            INIT_79 => X"0000000000000000000000680000000000000000000000000000005e00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000005200000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"000000bd00000000000000000000000000000009000000000000000000000000",
            INIT_7D => X"0000000b00000000000000000000000000000000000000000000002e00000000",
            INIT_7E => X"0000000000000000000000120000000000000000000000000000000d00000000",
            INIT_7F => X"0000000000000000000000230000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE1;


    MEM_IFMAP_LAYER1_INSTANCE2 : if BRAM_NAME = "ifmap_layer1_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000056000000000000000000000000",
            INIT_01 => X"0000008100000000000000000000000000000064000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000002900000000000000000000000000000044000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"00000000000000000000001400000000000000bd000000000000004500000000",
            INIT_06 => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000007000000000",
            INIT_08 => X"00000038000000000000008b0000000000000088000000000000000e00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000100000000000000000000000000000035000000000000000f00000000",
            INIT_0B => X"0000000000000000000000200000000000000178000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000005900000000000000000000000000000000000000000000001700000000",
            INIT_0F => X"0000000000000000000000120000000000000000000000000000009c00000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000f00000000000000000000000000000012000000000000001900000000",
            INIT_12 => X"0000000f00000000000000c70000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000020000000000000003000000000000000000000000",
            INIT_15 => X"00000000000000000000002a0000000000000098000000000000000000000000",
            INIT_16 => X"00000000000000000000002b0000000000000055000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_18 => X"0000000a00000000000000000000000000000000000000000000000900000000",
            INIT_19 => X"0000004f00000000000000560000000000000042000000000000005200000000",
            INIT_1A => X"0000005400000000000000450000000000000058000000000000005800000000",
            INIT_1B => X"0000003e0000000000000047000000000000005f000000000000005c00000000",
            INIT_1C => X"0000005a00000000000000510000000000000049000000000000003700000000",
            INIT_1D => X"0000005e00000000000000450000000000000050000000000000005700000000",
            INIT_1E => X"0000006800000000000000640000000000000097000000000000003c00000000",
            INIT_1F => X"000000320000000000000045000000000000001e000000000000004000000000",
            INIT_20 => X"0000007e00000000000000570000000000000023000000000000001400000000",
            INIT_21 => X"0000004800000000000000610000000000000056000000000000000000000000",
            INIT_22 => X"000000000000000000000017000000000000008d000000000000000000000000",
            INIT_23 => X"00000053000000000000001c000000000000001d000000000000000000000000",
            INIT_24 => X"0000000000000000000000b50000000000000031000000000000000000000000",
            INIT_25 => X"0000000500000000000000960000000000000047000000000000004b00000000",
            INIT_26 => X"0000000000000000000000280000000000000027000000000000004e00000000",
            INIT_27 => X"00000045000000000000004d0000000000000000000000000000008500000000",
            INIT_28 => X"0000007000000000000000000000000000000066000000000000000000000000",
            INIT_29 => X"0000005f000000000000000a0000000000000069000000000000000000000000",
            INIT_2A => X"0000001600000000000000000000000000000047000000000000006b00000000",
            INIT_2B => X"000000000000000000000063000000000000001e000000000000006400000000",
            INIT_2C => X"00000043000000000000008c000000000000000c000000000000000000000000",
            INIT_2D => X"0000003200000000000000a50000000000000000000000000000000000000000",
            INIT_2E => X"00000065000000000000006a000000000000000000000000000000a600000000",
            INIT_2F => X"00000000000000000000003d000000000000002e000000000000000000000000",
            INIT_30 => X"0000000000000000000000b80000000000000016000000000000007900000000",
            INIT_31 => X"000000720000000000000064000000000000001f000000000000000000000000",
            INIT_32 => X"000000010000000000000056000000000000006d000000000000000000000000",
            INIT_33 => X"000000400000000000000017000000000000003b000000000000000000000000",
            INIT_34 => X"000000000000000000000000000000000000006e000000000000000000000000",
            INIT_35 => X"0000000000000000000000530000000000000010000000000000008300000000",
            INIT_36 => X"0000000000000000000000000000000000000058000000000000006300000000",
            INIT_37 => X"000000a10000000000000000000000000000003b000000000000003200000000",
            INIT_38 => X"0000002700000000000000000000000000000049000000000000000000000000",
            INIT_39 => X"0000000000000000000000430000000000000000000000000000004d00000000",
            INIT_3A => X"0000003000000000000000030000000000000000000000000000006700000000",
            INIT_3B => X"0000000000000000000000c40000000000000000000000000000001a00000000",
            INIT_3C => X"0000005200000000000000000000000000000000000000000000002400000000",
            INIT_3D => X"000000000000000000000065000000000000001a000000000000000300000000",
            INIT_3E => X"00000000000000000000004f000000000000000d000000000000000000000000",
            INIT_3F => X"000000f800000000000000000000000000000098000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006e00000000000000090000000000000000000000000000001000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_42 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_43 => X"0000002500000000000000850000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"000000000000000000000000000000000000006d000000000000003e00000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"000000b800000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000040000000000000033000000000000003d00000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"000000000000000000000000000000000000005f000000000000000000000000",
            INIT_58 => X"0000000000000000000000340000000000000000000000000000000000000000",
            INIT_59 => X"00000000000000000000000000000000000000a8000000000000001000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"00000000000000000000001d0000000000000017000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000005b00000000",
            INIT_60 => X"000000000000000000000000000000000000004c000000000000000000000000",
            INIT_61 => X"000000000000000000000000000000000000004d000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"000000000000000000000054000000000000005a000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_68 => X"00000000000000000000004a0000000000000000000000000000000000000000",
            INIT_69 => X"00000000000000000000002d0000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"000000070000000000000016000000000000002b000000000000008000000000",
            INIT_6E => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_70 => X"0000002600000000000000000000000000000022000000000000000000000000",
            INIT_71 => X"0000000000000000000000280000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000029000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"000000000000000000000010000000000000001b000000000000000000000000",
            INIT_75 => X"0000005500000000000000a10000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000030000000000000002600000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_78 => X"000000b5000000000000006b0000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000008b00000000",
            INIT_7A => X"0000008500000000000000130000000000000017000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000043000000000000008700000000",
            INIT_7C => X"0000000300000000000000000000000000000000000000000000001e00000000",
            INIT_7D => X"0000000000000000000000000000000000000001000000000000000300000000",
            INIT_7E => X"0000003500000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000330000000000000000000000000000006500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE2;


    MEM_IFMAP_LAYER1_INSTANCE3 : if BRAM_NAME = "ifmap_layer1_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000001a00000000000000040000000000000000000000000000000000000000",
            INIT_02 => X"0000007200000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"000000000000000000000000000000000000001d000000000000004f00000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"000000170000000000000048000000000000000b000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000002300000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000024000000000000001400000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000003100000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"00000000000000000000001e0000000000000000000000000000001600000000",
            INIT_18 => X"0000003c0000000000000000000000000000000f000000000000001a00000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_1A => X"000000230000000000000017000000000000000d000000000000000000000000",
            INIT_1B => X"0000001000000000000000130000000000000005000000000000000000000000",
            INIT_1C => X"0000002c00000000000000180000000000000000000000000000002700000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"00000000000000000000004d0000000000000000000000000000002f00000000",
            INIT_1F => X"000000190000000000000000000000000000000e000000000000001900000000",
            INIT_20 => X"00000000000000000000007a0000000000000007000000000000001400000000",
            INIT_21 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"000000260000000000000000000000000000002e000000000000000d00000000",
            INIT_23 => X"0000000600000000000000100000000000000011000000000000002300000000",
            INIT_24 => X"0000000000000000000000000000000000000058000000000000002200000000",
            INIT_25 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_26 => X"0000002500000000000000200000000000000000000000000000000000000000",
            INIT_27 => X"0000005400000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"00000000000000000000000d0000000000000053000000000000004400000000",
            INIT_29 => X"0000000000000000000000270000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_2B => X"0000003800000000000000380000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000100000000000000029000000000000007900000000",
            INIT_2D => X"0000000000000000000000010000000000000049000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000004000000000000001300000000",
            INIT_2F => X"0000006700000000000000240000000000000044000000000000000000000000",
            INIT_30 => X"00000031000000000000004000000000000000a6000000000000000000000000",
            INIT_31 => X"000000560000000000000041000000000000004b000000000000003d00000000",
            INIT_32 => X"0000005000000000000000500000000000000079000000000000007300000000",
            INIT_33 => X"0000002600000000000000200000000000000043000000000000006a00000000",
            INIT_34 => X"0000007f00000000000000840000000000000081000000000000008d00000000",
            INIT_35 => X"000000ba00000000000000b10000000000000098000000000000009b00000000",
            INIT_36 => X"000000f900000000000000cc00000000000000cc00000000000000cc00000000",
            INIT_37 => X"0000007e00000000000000780000000000000000000000000000006900000000",
            INIT_38 => X"000000af00000000000000a800000000000000af00000000000000ae00000000",
            INIT_39 => X"000000cf00000000000000d300000000000000cd00000000000000ba00000000",
            INIT_3A => X"000000db000000000000010400000000000000e100000000000000ca00000000",
            INIT_3B => X"000000ac000000000000009600000000000000bf000000000000002200000000",
            INIT_3C => X"000000c200000000000000b000000000000000ae00000000000000bf00000000",
            INIT_3D => X"000000f200000000000000e700000000000000db00000000000000da00000000",
            INIT_3E => X"000000cd00000000000000f1000000000000010200000000000000fc00000000",
            INIT_3F => X"000000a600000000000000a600000000000000a6000000000000009100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d600000000000000d200000000000000b600000000000000ab00000000",
            INIT_41 => X"00000103000000000000011300000000000000cd00000000000000c800000000",
            INIT_42 => X"000000e200000000000000e100000000000000e300000000000000d500000000",
            INIT_43 => X"000000fd00000000000000eb00000000000000d500000000000000e100000000",
            INIT_44 => X"00000095000000000000008800000000000000a900000000000000e100000000",
            INIT_45 => X"000000dd00000000000000c400000000000000c700000000000000ae00000000",
            INIT_46 => X"000000df00000000000000ea00000000000000ee00000000000000f200000000",
            INIT_47 => X"0000008100000000000000b500000000000000c000000000000000e800000000",
            INIT_48 => X"0000004c00000000000000300000000000000027000000000000003d00000000",
            INIT_49 => X"00000090000000000000008400000000000000b4000000000000008400000000",
            INIT_4A => X"000000d600000000000000f300000000000000f200000000000000ea00000000",
            INIT_4B => X"0000003b00000000000000170000000000000033000000000000006f00000000",
            INIT_4C => X"0000002f000000000000002c0000000000000010000000000000001c00000000",
            INIT_4D => X"000000ce0000000000000066000000000000002f000000000000009600000000",
            INIT_4E => X"0000005a000000000000006e00000000000000c100000000000000e600000000",
            INIT_4F => X"0000003a000000000000002a000000000000001c000000000000001c00000000",
            INIT_50 => X"0000006800000000000000190000000000000012000000000000002f00000000",
            INIT_51 => X"0000007f00000000000000a7000000000000005d000000000000000000000000",
            INIT_52 => X"0000002200000000000000400000000000000067000000000000006e00000000",
            INIT_53 => X"0000002700000000000000370000000000000025000000000000002200000000",
            INIT_54 => X"00000000000000000000003a0000000000000018000000000000002200000000",
            INIT_55 => X"0000005100000000000000d40000000000000093000000000000002b00000000",
            INIT_56 => X"00000032000000000000002f000000000000005d000000000000003500000000",
            INIT_57 => X"000000160000000000000004000000000000002c000000000000003d00000000",
            INIT_58 => X"0000004c00000000000000000000000000000016000000000000000f00000000",
            INIT_59 => X"00000054000000000000008e00000000000000b7000000000000004800000000",
            INIT_5A => X"000000550000000000000019000000000000002d000000000000003d00000000",
            INIT_5B => X"00000015000000000000001b0000000000000010000000000000000f00000000",
            INIT_5C => X"00000008000000000000000e0000000000000000000000000000002800000000",
            INIT_5D => X"000000220000000000000042000000000000006b000000000000005900000000",
            INIT_5E => X"000000320000000000000082000000000000001d000000000000002a00000000",
            INIT_5F => X"000000680000000000000034000000000000000d000000000000001500000000",
            INIT_60 => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"00000037000000000000002d0000000000000033000000000000003f00000000",
            INIT_62 => X"0000000e00000000000000260000000000000083000000000000001200000000",
            INIT_63 => X"0000001600000000000000b90000000000000068000000000000002500000000",
            INIT_64 => X"0000000000000000000000200000000000000000000000000000000d00000000",
            INIT_65 => X"00000021000000000000003d000000000000001b000000000000001b00000000",
            INIT_66 => X"000000250000000000000000000000000000000d000000000000001400000000",
            INIT_67 => X"0000000b000000000000000500000000000000a200000000000000a300000000",
            INIT_68 => X"00000000000000000000001e0000000000000012000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000006a00000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000003b00000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000006700000000000000760000000000000066000000000000000000000000",
            INIT_7B => X"0000007300000000000000610000000000000064000000000000006300000000",
            INIT_7C => X"000000680000000000000070000000000000007e000000000000008f00000000",
            INIT_7D => X"0000005b000000000000004e000000000000004d000000000000006500000000",
            INIT_7E => X"0000006e00000000000000740000000000000075000000000000006200000000",
            INIT_7F => X"0000007500000000000000220000000000000000000000000000006600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE3;


    MEM_IFMAP_LAYER1_INSTANCE4 : if BRAM_NAME = "ifmap_layer1_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000009300000000",
            INIT_01 => X"0000006f00000000000000470000000000000050000000000000001400000000",
            INIT_02 => X"0000008000000000000000790000000000000070000000000000009a00000000",
            INIT_03 => X"00000000000000000000000c000000000000003400000000000000c200000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"000000000000000000000000000000000000003b000000000000000000000000",
            INIT_06 => X"00000004000000000000004b0000000000000077000000000000004b00000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000003d00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000002900000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000006d00000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000005200000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000002e000000000000004a0000000000000007000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_1A => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_1F => X"00000000000000000000003e0000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000002400000000000000230000000000000000000000000000000000000000",
            INIT_33 => X"0000001c00000000000000230000000000000024000000000000001900000000",
            INIT_34 => X"0000002c00000000000000250000000000000024000000000000002100000000",
            INIT_35 => X"0000001a00000000000000120000000000000011000000000000001800000000",
            INIT_36 => X"0000001c00000000000000260000000000000026000000000000002a00000000",
            INIT_37 => X"000000020000000000000050000000000000001e000000000000002800000000",
            INIT_38 => X"00000028000000000000001c0000000000000015000000000000001d00000000",
            INIT_39 => X"0000002e00000000000000270000000000000013000000000000001c00000000",
            INIT_3A => X"0000002800000000000000270000000000000026000000000000002f00000000",
            INIT_3B => X"00000011000000000000000f0000000000000060000000000000002d00000000",
            INIT_3C => X"000000000000000000000014000000000000002c000000000000000200000000",
            INIT_3D => X"0000004900000000000000380000000000000016000000000000002800000000",
            INIT_3E => X"0000002b00000000000000230000000000000035000000000000002e00000000",
            INIT_3F => X"0000001d00000000000000000000000000000042000000000000000600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000019000000000000000f000000000000000a000000000000000d00000000",
            INIT_41 => X"000000560000000000000000000000000000002d000000000000001c00000000",
            INIT_42 => X"0000000000000000000000350000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000290000000000000000000000000000000000000000",
            INIT_44 => X"0000002a00000000000000260000000000000000000000000000001800000000",
            INIT_45 => X"0000000000000000000000340000000000000000000000000000000000000000",
            INIT_46 => X"0000002800000000000000000000000000000049000000000000000000000000",
            INIT_47 => X"00000000000000000000000d000000000000004b000000000000000700000000",
            INIT_48 => X"000000000000000000000011000000000000001f000000000000000000000000",
            INIT_49 => X"000000420000000000000000000000000000006d000000000000000000000000",
            INIT_4A => X"0000000000000000000000440000000000000000000000000000004e00000000",
            INIT_4B => X"0000000300000000000000000000000000000044000000000000003600000000",
            INIT_4C => X"0000000000000000000000110000000000000025000000000000001100000000",
            INIT_4D => X"0000000d000000000000004b0000000000000000000000000000002b00000000",
            INIT_4E => X"0000001b00000000000000040000000000000000000000000000004000000000",
            INIT_4F => X"0000001100000000000000150000000000000009000000000000003800000000",
            INIT_50 => X"0000000100000000000000000000000000000000000000000000001a00000000",
            INIT_51 => X"0000000000000000000000000000000000000034000000000000000000000000",
            INIT_52 => X"0000003300000000000000070000000000000048000000000000001800000000",
            INIT_53 => X"0000002f00000000000000150000000000000000000000000000005300000000",
            INIT_54 => X"0000001200000000000000000000000000000000000000000000002900000000",
            INIT_55 => X"0000000000000000000000000000000000000009000000000000001900000000",
            INIT_56 => X"0000000a00000000000000030000000000000000000000000000006300000000",
            INIT_57 => X"0000001900000000000000340000000000000031000000000000001300000000",
            INIT_58 => X"0000000000000000000000170000000000000000000000000000006600000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000001700000000000000220000000000000000000000000000000000000000",
            INIT_5B => X"000000430000000000000034000000000000003d000000000000000b00000000",
            INIT_5C => X"0000002e00000000000000400000000000000000000000000000000000000000",
            INIT_5D => X"0000001a0000000000000016000000000000001d000000000000000000000000",
            INIT_5E => X"000000270000000000000023000000000000002b000000000000002300000000",
            INIT_5F => X"0000001a0000000000000027000000000000001d000000000000002300000000",
            INIT_60 => X"0000001200000000000000000000000000000068000000000000000000000000",
            INIT_61 => X"000000280000000000000025000000000000001a000000000000001900000000",
            INIT_62 => X"0000001400000000000000210000000000000023000000000000002800000000",
            INIT_63 => X"00000000000000000000001f0000000000000025000000000000001800000000",
            INIT_64 => X"0000001a0000000000000014000000000000000c000000000000008b00000000",
            INIT_65 => X"0000002000000000000000170000000000000014000000000000001d00000000",
            INIT_66 => X"0000003d00000000000000280000000000000021000000000000003100000000",
            INIT_67 => X"0000007300000000000000190000000000000023000000000000001800000000",
            INIT_68 => X"000000100000000000000023000000000000002c000000000000002f00000000",
            INIT_69 => X"0000001800000000000000260000000000000022000000000000001800000000",
            INIT_6A => X"0000004e0000000000000028000000000000003b000000000000001d00000000",
            INIT_6B => X"0000004d0000000000000052000000000000004f000000000000005900000000",
            INIT_6C => X"0000004b0000000000000056000000000000005a000000000000005400000000",
            INIT_6D => X"0000003d00000000000000410000000000000045000000000000004e00000000",
            INIT_6E => X"0000005600000000000000490000000000000033000000000000003f00000000",
            INIT_6F => X"00000082000000000000004b0000000000000059000000000000005300000000",
            INIT_70 => X"0000001d000000000000003c0000000000000060000000000000005900000000",
            INIT_71 => X"00000037000000000000002e000000000000002a000000000000002900000000",
            INIT_72 => X"00000057000000000000003c0000000000000063000000000000003d00000000",
            INIT_73 => X"0000003e00000000000000910000000000000056000000000000005400000000",
            INIT_74 => X"00000054000000000000003f0000000000000000000000000000000d00000000",
            INIT_75 => X"0000003f00000000000000180000000000000029000000000000002100000000",
            INIT_76 => X"00000054000000000000005d0000000000000029000000000000003900000000",
            INIT_77 => X"00000019000000000000005a0000000000000021000000000000006200000000",
            INIT_78 => X"0000003b00000000000000570000000000000046000000000000001d00000000",
            INIT_79 => X"0000003300000000000000250000000000000003000000000000001300000000",
            INIT_7A => X"000000ac00000000000000210000000000000059000000000000008c00000000",
            INIT_7B => X"00000024000000000000002d0000000000000071000000000000006200000000",
            INIT_7C => X"0000002100000000000000330000000000000062000000000000000000000000",
            INIT_7D => X"000000a900000000000000400000000000000004000000000000000800000000",
            INIT_7E => X"0000006400000000000000bb0000000000000055000000000000006000000000",
            INIT_7F => X"00000046000000000000002e000000000000003b000000000000009300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE4;


    MEM_IFMAP_LAYER1_INSTANCE5 : if BRAM_NAME = "ifmap_layer1_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001200000000000000290000000000000026000000000000008a00000000",
            INIT_01 => X"0000005300000000000000ca0000000000000023000000000000000000000000",
            INIT_02 => X"000000c60000000000000074000000000000006d000000000000004c00000000",
            INIT_03 => X"0000006c000000000000007e0000000000000041000000000000005500000000",
            INIT_04 => X"0000002a0000000000000027000000000000001a000000000000002c00000000",
            INIT_05 => X"00000054000000000000002e0000000000000090000000000000005f00000000",
            INIT_06 => X"00000060000000000000007b00000000000000cb000000000000002f00000000",
            INIT_07 => X"000000350000000000000066000000000000007a000000000000003100000000",
            INIT_08 => X"0000008d000000000000001e000000000000004b000000000000002100000000",
            INIT_09 => X"000000470000000000000067000000000000004b00000000000000a800000000",
            INIT_0A => X"0000002a000000000000004e0000000000000042000000000000004600000000",
            INIT_0B => X"0000000900000000000000170000000000000069000000000000005700000000",
            INIT_0C => X"0000009f00000000000000a00000000000000050000000000000002800000000",
            INIT_0D => X"00000012000000000000006a0000000000000053000000000000007000000000",
            INIT_0E => X"0000004d00000000000000480000000000000087000000000000002300000000",
            INIT_0F => X"0000005d00000000000000200000000000000000000000000000001a00000000",
            INIT_10 => X"00000073000000000000009b00000000000000b3000000000000005200000000",
            INIT_11 => X"00000094000000000000005e0000000000000096000000000000006f00000000",
            INIT_12 => X"000000000000000000000000000000000000004800000000000000a100000000",
            INIT_13 => X"00000030000000000000003e000000000000001e000000000000000000000000",
            INIT_14 => X"000000fb00000000000000640000000000000089000000000000008400000000",
            INIT_15 => X"000000280000000000000033000000000000002d00000000000000fb00000000",
            INIT_16 => X"000000150000000000000016000000000000000a000000000000001500000000",
            INIT_17 => X"00000020000000000000001d0000000000000025000000000000001a00000000",
            INIT_18 => X"00000026000000000000012e000000000000004e000000000000006000000000",
            INIT_19 => X"0000000900000000000000100000000000000018000000000000001500000000",
            INIT_1A => X"00000030000000000000001e000000000000000c000000000000000800000000",
            INIT_1B => X"0000001900000000000000170000000000000021000000000000001e00000000",
            INIT_1C => X"00000017000000000000001600000000000000dd000000000000006500000000",
            INIT_1D => X"00000015000000000000000d0000000000000014000000000000001400000000",
            INIT_1E => X"0000002600000000000000110000000000000026000000000000001b00000000",
            INIT_1F => X"0000002a00000000000000160000000000000021000000000000005700000000",
            INIT_20 => X"0000001b0000000000000015000000000000000d000000000000004800000000",
            INIT_21 => X"0000001e00000000000000210000000000000018000000000000000f00000000",
            INIT_22 => X"000000100000000000000051000000000000001b000000000000000700000000",
            INIT_23 => X"0000000300000000000000080000000000000007000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_26 => X"0000000a00000000000000010000000000000000000000000000000000000000",
            INIT_27 => X"000000080000000000000000000000000000000b000000000000001a00000000",
            INIT_28 => X"000000000000000000000021000000000000000000000000000000ac00000000",
            INIT_29 => X"00000000000000000000000e0000000000000020000000000000001e00000000",
            INIT_2A => X"000000000000000000000015000000000000000c000000000000000000000000",
            INIT_2B => X"00000000000000000000000e0000000000000000000000000000000b00000000",
            INIT_2C => X"0000005a000000000000001f0000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000a30000000000000000000000000000001e00000000",
            INIT_2F => X"0000004200000000000000000000000000000035000000000000001400000000",
            INIT_30 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_31 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"000000040000000000000000000000000000008e000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000008500000000",
            INIT_34 => X"0000000000000000000000000000000000000035000000000000000000000000",
            INIT_35 => X"0000000000000000000000110000000000000000000000000000001600000000",
            INIT_36 => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000012c00000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"00000069000000000000003c0000000000000000000000000000000000000000",
            INIT_3B => X"000000cc00000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000830000000000000011000000000000000000000000",
            INIT_3F => X"0000000000000000000000700000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_41 => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000003e00000000000000000000000000000000000000000000000d00000000",
            INIT_43 => X"0000000000000000000000270000000000000000000000000000000000000000",
            INIT_44 => X"00000000000000000000003f0000000000000008000000000000000000000000",
            INIT_45 => X"0000000000000000000000200000000000000000000000000000000000000000",
            INIT_46 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_47 => X"0000004a00000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000470000000000000000000000000000005500000000",
            INIT_49 => X"0000003d000000000000000000000000000000eb000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000006100000000",
            INIT_4B => X"000000000000000000000025000000000000005f000000000000002e00000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"000000000000000000000000000000000000000000000000000000ba00000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000025000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_62 => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000005400000000",
            INIT_64 => X"000000000000000000000000000000000000000000000000000000c500000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000002f00000000",
            INIT_66 => X"000000000000000000000000000000000000002d000000000000001300000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"000000af00000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"00000000000000000000000f0000000000000000000000000000009200000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000003b00000000",
            INIT_6C => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"000000000000000000000000000000000000002d000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000015a00000000",
            INIT_70 => X"0000000000000000000000000000000000000092000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000003600000000",
            INIT_72 => X"000000d700000000000000000000000000000004000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000059000000000000000000000000",
            INIT_74 => X"000000000000000000000000000000000000000000000000000000be00000000",
            INIT_75 => X"0000001900000000000000000000000000000000000000000000000400000000",
            INIT_76 => X"000000d4000000000000003e0000000000000000000000000000000000000000",
            INIT_77 => X"0000008700000000000000000000000000000007000000000000000000000000",
            INIT_78 => X"0000000700000000000000360000000000000000000000000000000000000000",
            INIT_79 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_7A => X"00000011000000000000005f0000000000000000000000000000006100000000",
            INIT_7B => X"000000b60000000000000000000000000000002d000000000000000000000000",
            INIT_7C => X"000000000000000000000043000000000000001d000000000000000000000000",
            INIT_7D => X"0000004d00000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"000000220000000000000000000000000000002a000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE5;


    MEM_IFMAP_LAYER1_INSTANCE6 : if BRAM_NAME = "ifmap_layer1_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b400000000000000000000000000000002000000000000004400000000",
            INIT_01 => X"0000000000000000000000850000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000003a00000000000001000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000051000000000000000000000000",
            INIT_06 => X"000000000000000000000007000000000000003d000000000000003c00000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"00000000000000000000008b0000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000004300000000000000820000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000001000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000030000000000000003200000000",
            INIT_12 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000009000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000009200000000000000970000000000000093000000000000008b00000000",
            INIT_4D => X"0000009b00000000000000ab000000000000009c000000000000008300000000",
            INIT_4E => X"000000710000000000000066000000000000005a000000000000007400000000",
            INIT_4F => X"00000099000000000000009a000000000000007f000000000000007900000000",
            INIT_50 => X"00000066000000000000009e0000000000000098000000000000009a00000000",
            INIT_51 => X"0000002a0000000000000039000000000000006e000000000000007600000000",
            INIT_52 => X"0000006e00000000000000200000000000000000000000000000000000000000",
            INIT_53 => X"000000a1000000000000007c0000000000000037000000000000007d00000000",
            INIT_54 => X"00000039000000000000004d000000000000009f00000000000000a000000000",
            INIT_55 => X"0000000000000000000000000000000000000022000000000000001500000000",
            INIT_56 => X"0000006200000000000000260000000000000000000000000000000000000000",
            INIT_57 => X"0000009f00000000000000910000000000000032000000000000000000000000",
            INIT_58 => X"000000000000000000000014000000000000005a000000000000006600000000",
            INIT_59 => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_5A => X"0000000000000000000000460000000000000000000000000000000000000000",
            INIT_5B => X"00000017000000000000009f0000000000000069000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_5E => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_5F => X"000000120000000000000006000000000000002f000000000000006e00000000",
            INIT_60 => X"0000002c00000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000005e00000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000250000000000000000000000000000006200000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_66 => X"0000003700000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000011000000000000003600000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_69 => X"0000000000000000000000470000000000000000000000000000000000000000",
            INIT_6A => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000002000000000000000000000000000000012000000000000000000000000",
            INIT_6C => X"000000000000000000000000000000000000002f000000000000000000000000",
            INIT_6D => X"000000000000000000000000000000000000005e000000000000003700000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000001a00000000000000000000000000000000000000000000000e00000000",
            INIT_70 => X"0000004b00000000000000020000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000006a00000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE6;


    MEM_IFMAP_LAYER1_INSTANCE7 : if BRAM_NAME = "ifmap_layer1_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE7;


    MEM_IFMAP_LAYER2_INSTANCE0 : if BRAM_NAME = "ifmap_layer2_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000019700000000000000550000000000000000000000000000011600000000",
            INIT_02 => X"00000000000000000000005200000000000000b7000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"000000f20000000000000026000000000000004700000000000000cc00000000",
            INIT_05 => X"0000000000000000000000170000000000000000000000000000002700000000",
            INIT_06 => X"0000002400000000000000000000000000000000000000000000005e00000000",
            INIT_07 => X"00000000000000000000006b000000000000007f000000000000000000000000",
            INIT_08 => X"00000000000000000000000000000000000001c4000000000000000000000000",
            INIT_09 => X"000000370000000000000059000000000000017d000000000000000000000000",
            INIT_0A => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"00000000000000000000009b0000000000000090000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000018000000000000001f00000000",
            INIT_12 => X"000000840000000000000000000000000000000f000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000d20000000000000000000000000000000000000000",
            INIT_15 => X"000001a900000000000000000000000000000000000000000000007400000000",
            INIT_16 => X"000000000000000000000018000000000000000500000000000000cc00000000",
            INIT_17 => X"0000001500000000000000270000000000000046000000000000023300000000",
            INIT_18 => X"0000000000000000000000000000000000000003000000000000001200000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000500000000000000000000000000000000000000000",
            INIT_21 => X"0000013200000000000000000000000000000087000000000000000000000000",
            INIT_22 => X"000000a300000000000000f5000000000000008800000000000000fb00000000",
            INIT_23 => X"000000f5000000000000015e000000000000013d000000000000000000000000",
            INIT_24 => X"000000db00000000000000b500000000000000d300000000000000da00000000",
            INIT_25 => X"000000000000000000000000000000000000003f000000000000015000000000",
            INIT_26 => X"0000001f0000000000000000000000000000006d000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000007500000000000000100000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000650000000000000000000000000000000000000000",
            INIT_2D => X"00000000000000000000000000000000000000ad000000000000000000000000",
            INIT_2E => X"000000b900000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"00000000000000000000002d0000000000000067000000000000001b00000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000c10000000000000000000000000000000000000000",
            INIT_34 => X"000000000000000000000000000000000000011b000000000000000000000000",
            INIT_35 => X"000000da00000000000000000000000000000053000000000000000000000000",
            INIT_36 => X"000000000000000000000058000000000000001b000000000000002e00000000",
            INIT_37 => X"0000000000000000000000aa0000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000052000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000001090000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000210000000000000000000000000000014300000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000040000000000000000000000000000002600000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"00000000000000000000000a0000000000000000000000000000000900000000",
            INIT_43 => X"0000001e0000000000000000000000000000002e000000000000000000000000",
            INIT_44 => X"0000000000000000000000390000000000000000000000000000002b00000000",
            INIT_45 => X"000000000000000000000000000000000000018b000000000000000000000000",
            INIT_46 => X"0000009e000000000000009b0000000000000000000000000000003900000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000010000000000000000000000000000011900000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"000001e4000000000000021c0000000000000258000000000000005300000000",
            INIT_4B => X"00000083000000000000000000000000000000a7000000000000011c00000000",
            INIT_4C => X"0000007f00000000000000000000000000000000000000000000001000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000057000000000000000000000000",
            INIT_4F => X"000000000000000000000056000000000000007c00000000000000d900000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000008300000000",
            INIT_51 => X"0000011c00000000000001150000000000000026000000000000003b00000000",
            INIT_52 => X"0000020f000000000000001b0000000000000007000000000000000000000000",
            INIT_53 => X"000000000000000000000000000000000000000b00000000000000a200000000",
            INIT_54 => X"00000000000000000000000800000000000000f7000000000000002200000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000780000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000042000000000000000000000000",
            INIT_5A => X"000000120000000000000000000000000000006e000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000570000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000bd0000000000000019000000000000004200000000",
            INIT_5E => X"000001bb00000000000000000000000000000042000000000000000400000000",
            INIT_5F => X"0000000100000000000000200000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000004900000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000004200000000000000290000000000000000000000000000000f00000000",
            INIT_63 => X"0000004f00000000000000000000000000000097000000000000000a00000000",
            INIT_64 => X"0000000000000000000000e10000000000000112000000000000000000000000",
            INIT_65 => X"0000000000000000000000390000000000000014000000000000000000000000",
            INIT_66 => X"0000000000000000000000a20000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000061000000000000000000000000",
            INIT_69 => X"000000ee000000000000007400000000000000cc000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000007300000000",
            INIT_6B => X"0000000000000000000000000000000000000111000000000000018700000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000150000000000000054000000000000006300000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000009100000000",
            INIT_72 => X"0000025b00000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000d80000000000000000000000000000000000000000",
            INIT_75 => X"0000000200000000000001a20000000000000000000000000000000000000000",
            INIT_76 => X"0000007100000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"000000000000000000000000000000000000008f000000000000000000000000",
            INIT_78 => X"000000000000000000000000000000000000003c000000000000002000000000",
            INIT_79 => X"0000000000000000000000000000000000000094000000000000000000000000",
            INIT_7A => X"0000002f00000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"000000e0000000000000014500000000000001de000000000000012700000000",
            INIT_7C => X"0000009900000000000000a6000000000000007c000000000000002f00000000",
            INIT_7D => X"00000000000000000000009b0000000000000000000000000000011600000000",
            INIT_7E => X"0000003000000000000000000000000000000000000000000000005900000000",
            INIT_7F => X"0000007c0000000000000000000000000000005f000000000000002700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE0;


    MEM_IFMAP_LAYER2_INSTANCE1 : if BRAM_NAME = "ifmap_layer2_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000006e0000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000003100000000000000d100000000000000e5000000000000002e00000000",
            INIT_03 => X"0000007600000000000001e90000000000000000000000000000009700000000",
            INIT_04 => X"0000009c00000000000000cc00000000000000dc00000000000000f900000000",
            INIT_05 => X"00000000000000000000005f000000000000003c000000000000000000000000",
            INIT_06 => X"0000004700000000000000f20000000000000002000000000000002c00000000",
            INIT_07 => X"00000000000000000000006a0000000000000036000000000000006900000000",
            INIT_08 => X"00000054000000000000009f00000000000000e4000000000000009f00000000",
            INIT_09 => X"000000000000000000000036000000000000000d000000000000000000000000",
            INIT_0A => X"0000009000000000000000f400000000000000aa000000000000000000000000",
            INIT_0B => X"0000008500000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000002200000000000000a300000000000000d4000000000000006a00000000",
            INIT_0D => X"0000000000000000000000ad000000000000000000000000000000e500000000",
            INIT_0E => X"000000e200000000000000fb0000000000000162000000000000000000000000",
            INIT_0F => X"0000004f00000000000000c900000000000000b4000000000000003c00000000",
            INIT_10 => X"00000067000000000000007b00000000000000f8000000000000000000000000",
            INIT_11 => X"00000000000000000000008e0000000000000031000000000000003900000000",
            INIT_12 => X"0000000000000000000000000000000000000004000000000000000500000000",
            INIT_13 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000680000000000000109000000000000004300000000",
            INIT_15 => X"0000000000000000000000e30000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000aa0000000000000000000000000000009b00000000",
            INIT_17 => X"000000da000000000000000000000000000001b1000000000000000000000000",
            INIT_18 => X"00000000000000000000005f0000000000000125000000000000004e00000000",
            INIT_19 => X"00000000000000000000008b0000000000000000000000000000011800000000",
            INIT_1A => X"000000d60000000000000000000000000000008a00000000000000a900000000",
            INIT_1B => X"0000000000000000000000000000000000000036000000000000004c00000000",
            INIT_1C => X"000000e2000000000000000000000000000001f5000000000000000000000000",
            INIT_1D => X"0000009a00000000000000000000000000000021000000000000000000000000",
            INIT_1E => X"00000008000000000000001a000000000000003b000000000000004e00000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"00000000000000000000001d0000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000860000000000000000000000000000015400000000",
            INIT_2D => X"00000000000000000000004b000000000000001a000000000000002b00000000",
            INIT_2E => X"000000000000000000000000000000000000007e000000000000000000000000",
            INIT_2F => X"00000000000000000000001d000000000000000000000000000001c300000000",
            INIT_30 => X"0000013b000000000000009d000000000000000000000000000000ac00000000",
            INIT_31 => X"000000f9000000000000004c0000000000000187000000000000014400000000",
            INIT_32 => X"00000000000000000000007600000000000000a8000000000000000000000000",
            INIT_33 => X"00000000000000000000002c0000000000000148000000000000000000000000",
            INIT_34 => X"000000000000000000000240000000000000003200000000000000a800000000",
            INIT_35 => X"000000000000000000000022000000000000002f000000000000000000000000",
            INIT_36 => X"0000000c000000000000002000000000000002fb000000000000000000000000",
            INIT_37 => X"0000000000000000000000600000000000000036000000000000002000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000006e0000000000000058000000000000002b000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000007e000000000000004f00000000000000e2000000000000005300000000",
            INIT_3D => X"0000001f00000000000000000000000000000099000000000000006b00000000",
            INIT_3E => X"0000009800000000000000170000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000005800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000010200000000000000c80000000000000000000000000000000000000000",
            INIT_42 => X"00000047000000000000002d000000000000000000000000000000fe00000000",
            INIT_43 => X"000000b40000000000000103000000000000012d00000000000000a500000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000004f00000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"000000000000000000000121000000000000008e000000000000004800000000",
            INIT_48 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_4A => X"0000015100000000000000000000000000000000000000000000007100000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000006a000000000000007700000000000000ca000000000000000000000000",
            INIT_4E => X"0000000000000000000000f0000000000000007a000000000000000000000000",
            INIT_4F => X"00000060000000000000001d0000000000000031000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000007300000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000003500000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"000000000000000000000000000000000000006f000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000af0000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000670000000000000000000000000000000000000000",
            INIT_72 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000115000000000000004f00000000",
            INIT_74 => X"000000c700000000000000b10000000000000086000000000000008900000000",
            INIT_75 => X"0000010d0000000000000080000000000000001a000000000000007900000000",
            INIT_76 => X"0000003b000000000000007e000000000000003200000000000000a200000000",
            INIT_77 => X"00000000000000000000000000000000000000b3000000000000011700000000",
            INIT_78 => X"000000000000000000000000000000000000005d000000000000002800000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000930000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000007b00000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_7D => X"0000000000000000000000f90000000000000043000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE1;


    MEM_IFMAP_LAYER2_INSTANCE2 : if BRAM_NAME = "ifmap_layer2_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000420000000000000000000000000000000000000000",
            INIT_02 => X"0000007900000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"000000000000000000000000000000000000002a000000000000007300000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000008600000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"000000bc00000000000000e600000000000000e6000000000000015100000000",
            INIT_18 => X"000000000000000000000000000000000000000000000000000000d500000000",
            INIT_19 => X"0000000000000000000000bd00000000000000a600000000000000b000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"000000380000000000000000000000000000006f000000000000000000000000",
            INIT_1D => X"000000c500000000000001080000000000000000000000000000004600000000",
            INIT_1E => X"0000000000000000000000330000000000000000000000000000001400000000",
            INIT_1F => X"00000020000000000000008e0000000000000000000000000000000000000000",
            INIT_20 => X"000000000000000000000066000000000000007e000000000000003900000000",
            INIT_21 => X"0000007300000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000003200000000000000c70000000000000000000000000000000000000000",
            INIT_23 => X"000000000000000000000000000000000000007b000000000000001a00000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000c90000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000008200000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000004000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000014b00000000000000310000000000000000000000000000000000000000",
            INIT_30 => X"00000000000000000000001200000000000000b100000000000000a000000000",
            INIT_31 => X"0000007300000000000000bf0000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000029000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000005200000000",
            INIT_39 => X"00000000000000000000000000000000000000b7000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"000000000000000000000000000000000000000000000000000000eb00000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000028000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000005000000000",
            INIT_43 => X"0000009500000000000000000000000000000000000000000000000f00000000",
            INIT_44 => X"0000004600000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000001000000000000000150000000000000000000000000000000000000000",
            INIT_46 => X"00000000000000000000007300000000000000a4000000000000000000000000",
            INIT_47 => X"0000000000000000000001810000000000000153000000000000000000000000",
            INIT_48 => X"0000014a00000000000001450000000000000115000000000000018300000000",
            INIT_49 => X"0000009700000000000000d0000000000000011b00000000000001c500000000",
            INIT_4A => X"00000108000000000000012f00000000000000de00000000000000c100000000",
            INIT_4B => X"0000000000000000000000a00000000000000000000000000000000000000000",
            INIT_4C => X"00000099000000000000000c00000000000001b1000000000000000800000000",
            INIT_4D => X"0000000000000000000000fb0000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000004000000000",
            INIT_4F => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_50 => X"00000000000000000000002e00000000000000b9000000000000000000000000",
            INIT_51 => X"00000000000000000000008f0000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"00000000000000000000011b00000000000000ef000000000000003e00000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000018000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"00000137000000000000021100000000000001db000000000000010f00000000",
            INIT_58 => X"0000000000000000000000380000000000000000000000000000003c00000000",
            INIT_59 => X"0000000900000000000000000000000000000000000000000000014a00000000",
            INIT_5A => X"0000012800000000000000000000000000000000000000000000005a00000000",
            INIT_5B => X"000000c2000000000000007d0000000000000067000000000000000000000000",
            INIT_5C => X"0000015100000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000400000000000000db00000000000000e9000000000000008800000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"000000cb00000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000009400000000000000300000000000000000000000000000000000000000",
            INIT_66 => X"000000000000000000000000000000000000001f000000000000000000000000",
            INIT_67 => X"0000007700000000000000e70000000000000023000000000000017c00000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000002e00000000",
            INIT_69 => X"000000b3000000000000007c0000000000000000000000000000003d00000000",
            INIT_6A => X"0000005300000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000005300000000",
            INIT_6C => X"0000000000000000000001080000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000067000000000000000000000000",
            INIT_6F => X"000000e7000000000000005d0000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000500000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000003100000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"000000000000000000000000000000000000002f000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000003000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"00000071000000000000005c00000000000000b0000000000000001200000000",
            INIT_7D => X"0000007b000000000000002c0000000000000000000000000000005000000000",
            INIT_7E => X"000000000000000000000008000000000000007a000000000000004e00000000",
            INIT_7F => X"0000000000000000000000660000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE2;


    MEM_IFMAP_LAYER2_INSTANCE3 : if BRAM_NAME = "ifmap_layer2_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003700000000000000000000000000000089000000000000000700000000",
            INIT_01 => X"00000024000000000000000000000000000000aa000000000000008600000000",
            INIT_02 => X"00000010000000000000004d0000000000000002000000000000004300000000",
            INIT_03 => X"00000034000000000000006200000000000000a000000000000000d000000000",
            INIT_04 => X"0000008200000000000000000000000000000000000000000000002a00000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE3;


    MEM_IFMAP_LAYER3_INSTANCE0 : if BRAM_NAME = "ifmap_layer3_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000dd0000000000000000000000000000000000000000",
            INIT_06 => X"0000018f00000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"000000000000000000000000000000000000007b000000000000000000000000",
            INIT_0B => X"000000f900000000000000850000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000fc0000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000017f00000000000001fa0000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_13 => X"0000000000000000000000000000000000000086000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000270000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000111000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"000002fe00000000000000810000000000000000000000000000017400000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"000000000000000000000000000000000000000000000000000000fb00000000",
            INIT_1C => X"000000000000000000000000000000000000035d000000000000000000000000",
            INIT_1D => X"00000126000000000000020600000000000002ba000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"000000000000000000000000000000000000000000000000000001f200000000",
            INIT_23 => X"0000009d00000000000003370000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"000001f500000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000a20000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"000001d400000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000007900000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000007b0000000000000000000000000000030d000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000010e00000000000000000000000000000108000000000000000000000000",
            INIT_2F => X"000000000000000000000000000000000000000000000000000003d700000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000003600000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"000000c100000000000000cf0000000000000000000000000000010b00000000",
            INIT_37 => X"0000000000000000000000c100000000000002bd000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"000001c50000000000000170000000000000023b000000000000000000000000",
            INIT_3A => X"0000008e000000000000000000000000000001f8000000000000000000000000",
            INIT_3B => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"000000b800000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"00000382000000000000023f000000000000015a000000000000008d00000000",
            INIT_3E => X"0000000000000000000002fd000000000000036300000000000003ed00000000",
            INIT_3F => X"0000013e000000000000000000000000000001c1000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000000000000000000000000000000000002b6000000000000029100000000",
            INIT_41 => X"0000000000000000000004730000000000000205000000000000000000000000",
            INIT_42 => X"0000031900000000000002ef0000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000061000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"000000000000000000000000000000000000000000000000000000c100000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"000000eb00000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"00000000000000000000000000000000000001e900000000000003c800000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000ce00000000000000000000000000000000000000000000009900000000",
            INIT_52 => X"000000000000000000000000000000000000022300000000000002f500000000",
            INIT_53 => X"00000000000000000000028c0000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"00000000000000000000000000000000000005cf000000000000033500000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"000001ea00000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"000000000000000000000000000000000000033b000000000000021300000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"00000090000000000000019f000000000000000000000000000000eb00000000",
            INIT_5B => X"000000000000000000000000000000000000000000000000000001cb00000000",
            INIT_5C => X"0000000000000000000002ff0000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000093000000000000006700000000",
            INIT_5E => X"000000000000000000000200000000000000019e000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000015e00000000",
            INIT_60 => X"0000000000000000000000d10000000000000000000000000000000000000000",
            INIT_61 => X"000001f900000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"00000000000000000000000000000000000002dc000000000000012c00000000",
            INIT_64 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_65 => X"000000000000000000000000000000000000011e00000000000001b500000000",
            INIT_66 => X"00000000000000000000021c0000000000000178000000000000034700000000",
            INIT_67 => X"0000004400000000000000ab0000000000000000000000000000000000000000",
            INIT_68 => X"000000000000000000000000000000000000000000000000000003db00000000",
            INIT_69 => X"0000000000000000000000bb0000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000031000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000db0000000000000000000000000000017e00000000",
            INIT_6D => X"00000000000000000000034f0000000000000000000000000000009a00000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"00000145000000000000028f0000000000000026000000000000000000000000",
            INIT_70 => X"0000000000000000000000b3000000000000016a000000000000004100000000",
            INIT_71 => X"0000036900000000000001b30000000000000000000000000000000000000000",
            INIT_72 => X"000000a900000000000000000000000000000000000000000000026e00000000",
            INIT_73 => X"0000008d00000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000001740000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000027b00000000",
            INIT_76 => X"00000000000000000000000000000000000001f9000000000000002700000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000033d00000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000010e00000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"000000000000000000000000000000000000001e000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER3_INSTANCE0;


    MEM_IFMAP_LAYER3_INSTANCE1 : if BRAM_NAME = "ifmap_layer3_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000043100000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000028400000000000000000000000000000000000000000000015700000000",
            INIT_02 => X"00000000000000000000000000000000000003e400000000000000d800000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000005a20000000000000559000000000000038300000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000011d00000000000001550000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000001670000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000007900000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"00000000000000000000036f0000000000000000000000000000000000000000",
            INIT_0C => X"000001ce000000000000019700000000000000c400000000000001ab00000000",
            INIT_0D => X"000001cc0000000000000000000000000000000000000000000001fb00000000",
            INIT_0E => X"0000030e00000000000000fa0000000000000345000000000000028b00000000",
            INIT_0F => X"000002f300000000000006ca0000000000000000000000000000043f00000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER3_INSTANCE1;


    MEM_GOLD_LAYER0_INSTANCE0 : if BRAM_NAME = "gold_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000021000000000000001f000000000000002f000000000000001800000000",
            INIT_01 => X"0000002c00000000000000240000000000000028000000000000001900000000",
            INIT_02 => X"0000001900000000000000080000000000000000000000000000001b00000000",
            INIT_03 => X"0000001c0000000000000027000000000000002a000000000000002800000000",
            INIT_04 => X"000000190000000000000021000000000000001d000000000000003b00000000",
            INIT_05 => X"0000001300000000000000100000000000000013000000000000001b00000000",
            INIT_06 => X"0000000b00000000000000080000000000000000000000000000000f00000000",
            INIT_07 => X"000000000000000000000000000000000000001b000000000000001000000000",
            INIT_08 => X"000000220000000000000014000000000000002b000000000000002100000000",
            INIT_09 => X"000000000000000000000009000000000000002c000000000000003400000000",
            INIT_0A => X"0000000000000000000000030000000000000012000000000000000700000000",
            INIT_0B => X"0000001b00000000000000000000000000000030000000000000002000000000",
            INIT_0C => X"0000000c000000000000000f0000000000000012000000000000001d00000000",
            INIT_0D => X"0000003200000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000100000000000000030000000000000000e00000000",
            INIT_0F => X"0000000000000000000000120000000000000000000000000000002000000000",
            INIT_10 => X"0000002a00000000000000370000000000000000000000000000000000000000",
            INIT_11 => X"0000001c000000000000001b0000000000000000000000000000001d00000000",
            INIT_12 => X"0000000000000000000000000000000000000021000000000000000e00000000",
            INIT_13 => X"0000002f000000000000000f0000000000000032000000000000000000000000",
            INIT_14 => X"00000034000000000000002b0000000000000041000000000000003000000000",
            INIT_15 => X"0000000000000000000000350000000000000005000000000000000000000000",
            INIT_16 => X"00000002000000000000000b0000000000000015000000000000001200000000",
            INIT_17 => X"000000000000000000000000000000000000005c000000000000001900000000",
            INIT_18 => X"0000000000000000000000380000000000000019000000000000000000000000",
            INIT_19 => X"0000000400000000000000080000000000000025000000000000002f00000000",
            INIT_1A => X"0000000000000000000000320000000000000000000000000000000f00000000",
            INIT_1B => X"0000001900000000000000000000000000000000000000000000002000000000",
            INIT_1C => X"000000260000000000000000000000000000003b000000000000001400000000",
            INIT_1D => X"0000003d00000000000000040000000000000000000000000000003700000000",
            INIT_1E => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_1F => X"0000000f00000000000000420000000000000028000000000000000000000000",
            INIT_20 => X"0000004200000000000000110000000000000019000000000000000000000000",
            INIT_21 => X"0000000c00000000000000020000000000000027000000000000001900000000",
            INIT_22 => X"0000000c0000000000000000000000000000003b000000000000000000000000",
            INIT_23 => X"0000000000000000000000190000000000000006000000000000000000000000",
            INIT_24 => X"00000000000000000000001e0000000000000023000000000000000300000000",
            INIT_25 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_26 => X"0000000000000000000000020000000000000000000000000000004000000000",
            INIT_27 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"00000008000000000000002b0000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_3F => X"0000001e00000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000100000000000000000000000000000000000000000000001300000000",
            INIT_41 => X"00000000000000000000000a000000000000000e00000000000000b700000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000022000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000023000000000000000000000000",
            INIT_4A => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000008700000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"000000000000000000000000000000000000001500000000000000a700000000",
            INIT_4D => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000004e00000000000000000000000000000000000000000000000b00000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"000000480000000000000000000000000000005a000000000000005f00000000",
            INIT_55 => X"0000002300000000000000000000000000000002000000000000000300000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_57 => X"0000000000000000000000990000000000000000000000000000000000000000",
            INIT_58 => X"0000003e00000000000000240000000000000000000000000000000000000000",
            INIT_59 => X"000000000000000000000000000000000000003a000000000000006d00000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"000000000000000000000047000000000000003f000000000000000c00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000860000000000000000000000000000000000000000",
            INIT_62 => X"0000007500000000000000bf0000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000050000000000000006300000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000740000000000000000000000000000000000000000",
            INIT_66 => X"000000000000000000000000000000000000005c000000000000002e00000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000005f00000000000000590000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000590000000000000000000000000000000000000000",
            INIT_6D => X"0000001a000000000000006e000000000000000d000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000013000000000000002100000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"00000020000000000000002e0000000000000000000000000000000000000000",
            INIT_71 => X"0000002700000000000000250000000000000023000000000000003600000000",
            INIT_72 => X"0000000d0000000000000025000000000000002d000000000000002800000000",
            INIT_73 => X"0000001700000000000000240000000000000028000000000000001100000000",
            INIT_74 => X"0000003a00000000000000240000000000000028000000000000001300000000",
            INIT_75 => X"0000000000000000000000000000000000000042000000000000001c00000000",
            INIT_76 => X"0000000000000000000000150000000000000001000000000000000000000000",
            INIT_77 => X"0000000c0000000000000025000000000000000d000000000000000000000000",
            INIT_78 => X"00000022000000000000002b0000000000000063000000000000000000000000",
            INIT_79 => X"000000000000000000000000000000000000000b000000000000003b00000000",
            INIT_7A => X"000000000000000000000000000000000000003d000000000000002100000000",
            INIT_7B => X"00000000000000000000001b0000000000000021000000000000000000000000",
            INIT_7C => X"0000000000000000000000360000000000000004000000000000006200000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000004800000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000009700000000",
            INIT_7F => X"000000000000000000000000000000000000006f000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE0;


    MEM_GOLD_LAYER0_INSTANCE1 : if BRAM_NAME = "gold_layer0_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001e000000000000000000000000000000f0000000000000000000000000",
            INIT_01 => X"000000e800000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000005100000000",
            INIT_04 => X"0000000000000000000000540000000000000044000000000000007000000000",
            INIT_05 => X"00000000000000000000012e0000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_07 => X"0000000000000000000000060000000000000000000000000000002b00000000",
            INIT_08 => X"0000000000000000000000000000000000000063000000000000005b00000000",
            INIT_09 => X"00000000000000000000000000000000000000bd000000000000000000000000",
            INIT_0A => X"0000001100000000000000000000000000000002000000000000000000000000",
            INIT_0B => X"0000008000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_0D => X"0000002800000000000000000000000000000000000000000000008700000000",
            INIT_0E => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_0F => X"0000003800000000000000070000000000000000000000000000000000000000",
            INIT_10 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_11 => X"0000001e000000000000002f0000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_13 => X"0000006d000000000000006a0000000000000000000000000000003d00000000",
            INIT_14 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_15 => X"00000004000000000000002d000000000000001a000000000000000000000000",
            INIT_16 => X"000000fb00000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"00000000000000000000003f0000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000002000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"00000000000000000000005d0000000000000000000000000000002a00000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000003f00000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"000000000000000000000000000000000000000000000000000000d800000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"000000fa00000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000100000000000000000000000000000000000000000000000700000000",
            INIT_29 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000700000000000000040000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000060000000000000001000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000003700000000000000000000000000000000000000000000000500000000",
            INIT_2F => X"0000000000000000000000560000000000000053000000000000001c00000000",
            INIT_30 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000003500000000000000500000000000000005000000000000000500000000",
            INIT_32 => X"000000000000000000000000000000000000002500000000000000a700000000",
            INIT_33 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_34 => X"00000008000000000000000c0000000000000052000000000000000f00000000",
            INIT_35 => X"000000000000000000000000000000000000003e000000000000000300000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000120000000000000000000000000000000800000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000023000000000000004100000000",
            INIT_3B => X"000000000000000000000000000000000000002a000000000000000000000000",
            INIT_3C => X"00000000000000000000004b0000000000000001000000000000000000000000",
            INIT_3D => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_3F => X"0000003900000000000000000000000000000015000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_41 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000020000000000000032000000000000002300000000",
            INIT_43 => X"0000001000000000000000190000000000000006000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000004a00000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"00000000000000000000001d0000000000000071000000000000006300000000",
            INIT_49 => X"000000310000000000000003000000000000003b000000000000008200000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_4B => X"0000000000000000000000000000000000000055000000000000000000000000",
            INIT_4C => X"0000000000000000000000170000000000000000000000000000003400000000",
            INIT_4D => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_4E => X"0000001f00000000000000050000000000000009000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_50 => X"00000034000000000000001d0000000000000000000000000000000000000000",
            INIT_51 => X"0000003300000000000000320000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_53 => X"000000aa00000000000000b1000000000000009c000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000003600000000",
            INIT_55 => X"0000000000000000000000000000000000000009000000000000000700000000",
            INIT_56 => X"0000006200000000000000000000000000000017000000000000002e00000000",
            INIT_57 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_5A => X"0000000200000000000000000000000000000000000000000000000b00000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_5D => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"000000000000000000000007000000000000001e000000000000009c00000000",
            INIT_5F => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000330000000000000023000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"000000a000000000000000060000000000000011000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"00000000000000000000004a0000000000000000000000000000000000000000",
            INIT_69 => X"0000007800000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"000000000000000000000000000000000000000a000000000000000900000000",
            INIT_6B => X"0000000000000000000000500000000000000000000000000000000c00000000",
            INIT_6C => X"0000000000000000000000000000000000000080000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000001900000000000000000000000000000002000000000000001400000000",
            INIT_6F => X"000000000000000000000000000000000000000d000000000000002600000000",
            INIT_70 => X"00000000000000000000001d0000000000000000000000000000004f00000000",
            INIT_71 => X"0000000000000000000000320000000000000015000000000000000000000000",
            INIT_72 => X"0000003400000000000000000000000000000000000000000000002a00000000",
            INIT_73 => X"0000004300000000000000000000000000000019000000000000000000000000",
            INIT_74 => X"0000000000000000000000190000000000000000000000000000000000000000",
            INIT_75 => X"0000002c000000000000000a0000000000000000000000000000000000000000",
            INIT_76 => X"00000000000000000000003d0000000000000062000000000000000000000000",
            INIT_77 => X"0000004b00000000000000000000000000000000000000000000000f00000000",
            INIT_78 => X"0000000000000000000000000000000000000039000000000000000000000000",
            INIT_79 => X"0000000000000000000000680000000000000000000000000000005e00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000005200000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"000000bd00000000000000000000000000000009000000000000000000000000",
            INIT_7D => X"0000000b00000000000000000000000000000000000000000000002e00000000",
            INIT_7E => X"0000000000000000000000120000000000000000000000000000000d00000000",
            INIT_7F => X"0000000000000000000000230000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE1;


    MEM_GOLD_LAYER0_INSTANCE2 : if BRAM_NAME = "gold_layer0_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000056000000000000000000000000",
            INIT_01 => X"0000008100000000000000000000000000000064000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000002900000000000000000000000000000044000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"00000000000000000000001400000000000000bd000000000000004500000000",
            INIT_06 => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000007000000000",
            INIT_08 => X"00000038000000000000008b0000000000000088000000000000000e00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000100000000000000000000000000000035000000000000000f00000000",
            INIT_0B => X"0000000000000000000000200000000000000178000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000005900000000000000000000000000000000000000000000001700000000",
            INIT_0F => X"0000000000000000000000120000000000000000000000000000009c00000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000f00000000000000000000000000000012000000000000001900000000",
            INIT_12 => X"0000000f00000000000000c70000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000020000000000000003000000000000000000000000",
            INIT_15 => X"00000000000000000000002a0000000000000098000000000000000000000000",
            INIT_16 => X"00000000000000000000002b0000000000000055000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_18 => X"0000000a00000000000000000000000000000000000000000000000900000000",
            INIT_19 => X"0000004f00000000000000560000000000000042000000000000005200000000",
            INIT_1A => X"0000005400000000000000450000000000000058000000000000005800000000",
            INIT_1B => X"0000003e0000000000000047000000000000005f000000000000005c00000000",
            INIT_1C => X"0000005a00000000000000510000000000000049000000000000003700000000",
            INIT_1D => X"0000005e00000000000000450000000000000050000000000000005700000000",
            INIT_1E => X"0000006800000000000000640000000000000097000000000000003c00000000",
            INIT_1F => X"000000320000000000000045000000000000001e000000000000004000000000",
            INIT_20 => X"0000007e00000000000000570000000000000023000000000000001400000000",
            INIT_21 => X"0000004800000000000000610000000000000056000000000000000000000000",
            INIT_22 => X"000000000000000000000017000000000000008d000000000000000000000000",
            INIT_23 => X"00000053000000000000001c000000000000001d000000000000000000000000",
            INIT_24 => X"0000000000000000000000b50000000000000031000000000000000000000000",
            INIT_25 => X"0000000500000000000000960000000000000047000000000000004b00000000",
            INIT_26 => X"0000000000000000000000280000000000000027000000000000004e00000000",
            INIT_27 => X"00000045000000000000004d0000000000000000000000000000008500000000",
            INIT_28 => X"0000007000000000000000000000000000000066000000000000000000000000",
            INIT_29 => X"0000005f000000000000000a0000000000000069000000000000000000000000",
            INIT_2A => X"0000001600000000000000000000000000000047000000000000006b00000000",
            INIT_2B => X"000000000000000000000063000000000000001e000000000000006400000000",
            INIT_2C => X"00000043000000000000008c000000000000000c000000000000000000000000",
            INIT_2D => X"0000003200000000000000a50000000000000000000000000000000000000000",
            INIT_2E => X"00000065000000000000006a000000000000000000000000000000a600000000",
            INIT_2F => X"00000000000000000000003d000000000000002e000000000000000000000000",
            INIT_30 => X"0000000000000000000000b80000000000000016000000000000007900000000",
            INIT_31 => X"000000720000000000000064000000000000001f000000000000000000000000",
            INIT_32 => X"000000010000000000000056000000000000006d000000000000000000000000",
            INIT_33 => X"000000400000000000000017000000000000003b000000000000000000000000",
            INIT_34 => X"000000000000000000000000000000000000006e000000000000000000000000",
            INIT_35 => X"0000000000000000000000530000000000000010000000000000008300000000",
            INIT_36 => X"0000000000000000000000000000000000000058000000000000006300000000",
            INIT_37 => X"000000a10000000000000000000000000000003b000000000000003200000000",
            INIT_38 => X"0000002700000000000000000000000000000049000000000000000000000000",
            INIT_39 => X"0000000000000000000000430000000000000000000000000000004d00000000",
            INIT_3A => X"0000003000000000000000030000000000000000000000000000006700000000",
            INIT_3B => X"0000000000000000000000c40000000000000000000000000000001a00000000",
            INIT_3C => X"0000005200000000000000000000000000000000000000000000002400000000",
            INIT_3D => X"000000000000000000000065000000000000001a000000000000000300000000",
            INIT_3E => X"00000000000000000000004f000000000000000d000000000000000000000000",
            INIT_3F => X"000000f800000000000000000000000000000098000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006e00000000000000090000000000000000000000000000001000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_42 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_43 => X"0000002500000000000000850000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"000000000000000000000000000000000000006d000000000000003e00000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"000000b800000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000040000000000000033000000000000003d00000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"000000000000000000000000000000000000005f000000000000000000000000",
            INIT_58 => X"0000000000000000000000340000000000000000000000000000000000000000",
            INIT_59 => X"00000000000000000000000000000000000000a8000000000000001000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"00000000000000000000001d0000000000000017000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000005b00000000",
            INIT_60 => X"000000000000000000000000000000000000004c000000000000000000000000",
            INIT_61 => X"000000000000000000000000000000000000004d000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"000000000000000000000054000000000000005a000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_68 => X"00000000000000000000004a0000000000000000000000000000000000000000",
            INIT_69 => X"00000000000000000000002d0000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"000000070000000000000016000000000000002b000000000000008000000000",
            INIT_6E => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_70 => X"0000002600000000000000000000000000000022000000000000000000000000",
            INIT_71 => X"0000000000000000000000280000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000029000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"000000000000000000000010000000000000001b000000000000000000000000",
            INIT_75 => X"0000005500000000000000a10000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000030000000000000002600000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_78 => X"000000b5000000000000006b0000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000008b00000000",
            INIT_7A => X"0000008500000000000000130000000000000017000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000043000000000000008700000000",
            INIT_7C => X"0000000300000000000000000000000000000000000000000000001e00000000",
            INIT_7D => X"0000000000000000000000000000000000000001000000000000000300000000",
            INIT_7E => X"0000003500000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000330000000000000000000000000000006500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE2;


    MEM_GOLD_LAYER0_INSTANCE3 : if BRAM_NAME = "gold_layer0_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000001a00000000000000040000000000000000000000000000000000000000",
            INIT_02 => X"0000007200000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"000000000000000000000000000000000000001d000000000000004f00000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"000000170000000000000048000000000000000b000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000002300000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000024000000000000001400000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000003100000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"00000000000000000000001e0000000000000000000000000000001600000000",
            INIT_18 => X"0000003c0000000000000000000000000000000f000000000000001a00000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_1A => X"000000230000000000000017000000000000000d000000000000000000000000",
            INIT_1B => X"0000001000000000000000130000000000000005000000000000000000000000",
            INIT_1C => X"0000002c00000000000000180000000000000000000000000000002700000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"00000000000000000000004d0000000000000000000000000000002f00000000",
            INIT_1F => X"000000190000000000000000000000000000000e000000000000001900000000",
            INIT_20 => X"00000000000000000000007a0000000000000007000000000000001400000000",
            INIT_21 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"000000260000000000000000000000000000002e000000000000000d00000000",
            INIT_23 => X"0000000600000000000000100000000000000011000000000000002300000000",
            INIT_24 => X"0000000000000000000000000000000000000058000000000000002200000000",
            INIT_25 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_26 => X"0000002500000000000000200000000000000000000000000000000000000000",
            INIT_27 => X"0000005400000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"00000000000000000000000d0000000000000053000000000000004400000000",
            INIT_29 => X"0000000000000000000000270000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_2B => X"0000003800000000000000380000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000100000000000000029000000000000007900000000",
            INIT_2D => X"0000000000000000000000010000000000000049000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000004000000000000001300000000",
            INIT_2F => X"0000006700000000000000240000000000000044000000000000000000000000",
            INIT_30 => X"00000031000000000000004000000000000000a6000000000000000000000000",
            INIT_31 => X"000000560000000000000041000000000000004b000000000000003d00000000",
            INIT_32 => X"0000005000000000000000500000000000000079000000000000007300000000",
            INIT_33 => X"0000002600000000000000200000000000000043000000000000006a00000000",
            INIT_34 => X"0000007f00000000000000840000000000000081000000000000008d00000000",
            INIT_35 => X"000000ba00000000000000b10000000000000098000000000000009b00000000",
            INIT_36 => X"000000f900000000000000cc00000000000000cc00000000000000cc00000000",
            INIT_37 => X"0000007e00000000000000780000000000000000000000000000006900000000",
            INIT_38 => X"000000af00000000000000a800000000000000af00000000000000ae00000000",
            INIT_39 => X"000000cf00000000000000d300000000000000cd00000000000000ba00000000",
            INIT_3A => X"000000db000000000000010400000000000000e100000000000000ca00000000",
            INIT_3B => X"000000ac000000000000009600000000000000bf000000000000002200000000",
            INIT_3C => X"000000c200000000000000b000000000000000ae00000000000000bf00000000",
            INIT_3D => X"000000f200000000000000e700000000000000db00000000000000da00000000",
            INIT_3E => X"000000cd00000000000000f1000000000000010200000000000000fc00000000",
            INIT_3F => X"000000a600000000000000a600000000000000a6000000000000009100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d600000000000000d200000000000000b600000000000000ab00000000",
            INIT_41 => X"00000103000000000000011300000000000000cd00000000000000c800000000",
            INIT_42 => X"000000e200000000000000e100000000000000e300000000000000d500000000",
            INIT_43 => X"000000fd00000000000000eb00000000000000d500000000000000e100000000",
            INIT_44 => X"00000095000000000000008800000000000000a900000000000000e100000000",
            INIT_45 => X"000000dd00000000000000c400000000000000c700000000000000ae00000000",
            INIT_46 => X"000000df00000000000000ea00000000000000ee00000000000000f200000000",
            INIT_47 => X"0000008100000000000000b500000000000000c000000000000000e800000000",
            INIT_48 => X"0000004c00000000000000300000000000000027000000000000003d00000000",
            INIT_49 => X"00000090000000000000008400000000000000b4000000000000008400000000",
            INIT_4A => X"000000d600000000000000f300000000000000f200000000000000ea00000000",
            INIT_4B => X"0000003b00000000000000170000000000000033000000000000006f00000000",
            INIT_4C => X"0000002f000000000000002c0000000000000010000000000000001c00000000",
            INIT_4D => X"000000ce0000000000000066000000000000002f000000000000009600000000",
            INIT_4E => X"0000005a000000000000006e00000000000000c100000000000000e600000000",
            INIT_4F => X"0000003a000000000000002a000000000000001c000000000000001c00000000",
            INIT_50 => X"0000006800000000000000190000000000000012000000000000002f00000000",
            INIT_51 => X"0000007f00000000000000a7000000000000005d000000000000000000000000",
            INIT_52 => X"0000002200000000000000400000000000000067000000000000006e00000000",
            INIT_53 => X"0000002700000000000000370000000000000025000000000000002200000000",
            INIT_54 => X"00000000000000000000003a0000000000000018000000000000002200000000",
            INIT_55 => X"0000005100000000000000d40000000000000093000000000000002b00000000",
            INIT_56 => X"00000032000000000000002f000000000000005d000000000000003500000000",
            INIT_57 => X"000000160000000000000004000000000000002c000000000000003d00000000",
            INIT_58 => X"0000004c00000000000000000000000000000016000000000000000f00000000",
            INIT_59 => X"00000054000000000000008e00000000000000b7000000000000004800000000",
            INIT_5A => X"000000550000000000000019000000000000002d000000000000003d00000000",
            INIT_5B => X"00000015000000000000001b0000000000000010000000000000000f00000000",
            INIT_5C => X"00000008000000000000000e0000000000000000000000000000002800000000",
            INIT_5D => X"000000220000000000000042000000000000006b000000000000005900000000",
            INIT_5E => X"000000320000000000000082000000000000001d000000000000002a00000000",
            INIT_5F => X"000000680000000000000034000000000000000d000000000000001500000000",
            INIT_60 => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"00000037000000000000002d0000000000000033000000000000003f00000000",
            INIT_62 => X"0000000e00000000000000260000000000000083000000000000001200000000",
            INIT_63 => X"0000001600000000000000b90000000000000068000000000000002500000000",
            INIT_64 => X"0000000000000000000000200000000000000000000000000000000d00000000",
            INIT_65 => X"00000021000000000000003d000000000000001b000000000000001b00000000",
            INIT_66 => X"000000250000000000000000000000000000000d000000000000001400000000",
            INIT_67 => X"0000000b000000000000000500000000000000a200000000000000a300000000",
            INIT_68 => X"00000000000000000000001e0000000000000012000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000006a00000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000003b00000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000006700000000000000760000000000000066000000000000000000000000",
            INIT_7B => X"0000007300000000000000610000000000000064000000000000006300000000",
            INIT_7C => X"000000680000000000000070000000000000007e000000000000008f00000000",
            INIT_7D => X"0000005b000000000000004e000000000000004d000000000000006500000000",
            INIT_7E => X"0000006e00000000000000740000000000000075000000000000006200000000",
            INIT_7F => X"0000007500000000000000220000000000000000000000000000006600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE3;


    MEM_GOLD_LAYER0_INSTANCE4 : if BRAM_NAME = "gold_layer0_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000009300000000",
            INIT_01 => X"0000006f00000000000000470000000000000050000000000000001400000000",
            INIT_02 => X"0000008000000000000000790000000000000070000000000000009a00000000",
            INIT_03 => X"00000000000000000000000c000000000000003400000000000000c200000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"000000000000000000000000000000000000003b000000000000000000000000",
            INIT_06 => X"00000004000000000000004b0000000000000077000000000000004b00000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000003d00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000002900000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000006d00000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000005200000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000002e000000000000004a0000000000000007000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_1A => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_1F => X"00000000000000000000003e0000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000002400000000000000230000000000000000000000000000000000000000",
            INIT_33 => X"0000001c00000000000000230000000000000024000000000000001900000000",
            INIT_34 => X"0000002c00000000000000250000000000000024000000000000002100000000",
            INIT_35 => X"0000001a00000000000000120000000000000011000000000000001800000000",
            INIT_36 => X"0000001c00000000000000260000000000000026000000000000002a00000000",
            INIT_37 => X"000000020000000000000050000000000000001e000000000000002800000000",
            INIT_38 => X"00000028000000000000001c0000000000000015000000000000001d00000000",
            INIT_39 => X"0000002e00000000000000270000000000000013000000000000001c00000000",
            INIT_3A => X"0000002800000000000000270000000000000026000000000000002f00000000",
            INIT_3B => X"00000011000000000000000f0000000000000060000000000000002d00000000",
            INIT_3C => X"000000000000000000000014000000000000002c000000000000000200000000",
            INIT_3D => X"0000004900000000000000380000000000000016000000000000002800000000",
            INIT_3E => X"0000002b00000000000000230000000000000035000000000000002e00000000",
            INIT_3F => X"0000001d00000000000000000000000000000042000000000000000600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000019000000000000000f000000000000000a000000000000000d00000000",
            INIT_41 => X"000000560000000000000000000000000000002d000000000000001c00000000",
            INIT_42 => X"0000000000000000000000350000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000290000000000000000000000000000000000000000",
            INIT_44 => X"0000002a00000000000000260000000000000000000000000000001800000000",
            INIT_45 => X"0000000000000000000000340000000000000000000000000000000000000000",
            INIT_46 => X"0000002800000000000000000000000000000049000000000000000000000000",
            INIT_47 => X"00000000000000000000000d000000000000004b000000000000000700000000",
            INIT_48 => X"000000000000000000000011000000000000001f000000000000000000000000",
            INIT_49 => X"000000420000000000000000000000000000006d000000000000000000000000",
            INIT_4A => X"0000000000000000000000440000000000000000000000000000004e00000000",
            INIT_4B => X"0000000300000000000000000000000000000044000000000000003600000000",
            INIT_4C => X"0000000000000000000000110000000000000025000000000000001100000000",
            INIT_4D => X"0000000d000000000000004b0000000000000000000000000000002b00000000",
            INIT_4E => X"0000001b00000000000000040000000000000000000000000000004000000000",
            INIT_4F => X"0000001100000000000000150000000000000009000000000000003800000000",
            INIT_50 => X"0000000100000000000000000000000000000000000000000000001a00000000",
            INIT_51 => X"0000000000000000000000000000000000000034000000000000000000000000",
            INIT_52 => X"0000003300000000000000070000000000000048000000000000001800000000",
            INIT_53 => X"0000002f00000000000000150000000000000000000000000000005300000000",
            INIT_54 => X"0000001200000000000000000000000000000000000000000000002900000000",
            INIT_55 => X"0000000000000000000000000000000000000009000000000000001900000000",
            INIT_56 => X"0000000a00000000000000030000000000000000000000000000006300000000",
            INIT_57 => X"0000001900000000000000340000000000000031000000000000001300000000",
            INIT_58 => X"0000000000000000000000170000000000000000000000000000006600000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000001700000000000000220000000000000000000000000000000000000000",
            INIT_5B => X"000000430000000000000034000000000000003d000000000000000b00000000",
            INIT_5C => X"0000002e00000000000000400000000000000000000000000000000000000000",
            INIT_5D => X"0000001a0000000000000016000000000000001d000000000000000000000000",
            INIT_5E => X"000000270000000000000023000000000000002b000000000000002300000000",
            INIT_5F => X"0000001a0000000000000027000000000000001d000000000000002300000000",
            INIT_60 => X"0000001200000000000000000000000000000068000000000000000000000000",
            INIT_61 => X"000000280000000000000025000000000000001a000000000000001900000000",
            INIT_62 => X"0000001400000000000000210000000000000023000000000000002800000000",
            INIT_63 => X"00000000000000000000001f0000000000000025000000000000001800000000",
            INIT_64 => X"0000001a0000000000000014000000000000000c000000000000008b00000000",
            INIT_65 => X"0000002000000000000000170000000000000014000000000000001d00000000",
            INIT_66 => X"0000003d00000000000000280000000000000021000000000000003100000000",
            INIT_67 => X"0000007300000000000000190000000000000023000000000000001800000000",
            INIT_68 => X"000000100000000000000023000000000000002c000000000000002f00000000",
            INIT_69 => X"0000001800000000000000260000000000000022000000000000001800000000",
            INIT_6A => X"0000004e0000000000000028000000000000003b000000000000001d00000000",
            INIT_6B => X"0000004d0000000000000052000000000000004f000000000000005900000000",
            INIT_6C => X"0000004b0000000000000056000000000000005a000000000000005400000000",
            INIT_6D => X"0000003d00000000000000410000000000000045000000000000004e00000000",
            INIT_6E => X"0000005600000000000000490000000000000033000000000000003f00000000",
            INIT_6F => X"00000082000000000000004b0000000000000059000000000000005300000000",
            INIT_70 => X"0000001d000000000000003c0000000000000060000000000000005900000000",
            INIT_71 => X"00000037000000000000002e000000000000002a000000000000002900000000",
            INIT_72 => X"00000057000000000000003c0000000000000063000000000000003d00000000",
            INIT_73 => X"0000003e00000000000000910000000000000056000000000000005400000000",
            INIT_74 => X"00000054000000000000003f0000000000000000000000000000000d00000000",
            INIT_75 => X"0000003f00000000000000180000000000000029000000000000002100000000",
            INIT_76 => X"00000054000000000000005d0000000000000029000000000000003900000000",
            INIT_77 => X"00000019000000000000005a0000000000000021000000000000006200000000",
            INIT_78 => X"0000003b00000000000000570000000000000046000000000000001d00000000",
            INIT_79 => X"0000003300000000000000250000000000000003000000000000001300000000",
            INIT_7A => X"000000ac00000000000000210000000000000059000000000000008c00000000",
            INIT_7B => X"00000024000000000000002d0000000000000071000000000000006200000000",
            INIT_7C => X"0000002100000000000000330000000000000062000000000000000000000000",
            INIT_7D => X"000000a900000000000000400000000000000004000000000000000800000000",
            INIT_7E => X"0000006400000000000000bb0000000000000055000000000000006000000000",
            INIT_7F => X"00000046000000000000002e000000000000003b000000000000009300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE4;


    MEM_GOLD_LAYER0_INSTANCE5 : if BRAM_NAME = "gold_layer0_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001200000000000000290000000000000026000000000000008a00000000",
            INIT_01 => X"0000005300000000000000ca0000000000000023000000000000000000000000",
            INIT_02 => X"000000c60000000000000074000000000000006d000000000000004c00000000",
            INIT_03 => X"0000006c000000000000007e0000000000000041000000000000005500000000",
            INIT_04 => X"0000002a0000000000000027000000000000001a000000000000002c00000000",
            INIT_05 => X"00000054000000000000002e0000000000000090000000000000005f00000000",
            INIT_06 => X"00000060000000000000007b00000000000000cb000000000000002f00000000",
            INIT_07 => X"000000350000000000000066000000000000007a000000000000003100000000",
            INIT_08 => X"0000008d000000000000001e000000000000004b000000000000002100000000",
            INIT_09 => X"000000470000000000000067000000000000004b00000000000000a800000000",
            INIT_0A => X"0000002a000000000000004e0000000000000042000000000000004600000000",
            INIT_0B => X"0000000900000000000000170000000000000069000000000000005700000000",
            INIT_0C => X"0000009f00000000000000a00000000000000050000000000000002800000000",
            INIT_0D => X"00000012000000000000006a0000000000000053000000000000007000000000",
            INIT_0E => X"0000004d00000000000000480000000000000087000000000000002300000000",
            INIT_0F => X"0000005d00000000000000200000000000000000000000000000001a00000000",
            INIT_10 => X"00000073000000000000009b00000000000000b3000000000000005200000000",
            INIT_11 => X"00000094000000000000005e0000000000000096000000000000006f00000000",
            INIT_12 => X"000000000000000000000000000000000000004800000000000000a100000000",
            INIT_13 => X"00000030000000000000003e000000000000001e000000000000000000000000",
            INIT_14 => X"000000fb00000000000000640000000000000089000000000000008400000000",
            INIT_15 => X"000000280000000000000033000000000000002d00000000000000fb00000000",
            INIT_16 => X"000000150000000000000016000000000000000a000000000000001500000000",
            INIT_17 => X"00000020000000000000001d0000000000000025000000000000001a00000000",
            INIT_18 => X"00000026000000000000012e000000000000004e000000000000006000000000",
            INIT_19 => X"0000000900000000000000100000000000000018000000000000001500000000",
            INIT_1A => X"00000030000000000000001e000000000000000c000000000000000800000000",
            INIT_1B => X"0000001900000000000000170000000000000021000000000000001e00000000",
            INIT_1C => X"00000017000000000000001600000000000000dd000000000000006500000000",
            INIT_1D => X"00000015000000000000000d0000000000000014000000000000001400000000",
            INIT_1E => X"0000002600000000000000110000000000000026000000000000001b00000000",
            INIT_1F => X"0000002a00000000000000160000000000000021000000000000005700000000",
            INIT_20 => X"0000001b0000000000000015000000000000000d000000000000004800000000",
            INIT_21 => X"0000001e00000000000000210000000000000018000000000000000f00000000",
            INIT_22 => X"000000100000000000000051000000000000001b000000000000000700000000",
            INIT_23 => X"0000000300000000000000080000000000000007000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_26 => X"0000000a00000000000000010000000000000000000000000000000000000000",
            INIT_27 => X"000000080000000000000000000000000000000b000000000000001a00000000",
            INIT_28 => X"000000000000000000000021000000000000000000000000000000ac00000000",
            INIT_29 => X"00000000000000000000000e0000000000000020000000000000001e00000000",
            INIT_2A => X"000000000000000000000015000000000000000c000000000000000000000000",
            INIT_2B => X"00000000000000000000000e0000000000000000000000000000000b00000000",
            INIT_2C => X"0000005a000000000000001f0000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000a30000000000000000000000000000001e00000000",
            INIT_2F => X"0000004200000000000000000000000000000035000000000000001400000000",
            INIT_30 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_31 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"000000040000000000000000000000000000008e000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000008500000000",
            INIT_34 => X"0000000000000000000000000000000000000035000000000000000000000000",
            INIT_35 => X"0000000000000000000000110000000000000000000000000000001600000000",
            INIT_36 => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000012c00000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"00000069000000000000003c0000000000000000000000000000000000000000",
            INIT_3B => X"000000cc00000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000830000000000000011000000000000000000000000",
            INIT_3F => X"0000000000000000000000700000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_41 => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000003e00000000000000000000000000000000000000000000000d00000000",
            INIT_43 => X"0000000000000000000000270000000000000000000000000000000000000000",
            INIT_44 => X"00000000000000000000003f0000000000000008000000000000000000000000",
            INIT_45 => X"0000000000000000000000200000000000000000000000000000000000000000",
            INIT_46 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_47 => X"0000004a00000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000470000000000000000000000000000005500000000",
            INIT_49 => X"0000003d000000000000000000000000000000eb000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000006100000000",
            INIT_4B => X"000000000000000000000025000000000000005f000000000000002e00000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"000000000000000000000000000000000000000000000000000000ba00000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000025000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_62 => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000005400000000",
            INIT_64 => X"000000000000000000000000000000000000000000000000000000c500000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000002f00000000",
            INIT_66 => X"000000000000000000000000000000000000002d000000000000001300000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"000000af00000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"00000000000000000000000f0000000000000000000000000000009200000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000003b00000000",
            INIT_6C => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"000000000000000000000000000000000000002d000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000015a00000000",
            INIT_70 => X"0000000000000000000000000000000000000092000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000003600000000",
            INIT_72 => X"000000d700000000000000000000000000000004000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000059000000000000000000000000",
            INIT_74 => X"000000000000000000000000000000000000000000000000000000be00000000",
            INIT_75 => X"0000001900000000000000000000000000000000000000000000000400000000",
            INIT_76 => X"000000d4000000000000003e0000000000000000000000000000000000000000",
            INIT_77 => X"0000008700000000000000000000000000000007000000000000000000000000",
            INIT_78 => X"0000000700000000000000360000000000000000000000000000000000000000",
            INIT_79 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_7A => X"00000011000000000000005f0000000000000000000000000000006100000000",
            INIT_7B => X"000000b60000000000000000000000000000002d000000000000000000000000",
            INIT_7C => X"000000000000000000000043000000000000001d000000000000000000000000",
            INIT_7D => X"0000004d00000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"000000220000000000000000000000000000002a000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE5;


    MEM_GOLD_LAYER0_INSTANCE6 : if BRAM_NAME = "gold_layer0_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b400000000000000000000000000000002000000000000004400000000",
            INIT_01 => X"0000000000000000000000850000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000003a00000000000001000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000051000000000000000000000000",
            INIT_06 => X"000000000000000000000007000000000000003d000000000000003c00000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"00000000000000000000008b0000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000004300000000000000820000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000001000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000030000000000000003200000000",
            INIT_12 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000009000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000009200000000000000970000000000000093000000000000008b00000000",
            INIT_4D => X"0000009b00000000000000ab000000000000009c000000000000008300000000",
            INIT_4E => X"000000710000000000000066000000000000005a000000000000007400000000",
            INIT_4F => X"00000099000000000000009a000000000000007f000000000000007900000000",
            INIT_50 => X"00000066000000000000009e0000000000000098000000000000009a00000000",
            INIT_51 => X"0000002a0000000000000039000000000000006e000000000000007600000000",
            INIT_52 => X"0000006e00000000000000200000000000000000000000000000000000000000",
            INIT_53 => X"000000a1000000000000007c0000000000000037000000000000007d00000000",
            INIT_54 => X"00000039000000000000004d000000000000009f00000000000000a000000000",
            INIT_55 => X"0000000000000000000000000000000000000022000000000000001500000000",
            INIT_56 => X"0000006200000000000000260000000000000000000000000000000000000000",
            INIT_57 => X"0000009f00000000000000910000000000000032000000000000000000000000",
            INIT_58 => X"000000000000000000000014000000000000005a000000000000006600000000",
            INIT_59 => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_5A => X"0000000000000000000000460000000000000000000000000000000000000000",
            INIT_5B => X"00000017000000000000009f0000000000000069000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_5E => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_5F => X"000000120000000000000006000000000000002f000000000000006e00000000",
            INIT_60 => X"0000002c00000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000005e00000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000250000000000000000000000000000006200000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_66 => X"0000003700000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000011000000000000003600000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_69 => X"0000000000000000000000470000000000000000000000000000000000000000",
            INIT_6A => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000002000000000000000000000000000000012000000000000000000000000",
            INIT_6C => X"000000000000000000000000000000000000002f000000000000000000000000",
            INIT_6D => X"000000000000000000000000000000000000005e000000000000003700000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000001a00000000000000000000000000000000000000000000000e00000000",
            INIT_70 => X"0000004b00000000000000020000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000006a00000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE6;


    MEM_GOLD_LAYER0_INSTANCE7 : if BRAM_NAME = "gold_layer0_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE7;


    MEM_GOLD_LAYER1_INSTANCE0 : if BRAM_NAME = "gold_layer1_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000019700000000000000550000000000000000000000000000011600000000",
            INIT_02 => X"00000000000000000000005200000000000000b7000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"000000f20000000000000026000000000000004700000000000000cc00000000",
            INIT_05 => X"0000000000000000000000170000000000000000000000000000002700000000",
            INIT_06 => X"0000002400000000000000000000000000000000000000000000005e00000000",
            INIT_07 => X"00000000000000000000006b000000000000007f000000000000000000000000",
            INIT_08 => X"00000000000000000000000000000000000001c4000000000000000000000000",
            INIT_09 => X"000000370000000000000059000000000000017d000000000000000000000000",
            INIT_0A => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"00000000000000000000009b0000000000000090000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000018000000000000001f00000000",
            INIT_12 => X"000000840000000000000000000000000000000f000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000d20000000000000000000000000000000000000000",
            INIT_15 => X"000001a900000000000000000000000000000000000000000000007400000000",
            INIT_16 => X"000000000000000000000018000000000000000500000000000000cc00000000",
            INIT_17 => X"0000001500000000000000270000000000000046000000000000023300000000",
            INIT_18 => X"0000000000000000000000000000000000000003000000000000001200000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000500000000000000000000000000000000000000000",
            INIT_21 => X"0000013200000000000000000000000000000087000000000000000000000000",
            INIT_22 => X"000000a300000000000000f5000000000000008800000000000000fb00000000",
            INIT_23 => X"000000f5000000000000015e000000000000013d000000000000000000000000",
            INIT_24 => X"000000db00000000000000b500000000000000d300000000000000da00000000",
            INIT_25 => X"000000000000000000000000000000000000003f000000000000015000000000",
            INIT_26 => X"0000001f0000000000000000000000000000006d000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000007500000000000000100000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000650000000000000000000000000000000000000000",
            INIT_2D => X"00000000000000000000000000000000000000ad000000000000000000000000",
            INIT_2E => X"000000b900000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"00000000000000000000002d0000000000000067000000000000001b00000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000c10000000000000000000000000000000000000000",
            INIT_34 => X"000000000000000000000000000000000000011b000000000000000000000000",
            INIT_35 => X"000000da00000000000000000000000000000053000000000000000000000000",
            INIT_36 => X"000000000000000000000058000000000000001b000000000000002e00000000",
            INIT_37 => X"0000000000000000000000aa0000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000052000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000001090000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000210000000000000000000000000000014300000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000040000000000000000000000000000002600000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"00000000000000000000000a0000000000000000000000000000000900000000",
            INIT_43 => X"0000001e0000000000000000000000000000002e000000000000000000000000",
            INIT_44 => X"0000000000000000000000390000000000000000000000000000002b00000000",
            INIT_45 => X"000000000000000000000000000000000000018b000000000000000000000000",
            INIT_46 => X"0000009e000000000000009b0000000000000000000000000000003900000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000010000000000000000000000000000011900000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"000001e4000000000000021c0000000000000258000000000000005300000000",
            INIT_4B => X"00000083000000000000000000000000000000a7000000000000011c00000000",
            INIT_4C => X"0000007f00000000000000000000000000000000000000000000001000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000057000000000000000000000000",
            INIT_4F => X"000000000000000000000056000000000000007c00000000000000d900000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000008300000000",
            INIT_51 => X"0000011c00000000000001150000000000000026000000000000003b00000000",
            INIT_52 => X"0000020f000000000000001b0000000000000007000000000000000000000000",
            INIT_53 => X"000000000000000000000000000000000000000b00000000000000a200000000",
            INIT_54 => X"00000000000000000000000800000000000000f7000000000000002200000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000780000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000042000000000000000000000000",
            INIT_5A => X"000000120000000000000000000000000000006e000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000570000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000bd0000000000000019000000000000004200000000",
            INIT_5E => X"000001bb00000000000000000000000000000042000000000000000400000000",
            INIT_5F => X"0000000100000000000000200000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000004900000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000004200000000000000290000000000000000000000000000000f00000000",
            INIT_63 => X"0000004f00000000000000000000000000000097000000000000000a00000000",
            INIT_64 => X"0000000000000000000000e10000000000000112000000000000000000000000",
            INIT_65 => X"0000000000000000000000390000000000000014000000000000000000000000",
            INIT_66 => X"0000000000000000000000a20000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000061000000000000000000000000",
            INIT_69 => X"000000ee000000000000007400000000000000cc000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000007300000000",
            INIT_6B => X"0000000000000000000000000000000000000111000000000000018700000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000150000000000000054000000000000006300000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000009100000000",
            INIT_72 => X"0000025b00000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000d80000000000000000000000000000000000000000",
            INIT_75 => X"0000000200000000000001a20000000000000000000000000000000000000000",
            INIT_76 => X"0000007100000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"000000000000000000000000000000000000008f000000000000000000000000",
            INIT_78 => X"000000000000000000000000000000000000003c000000000000002000000000",
            INIT_79 => X"0000000000000000000000000000000000000094000000000000000000000000",
            INIT_7A => X"0000002f00000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"000000e0000000000000014500000000000001de000000000000012700000000",
            INIT_7C => X"0000009900000000000000a6000000000000007c000000000000002f00000000",
            INIT_7D => X"00000000000000000000009b0000000000000000000000000000011600000000",
            INIT_7E => X"0000003000000000000000000000000000000000000000000000005900000000",
            INIT_7F => X"0000007c0000000000000000000000000000005f000000000000002700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE0;


    MEM_GOLD_LAYER1_INSTANCE1 : if BRAM_NAME = "gold_layer1_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000006e0000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000003100000000000000d100000000000000e5000000000000002e00000000",
            INIT_03 => X"0000007600000000000001e90000000000000000000000000000009700000000",
            INIT_04 => X"0000009c00000000000000cc00000000000000dc00000000000000f900000000",
            INIT_05 => X"00000000000000000000005f000000000000003c000000000000000000000000",
            INIT_06 => X"0000004700000000000000f20000000000000002000000000000002c00000000",
            INIT_07 => X"00000000000000000000006a0000000000000036000000000000006900000000",
            INIT_08 => X"00000054000000000000009f00000000000000e4000000000000009f00000000",
            INIT_09 => X"000000000000000000000036000000000000000d000000000000000000000000",
            INIT_0A => X"0000009000000000000000f400000000000000aa000000000000000000000000",
            INIT_0B => X"0000008500000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000002200000000000000a300000000000000d4000000000000006a00000000",
            INIT_0D => X"0000000000000000000000ad000000000000000000000000000000e500000000",
            INIT_0E => X"000000e200000000000000fb0000000000000162000000000000000000000000",
            INIT_0F => X"0000004f00000000000000c900000000000000b4000000000000003c00000000",
            INIT_10 => X"00000067000000000000007b00000000000000f8000000000000000000000000",
            INIT_11 => X"00000000000000000000008e0000000000000031000000000000003900000000",
            INIT_12 => X"0000000000000000000000000000000000000004000000000000000500000000",
            INIT_13 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000680000000000000109000000000000004300000000",
            INIT_15 => X"0000000000000000000000e30000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000aa0000000000000000000000000000009b00000000",
            INIT_17 => X"000000da000000000000000000000000000001b1000000000000000000000000",
            INIT_18 => X"00000000000000000000005f0000000000000125000000000000004e00000000",
            INIT_19 => X"00000000000000000000008b0000000000000000000000000000011800000000",
            INIT_1A => X"000000d60000000000000000000000000000008a00000000000000a900000000",
            INIT_1B => X"0000000000000000000000000000000000000036000000000000004c00000000",
            INIT_1C => X"000000e2000000000000000000000000000001f5000000000000000000000000",
            INIT_1D => X"0000009a00000000000000000000000000000021000000000000000000000000",
            INIT_1E => X"00000008000000000000001a000000000000003b000000000000004e00000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"00000000000000000000001d0000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000860000000000000000000000000000015400000000",
            INIT_2D => X"00000000000000000000004b000000000000001a000000000000002b00000000",
            INIT_2E => X"000000000000000000000000000000000000007e000000000000000000000000",
            INIT_2F => X"00000000000000000000001d000000000000000000000000000001c300000000",
            INIT_30 => X"0000013b000000000000009d000000000000000000000000000000ac00000000",
            INIT_31 => X"000000f9000000000000004c0000000000000187000000000000014400000000",
            INIT_32 => X"00000000000000000000007600000000000000a8000000000000000000000000",
            INIT_33 => X"00000000000000000000002c0000000000000148000000000000000000000000",
            INIT_34 => X"000000000000000000000240000000000000003200000000000000a800000000",
            INIT_35 => X"000000000000000000000022000000000000002f000000000000000000000000",
            INIT_36 => X"0000000c000000000000002000000000000002fb000000000000000000000000",
            INIT_37 => X"0000000000000000000000600000000000000036000000000000002000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000006e0000000000000058000000000000002b000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000007e000000000000004f00000000000000e2000000000000005300000000",
            INIT_3D => X"0000001f00000000000000000000000000000099000000000000006b00000000",
            INIT_3E => X"0000009800000000000000170000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000005800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000010200000000000000c80000000000000000000000000000000000000000",
            INIT_42 => X"00000047000000000000002d000000000000000000000000000000fe00000000",
            INIT_43 => X"000000b40000000000000103000000000000012d00000000000000a500000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000004f00000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"000000000000000000000121000000000000008e000000000000004800000000",
            INIT_48 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_4A => X"0000015100000000000000000000000000000000000000000000007100000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000006a000000000000007700000000000000ca000000000000000000000000",
            INIT_4E => X"0000000000000000000000f0000000000000007a000000000000000000000000",
            INIT_4F => X"00000060000000000000001d0000000000000031000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000007300000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000003500000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"000000000000000000000000000000000000006f000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000af0000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000670000000000000000000000000000000000000000",
            INIT_72 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000115000000000000004f00000000",
            INIT_74 => X"000000c700000000000000b10000000000000086000000000000008900000000",
            INIT_75 => X"0000010d0000000000000080000000000000001a000000000000007900000000",
            INIT_76 => X"0000003b000000000000007e000000000000003200000000000000a200000000",
            INIT_77 => X"00000000000000000000000000000000000000b3000000000000011700000000",
            INIT_78 => X"000000000000000000000000000000000000005d000000000000002800000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000930000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000007b00000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_7D => X"0000000000000000000000f90000000000000043000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE1;


    MEM_GOLD_LAYER1_INSTANCE2 : if BRAM_NAME = "gold_layer1_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000420000000000000000000000000000000000000000",
            INIT_02 => X"0000007900000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"000000000000000000000000000000000000002a000000000000007300000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000008600000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"000000bc00000000000000e600000000000000e6000000000000015100000000",
            INIT_18 => X"000000000000000000000000000000000000000000000000000000d500000000",
            INIT_19 => X"0000000000000000000000bd00000000000000a600000000000000b000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"000000380000000000000000000000000000006f000000000000000000000000",
            INIT_1D => X"000000c500000000000001080000000000000000000000000000004600000000",
            INIT_1E => X"0000000000000000000000330000000000000000000000000000001400000000",
            INIT_1F => X"00000020000000000000008e0000000000000000000000000000000000000000",
            INIT_20 => X"000000000000000000000066000000000000007e000000000000003900000000",
            INIT_21 => X"0000007300000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000003200000000000000c70000000000000000000000000000000000000000",
            INIT_23 => X"000000000000000000000000000000000000007b000000000000001a00000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000c90000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000008200000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000004000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000014b00000000000000310000000000000000000000000000000000000000",
            INIT_30 => X"00000000000000000000001200000000000000b100000000000000a000000000",
            INIT_31 => X"0000007300000000000000bf0000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000029000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000005200000000",
            INIT_39 => X"00000000000000000000000000000000000000b7000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"000000000000000000000000000000000000000000000000000000eb00000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000028000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000005000000000",
            INIT_43 => X"0000009500000000000000000000000000000000000000000000000f00000000",
            INIT_44 => X"0000004600000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000001000000000000000150000000000000000000000000000000000000000",
            INIT_46 => X"00000000000000000000007300000000000000a4000000000000000000000000",
            INIT_47 => X"0000000000000000000001810000000000000153000000000000000000000000",
            INIT_48 => X"0000014a00000000000001450000000000000115000000000000018300000000",
            INIT_49 => X"0000009700000000000000d0000000000000011b00000000000001c500000000",
            INIT_4A => X"00000108000000000000012f00000000000000de00000000000000c100000000",
            INIT_4B => X"0000000000000000000000a00000000000000000000000000000000000000000",
            INIT_4C => X"00000099000000000000000c00000000000001b1000000000000000800000000",
            INIT_4D => X"0000000000000000000000fb0000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000004000000000",
            INIT_4F => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_50 => X"00000000000000000000002e00000000000000b9000000000000000000000000",
            INIT_51 => X"00000000000000000000008f0000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"00000000000000000000011b00000000000000ef000000000000003e00000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000018000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"00000137000000000000021100000000000001db000000000000010f00000000",
            INIT_58 => X"0000000000000000000000380000000000000000000000000000003c00000000",
            INIT_59 => X"0000000900000000000000000000000000000000000000000000014a00000000",
            INIT_5A => X"0000012800000000000000000000000000000000000000000000005a00000000",
            INIT_5B => X"000000c2000000000000007d0000000000000067000000000000000000000000",
            INIT_5C => X"0000015100000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000400000000000000db00000000000000e9000000000000008800000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"000000cb00000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000009400000000000000300000000000000000000000000000000000000000",
            INIT_66 => X"000000000000000000000000000000000000001f000000000000000000000000",
            INIT_67 => X"0000007700000000000000e70000000000000023000000000000017c00000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000002e00000000",
            INIT_69 => X"000000b3000000000000007c0000000000000000000000000000003d00000000",
            INIT_6A => X"0000005300000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000005300000000",
            INIT_6C => X"0000000000000000000001080000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000067000000000000000000000000",
            INIT_6F => X"000000e7000000000000005d0000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000500000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000003100000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"000000000000000000000000000000000000002f000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000003000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"00000071000000000000005c00000000000000b0000000000000001200000000",
            INIT_7D => X"0000007b000000000000002c0000000000000000000000000000005000000000",
            INIT_7E => X"000000000000000000000008000000000000007a000000000000004e00000000",
            INIT_7F => X"0000000000000000000000660000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE2;


    MEM_GOLD_LAYER1_INSTANCE3 : if BRAM_NAME = "gold_layer1_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003700000000000000000000000000000089000000000000000700000000",
            INIT_01 => X"00000024000000000000000000000000000000aa000000000000008600000000",
            INIT_02 => X"00000010000000000000004d0000000000000002000000000000004300000000",
            INIT_03 => X"00000034000000000000006200000000000000a000000000000000d000000000",
            INIT_04 => X"0000008200000000000000000000000000000000000000000000002a00000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE3;


    MEM_GOLD_LAYER2_INSTANCE0 : if BRAM_NAME = "gold_layer2_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000dd0000000000000000000000000000000000000000",
            INIT_06 => X"0000018f00000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"000000000000000000000000000000000000007b000000000000000000000000",
            INIT_0B => X"000000f900000000000000850000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000fc0000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000017f00000000000001fa0000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_13 => X"0000000000000000000000000000000000000086000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000270000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000111000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"000002fe00000000000000810000000000000000000000000000017400000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"000000000000000000000000000000000000000000000000000000fb00000000",
            INIT_1C => X"000000000000000000000000000000000000035d000000000000000000000000",
            INIT_1D => X"00000126000000000000020600000000000002ba000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"000000000000000000000000000000000000000000000000000001f200000000",
            INIT_23 => X"0000009d00000000000003370000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"000001f500000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000a20000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"000001d400000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000007900000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000007b0000000000000000000000000000030d000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000010e00000000000000000000000000000108000000000000000000000000",
            INIT_2F => X"000000000000000000000000000000000000000000000000000003d700000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000003600000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"000000c100000000000000cf0000000000000000000000000000010b00000000",
            INIT_37 => X"0000000000000000000000c100000000000002bd000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"000001c50000000000000170000000000000023b000000000000000000000000",
            INIT_3A => X"0000008e000000000000000000000000000001f8000000000000000000000000",
            INIT_3B => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"000000b800000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"00000382000000000000023f000000000000015a000000000000008d00000000",
            INIT_3E => X"0000000000000000000002fd000000000000036300000000000003ed00000000",
            INIT_3F => X"0000013e000000000000000000000000000001c1000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000000000000000000000000000000000002b6000000000000029100000000",
            INIT_41 => X"0000000000000000000004730000000000000205000000000000000000000000",
            INIT_42 => X"0000031900000000000002ef0000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000061000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"000000000000000000000000000000000000000000000000000000c100000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"000000eb00000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"00000000000000000000000000000000000001e900000000000003c800000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000ce00000000000000000000000000000000000000000000009900000000",
            INIT_52 => X"000000000000000000000000000000000000022300000000000002f500000000",
            INIT_53 => X"00000000000000000000028c0000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"00000000000000000000000000000000000005cf000000000000033500000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"000001ea00000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"000000000000000000000000000000000000033b000000000000021300000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"00000090000000000000019f000000000000000000000000000000eb00000000",
            INIT_5B => X"000000000000000000000000000000000000000000000000000001cb00000000",
            INIT_5C => X"0000000000000000000002ff0000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000093000000000000006700000000",
            INIT_5E => X"000000000000000000000200000000000000019e000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000015e00000000",
            INIT_60 => X"0000000000000000000000d10000000000000000000000000000000000000000",
            INIT_61 => X"000001f900000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"00000000000000000000000000000000000002dc000000000000012c00000000",
            INIT_64 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_65 => X"000000000000000000000000000000000000011e00000000000001b500000000",
            INIT_66 => X"00000000000000000000021c0000000000000178000000000000034700000000",
            INIT_67 => X"0000004400000000000000ab0000000000000000000000000000000000000000",
            INIT_68 => X"000000000000000000000000000000000000000000000000000003db00000000",
            INIT_69 => X"0000000000000000000000bb0000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000031000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000db0000000000000000000000000000017e00000000",
            INIT_6D => X"00000000000000000000034f0000000000000000000000000000009a00000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"00000145000000000000028f0000000000000026000000000000000000000000",
            INIT_70 => X"0000000000000000000000b3000000000000016a000000000000004100000000",
            INIT_71 => X"0000036900000000000001b30000000000000000000000000000000000000000",
            INIT_72 => X"000000a900000000000000000000000000000000000000000000026e00000000",
            INIT_73 => X"0000008d00000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000001740000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000027b00000000",
            INIT_76 => X"00000000000000000000000000000000000001f9000000000000002700000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000033d00000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000010e00000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"000000000000000000000000000000000000001e000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER2_INSTANCE0;


    MEM_GOLD_LAYER2_INSTANCE1 : if BRAM_NAME = "gold_layer2_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000043100000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000028400000000000000000000000000000000000000000000015700000000",
            INIT_02 => X"00000000000000000000000000000000000003e400000000000000d800000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000005a20000000000000559000000000000038300000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000011d00000000000001550000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000001670000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000007900000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"00000000000000000000036f0000000000000000000000000000000000000000",
            INIT_0C => X"000001ce000000000000019700000000000000c400000000000001ab00000000",
            INIT_0D => X"000001cc0000000000000000000000000000000000000000000001fb00000000",
            INIT_0E => X"0000030e00000000000000fa0000000000000345000000000000028b00000000",
            INIT_0F => X"000002f300000000000006ca0000000000000000000000000000043f00000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER2_INSTANCE1;


    MEM_GOLD_LAYER3_INSTANCE0 : if BRAM_NAME = "gold_layer3_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffe2bf70fffffffffff41a5dffffffffffe87547fffffffffffdee13ffffffff",
            INIT_01 => X"ffe17153ffffffffffded97affffffffffe27f99ffffffffffe9d569ffffffff",
            INIT_02 => X"fff1648cffffffffffddd902ffffffff",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER3_INSTANCE0;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE0 : if BRAM_NAME = "sampleifmap_layersamples_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a600000000000000a5000000000000009f000000000000009e00000000",
            INIT_01 => X"0000009f00000000000000a2000000000000009c00000000000000a000000000",
            INIT_02 => X"000000a000000000000000a1000000000000009f000000000000009e00000000",
            INIT_03 => X"000000aa00000000000000a900000000000000a600000000000000a100000000",
            INIT_04 => X"000000a000000000000000a000000000000000a200000000000000a700000000",
            INIT_05 => X"0000009400000000000000960000000000000095000000000000009c00000000",
            INIT_06 => X"0000008d000000000000008c000000000000008f000000000000009500000000",
            INIT_07 => X"00000074000000000000007e0000000000000089000000000000008f00000000",
            INIT_08 => X"000000a6000000000000009f0000000000000097000000000000009800000000",
            INIT_09 => X"000000a200000000000000a400000000000000a000000000000000a200000000",
            INIT_0A => X"0000009f000000000000009b000000000000009c00000000000000a300000000",
            INIT_0B => X"000000ab00000000000000ab00000000000000aa00000000000000a300000000",
            INIT_0C => X"00000097000000000000009a00000000000000a000000000000000a900000000",
            INIT_0D => X"0000008d000000000000008c000000000000008b000000000000009100000000",
            INIT_0E => X"0000008e00000000000000910000000000000093000000000000009500000000",
            INIT_0F => X"00000077000000000000007d0000000000000088000000000000008f00000000",
            INIT_10 => X"000000a7000000000000009e0000000000000097000000000000009700000000",
            INIT_11 => X"000000a500000000000000a500000000000000a300000000000000a000000000",
            INIT_12 => X"0000009d000000000000009e00000000000000a200000000000000a300000000",
            INIT_13 => X"000000a900000000000000a700000000000000a600000000000000a100000000",
            INIT_14 => X"000000790000000000000091000000000000009f00000000000000aa00000000",
            INIT_15 => X"0000007200000000000000650000000000000062000000000000006e00000000",
            INIT_16 => X"0000008c000000000000008f0000000000000086000000000000007800000000",
            INIT_17 => X"000000780000000000000082000000000000008b000000000000008e00000000",
            INIT_18 => X"000000ae00000000000000a0000000000000009b000000000000009b00000000",
            INIT_19 => X"000000a900000000000000a900000000000000a700000000000000a700000000",
            INIT_1A => X"000000bf00000000000000a700000000000000a500000000000000a500000000",
            INIT_1B => X"000000a400000000000000a2000000000000009d00000000000000b100000000",
            INIT_1C => X"0000006700000000000000680000000000000095000000000000009e00000000",
            INIT_1D => X"0000004a0000000000000050000000000000005c000000000000006200000000",
            INIT_1E => X"0000008400000000000000710000000000000053000000000000005600000000",
            INIT_1F => X"0000007f0000000000000088000000000000008c000000000000008c00000000",
            INIT_20 => X"000000aa00000000000000a1000000000000009c000000000000009b00000000",
            INIT_21 => X"000000a600000000000000a900000000000000a300000000000000a900000000",
            INIT_22 => X"000000f600000000000000ad00000000000000a400000000000000a400000000",
            INIT_23 => X"0000008e0000000000000092000000000000009700000000000000c300000000",
            INIT_24 => X"000000710000000000000055000000000000004e000000000000006f00000000",
            INIT_25 => X"0000005d0000000000000061000000000000006a000000000000007000000000",
            INIT_26 => X"0000006900000000000000550000000000000054000000000000004a00000000",
            INIT_27 => X"000000810000000000000085000000000000008a000000000000008000000000",
            INIT_28 => X"0000009300000000000000820000000000000085000000000000009400000000",
            INIT_29 => X"000000a700000000000000a700000000000000a500000000000000a100000000",
            INIT_2A => X"000000b400000000000000a300000000000000a500000000000000a300000000",
            INIT_2B => X"0000004200000000000000610000000000000080000000000000009d00000000",
            INIT_2C => X"0000007600000000000000590000000000000042000000000000004500000000",
            INIT_2D => X"0000005e00000000000000720000000000000077000000000000007a00000000",
            INIT_2E => X"00000043000000000000003a000000000000005b000000000000006300000000",
            INIT_2F => X"00000086000000000000008a000000000000008c000000000000006c00000000",
            INIT_30 => X"00000058000000000000002f000000000000006d000000000000007f00000000",
            INIT_31 => X"000000aa00000000000000a800000000000000aa000000000000009900000000",
            INIT_32 => X"0000009300000000000000a400000000000000a600000000000000a900000000",
            INIT_33 => X"000000440000000000000064000000000000007f000000000000008100000000",
            INIT_34 => X"0000008400000000000000530000000000000048000000000000004e00000000",
            INIT_35 => X"0000006b0000000000000069000000000000007c000000000000009200000000",
            INIT_36 => X"0000002e000000000000003f0000000000000055000000000000007300000000",
            INIT_37 => X"00000086000000000000008d0000000000000084000000000000004f00000000",
            INIT_38 => X"00000046000000000000002a0000000000000063000000000000008300000000",
            INIT_39 => X"000000a800000000000000a500000000000000a7000000000000008f00000000",
            INIT_3A => X"00000078000000000000008c00000000000000a100000000000000ab00000000",
            INIT_3B => X"0000005800000000000000740000000000000090000000000000008200000000",
            INIT_3C => X"0000007c000000000000004d0000000000000055000000000000005b00000000",
            INIT_3D => X"0000006a0000000000000066000000000000008800000000000000a300000000",
            INIT_3E => X"0000003100000000000000360000000000000055000000000000006400000000",
            INIT_3F => X"00000088000000000000008a000000000000006b000000000000003900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007c0000000000000036000000000000006700000000000000aa00000000",
            INIT_41 => X"000000a600000000000000a300000000000000a1000000000000009900000000",
            INIT_42 => X"0000007d000000000000007100000000000000ae00000000000000a500000000",
            INIT_43 => X"000000560000000000000079000000000000009c000000000000009d00000000",
            INIT_44 => X"0000005100000000000000500000000000000054000000000000005200000000",
            INIT_45 => X"0000005700000000000000710000000000000092000000000000008a00000000",
            INIT_46 => X"0000003800000000000000470000000000000056000000000000005300000000",
            INIT_47 => X"000000890000000000000085000000000000004a000000000000002800000000",
            INIT_48 => X"0000009a000000000000005e000000000000008600000000000000b400000000",
            INIT_49 => X"00000099000000000000009c000000000000009e00000000000000ae00000000",
            INIT_4A => X"0000009c00000000000000cf00000000000000ed00000000000000cf00000000",
            INIT_4B => X"0000005d000000000000007d000000000000009400000000000000ae00000000",
            INIT_4C => X"0000004c000000000000003b000000000000004a000000000000005600000000",
            INIT_4D => X"0000006a0000000000000085000000000000008f000000000000008900000000",
            INIT_4E => X"0000004b00000000000000540000000000000057000000000000005600000000",
            INIT_4F => X"00000084000000000000005f0000000000000028000000000000003200000000",
            INIT_50 => X"000000a5000000000000008e000000000000006c00000000000000b700000000",
            INIT_51 => X"0000007a000000000000009f000000000000009b00000000000000b100000000",
            INIT_52 => X"000000a400000000000000dc00000000000000ed00000000000000d500000000",
            INIT_53 => X"00000078000000000000007d000000000000009c00000000000000b700000000",
            INIT_54 => X"0000005b000000000000002d0000000000000050000000000000004e00000000",
            INIT_55 => X"0000006b000000000000009b000000000000009d00000000000000af00000000",
            INIT_56 => X"0000004e00000000000000580000000000000067000000000000005700000000",
            INIT_57 => X"00000068000000000000003b0000000000000029000000000000003b00000000",
            INIT_58 => X"000000aa0000000000000087000000000000006400000000000000bc00000000",
            INIT_59 => X"0000008600000000000000ad00000000000000a600000000000000bb00000000",
            INIT_5A => X"000000aa00000000000000c700000000000000c2000000000000007500000000",
            INIT_5B => X"00000075000000000000008600000000000000bd00000000000000b900000000",
            INIT_5C => X"0000007d00000000000000260000000000000054000000000000006600000000",
            INIT_5D => X"0000005d000000000000009200000000000000a000000000000000d200000000",
            INIT_5E => X"000000550000000000000068000000000000005e000000000000005300000000",
            INIT_5F => X"0000004c000000000000003e0000000000000037000000000000004900000000",
            INIT_60 => X"000000af000000000000007f000000000000005a00000000000000bd00000000",
            INIT_61 => X"0000009f00000000000000b200000000000000a600000000000000ae00000000",
            INIT_62 => X"0000008900000000000000a800000000000000a8000000000000006100000000",
            INIT_63 => X"0000007b00000000000000a000000000000000d800000000000000ba00000000",
            INIT_64 => X"0000009600000000000000320000000000000073000000000000007800000000",
            INIT_65 => X"0000005b000000000000007b000000000000009b00000000000000c200000000",
            INIT_66 => X"00000056000000000000005f0000000000000054000000000000005400000000",
            INIT_67 => X"00000049000000000000004f0000000000000049000000000000005400000000",
            INIT_68 => X"000000b90000000000000098000000000000005d00000000000000bd00000000",
            INIT_69 => X"000000a700000000000000ad0000000000000088000000000000007700000000",
            INIT_6A => X"000000a700000000000000910000000000000093000000000000006700000000",
            INIT_6B => X"0000008d00000000000000b400000000000000e200000000000000bd00000000",
            INIT_6C => X"0000009a00000000000000470000000000000075000000000000007e00000000",
            INIT_6D => X"000000570000000000000072000000000000009500000000000000ba00000000",
            INIT_6E => X"0000006300000000000000500000000000000048000000000000005000000000",
            INIT_6F => X"0000005e0000000000000061000000000000005a000000000000006400000000",
            INIT_70 => X"000000ba00000000000000a8000000000000006c00000000000000c200000000",
            INIT_71 => X"000000a7000000000000009c0000000000000063000000000000006900000000",
            INIT_72 => X"000000c6000000000000008a0000000000000073000000000000006400000000",
            INIT_73 => X"0000009a000000000000009100000000000000ac00000000000000be00000000",
            INIT_74 => X"0000009800000000000000470000000000000067000000000000009200000000",
            INIT_75 => X"0000006e0000000000000082000000000000008900000000000000b300000000",
            INIT_76 => X"0000006d000000000000005f000000000000005b000000000000005500000000",
            INIT_77 => X"0000007500000000000000610000000000000064000000000000007300000000",
            INIT_78 => X"000000b800000000000000ac000000000000008400000000000000c500000000",
            INIT_79 => X"0000009b000000000000008c000000000000004e000000000000008200000000",
            INIT_7A => X"000000e6000000000000008f0000000000000082000000000000007300000000",
            INIT_7B => X"000000830000000000000087000000000000009100000000000000f200000000",
            INIT_7C => X"00000090000000000000005f000000000000006c000000000000007900000000",
            INIT_7D => X"000000570000000000000070000000000000009800000000000000a800000000",
            INIT_7E => X"0000007000000000000000690000000000000057000000000000004700000000",
            INIT_7F => X"0000008800000000000000790000000000000067000000000000007800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE0;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE1 : if BRAM_NAME = "sampleifmap_layersamples_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bf00000000000000a8000000000000009200000000000000cb00000000",
            INIT_01 => X"0000008a000000000000007e000000000000004e00000000000000a800000000",
            INIT_02 => X"000000ad000000000000009a0000000000000060000000000000008a00000000",
            INIT_03 => X"000000710000000000000071000000000000008c00000000000000a200000000",
            INIT_04 => X"000000ab00000000000000700000000000000069000000000000006500000000",
            INIT_05 => X"0000006d00000000000000870000000000000094000000000000009c00000000",
            INIT_06 => X"00000065000000000000005e000000000000004f000000000000004e00000000",
            INIT_07 => X"000000900000000000000097000000000000007d000000000000006b00000000",
            INIT_08 => X"000000b700000000000000a400000000000000a300000000000000d600000000",
            INIT_09 => X"0000009c0000000000000060000000000000005e00000000000000b000000000",
            INIT_0A => X"000000760000000000000081000000000000006a000000000000009400000000",
            INIT_0B => X"0000007300000000000000660000000000000074000000000000007200000000",
            INIT_0C => X"0000007600000000000000900000000000000065000000000000005600000000",
            INIT_0D => X"0000004b00000000000000850000000000000080000000000000004400000000",
            INIT_0E => X"000000660000000000000047000000000000003a000000000000003c00000000",
            INIT_0F => X"0000008c0000000000000096000000000000008f000000000000007400000000",
            INIT_10 => X"000000ad00000000000000a700000000000000b200000000000000d400000000",
            INIT_11 => X"0000008d0000000000000056000000000000007c00000000000000b000000000",
            INIT_12 => X"0000004d00000000000000680000000000000087000000000000009900000000",
            INIT_13 => X"000000930000000000000081000000000000007c000000000000008600000000",
            INIT_14 => X"000000840000000000000096000000000000005c000000000000005500000000",
            INIT_15 => X"00000040000000000000004b000000000000006b000000000000007500000000",
            INIT_16 => X"0000008500000000000000560000000000000041000000000000002c00000000",
            INIT_17 => X"00000097000000000000009a00000000000000a0000000000000009b00000000",
            INIT_18 => X"000000ae00000000000000ab00000000000000bb00000000000000c700000000",
            INIT_19 => X"000000770000000000000056000000000000009000000000000000b100000000",
            INIT_1A => X"0000004600000000000000900000000000000089000000000000007a00000000",
            INIT_1B => X"000000b80000000000000091000000000000006c000000000000008100000000",
            INIT_1C => X"0000008900000000000000830000000000000049000000000000007400000000",
            INIT_1D => X"0000003400000000000000330000000000000059000000000000008600000000",
            INIT_1E => X"000000a30000000000000079000000000000005a000000000000002f00000000",
            INIT_1F => X"00000095000000000000009e00000000000000a400000000000000ab00000000",
            INIT_20 => X"000000b100000000000000b300000000000000c300000000000000a500000000",
            INIT_21 => X"000000830000000000000063000000000000009800000000000000b500000000",
            INIT_22 => X"00000050000000000000005d000000000000006700000000000000ab00000000",
            INIT_23 => X"000000bf00000000000000b2000000000000007a000000000000005d00000000",
            INIT_24 => X"0000005700000000000000590000000000000064000000000000009600000000",
            INIT_25 => X"000000180000000000000026000000000000002e000000000000003c00000000",
            INIT_26 => X"00000090000000000000006c000000000000003c000000000000002e00000000",
            INIT_27 => X"00000078000000000000007f0000000000000080000000000000009000000000",
            INIT_28 => X"000000b200000000000000b100000000000000c3000000000000007500000000",
            INIT_29 => X"000000960000000000000053000000000000008a00000000000000b500000000",
            INIT_2A => X"00000086000000000000008500000000000000db00000000000000f500000000",
            INIT_2B => X"000000c200000000000000be00000000000000b0000000000000009500000000",
            INIT_2C => X"0000003d000000000000006e000000000000007d00000000000000a800000000",
            INIT_2D => X"0000003a00000000000000310000000000000022000000000000002300000000",
            INIT_2E => X"000000480000000000000045000000000000003a000000000000003d00000000",
            INIT_2F => X"00000037000000000000003b0000000000000045000000000000004e00000000",
            INIT_30 => X"000000b000000000000000ae00000000000000af000000000000004f00000000",
            INIT_31 => X"000000d3000000000000006d000000000000008c00000000000000b100000000",
            INIT_32 => X"0000007c00000000000000d000000000000000fc00000000000000fd00000000",
            INIT_33 => X"0000007a0000000000000074000000000000007c000000000000007200000000",
            INIT_34 => X"0000003c00000000000000440000000000000044000000000000006800000000",
            INIT_35 => X"0000003800000000000000330000000000000032000000000000003400000000",
            INIT_36 => X"00000033000000000000002b0000000000000033000000000000003800000000",
            INIT_37 => X"0000002a000000000000002b0000000000000030000000000000003b00000000",
            INIT_38 => X"000000a800000000000000900000000000000060000000000000002900000000",
            INIT_39 => X"000000f600000000000000a500000000000000a500000000000000b200000000",
            INIT_3A => X"0000003c000000000000006e00000000000000e300000000000000fd00000000",
            INIT_3B => X"0000003000000000000000310000000000000031000000000000003500000000",
            INIT_3C => X"0000002a000000000000002e000000000000002a000000000000002d00000000",
            INIT_3D => X"0000002b000000000000002e000000000000002e000000000000002600000000",
            INIT_3E => X"00000032000000000000002e000000000000002e000000000000002a00000000",
            INIT_3F => X"0000002d00000000000000330000000000000035000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000083000000000000003b000000000000001d000000000000001d00000000",
            INIT_41 => X"000000fe00000000000000c2000000000000008400000000000000a600000000",
            INIT_42 => X"00000032000000000000003d000000000000008d00000000000000f100000000",
            INIT_43 => X"0000003200000000000000310000000000000033000000000000003200000000",
            INIT_44 => X"000000220000000000000027000000000000002a000000000000002f00000000",
            INIT_45 => X"0000002a00000000000000260000000000000027000000000000002300000000",
            INIT_46 => X"0000003b000000000000003e0000000000000038000000000000002d00000000",
            INIT_47 => X"00000033000000000000002e0000000000000032000000000000003800000000",
            INIT_48 => X"000000490000000000000022000000000000001e000000000000003000000000",
            INIT_49 => X"0000010000000000000000d70000000000000080000000000000008000000000",
            INIT_4A => X"000000320000000000000036000000000000004200000000000000bb00000000",
            INIT_4B => X"0000002d000000000000002e0000000000000034000000000000003400000000",
            INIT_4C => X"0000002700000000000000240000000000000029000000000000002b00000000",
            INIT_4D => X"0000002e000000000000002b0000000000000028000000000000002800000000",
            INIT_4E => X"0000003b0000000000000040000000000000003e000000000000003b00000000",
            INIT_4F => X"0000005300000000000000460000000000000032000000000000003600000000",
            INIT_50 => X"00000029000000000000001f0000000000000023000000000000003400000000",
            INIT_51 => X"000000f000000000000000e00000000000000080000000000000004200000000",
            INIT_52 => X"000000380000000000000031000000000000003a000000000000007c00000000",
            INIT_53 => X"0000002f000000000000002c000000000000002c000000000000003600000000",
            INIT_54 => X"0000002c000000000000002b000000000000002b000000000000002e00000000",
            INIT_55 => X"0000003a0000000000000036000000000000002d000000000000002c00000000",
            INIT_56 => X"00000024000000000000002b000000000000002e000000000000003600000000",
            INIT_57 => X"0000004c00000000000000550000000000000049000000000000003300000000",
            INIT_58 => X"00000023000000000000001d0000000000000023000000000000003200000000",
            INIT_59 => X"000000d300000000000000ca000000000000004e000000000000002c00000000",
            INIT_5A => X"0000003000000000000000360000000000000041000000000000006100000000",
            INIT_5B => X"0000002d00000000000000280000000000000030000000000000003a00000000",
            INIT_5C => X"0000002e000000000000002f0000000000000030000000000000002f00000000",
            INIT_5D => X"0000003000000000000000270000000000000027000000000000003300000000",
            INIT_5E => X"00000028000000000000001c0000000000000027000000000000002f00000000",
            INIT_5F => X"00000033000000000000002e0000000000000043000000000000004300000000",
            INIT_60 => X"0000002100000000000000200000000000000023000000000000003200000000",
            INIT_61 => X"000000aa0000000000000068000000000000002e000000000000002900000000",
            INIT_62 => X"0000003500000000000000340000000000000036000000000000004000000000",
            INIT_63 => X"0000002d0000000000000036000000000000003a000000000000003d00000000",
            INIT_64 => X"00000031000000000000002e0000000000000029000000000000002a00000000",
            INIT_65 => X"000000270000000000000028000000000000002a000000000000002e00000000",
            INIT_66 => X"0000003f000000000000002c0000000000000028000000000000002500000000",
            INIT_67 => X"00000033000000000000000f000000000000001f000000000000002f00000000",
            INIT_68 => X"00000026000000000000001f000000000000002a000000000000004400000000",
            INIT_69 => X"00000047000000000000002a000000000000002b000000000000002500000000",
            INIT_6A => X"00000026000000000000001b000000000000001f000000000000003100000000",
            INIT_6B => X"00000035000000000000003a0000000000000038000000000000003100000000",
            INIT_6C => X"000000350000000000000039000000000000003c000000000000003800000000",
            INIT_6D => X"000000210000000000000027000000000000002d000000000000003200000000",
            INIT_6E => X"00000049000000000000004f000000000000003e000000000000002a00000000",
            INIT_6F => X"00000028000000000000000d0000000000000026000000000000003800000000",
            INIT_70 => X"0000002b00000000000000230000000000000031000000000000003d00000000",
            INIT_71 => X"00000028000000000000002c000000000000002a000000000000002700000000",
            INIT_72 => X"0000001e0000000000000017000000000000001b000000000000002a00000000",
            INIT_73 => X"0000002f0000000000000024000000000000001d000000000000001b00000000",
            INIT_74 => X"0000004b0000000000000042000000000000003e000000000000003800000000",
            INIT_75 => X"0000002b000000000000002b0000000000000031000000000000004500000000",
            INIT_76 => X"0000005d000000000000006d0000000000000055000000000000003c00000000",
            INIT_77 => X"00000014000000000000001d000000000000001a000000000000003c00000000",
            INIT_78 => X"0000002b000000000000002d0000000000000038000000000000003600000000",
            INIT_79 => X"0000002600000000000000280000000000000028000000000000002800000000",
            INIT_7A => X"0000001d0000000000000016000000000000001a000000000000002400000000",
            INIT_7B => X"000000120000000000000013000000000000001d000000000000001900000000",
            INIT_7C => X"0000004a000000000000003d000000000000002f000000000000002000000000",
            INIT_7D => X"0000002d00000000000000340000000000000035000000000000004200000000",
            INIT_7E => X"0000005900000000000000690000000000000059000000000000004300000000",
            INIT_7F => X"0000001500000000000000220000000000000018000000000000003000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE1;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE2 : if BRAM_NAME = "sampleifmap_layersamples_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000760000000000000074000000000000006f000000000000007000000000",
            INIT_01 => X"000000710000000000000073000000000000006d000000000000007000000000",
            INIT_02 => X"0000006f00000000000000740000000000000071000000000000006f00000000",
            INIT_03 => X"0000007700000000000000750000000000000075000000000000006f00000000",
            INIT_04 => X"00000070000000000000006f0000000000000071000000000000007500000000",
            INIT_05 => X"0000006a000000000000006b000000000000006b000000000000006d00000000",
            INIT_06 => X"0000006100000000000000620000000000000065000000000000006b00000000",
            INIT_07 => X"00000055000000000000005b000000000000005f000000000000006100000000",
            INIT_08 => X"000000740000000000000072000000000000006e000000000000007000000000",
            INIT_09 => X"0000007200000000000000750000000000000071000000000000007000000000",
            INIT_0A => X"0000006e000000000000006f000000000000006e000000000000007400000000",
            INIT_0B => X"0000007300000000000000750000000000000077000000000000007100000000",
            INIT_0C => X"000000730000000000000070000000000000006f000000000000007300000000",
            INIT_0D => X"0000006400000000000000660000000000000068000000000000006e00000000",
            INIT_0E => X"0000006100000000000000660000000000000066000000000000006900000000",
            INIT_0F => X"00000058000000000000005b000000000000005f000000000000006200000000",
            INIT_10 => X"0000006f000000000000006f000000000000006d000000000000006e00000000",
            INIT_11 => X"0000007500000000000000750000000000000073000000000000006a00000000",
            INIT_12 => X"0000006d00000000000000720000000000000073000000000000007300000000",
            INIT_13 => X"0000007100000000000000720000000000000073000000000000006f00000000",
            INIT_14 => X"00000060000000000000006f0000000000000072000000000000007400000000",
            INIT_15 => X"00000055000000000000004d000000000000004e000000000000005a00000000",
            INIT_16 => X"0000006300000000000000670000000000000060000000000000005600000000",
            INIT_17 => X"00000059000000000000005f0000000000000062000000000000006300000000",
            INIT_18 => X"00000070000000000000006d000000000000006e000000000000006b00000000",
            INIT_19 => X"0000007700000000000000780000000000000075000000000000006e00000000",
            INIT_1A => X"00000092000000000000007b0000000000000075000000000000007300000000",
            INIT_1B => X"000000720000000000000073000000000000006f000000000000008200000000",
            INIT_1C => X"000000570000000000000050000000000000006f000000000000007000000000",
            INIT_1D => X"0000003f000000000000004b000000000000005a000000000000005a00000000",
            INIT_1E => X"000000620000000000000055000000000000003e000000000000004600000000",
            INIT_1F => X"0000005e00000000000000630000000000000065000000000000006600000000",
            INIT_20 => X"0000007200000000000000730000000000000072000000000000006b00000000",
            INIT_21 => X"0000007400000000000000780000000000000071000000000000007200000000",
            INIT_22 => X"000000d600000000000000800000000000000074000000000000007100000000",
            INIT_23 => X"0000006c000000000000006f0000000000000072000000000000009c00000000",
            INIT_24 => X"0000006700000000000000450000000000000035000000000000005000000000",
            INIT_25 => X"0000005e00000000000000660000000000000072000000000000006e00000000",
            INIT_26 => X"000000530000000000000049000000000000004e000000000000004800000000",
            INIT_27 => X"0000005d000000000000005e0000000000000065000000000000006000000000",
            INIT_28 => X"0000007000000000000000640000000000000068000000000000006d00000000",
            INIT_29 => X"0000007300000000000000740000000000000071000000000000007300000000",
            INIT_2A => X"0000008a00000000000000760000000000000074000000000000006f00000000",
            INIT_2B => X"00000032000000000000004b0000000000000066000000000000007a00000000",
            INIT_2C => X"0000007100000000000000530000000000000038000000000000003a00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007900000000",
            INIT_2E => X"0000003a000000000000003a000000000000005b000000000000006400000000",
            INIT_2F => X"0000005f00000000000000620000000000000069000000000000005400000000",
            INIT_30 => X"0000004a0000000000000025000000000000005f000000000000006400000000",
            INIT_31 => X"0000007600000000000000730000000000000076000000000000007500000000",
            INIT_32 => X"0000006b00000000000000780000000000000074000000000000007500000000",
            INIT_33 => X"000000430000000000000057000000000000006c000000000000006200000000",
            INIT_34 => X"000000820000000000000054000000000000004b000000000000005300000000",
            INIT_35 => X"0000006600000000000000630000000000000076000000000000008e00000000",
            INIT_36 => X"0000002f00000000000000470000000000000053000000000000006f00000000",
            INIT_37 => X"0000005d00000000000000630000000000000062000000000000003d00000000",
            INIT_38 => X"00000040000000000000002b0000000000000060000000000000007300000000",
            INIT_39 => X"0000007400000000000000720000000000000075000000000000006f00000000",
            INIT_3A => X"0000005e000000000000006d0000000000000071000000000000007700000000",
            INIT_3B => X"00000057000000000000006a0000000000000083000000000000006e00000000",
            INIT_3C => X"00000076000000000000004d0000000000000058000000000000005f00000000",
            INIT_3D => X"00000062000000000000005d000000000000007c000000000000009900000000",
            INIT_3E => X"00000035000000000000003c0000000000000051000000000000005d00000000",
            INIT_3F => X"0000006100000000000000670000000000000053000000000000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000079000000000000003a000000000000006900000000000000a100000000",
            INIT_41 => X"0000007a00000000000000750000000000000071000000000000007c00000000",
            INIT_42 => X"0000006900000000000000590000000000000087000000000000007900000000",
            INIT_43 => X"00000050000000000000006f000000000000008f000000000000008d00000000",
            INIT_44 => X"00000047000000000000004e0000000000000055000000000000005100000000",
            INIT_45 => X"0000004f00000000000000670000000000000087000000000000007d00000000",
            INIT_46 => X"0000003900000000000000490000000000000052000000000000004d00000000",
            INIT_47 => X"00000067000000000000006a000000000000003b000000000000002300000000",
            INIT_48 => X"0000009a0000000000000064000000000000008b00000000000000b000000000",
            INIT_49 => X"0000007600000000000000740000000000000074000000000000009500000000",
            INIT_4A => X"0000008300000000000000b400000000000000d600000000000000b400000000",
            INIT_4B => X"00000055000000000000006e0000000000000083000000000000009900000000",
            INIT_4C => X"000000440000000000000039000000000000004a000000000000005400000000",
            INIT_4D => X"00000062000000000000007c0000000000000085000000000000007d00000000",
            INIT_4E => X"0000004c00000000000000550000000000000055000000000000005100000000",
            INIT_4F => X"00000067000000000000004b000000000000001e000000000000003100000000",
            INIT_50 => X"000000a90000000000000097000000000000007400000000000000b700000000",
            INIT_51 => X"0000005900000000000000760000000000000070000000000000009c00000000",
            INIT_52 => X"0000008700000000000000bf00000000000000e000000000000000c500000000",
            INIT_53 => X"0000006f000000000000006c0000000000000089000000000000009f00000000",
            INIT_54 => X"00000055000000000000002c0000000000000050000000000000004c00000000",
            INIT_55 => X"000000640000000000000093000000000000009300000000000000a500000000",
            INIT_56 => X"0000004f00000000000000580000000000000066000000000000005300000000",
            INIT_57 => X"00000051000000000000002e0000000000000024000000000000003b00000000",
            INIT_58 => X"000000af0000000000000090000000000000006c00000000000000bf00000000",
            INIT_59 => X"0000005d000000000000007b000000000000007800000000000000a700000000",
            INIT_5A => X"0000008e00000000000000ab00000000000000b6000000000000005f00000000",
            INIT_5B => X"0000006b000000000000007700000000000000ab00000000000000a100000000",
            INIT_5C => X"0000007900000000000000260000000000000054000000000000006200000000",
            INIT_5D => X"00000059000000000000008b000000000000009800000000000000c900000000",
            INIT_5E => X"000000570000000000000068000000000000005d000000000000005000000000",
            INIT_5F => X"0000003800000000000000370000000000000035000000000000004b00000000",
            INIT_60 => X"000000b40000000000000086000000000000006000000000000000c200000000",
            INIT_61 => X"0000006d000000000000007b000000000000007b000000000000009c00000000",
            INIT_62 => X"000000720000000000000090000000000000009a000000000000004400000000",
            INIT_63 => X"00000071000000000000009500000000000000ca00000000000000a600000000",
            INIT_64 => X"0000009300000000000000320000000000000072000000000000007200000000",
            INIT_65 => X"000000580000000000000076000000000000009500000000000000bb00000000",
            INIT_66 => X"00000057000000000000005f0000000000000054000000000000005300000000",
            INIT_67 => X"00000037000000000000004a0000000000000049000000000000005700000000",
            INIT_68 => X"000000bc000000000000009a000000000000005f00000000000000c000000000",
            INIT_69 => X"00000074000000000000007c000000000000006a000000000000006e00000000",
            INIT_6A => X"00000095000000000000007d0000000000000084000000000000004800000000",
            INIT_6B => X"0000008300000000000000ac00000000000000d800000000000000ae00000000",
            INIT_6C => X"0000009800000000000000470000000000000072000000000000007500000000",
            INIT_6D => X"00000055000000000000006e000000000000009000000000000000b500000000",
            INIT_6E => X"0000006400000000000000500000000000000049000000000000005000000000",
            INIT_6F => X"0000004900000000000000590000000000000058000000000000006500000000",
            INIT_70 => X"000000ba00000000000000a7000000000000006b00000000000000c400000000",
            INIT_71 => X"0000007a00000000000000770000000000000059000000000000006d00000000",
            INIT_72 => X"000000b9000000000000007b000000000000006a000000000000004a00000000",
            INIT_73 => X"0000008f000000000000008c00000000000000a500000000000000b400000000",
            INIT_74 => X"0000009800000000000000470000000000000064000000000000008800000000",
            INIT_75 => X"0000006d0000000000000080000000000000008500000000000000af00000000",
            INIT_76 => X"0000006e0000000000000060000000000000005d000000000000005600000000",
            INIT_77 => X"0000005f00000000000000550000000000000060000000000000007400000000",
            INIT_78 => X"000000b200000000000000a7000000000000008100000000000000c500000000",
            INIT_79 => X"0000007d00000000000000780000000000000053000000000000008900000000",
            INIT_7A => X"000000dd00000000000000830000000000000078000000000000005e00000000",
            INIT_7B => X"000000790000000000000082000000000000008a00000000000000ec00000000",
            INIT_7C => X"0000008600000000000000580000000000000068000000000000007000000000",
            INIT_7D => X"00000055000000000000006c0000000000000093000000000000009f00000000",
            INIT_7E => X"0000006d00000000000000680000000000000058000000000000004800000000",
            INIT_7F => X"0000006800000000000000600000000000000056000000000000006e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE2;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE3 : if BRAM_NAME = "sampleifmap_layersamples_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b600000000000000a4000000000000009200000000000000cb00000000",
            INIT_01 => X"0000007e000000000000007d000000000000005600000000000000aa00000000",
            INIT_02 => X"000000a3000000000000008f0000000000000050000000000000007900000000",
            INIT_03 => X"0000006a000000000000006a0000000000000084000000000000009800000000",
            INIT_04 => X"0000008f000000000000005a0000000000000065000000000000006500000000",
            INIT_05 => X"000000690000000000000082000000000000008d000000000000008a00000000",
            INIT_06 => X"0000005b000000000000005d000000000000004f000000000000004c00000000",
            INIT_07 => X"00000068000000000000006c0000000000000058000000000000005300000000",
            INIT_08 => X"000000b800000000000000a700000000000000a600000000000000d700000000",
            INIT_09 => X"000000950000000000000060000000000000006600000000000000b600000000",
            INIT_0A => X"000000690000000000000074000000000000005d000000000000008900000000",
            INIT_0B => X"0000006e000000000000005b0000000000000069000000000000006600000000",
            INIT_0C => X"0000006000000000000000800000000000000067000000000000005b00000000",
            INIT_0D => X"00000045000000000000007e0000000000000078000000000000003800000000",
            INIT_0E => X"0000005d00000000000000460000000000000038000000000000003800000000",
            INIT_0F => X"0000006e00000000000000740000000000000070000000000000005e00000000",
            INIT_10 => X"000000b500000000000000af00000000000000b800000000000000d300000000",
            INIT_11 => X"0000008b0000000000000058000000000000008300000000000000b800000000",
            INIT_12 => X"00000040000000000000005a0000000000000080000000000000009400000000",
            INIT_13 => X"0000008f0000000000000075000000000000006f000000000000007900000000",
            INIT_14 => X"00000075000000000000008b0000000000000060000000000000005c00000000",
            INIT_15 => X"0000003b00000000000000440000000000000063000000000000006d00000000",
            INIT_16 => X"000000690000000000000045000000000000003e000000000000002900000000",
            INIT_17 => X"0000006f00000000000000730000000000000078000000000000007700000000",
            INIT_18 => X"000000b300000000000000b000000000000000bd00000000000000c000000000",
            INIT_19 => X"00000079000000000000005a000000000000009500000000000000b600000000",
            INIT_1A => X"0000003b00000000000000860000000000000088000000000000007c00000000",
            INIT_1B => X"000000b000000000000000860000000000000061000000000000007600000000",
            INIT_1C => X"0000007c0000000000000077000000000000004b000000000000007600000000",
            INIT_1D => X"0000003300000000000000310000000000000056000000000000008100000000",
            INIT_1E => X"00000076000000000000005b000000000000005a000000000000003100000000",
            INIT_1F => X"0000006b000000000000006f0000000000000071000000000000007900000000",
            INIT_20 => X"000000ad00000000000000b200000000000000c1000000000000009c00000000",
            INIT_21 => X"000000870000000000000067000000000000009d00000000000000b500000000",
            INIT_22 => X"0000004d000000000000005a000000000000006900000000000000af00000000",
            INIT_23 => X"000000b600000000000000ad0000000000000076000000000000005a00000000",
            INIT_24 => X"0000004d000000000000004e0000000000000064000000000000009400000000",
            INIT_25 => X"00000021000000000000002e0000000000000034000000000000003d00000000",
            INIT_26 => X"0000007d00000000000000640000000000000047000000000000003900000000",
            INIT_27 => X"000000690000000000000071000000000000006d000000000000007b00000000",
            INIT_28 => X"000000a900000000000000b200000000000000c8000000000000007800000000",
            INIT_29 => X"000000990000000000000057000000000000009000000000000000b300000000",
            INIT_2A => X"0000008d000000000000008c00000000000000de00000000000000f700000000",
            INIT_2B => X"000000c000000000000000c400000000000000b6000000000000009c00000000",
            INIT_2C => X"0000003e000000000000006d000000000000008500000000000000ac00000000",
            INIT_2D => X"0000005100000000000000460000000000000036000000000000003100000000",
            INIT_2E => X"0000006500000000000000630000000000000054000000000000005500000000",
            INIT_2F => X"0000005a000000000000005c0000000000000060000000000000006800000000",
            INIT_30 => X"000000ac00000000000000b700000000000000c5000000000000006900000000",
            INIT_31 => X"000000d30000000000000070000000000000009200000000000000b100000000",
            INIT_32 => X"0000008f00000000000000e000000000000000fd00000000000000fc00000000",
            INIT_33 => X"000000850000000000000085000000000000008d000000000000008400000000",
            INIT_34 => X"000000520000000000000057000000000000005d000000000000007c00000000",
            INIT_35 => X"0000005d00000000000000550000000000000054000000000000005400000000",
            INIT_36 => X"000000680000000000000060000000000000005b000000000000005e00000000",
            INIT_37 => X"0000005f00000000000000610000000000000061000000000000006c00000000",
            INIT_38 => X"000000ae00000000000000a80000000000000089000000000000005900000000",
            INIT_39 => X"000000f500000000000000a600000000000000aa00000000000000b600000000",
            INIT_3A => X"00000058000000000000008800000000000000e700000000000000fb00000000",
            INIT_3B => X"00000048000000000000004b000000000000004c000000000000005000000000",
            INIT_3C => X"0000005200000000000000510000000000000051000000000000004f00000000",
            INIT_3D => X"000000570000000000000059000000000000005a000000000000005600000000",
            INIT_3E => X"00000060000000000000005e000000000000005d000000000000005900000000",
            INIT_3F => X"0000005a000000000000005f000000000000005e000000000000006000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009900000000000000660000000000000057000000000000005b00000000",
            INIT_41 => X"000000fa00000000000000bd000000000000008800000000000000b300000000",
            INIT_42 => X"00000054000000000000005e000000000000009f00000000000000f500000000",
            INIT_43 => X"0000005400000000000000530000000000000055000000000000005400000000",
            INIT_44 => X"0000004f00000000000000520000000000000054000000000000005600000000",
            INIT_45 => X"0000005900000000000000550000000000000056000000000000005300000000",
            INIT_46 => X"0000006500000000000000670000000000000067000000000000005c00000000",
            INIT_47 => X"00000067000000000000005e0000000000000063000000000000006600000000",
            INIT_48 => X"0000006a0000000000000055000000000000005e000000000000006f00000000",
            INIT_49 => X"000000fd00000000000000d50000000000000088000000000000009400000000",
            INIT_4A => X"00000058000000000000005b000000000000005d00000000000000c600000000",
            INIT_4B => X"000000520000000000000053000000000000005a000000000000005a00000000",
            INIT_4C => X"0000005300000000000000500000000000000051000000000000005200000000",
            INIT_4D => X"0000005f000000000000005c0000000000000059000000000000005600000000",
            INIT_4E => X"0000006c000000000000006d000000000000006e000000000000006c00000000",
            INIT_4F => X"00000089000000000000007b0000000000000069000000000000006c00000000",
            INIT_50 => X"0000005300000000000000560000000000000063000000000000007200000000",
            INIT_51 => X"000000f500000000000000e50000000000000091000000000000005f00000000",
            INIT_52 => X"0000005e0000000000000057000000000000005c000000000000008f00000000",
            INIT_53 => X"0000005300000000000000520000000000000052000000000000005c00000000",
            INIT_54 => X"0000005800000000000000560000000000000053000000000000005400000000",
            INIT_55 => X"0000006e000000000000006a0000000000000061000000000000005a00000000",
            INIT_56 => X"0000005b000000000000005f0000000000000061000000000000006900000000",
            INIT_57 => X"0000007d000000000000008a0000000000000082000000000000006c00000000",
            INIT_58 => X"0000005600000000000000590000000000000062000000000000006e00000000",
            INIT_59 => X"000000e400000000000000db000000000000006a000000000000005300000000",
            INIT_5A => X"00000057000000000000005e0000000000000068000000000000007e00000000",
            INIT_5B => X"0000005200000000000000500000000000000057000000000000006100000000",
            INIT_5C => X"0000005900000000000000590000000000000057000000000000005400000000",
            INIT_5D => X"00000066000000000000005d000000000000005c000000000000006100000000",
            INIT_5E => X"000000650000000000000055000000000000005d000000000000006500000000",
            INIT_5F => X"000000600000000000000062000000000000007e000000000000008100000000",
            INIT_60 => X"00000058000000000000005c0000000000000061000000000000006c00000000",
            INIT_61 => X"000000c500000000000000850000000000000054000000000000005800000000",
            INIT_62 => X"0000005f000000000000005e0000000000000061000000000000006400000000",
            INIT_63 => X"0000005300000000000000600000000000000064000000000000006700000000",
            INIT_64 => X"0000005c00000000000000580000000000000050000000000000004f00000000",
            INIT_65 => X"0000005c000000000000005d000000000000005f000000000000005c00000000",
            INIT_66 => X"0000007d0000000000000066000000000000005d000000000000005a00000000",
            INIT_67 => X"0000005d000000000000003c000000000000005a000000000000006e00000000",
            INIT_68 => X"0000005b00000000000000580000000000000064000000000000007c00000000",
            INIT_69 => X"0000006b000000000000004f0000000000000059000000000000005700000000",
            INIT_6A => X"000000520000000000000047000000000000004d000000000000005900000000",
            INIT_6B => X"0000005c00000000000000660000000000000064000000000000005d00000000",
            INIT_6C => X"0000006100000000000000630000000000000063000000000000005e00000000",
            INIT_6D => X"000000530000000000000058000000000000005e000000000000005f00000000",
            INIT_6E => X"0000008300000000000000840000000000000070000000000000005b00000000",
            INIT_6F => X"0000005500000000000000400000000000000061000000000000007400000000",
            INIT_70 => X"0000005b00000000000000550000000000000066000000000000007400000000",
            INIT_71 => X"000000510000000000000058000000000000005c000000000000005a00000000",
            INIT_72 => X"0000004a00000000000000430000000000000048000000000000005500000000",
            INIT_73 => X"0000005600000000000000500000000000000049000000000000004700000000",
            INIT_74 => X"00000077000000000000006d0000000000000065000000000000005f00000000",
            INIT_75 => X"000000580000000000000058000000000000005f000000000000007100000000",
            INIT_76 => X"00000091000000000000009c0000000000000082000000000000006900000000",
            INIT_77 => X"0000004000000000000000520000000000000052000000000000007300000000",
            INIT_78 => X"0000005600000000000000590000000000000069000000000000006b00000000",
            INIT_79 => X"000000510000000000000057000000000000005c000000000000005900000000",
            INIT_7A => X"0000004900000000000000420000000000000045000000000000004f00000000",
            INIT_7B => X"0000003a000000000000003f0000000000000049000000000000004500000000",
            INIT_7C => X"0000007700000000000000680000000000000057000000000000004600000000",
            INIT_7D => X"00000057000000000000005f0000000000000060000000000000006f00000000",
            INIT_7E => X"0000008700000000000000920000000000000083000000000000006d00000000",
            INIT_7F => X"000000430000000000000054000000000000004d000000000000006300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE3;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE4 : if BRAM_NAME = "sampleifmap_layersamples_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000350000000000000033000000000000002f000000000000003100000000",
            INIT_01 => X"0000002d000000000000002f0000000000000029000000000000002e00000000",
            INIT_02 => X"0000003400000000000000290000000000000029000000000000002c00000000",
            INIT_03 => X"0000002c000000000000002d0000000000000029000000000000003100000000",
            INIT_04 => X"0000002b00000000000000270000000000000026000000000000002800000000",
            INIT_05 => X"0000002b000000000000002d000000000000002d000000000000002c00000000",
            INIT_06 => X"00000029000000000000002b0000000000000027000000000000002c00000000",
            INIT_07 => X"0000002100000000000000240000000000000024000000000000002600000000",
            INIT_08 => X"00000038000000000000002d0000000000000028000000000000003300000000",
            INIT_09 => X"0000002d000000000000002f000000000000002b000000000000003100000000",
            INIT_0A => X"0000003600000000000000290000000000000026000000000000002e00000000",
            INIT_0B => X"0000002100000000000000280000000000000029000000000000003400000000",
            INIT_0C => X"0000003200000000000000290000000000000021000000000000001e00000000",
            INIT_0D => X"0000003000000000000000340000000000000037000000000000003500000000",
            INIT_0E => X"00000026000000000000002d000000000000002e000000000000003200000000",
            INIT_0F => X"000000220000000000000020000000000000001f000000000000002200000000",
            INIT_10 => X"0000003000000000000000240000000000000021000000000000002f00000000",
            INIT_11 => X"0000002d000000000000002d000000000000002c000000000000002a00000000",
            INIT_12 => X"000000390000000000000030000000000000002b000000000000002b00000000",
            INIT_13 => X"0000002300000000000000250000000000000026000000000000003300000000",
            INIT_14 => X"000000310000000000000036000000000000002f000000000000002700000000",
            INIT_15 => X"00000032000000000000002f0000000000000032000000000000003400000000",
            INIT_16 => X"0000002700000000000000330000000000000037000000000000003000000000",
            INIT_17 => X"0000002100000000000000220000000000000022000000000000002300000000",
            INIT_18 => X"0000002c000000000000001f0000000000000020000000000000002800000000",
            INIT_19 => X"000000300000000000000030000000000000002e000000000000002b00000000",
            INIT_1A => X"0000005f0000000000000039000000000000002d000000000000002c00000000",
            INIT_1B => X"00000036000000000000002f0000000000000029000000000000004b00000000",
            INIT_1C => X"00000041000000000000002f0000000000000043000000000000003a00000000",
            INIT_1D => X"0000003200000000000000420000000000000054000000000000004c00000000",
            INIT_1E => X"0000002e000000000000002d0000000000000027000000000000003400000000",
            INIT_1F => X"0000002400000000000000270000000000000027000000000000002b00000000",
            INIT_20 => X"0000002f00000000000000310000000000000030000000000000002900000000",
            INIT_21 => X"0000002c000000000000002f0000000000000028000000000000002b00000000",
            INIT_22 => X"000000a4000000000000003b000000000000002a000000000000002900000000",
            INIT_23 => X"00000047000000000000003c0000000000000038000000000000006b00000000",
            INIT_24 => X"000000620000000000000038000000000000001f000000000000003200000000",
            INIT_25 => X"0000005d00000000000000690000000000000076000000000000006f00000000",
            INIT_26 => X"0000002d000000000000002f0000000000000046000000000000004300000000",
            INIT_27 => X"000000240000000000000024000000000000002e000000000000003000000000",
            INIT_28 => X"0000003500000000000000390000000000000040000000000000003600000000",
            INIT_29 => X"0000002900000000000000290000000000000027000000000000002c00000000",
            INIT_2A => X"00000055000000000000002a0000000000000027000000000000002500000000",
            INIT_2B => X"0000001f000000000000002b000000000000003a000000000000004e00000000",
            INIT_2C => X"0000006e000000000000004c000000000000002d000000000000002b00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007800000000",
            INIT_2E => X"00000025000000000000002f0000000000000056000000000000006100000000",
            INIT_2F => X"00000028000000000000002c000000000000003a000000000000003100000000",
            INIT_30 => X"0000001c00000000000000110000000000000050000000000000003900000000",
            INIT_31 => X"0000002b0000000000000028000000000000002b000000000000003000000000",
            INIT_32 => X"0000003400000000000000270000000000000025000000000000002a00000000",
            INIT_33 => X"000000390000000000000046000000000000004b000000000000003b00000000",
            INIT_34 => X"00000079000000000000004a0000000000000040000000000000004800000000",
            INIT_35 => X"0000005e000000000000005a000000000000006c000000000000008400000000",
            INIT_36 => X"000000270000000000000045000000000000004d000000000000006700000000",
            INIT_37 => X"000000270000000000000030000000000000003a000000000000002400000000",
            INIT_38 => X"000000290000000000000026000000000000005c000000000000005a00000000",
            INIT_39 => X"000000270000000000000024000000000000002a000000000000003800000000",
            INIT_3A => X"0000003100000000000000330000000000000033000000000000003100000000",
            INIT_3B => X"0000004f000000000000005d000000000000006b000000000000004d00000000",
            INIT_3C => X"0000006b00000000000000450000000000000052000000000000005800000000",
            INIT_3D => X"0000005800000000000000510000000000000070000000000000008c00000000",
            INIT_3E => X"00000031000000000000003a000000000000004a000000000000005400000000",
            INIT_3F => X"0000002700000000000000330000000000000032000000000000002000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000071000000000000003b0000000000000069000000000000009000000000",
            INIT_41 => X"000000320000000000000029000000000000002b000000000000005200000000",
            INIT_42 => X"0000004e000000000000003b000000000000005f000000000000004200000000",
            INIT_43 => X"0000004a00000000000000650000000000000080000000000000007900000000",
            INIT_44 => X"0000003d00000000000000490000000000000052000000000000004d00000000",
            INIT_45 => X"00000046000000000000005d000000000000007b000000000000007000000000",
            INIT_46 => X"000000350000000000000043000000000000004c000000000000004500000000",
            INIT_47 => X"0000002d000000000000003b0000000000000023000000000000001b00000000",
            INIT_48 => X"000000950000000000000069000000000000008f00000000000000a300000000",
            INIT_49 => X"0000003c000000000000002f0000000000000033000000000000007000000000",
            INIT_4A => X"0000007700000000000000a600000000000000c6000000000000009200000000",
            INIT_4B => X"0000004f000000000000006b000000000000007d000000000000009100000000",
            INIT_4C => X"0000003a00000000000000350000000000000047000000000000004f00000000",
            INIT_4D => X"000000590000000000000072000000000000007a000000000000007000000000",
            INIT_4E => X"00000047000000000000004e000000000000004e000000000000004a00000000",
            INIT_4F => X"00000039000000000000002c000000000000000f000000000000002b00000000",
            INIT_50 => X"000000a8000000000000009e000000000000007a00000000000000af00000000",
            INIT_51 => X"0000002f00000000000000330000000000000032000000000000007a00000000",
            INIT_52 => X"0000008300000000000000bc00000000000000e200000000000000b300000000",
            INIT_53 => X"0000006800000000000000680000000000000084000000000000009b00000000",
            INIT_54 => X"0000004d0000000000000028000000000000004d000000000000004500000000",
            INIT_55 => X"0000005c000000000000008a0000000000000089000000000000009a00000000",
            INIT_56 => X"00000049000000000000004f0000000000000060000000000000004d00000000",
            INIT_57 => X"0000002e000000000000001f0000000000000021000000000000003b00000000",
            INIT_58 => X"000000b20000000000000099000000000000007400000000000000bd00000000",
            INIT_59 => X"0000002c0000000000000037000000000000003b000000000000008800000000",
            INIT_5A => X"0000008500000000000000a400000000000000bc000000000000005000000000",
            INIT_5B => X"0000005f000000000000006a000000000000009f000000000000009700000000",
            INIT_5C => X"000000710000000000000022000000000000004f000000000000005900000000",
            INIT_5D => X"000000520000000000000082000000000000008e00000000000000c000000000",
            INIT_5E => X"00000051000000000000005e0000000000000058000000000000004b00000000",
            INIT_5F => X"0000001a00000000000000300000000000000037000000000000004e00000000",
            INIT_60 => X"000000b90000000000000090000000000000006900000000000000c200000000",
            INIT_61 => X"0000002f00000000000000350000000000000044000000000000008500000000",
            INIT_62 => X"0000005e000000000000007e0000000000000098000000000000002c00000000",
            INIT_63 => X"00000062000000000000008100000000000000b7000000000000009400000000",
            INIT_64 => X"0000008c000000000000002f000000000000006d000000000000006900000000",
            INIT_65 => X"00000053000000000000006f000000000000008c00000000000000b200000000",
            INIT_66 => X"0000005100000000000000550000000000000050000000000000004f00000000",
            INIT_67 => X"0000001800000000000000400000000000000049000000000000005900000000",
            INIT_68 => X"000000c000000000000000a3000000000000006700000000000000c100000000",
            INIT_69 => X"00000032000000000000003a0000000000000042000000000000006200000000",
            INIT_6A => X"0000007f00000000000000670000000000000078000000000000002700000000",
            INIT_6B => X"00000075000000000000009d00000000000000c8000000000000009b00000000",
            INIT_6C => X"000000930000000000000044000000000000006d000000000000006b00000000",
            INIT_6D => X"000000500000000000000068000000000000008800000000000000ae00000000",
            INIT_6E => X"0000005e00000000000000480000000000000046000000000000004c00000000",
            INIT_6F => X"0000002200000000000000450000000000000051000000000000006300000000",
            INIT_70 => X"000000bc00000000000000ac000000000000007000000000000000c400000000",
            INIT_71 => X"00000037000000000000003e0000000000000043000000000000006d00000000",
            INIT_72 => X"000000a900000000000000670000000000000058000000000000002200000000",
            INIT_73 => X"00000086000000000000008c000000000000009f00000000000000a900000000",
            INIT_74 => X"000000950000000000000046000000000000005f000000000000007d00000000",
            INIT_75 => X"00000069000000000000007a000000000000007f00000000000000aa00000000",
            INIT_76 => X"00000068000000000000005a000000000000005b000000000000005300000000",
            INIT_77 => X"0000002f00000000000000350000000000000050000000000000006f00000000",
            INIT_78 => X"000000b500000000000000ae000000000000008800000000000000c500000000",
            INIT_79 => X"0000004d0000000000000058000000000000004d000000000000008e00000000",
            INIT_7A => X"000000d30000000000000074000000000000005d000000000000003400000000",
            INIT_7B => X"000000700000000000000082000000000000008900000000000000e600000000",
            INIT_7C => X"00000076000000000000004b000000000000005f000000000000006500000000",
            INIT_7D => X"000000500000000000000065000000000000008a000000000000009200000000",
            INIT_7E => X"0000006300000000000000630000000000000057000000000000004400000000",
            INIT_7F => X"0000003000000000000000300000000000000036000000000000005d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE4;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE5 : if BRAM_NAME = "sampleifmap_layersamples_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bc00000000000000b200000000000000a000000000000000cc00000000",
            INIT_01 => X"00000071000000000000007e000000000000005a00000000000000ac00000000",
            INIT_02 => X"0000009b00000000000000850000000000000025000000000000005200000000",
            INIT_03 => X"0000005a00000000000000580000000000000075000000000000008d00000000",
            INIT_04 => X"00000068000000000000003a0000000000000057000000000000005c00000000",
            INIT_05 => X"000000610000000000000076000000000000007e000000000000006d00000000",
            INIT_06 => X"00000052000000000000005e000000000000004d000000000000004800000000",
            INIT_07 => X"0000002e0000000000000037000000000000002d000000000000003700000000",
            INIT_08 => X"000000c200000000000000b800000000000000b400000000000000d700000000",
            INIT_09 => X"000000910000000000000066000000000000006900000000000000ba00000000",
            INIT_0A => X"0000005f0000000000000069000000000000003d000000000000006f00000000",
            INIT_0B => X"0000006200000000000000490000000000000059000000000000005900000000",
            INIT_0C => X"000000400000000000000066000000000000005f000000000000005800000000",
            INIT_0D => X"0000003d00000000000000730000000000000069000000000000002000000000",
            INIT_0E => X"0000004e00000000000000410000000000000035000000000000003300000000",
            INIT_0F => X"0000003600000000000000400000000000000044000000000000004000000000",
            INIT_10 => X"000000c100000000000000bd00000000000000c000000000000000cd00000000",
            INIT_11 => X"0000008f0000000000000060000000000000008500000000000000bc00000000",
            INIT_12 => X"000000370000000000000050000000000000006f000000000000008d00000000",
            INIT_13 => X"0000008500000000000000640000000000000060000000000000006c00000000",
            INIT_14 => X"0000005d0000000000000078000000000000005d000000000000005d00000000",
            INIT_15 => X"00000034000000000000003a0000000000000056000000000000005c00000000",
            INIT_16 => X"0000003b0000000000000028000000000000003c000000000000002700000000",
            INIT_17 => X"0000002e000000000000002d0000000000000036000000000000003e00000000",
            INIT_18 => X"000000b900000000000000b500000000000000bb00000000000000b400000000",
            INIT_19 => X"000000840000000000000063000000000000009800000000000000b800000000",
            INIT_1A => X"00000033000000000000007e0000000000000087000000000000008200000000",
            INIT_1B => X"000000a8000000000000007b0000000000000056000000000000006c00000000",
            INIT_1C => X"0000006900000000000000670000000000000049000000000000007600000000",
            INIT_1D => X"00000032000000000000002c000000000000004e000000000000007600000000",
            INIT_1E => X"00000044000000000000003c000000000000005d000000000000003400000000",
            INIT_1F => X"0000002e00000000000000320000000000000034000000000000004000000000",
            INIT_20 => X"000000ac00000000000000af00000000000000bb000000000000009200000000",
            INIT_21 => X"00000092000000000000006f00000000000000a000000000000000b400000000",
            INIT_22 => X"000000490000000000000057000000000000006f00000000000000b900000000",
            INIT_23 => X"000000b100000000000000ad0000000000000074000000000000005600000000",
            INIT_24 => X"0000003f00000000000000420000000000000065000000000000009400000000",
            INIT_25 => X"0000002900000000000000330000000000000036000000000000003900000000",
            INIT_26 => X"00000052000000000000004b0000000000000053000000000000004500000000",
            INIT_27 => X"0000003f0000000000000045000000000000003d000000000000004c00000000",
            INIT_28 => X"000000a800000000000000b000000000000000c8000000000000007c00000000",
            INIT_29 => X"0000009f000000000000005b000000000000009300000000000000b300000000",
            INIT_2A => X"00000093000000000000009000000000000000e100000000000000fa00000000",
            INIT_2B => X"000000c500000000000000d000000000000000c000000000000000a400000000",
            INIT_2C => X"0000003e000000000000006d000000000000008f00000000000000b500000000",
            INIT_2D => X"0000006600000000000000570000000000000044000000000000003a00000000",
            INIT_2E => X"00000077000000000000007a000000000000006f000000000000006e00000000",
            INIT_2F => X"0000007300000000000000700000000000000070000000000000007800000000",
            INIT_30 => X"000000b100000000000000c000000000000000d5000000000000008500000000",
            INIT_31 => X"000000d10000000000000071000000000000009600000000000000b600000000",
            INIT_32 => X"0000009d00000000000000e800000000000000fc00000000000000f700000000",
            INIT_33 => X"00000098000000000000009c00000000000000a2000000000000009500000000",
            INIT_34 => X"0000006500000000000000680000000000000077000000000000009400000000",
            INIT_35 => X"0000007d0000000000000073000000000000006e000000000000006f00000000",
            INIT_36 => X"0000008d00000000000000870000000000000082000000000000008300000000",
            INIT_37 => X"0000008400000000000000890000000000000084000000000000008e00000000",
            INIT_38 => X"000000bc00000000000000bc00000000000000a8000000000000008700000000",
            INIT_39 => X"000000ed00000000000000a400000000000000ae00000000000000c000000000",
            INIT_3A => X"0000006f000000000000009900000000000000e400000000000000f100000000",
            INIT_3B => X"00000065000000000000006b0000000000000069000000000000006900000000",
            INIT_3C => X"0000007400000000000000710000000000000078000000000000007300000000",
            INIT_3D => X"00000080000000000000007e000000000000007d000000000000007d00000000",
            INIT_3E => X"000000890000000000000089000000000000008b000000000000008400000000",
            INIT_3F => X"00000085000000000000008b0000000000000086000000000000008700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b000000000000000860000000000000082000000000000008d00000000",
            INIT_41 => X"000000f200000000000000b5000000000000008900000000000000bf00000000",
            INIT_42 => X"00000076000000000000007f00000000000000af00000000000000f500000000",
            INIT_43 => X"0000007400000000000000780000000000000079000000000000007700000000",
            INIT_44 => X"0000007100000000000000730000000000000075000000000000007500000000",
            INIT_45 => X"00000082000000000000007d000000000000007d000000000000007800000000",
            INIT_46 => X"0000008e000000000000008e0000000000000091000000000000008600000000",
            INIT_47 => X"00000095000000000000008c0000000000000090000000000000009200000000",
            INIT_48 => X"00000088000000000000007c000000000000008c00000000000000a200000000",
            INIT_49 => X"000000f900000000000000d1000000000000008f00000000000000a700000000",
            INIT_4A => X"0000007d0000000000000080000000000000007600000000000000cd00000000",
            INIT_4B => X"000000730000000000000079000000000000007f000000000000007f00000000",
            INIT_4C => X"0000007500000000000000710000000000000070000000000000007100000000",
            INIT_4D => X"0000008a00000000000000860000000000000083000000000000007b00000000",
            INIT_4E => X"0000009500000000000000930000000000000098000000000000009600000000",
            INIT_4F => X"000000b600000000000000a70000000000000098000000000000009a00000000",
            INIT_50 => X"0000007a0000000000000082000000000000009300000000000000a500000000",
            INIT_51 => X"000000f700000000000000ea00000000000000a4000000000000007e00000000",
            INIT_52 => X"00000083000000000000007b0000000000000072000000000000009900000000",
            INIT_53 => X"0000007700000000000000770000000000000077000000000000008100000000",
            INIT_54 => X"0000007f000000000000007b0000000000000077000000000000007700000000",
            INIT_55 => X"0000009a0000000000000096000000000000008d000000000000008300000000",
            INIT_56 => X"0000008a000000000000008c000000000000008d000000000000009600000000",
            INIT_57 => X"000000a900000000000000b600000000000000b2000000000000009e00000000",
            INIT_58 => X"00000085000000000000008a000000000000009500000000000000a200000000",
            INIT_59 => X"000000ea00000000000000e9000000000000008a000000000000007e00000000",
            INIT_5A => X"0000007c0000000000000081000000000000007e000000000000008c00000000",
            INIT_5B => X"000000770000000000000074000000000000007b000000000000008500000000",
            INIT_5C => X"000000840000000000000082000000000000007e000000000000007a00000000",
            INIT_5D => X"00000094000000000000008b000000000000008a000000000000008c00000000",
            INIT_5E => X"000000990000000000000085000000000000008b000000000000009300000000",
            INIT_5F => X"0000008b000000000000008e00000000000000b000000000000000b600000000",
            INIT_60 => X"0000008d000000000000008f000000000000009300000000000000a100000000",
            INIT_61 => X"000000d3000000000000009f000000000000007d000000000000008a00000000",
            INIT_62 => X"0000008200000000000000800000000000000079000000000000007700000000",
            INIT_63 => X"0000007800000000000000830000000000000087000000000000008b00000000",
            INIT_64 => X"0000008700000000000000820000000000000078000000000000007600000000",
            INIT_65 => X"00000088000000000000008a000000000000008b000000000000008800000000",
            INIT_66 => X"000000b20000000000000097000000000000008a000000000000008700000000",
            INIT_67 => X"000000880000000000000067000000000000008c00000000000000a400000000",
            INIT_68 => X"000000920000000000000089000000000000009400000000000000b100000000",
            INIT_69 => X"0000008500000000000000710000000000000084000000000000008b00000000",
            INIT_6A => X"0000007500000000000000690000000000000069000000000000007200000000",
            INIT_6B => X"0000008000000000000000890000000000000087000000000000008000000000",
            INIT_6C => X"0000008a000000000000008b0000000000000089000000000000008300000000",
            INIT_6D => X"0000007d00000000000000830000000000000088000000000000008900000000",
            INIT_6E => X"000000b500000000000000b3000000000000009a000000000000008500000000",
            INIT_6F => X"0000007f000000000000006c000000000000009200000000000000a800000000",
            INIT_70 => X"0000008f0000000000000084000000000000009400000000000000a800000000",
            INIT_71 => X"00000070000000000000007d0000000000000086000000000000008b00000000",
            INIT_72 => X"0000006d00000000000000660000000000000068000000000000007300000000",
            INIT_73 => X"000000780000000000000073000000000000006c000000000000006a00000000",
            INIT_74 => X"0000009c00000000000000900000000000000087000000000000008000000000",
            INIT_75 => X"0000007f000000000000007f0000000000000086000000000000009800000000",
            INIT_76 => X"000000be00000000000000c500000000000000aa000000000000009000000000",
            INIT_77 => X"0000006b000000000000007e000000000000008200000000000000a400000000",
            INIT_78 => X"000000860000000000000084000000000000009500000000000000a000000000",
            INIT_79 => X"00000073000000000000007b0000000000000084000000000000008600000000",
            INIT_7A => X"0000006c00000000000000650000000000000069000000000000007200000000",
            INIT_7B => X"000000590000000000000062000000000000006c000000000000006800000000",
            INIT_7C => X"0000009800000000000000890000000000000076000000000000006400000000",
            INIT_7D => X"0000007b00000000000000820000000000000083000000000000009100000000",
            INIT_7E => X"000000af00000000000000b600000000000000a7000000000000009100000000",
            INIT_7F => X"0000006e0000000000000081000000000000007c000000000000009100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE5;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE6 : if BRAM_NAME = "sampleifmap_layersamples_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e800000000000000e800000000000000e700000000000000eb00000000",
            INIT_01 => X"000000e800000000000000e800000000000000e800000000000000e800000000",
            INIT_02 => X"000000e900000000000000e900000000000000e800000000000000e800000000",
            INIT_03 => X"000000e900000000000000e900000000000000e900000000000000e900000000",
            INIT_04 => X"000000e600000000000000e700000000000000e800000000000000e900000000",
            INIT_05 => X"000000e900000000000000e800000000000000e800000000000000e800000000",
            INIT_06 => X"000000e800000000000000e800000000000000e900000000000000e800000000",
            INIT_07 => X"000000e800000000000000e900000000000000e900000000000000e800000000",
            INIT_08 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_09 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_0A => X"000000ec00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_0B => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_0C => X"000000ea00000000000000ec00000000000000ec00000000000000ed00000000",
            INIT_0D => X"000000ec00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_0E => X"000000eb00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_0F => X"000000eb00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_10 => X"000000ea00000000000000ea00000000000000ea00000000000000ed00000000",
            INIT_11 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_12 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_13 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_14 => X"000000ea00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_15 => X"000000ea00000000000000e700000000000000e700000000000000e300000000",
            INIT_16 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_17 => X"000000ea00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_18 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_19 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_1A => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_1B => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_1C => X"000000df00000000000000e400000000000000e800000000000000e900000000",
            INIT_1D => X"000000e400000000000000cf00000000000000d100000000000000ba00000000",
            INIT_1E => X"000000ea00000000000000ea00000000000000ea00000000000000ec00000000",
            INIT_1F => X"000000eb00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_20 => X"000000eb00000000000000eb00000000000000ea00000000000000ed00000000",
            INIT_21 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_22 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_23 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_24 => X"000000cb00000000000000db00000000000000e900000000000000ec00000000",
            INIT_25 => X"000000e600000000000000d600000000000000c300000000000000a300000000",
            INIT_26 => X"000000eb00000000000000eb00000000000000eb00000000000000ed00000000",
            INIT_27 => X"000000ec00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_28 => X"000000ec00000000000000ec00000000000000ec00000000000000ef00000000",
            INIT_29 => X"000000eb00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_2A => X"000000ed00000000000000ed00000000000000eb00000000000000ea00000000",
            INIT_2B => X"000000e500000000000000eb00000000000000e800000000000000ea00000000",
            INIT_2C => X"000000ae00000000000000b900000000000000c200000000000000d000000000",
            INIT_2D => X"000000e200000000000000cf00000000000000b800000000000000a500000000",
            INIT_2E => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_2F => X"000000ed00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_30 => X"000000e700000000000000e800000000000000e400000000000000e400000000",
            INIT_31 => X"000000ec00000000000000ed00000000000000ed00000000000000ea00000000",
            INIT_32 => X"000000ef00000000000000ef00000000000000ed00000000000000ed00000000",
            INIT_33 => X"000000dd00000000000000e900000000000000e000000000000000e100000000",
            INIT_34 => X"0000009a000000000000009f00000000000000a100000000000000b700000000",
            INIT_35 => X"000000c6000000000000009c000000000000008f000000000000009000000000",
            INIT_36 => X"000000eb00000000000000eb00000000000000ec00000000000000e900000000",
            INIT_37 => X"000000ef00000000000000ed00000000000000ec00000000000000eb00000000",
            INIT_38 => X"000000e300000000000000e600000000000000e000000000000000d400000000",
            INIT_39 => X"000000ee00000000000000ed00000000000000ea00000000000000e500000000",
            INIT_3A => X"000000f000000000000000ef00000000000000ef00000000000000ef00000000",
            INIT_3B => X"000000d600000000000000e900000000000000db00000000000000c900000000",
            INIT_3C => X"000000ad00000000000000b800000000000000b900000000000000c100000000",
            INIT_3D => X"000000ba00000000000000a2000000000000009f00000000000000a500000000",
            INIT_3E => X"000000e900000000000000e900000000000000ea00000000000000e500000000",
            INIT_3F => X"000000ee00000000000000ed00000000000000ec00000000000000ea00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000e100000000000000e100000000000000dd00000000000000d800000000",
            INIT_41 => X"000000ee00000000000000ec00000000000000e700000000000000e300000000",
            INIT_42 => X"000000ef00000000000000ed00000000000000ee00000000000000ee00000000",
            INIT_43 => X"000000e600000000000000e900000000000000dc00000000000000c500000000",
            INIT_44 => X"000000d000000000000000db00000000000000d100000000000000d100000000",
            INIT_45 => X"000000da00000000000000d900000000000000d200000000000000d100000000",
            INIT_46 => X"000000e600000000000000e400000000000000e400000000000000e100000000",
            INIT_47 => X"000000ee00000000000000ed00000000000000eb00000000000000e600000000",
            INIT_48 => X"00000088000000000000007c0000000000000077000000000000007600000000",
            INIT_49 => X"000000ed00000000000000eb00000000000000e100000000000000ac00000000",
            INIT_4A => X"000000e900000000000000eb00000000000000eb00000000000000ec00000000",
            INIT_4B => X"000000ec00000000000000e800000000000000e200000000000000d600000000",
            INIT_4C => X"000000e100000000000000e700000000000000e300000000000000e400000000",
            INIT_4D => X"000000b900000000000000c900000000000000d900000000000000e100000000",
            INIT_4E => X"000000ba00000000000000a700000000000000a700000000000000ac00000000",
            INIT_4F => X"000000ee00000000000000ec00000000000000eb00000000000000df00000000",
            INIT_50 => X"0000006f000000000000006c0000000000000067000000000000006d00000000",
            INIT_51 => X"000000e500000000000000e300000000000000de000000000000009200000000",
            INIT_52 => X"000000e600000000000000e700000000000000ea00000000000000ec00000000",
            INIT_53 => X"000000e600000000000000e800000000000000e700000000000000e500000000",
            INIT_54 => X"000000df00000000000000e500000000000000e700000000000000e700000000",
            INIT_55 => X"00000089000000000000009200000000000000a400000000000000bf00000000",
            INIT_56 => X"0000009500000000000000790000000000000080000000000000008600000000",
            INIT_57 => X"000000ed00000000000000eb00000000000000ea00000000000000d800000000",
            INIT_58 => X"000000c800000000000000c700000000000000bc00000000000000c300000000",
            INIT_59 => X"000000d300000000000000d500000000000000df00000000000000d100000000",
            INIT_5A => X"000000d200000000000000db00000000000000dc00000000000000d800000000",
            INIT_5B => X"000000dc00000000000000d800000000000000d300000000000000d100000000",
            INIT_5C => X"000000da00000000000000e100000000000000e200000000000000e100000000",
            INIT_5D => X"000000b200000000000000b500000000000000af00000000000000b700000000",
            INIT_5E => X"000000b9000000000000008e00000000000000aa00000000000000ba00000000",
            INIT_5F => X"000000ec00000000000000ea00000000000000e700000000000000db00000000",
            INIT_60 => X"000000d600000000000000ca00000000000000bf00000000000000c100000000",
            INIT_61 => X"000000ab00000000000000cb00000000000000d600000000000000df00000000",
            INIT_62 => X"0000006200000000000000ae00000000000000cf00000000000000b100000000",
            INIT_63 => X"0000007a000000000000006f0000000000000065000000000000005d00000000",
            INIT_64 => X"000000df00000000000000ca0000000000000099000000000000008900000000",
            INIT_65 => X"000000d900000000000000df00000000000000dc00000000000000da00000000",
            INIT_66 => X"000000de00000000000000c400000000000000d400000000000000dd00000000",
            INIT_67 => X"000000eb00000000000000e800000000000000dd00000000000000db00000000",
            INIT_68 => X"0000007d0000000000000071000000000000006f000000000000007100000000",
            INIT_69 => X"000000be00000000000000bf00000000000000aa000000000000008a00000000",
            INIT_6A => X"00000036000000000000009e00000000000000d800000000000000d000000000",
            INIT_6B => X"0000004200000000000000350000000000000031000000000000002d00000000",
            INIT_6C => X"000000ea00000000000000dd000000000000009f000000000000006600000000",
            INIT_6D => X"000000cf00000000000000df00000000000000e300000000000000e900000000",
            INIT_6E => X"000000c700000000000000d400000000000000d300000000000000ca00000000",
            INIT_6F => X"000000dd00000000000000d300000000000000bc00000000000000b300000000",
            INIT_70 => X"00000044000000000000003f0000000000000045000000000000003d00000000",
            INIT_71 => X"000000c30000000000000097000000000000008b000000000000007b00000000",
            INIT_72 => X"0000006700000000000000a300000000000000ce00000000000000d600000000",
            INIT_73 => X"000000b5000000000000008a0000000000000065000000000000005f00000000",
            INIT_74 => X"000000cd00000000000000db00000000000000dd00000000000000cf00000000",
            INIT_75 => X"000000830000000000000093000000000000009e00000000000000b700000000",
            INIT_76 => X"0000008500000000000000880000000000000082000000000000007d00000000",
            INIT_77 => X"000000c500000000000000b6000000000000008a000000000000008000000000",
            INIT_78 => X"0000007f0000000000000055000000000000003a000000000000002800000000",
            INIT_79 => X"000000a300000000000000770000000000000060000000000000008400000000",
            INIT_7A => X"000000b500000000000000b600000000000000b800000000000000ad00000000",
            INIT_7B => X"000000c800000000000000da00000000000000c600000000000000b700000000",
            INIT_7C => X"000000840000000000000091000000000000009f00000000000000ae00000000",
            INIT_7D => X"00000063000000000000005e0000000000000062000000000000007400000000",
            INIT_7E => X"0000008a000000000000007a000000000000006b000000000000006900000000",
            INIT_7F => X"000000b900000000000000bc000000000000009d000000000000009600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE6;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE7 : if BRAM_NAME = "sampleifmap_layersamples_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ce0000000000000086000000000000001a000000000000000d00000000",
            INIT_01 => X"000000ac000000000000008d0000000000000076000000000000008a00000000",
            INIT_02 => X"000000e400000000000000dc00000000000000cf00000000000000b500000000",
            INIT_03 => X"000000b000000000000000e200000000000000e600000000000000e000000000",
            INIT_04 => X"00000091000000000000008e000000000000008a000000000000009000000000",
            INIT_05 => X"0000009a00000000000000950000000000000095000000000000009a00000000",
            INIT_06 => X"000000bb00000000000000ad00000000000000a0000000000000009d00000000",
            INIT_07 => X"0000009d00000000000000a500000000000000b200000000000000be00000000",
            INIT_08 => X"000000e100000000000000c8000000000000003a000000000000000500000000",
            INIT_09 => X"000000e200000000000000d400000000000000c700000000000000c500000000",
            INIT_0A => X"000000e600000000000000e800000000000000e900000000000000e500000000",
            INIT_0B => X"000000d200000000000000dd00000000000000df00000000000000d100000000",
            INIT_0C => X"000000bc00000000000000c100000000000000b400000000000000c600000000",
            INIT_0D => X"000000b800000000000000c000000000000000c200000000000000bd00000000",
            INIT_0E => X"0000009000000000000000a100000000000000ab00000000000000ac00000000",
            INIT_0F => X"0000008a00000000000000800000000000000083000000000000008800000000",
            INIT_10 => X"000000ba00000000000000be0000000000000091000000000000002700000000",
            INIT_11 => X"000000c200000000000000c200000000000000c000000000000000b800000000",
            INIT_12 => X"000000be00000000000000c000000000000000bf00000000000000c200000000",
            INIT_13 => X"00000093000000000000009a00000000000000b400000000000000b100000000",
            INIT_14 => X"000000710000000000000092000000000000009c000000000000009100000000",
            INIT_15 => X"0000006f000000000000007e0000000000000084000000000000007200000000",
            INIT_16 => X"0000005e000000000000005d000000000000005b000000000000005c00000000",
            INIT_17 => X"0000008100000000000000810000000000000079000000000000006900000000",
            INIT_18 => X"00000089000000000000008f00000000000000a2000000000000007a00000000",
            INIT_19 => X"00000082000000000000007f0000000000000080000000000000008300000000",
            INIT_1A => X"00000081000000000000007f0000000000000080000000000000008300000000",
            INIT_1B => X"000000640000000000000068000000000000007c000000000000008100000000",
            INIT_1C => X"0000005e00000000000000700000000000000076000000000000006600000000",
            INIT_1D => X"000000530000000000000057000000000000005e000000000000005e00000000",
            INIT_1E => X"00000065000000000000005d0000000000000053000000000000005000000000",
            INIT_1F => X"0000008200000000000000790000000000000073000000000000006c00000000",
            INIT_20 => X"00000050000000000000004d000000000000004c000000000000004900000000",
            INIT_21 => X"0000005a00000000000000570000000000000057000000000000005400000000",
            INIT_22 => X"00000071000000000000006b0000000000000066000000000000005e00000000",
            INIT_23 => X"0000007800000000000000760000000000000076000000000000007300000000",
            INIT_24 => X"00000064000000000000006a000000000000006e000000000000007300000000",
            INIT_25 => X"00000050000000000000004f0000000000000055000000000000005f00000000",
            INIT_26 => X"000000520000000000000050000000000000004d000000000000005000000000",
            INIT_27 => X"00000088000000000000007d0000000000000071000000000000005c00000000",
            INIT_28 => X"0000001200000000000000090000000000000003000000000000000d00000000",
            INIT_29 => X"0000001600000000000000140000000000000015000000000000001200000000",
            INIT_2A => X"00000030000000000000002a0000000000000022000000000000001a00000000",
            INIT_2B => X"000000460000000000000042000000000000003c000000000000003400000000",
            INIT_2C => X"0000003c00000000000000430000000000000048000000000000004700000000",
            INIT_2D => X"0000003900000000000000350000000000000035000000000000003700000000",
            INIT_2E => X"0000005700000000000000480000000000000039000000000000003900000000",
            INIT_2F => X"0000008900000000000000820000000000000078000000000000006800000000",
            INIT_30 => X"000000200000000000000008000000000000000b000000000000002400000000",
            INIT_31 => X"0000000300000000000000080000000000000016000000000000002400000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_33 => X"0000000300000000000000010000000000000005000000000000000600000000",
            INIT_34 => X"0000001500000000000000150000000000000018000000000000000d00000000",
            INIT_35 => X"00000027000000000000001e0000000000000016000000000000001500000000",
            INIT_36 => X"0000007b00000000000000710000000000000055000000000000003900000000",
            INIT_37 => X"000000990000000000000086000000000000007a000000000000007400000000",
            INIT_38 => X"0000001b000000000000000d000000000000001a000000000000002300000000",
            INIT_39 => X"0000001b00000000000000310000000000000046000000000000004700000000",
            INIT_3A => X"0000000000000000000000020000000000000005000000000000000f00000000",
            INIT_3B => X"0000000a000000000000001f0000000000000039000000000000001100000000",
            INIT_3C => X"0000000e00000000000000070000000000000004000000000000000400000000",
            INIT_3D => X"00000056000000000000003e0000000000000029000000000000001900000000",
            INIT_3E => X"0000007200000000000000840000000000000090000000000000007a00000000",
            INIT_3F => X"000000ac00000000000000920000000000000084000000000000007500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000030000000000000004000000000000000d000000000000001000000000",
            INIT_41 => X"0000002400000000000000360000000000000041000000000000002d00000000",
            INIT_42 => X"0000000000000000000000020000000000000004000000000000001200000000",
            INIT_43 => X"0000008300000000000000a10000000000000076000000000000000700000000",
            INIT_44 => X"0000006d00000000000000690000000000000069000000000000007000000000",
            INIT_45 => X"00000097000000000000009a000000000000008a000000000000007600000000",
            INIT_46 => X"00000078000000000000006a0000000000000069000000000000007f00000000",
            INIT_47 => X"000000b800000000000000a4000000000000008e000000000000008100000000",
            INIT_48 => X"000000000000000000000000000000000000000c000000000000002800000000",
            INIT_49 => X"000000150000000000000020000000000000001e000000000000000c00000000",
            INIT_4A => X"0000000300000000000000020000000000000002000000000000000700000000",
            INIT_4B => X"000000cd00000000000000b60000000000000044000000000000000000000000",
            INIT_4C => X"000000bb00000000000000c300000000000000c200000000000000c400000000",
            INIT_4D => X"00000067000000000000007b000000000000009600000000000000ac00000000",
            INIT_4E => X"00000081000000000000007a0000000000000068000000000000005f00000000",
            INIT_4F => X"000000b900000000000000ab0000000000000098000000000000008400000000",
            INIT_50 => X"000000010000000000000001000000000000001a000000000000004500000000",
            INIT_51 => X"0000000c0000000000000012000000000000000c000000000000000400000000",
            INIT_52 => X"0000000400000000000000020000000000000002000000000000000400000000",
            INIT_53 => X"000000cb00000000000000990000000000000020000000000000000100000000",
            INIT_54 => X"0000009b00000000000000b300000000000000bf00000000000000c300000000",
            INIT_55 => X"0000005e0000000000000051000000000000005b000000000000007700000000",
            INIT_56 => X"00000081000000000000007d000000000000007d000000000000007500000000",
            INIT_57 => X"000000b800000000000000ad00000000000000a2000000000000009000000000",
            INIT_58 => X"000000020000000000000001000000000000002f000000000000005300000000",
            INIT_59 => X"0000000400000000000000070000000000000005000000000000000200000000",
            INIT_5A => X"0000000300000000000000010000000000000001000000000000000100000000",
            INIT_5B => X"000000cd000000000000008e000000000000001b000000000000000100000000",
            INIT_5C => X"00000055000000000000007900000000000000a900000000000000c600000000",
            INIT_5D => X"0000007900000000000000660000000000000055000000000000004a00000000",
            INIT_5E => X"000000840000000000000079000000000000007a000000000000008000000000",
            INIT_5F => X"000000ba00000000000000b000000000000000a5000000000000009300000000",
            INIT_60 => X"0000000300000000000000060000000000000036000000000000005c00000000",
            INIT_61 => X"0000000100000000000000010000000000000001000000000000000200000000",
            INIT_62 => X"0000000100000000000000010000000000000001000000000000000100000000",
            INIT_63 => X"0000009d0000000000000066000000000000000f000000000000000000000000",
            INIT_64 => X"0000004a0000000000000038000000000000004a000000000000007500000000",
            INIT_65 => X"0000007c000000000000007a0000000000000073000000000000006300000000",
            INIT_66 => X"000000880000000000000080000000000000007d000000000000007b00000000",
            INIT_67 => X"000000bc00000000000000b100000000000000a2000000000000009400000000",
            INIT_68 => X"0000000b0000000000000013000000000000002b000000000000005700000000",
            INIT_69 => X"0000000200000000000000020000000000000005000000000000000800000000",
            INIT_6A => X"0000000200000000000000030000000000000003000000000000000300000000",
            INIT_6B => X"00000047000000000000002a0000000000000004000000000000000000000000",
            INIT_6C => X"0000007100000000000000500000000000000039000000000000003500000000",
            INIT_6D => X"00000074000000000000007b0000000000000086000000000000008400000000",
            INIT_6E => X"0000008f000000000000008b0000000000000083000000000000007800000000",
            INIT_6F => X"000000bc00000000000000b600000000000000a9000000000000009c00000000",
            INIT_70 => X"0000001f0000000000000024000000000000002e000000000000005200000000",
            INIT_71 => X"0000001000000000000000110000000000000016000000000000001b00000000",
            INIT_72 => X"0000001300000000000000140000000000000013000000000000001200000000",
            INIT_73 => X"0000004000000000000000250000000000000017000000000000001300000000",
            INIT_74 => X"0000008000000000000000740000000000000068000000000000005700000000",
            INIT_75 => X"0000007300000000000000750000000000000083000000000000008b00000000",
            INIT_76 => X"00000094000000000000008b0000000000000083000000000000007b00000000",
            INIT_77 => X"000000bb00000000000000b900000000000000ae000000000000009f00000000",
            INIT_78 => X"00000037000000000000003a000000000000003e000000000000005500000000",
            INIT_79 => X"00000030000000000000002e000000000000002f000000000000003300000000",
            INIT_7A => X"0000003700000000000000350000000000000033000000000000003100000000",
            INIT_7B => X"0000006800000000000000510000000000000044000000000000003b00000000",
            INIT_7C => X"0000007f0000000000000085000000000000007f000000000000007400000000",
            INIT_7D => X"0000007a00000000000000720000000000000076000000000000007f00000000",
            INIT_7E => X"00000095000000000000008d0000000000000088000000000000008100000000",
            INIT_7F => X"000000ba00000000000000b400000000000000a8000000000000009e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE7;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE8 : if BRAM_NAME = "sampleifmap_layersamples_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e800000000000000e800000000000000e700000000000000eb00000000",
            INIT_01 => X"000000e800000000000000e800000000000000e800000000000000e800000000",
            INIT_02 => X"000000e900000000000000e900000000000000e800000000000000e800000000",
            INIT_03 => X"000000e800000000000000e900000000000000e900000000000000e900000000",
            INIT_04 => X"000000e900000000000000e900000000000000e700000000000000e700000000",
            INIT_05 => X"000000e900000000000000e800000000000000e700000000000000e800000000",
            INIT_06 => X"000000e800000000000000e800000000000000e900000000000000e900000000",
            INIT_07 => X"000000e800000000000000e900000000000000e900000000000000e800000000",
            INIT_08 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_09 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_0A => X"000000ec00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_0B => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_0C => X"000000ec00000000000000ec00000000000000ea00000000000000ea00000000",
            INIT_0D => X"000000ec00000000000000ec00000000000000ea00000000000000eb00000000",
            INIT_0E => X"000000eb00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_0F => X"000000eb00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_10 => X"000000ea00000000000000ea00000000000000ea00000000000000ed00000000",
            INIT_11 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_12 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_13 => X"000000ea00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_14 => X"000000eb00000000000000eb00000000000000ea00000000000000e900000000",
            INIT_15 => X"000000ea00000000000000e900000000000000eb00000000000000e600000000",
            INIT_16 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_17 => X"000000ea00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_18 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_19 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_1A => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_1B => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_1C => X"000000e200000000000000e600000000000000e800000000000000e900000000",
            INIT_1D => X"000000e400000000000000d200000000000000d800000000000000c000000000",
            INIT_1E => X"000000ea00000000000000ea00000000000000ea00000000000000eb00000000",
            INIT_1F => X"000000eb00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_20 => X"000000eb00000000000000eb00000000000000ea00000000000000ed00000000",
            INIT_21 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_22 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_23 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_24 => X"000000d200000000000000e100000000000000ed00000000000000ee00000000",
            INIT_25 => X"000000e500000000000000da00000000000000cd00000000000000ac00000000",
            INIT_26 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_27 => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_28 => X"000000eb00000000000000eb00000000000000eb00000000000000ef00000000",
            INIT_29 => X"000000eb00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_2A => X"000000ec00000000000000ec00000000000000eb00000000000000ea00000000",
            INIT_2B => X"000000e700000000000000ed00000000000000e900000000000000eb00000000",
            INIT_2C => X"000000bc00000000000000c600000000000000cd00000000000000d800000000",
            INIT_2D => X"000000e400000000000000d700000000000000c400000000000000b300000000",
            INIT_2E => X"000000ec00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_2F => X"000000ed00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_30 => X"000000e400000000000000e600000000000000e300000000000000e500000000",
            INIT_31 => X"000000ed00000000000000ed00000000000000ec00000000000000e800000000",
            INIT_32 => X"000000ed00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_33 => X"000000e200000000000000ed00000000000000e400000000000000e500000000",
            INIT_34 => X"000000b000000000000000b400000000000000b400000000000000c500000000",
            INIT_35 => X"000000ce00000000000000a9000000000000009f00000000000000a300000000",
            INIT_36 => X"000000eb00000000000000ec00000000000000ed00000000000000ee00000000",
            INIT_37 => X"000000ed00000000000000ed00000000000000ee00000000000000ec00000000",
            INIT_38 => X"000000e800000000000000ea00000000000000e600000000000000dc00000000",
            INIT_39 => X"000000ed00000000000000ee00000000000000ed00000000000000ea00000000",
            INIT_3A => X"000000ee00000000000000ec00000000000000ed00000000000000ed00000000",
            INIT_3B => X"000000da00000000000000ec00000000000000de00000000000000cc00000000",
            INIT_3C => X"000000bf00000000000000c900000000000000c900000000000000cc00000000",
            INIT_3D => X"000000c700000000000000b000000000000000ae00000000000000b600000000",
            INIT_3E => X"000000ee00000000000000ee00000000000000ef00000000000000ef00000000",
            INIT_3F => X"000000ee00000000000000ef00000000000000ef00000000000000ef00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ef00000000000000ee00000000000000ec00000000000000ea00000000",
            INIT_41 => X"000000ec00000000000000ed00000000000000ee00000000000000f000000000",
            INIT_42 => X"000000ef00000000000000ed00000000000000ec00000000000000ec00000000",
            INIT_43 => X"000000e700000000000000ea00000000000000dd00000000000000c600000000",
            INIT_44 => X"000000da00000000000000e400000000000000d800000000000000d500000000",
            INIT_45 => X"000000eb00000000000000e900000000000000e000000000000000dd00000000",
            INIT_46 => X"000000f000000000000000ef00000000000000ee00000000000000f000000000",
            INIT_47 => X"000000ee00000000000000f000000000000000f000000000000000f000000000",
            INIT_48 => X"0000009b000000000000008e000000000000008a000000000000008c00000000",
            INIT_49 => X"000000ea00000000000000ec00000000000000ea00000000000000bc00000000",
            INIT_4A => X"000000ed00000000000000ed00000000000000eb00000000000000e900000000",
            INIT_4B => X"000000ed00000000000000ea00000000000000e400000000000000d800000000",
            INIT_4C => X"000000e800000000000000ec00000000000000e600000000000000e600000000",
            INIT_4D => X"000000cc00000000000000db00000000000000e900000000000000ed00000000",
            INIT_4E => X"000000c700000000000000b400000000000000b300000000000000bd00000000",
            INIT_4F => X"000000f000000000000000f000000000000000f100000000000000eb00000000",
            INIT_50 => X"0000007f000000000000007d0000000000000079000000000000008200000000",
            INIT_51 => X"000000e200000000000000e400000000000000e5000000000000009f00000000",
            INIT_52 => X"000000ed00000000000000ec00000000000000ea00000000000000e800000000",
            INIT_53 => X"000000eb00000000000000ed00000000000000eb00000000000000ea00000000",
            INIT_54 => X"000000e800000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_55 => X"0000009c00000000000000a500000000000000b800000000000000ce00000000",
            INIT_56 => X"000000a20000000000000085000000000000008c000000000000009500000000",
            INIT_57 => X"000000f000000000000000f000000000000000f100000000000000e400000000",
            INIT_58 => X"000000d300000000000000d300000000000000ca00000000000000d400000000",
            INIT_59 => X"000000d100000000000000d500000000000000e300000000000000d900000000",
            INIT_5A => X"000000dd00000000000000e200000000000000de00000000000000d500000000",
            INIT_5B => X"000000e500000000000000e100000000000000dd00000000000000db00000000",
            INIT_5C => X"000000e700000000000000ed00000000000000ec00000000000000ea00000000",
            INIT_5D => X"000000c200000000000000c800000000000000c600000000000000cc00000000",
            INIT_5E => X"000000c3000000000000009700000000000000b200000000000000c500000000",
            INIT_5F => X"000000f000000000000000f100000000000000f000000000000000e600000000",
            INIT_60 => X"000000d900000000000000d300000000000000ca00000000000000cf00000000",
            INIT_61 => X"000000ae00000000000000d000000000000000db00000000000000e100000000",
            INIT_62 => X"0000007000000000000000b800000000000000d500000000000000b400000000",
            INIT_63 => X"0000008a00000000000000810000000000000079000000000000007200000000",
            INIT_64 => X"000000ec00000000000000d800000000000000a7000000000000009800000000",
            INIT_65 => X"000000e200000000000000ea00000000000000e900000000000000e800000000",
            INIT_66 => X"000000e600000000000000cb00000000000000db00000000000000e400000000",
            INIT_67 => X"000000f100000000000000ef00000000000000e600000000000000e300000000",
            INIT_68 => X"00000083000000000000007d000000000000007d000000000000008200000000",
            INIT_69 => X"000000c700000000000000c900000000000000b6000000000000009100000000",
            INIT_6A => X"0000004700000000000000ac00000000000000e600000000000000db00000000",
            INIT_6B => X"0000005400000000000000490000000000000049000000000000004600000000",
            INIT_6C => X"000000ef00000000000000e300000000000000a8000000000000007200000000",
            INIT_6D => X"000000d300000000000000e400000000000000e700000000000000ed00000000",
            INIT_6E => X"000000ce00000000000000db00000000000000da00000000000000d000000000",
            INIT_6F => X"000000e700000000000000dd00000000000000c500000000000000ba00000000",
            INIT_70 => X"00000055000000000000004f0000000000000056000000000000005100000000",
            INIT_71 => X"000000c8000000000000009d000000000000009b000000000000008d00000000",
            INIT_72 => X"0000007900000000000000b400000000000000df00000000000000e400000000",
            INIT_73 => X"000000c000000000000000970000000000000075000000000000007000000000",
            INIT_74 => X"000000cb00000000000000db00000000000000de00000000000000d400000000",
            INIT_75 => X"0000008a000000000000009a00000000000000a600000000000000ba00000000",
            INIT_76 => X"0000008e0000000000000092000000000000008b000000000000008500000000",
            INIT_77 => X"000000d400000000000000c50000000000000099000000000000008900000000",
            INIT_78 => X"0000009000000000000000620000000000000046000000000000003500000000",
            INIT_79 => X"0000009e0000000000000073000000000000006b000000000000009700000000",
            INIT_7A => X"000000c100000000000000c200000000000000c200000000000000b400000000",
            INIT_7B => X"000000d200000000000000e400000000000000d100000000000000c200000000",
            INIT_7C => X"00000088000000000000009600000000000000a500000000000000b500000000",
            INIT_7D => X"0000006f000000000000006a000000000000006f000000000000007d00000000",
            INIT_7E => X"0000009700000000000000870000000000000079000000000000007600000000",
            INIT_7F => X"000000cb00000000000000ce00000000000000ae00000000000000a400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE8;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE9 : if BRAM_NAME = "sampleifmap_layersamples_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d8000000000000008c000000000000001d000000000000000f00000000",
            INIT_01 => X"000000a20000000000000085000000000000007b000000000000009600000000",
            INIT_02 => X"000000ea00000000000000e000000000000000d100000000000000b500000000",
            INIT_03 => X"000000bd00000000000000ee00000000000000f100000000000000ea00000000",
            INIT_04 => X"000000a3000000000000009e000000000000009a000000000000009f00000000",
            INIT_05 => X"000000ab00000000000000a500000000000000a500000000000000ab00000000",
            INIT_06 => X"000000cc00000000000000be00000000000000b100000000000000ae00000000",
            INIT_07 => X"000000af00000000000000b700000000000000c400000000000000cf00000000",
            INIT_08 => X"000000e800000000000000cf000000000000003e000000000000000500000000",
            INIT_09 => X"000000e000000000000000d400000000000000cf00000000000000cd00000000",
            INIT_0A => X"000000ee00000000000000ee00000000000000ec00000000000000e600000000",
            INIT_0B => X"000000e400000000000000ee00000000000000ee00000000000000dd00000000",
            INIT_0C => X"000000d500000000000000d800000000000000c800000000000000d900000000",
            INIT_0D => X"000000cc00000000000000d400000000000000d600000000000000d400000000",
            INIT_0E => X"000000a500000000000000b500000000000000bf00000000000000c100000000",
            INIT_0F => X"0000009a000000000000008f0000000000000092000000000000009c00000000",
            INIT_10 => X"000000c400000000000000cc000000000000009b000000000000002d00000000",
            INIT_11 => X"000000d000000000000000d300000000000000d300000000000000c500000000",
            INIT_12 => X"000000cf00000000000000cf00000000000000cb00000000000000ce00000000",
            INIT_13 => X"000000a900000000000000b000000000000000c600000000000000c100000000",
            INIT_14 => X"0000008500000000000000a300000000000000ab00000000000000a100000000",
            INIT_15 => X"000000870000000000000096000000000000009d000000000000008900000000",
            INIT_16 => X"0000007400000000000000720000000000000070000000000000007300000000",
            INIT_17 => X"0000008e000000000000008d0000000000000085000000000000007d00000000",
            INIT_18 => X"0000009a00000000000000a000000000000000b3000000000000008700000000",
            INIT_19 => X"0000009600000000000000960000000000000098000000000000009800000000",
            INIT_1A => X"0000009500000000000000930000000000000093000000000000009600000000",
            INIT_1B => X"0000007a000000000000007e0000000000000091000000000000009500000000",
            INIT_1C => X"0000006d00000000000000800000000000000086000000000000007800000000",
            INIT_1D => X"0000006700000000000000700000000000000075000000000000007000000000",
            INIT_1E => X"00000075000000000000006f0000000000000067000000000000006100000000",
            INIT_1F => X"000000900000000000000085000000000000007d000000000000007900000000",
            INIT_20 => X"0000005d000000000000005a000000000000005a000000000000005700000000",
            INIT_21 => X"0000006900000000000000660000000000000066000000000000006200000000",
            INIT_22 => X"00000083000000000000007c0000000000000077000000000000006f00000000",
            INIT_23 => X"0000008500000000000000840000000000000088000000000000008900000000",
            INIT_24 => X"00000077000000000000007f0000000000000085000000000000008800000000",
            INIT_25 => X"0000005c00000000000000610000000000000065000000000000006d00000000",
            INIT_26 => X"0000006200000000000000640000000000000064000000000000005e00000000",
            INIT_27 => X"0000009500000000000000870000000000000077000000000000006800000000",
            INIT_28 => X"0000001a0000000000000010000000000000000b000000000000001900000000",
            INIT_29 => X"0000001e00000000000000190000000000000019000000000000001a00000000",
            INIT_2A => X"0000003b0000000000000033000000000000002b000000000000002400000000",
            INIT_2B => X"0000004f000000000000004d000000000000004b000000000000004500000000",
            INIT_2C => X"0000004800000000000000510000000000000058000000000000005700000000",
            INIT_2D => X"0000004500000000000000450000000000000044000000000000004300000000",
            INIT_2E => X"000000640000000000000059000000000000004e000000000000004700000000",
            INIT_2F => X"000000920000000000000088000000000000007c000000000000007100000000",
            INIT_30 => X"0000002c000000000000000d0000000000000010000000000000002e00000000",
            INIT_31 => X"00000008000000000000000b0000000000000019000000000000002d00000000",
            INIT_32 => X"0000000400000000000000020000000000000002000000000000000400000000",
            INIT_33 => X"0000001700000000000000130000000000000012000000000000000d00000000",
            INIT_34 => X"0000001f00000000000000210000000000000026000000000000001d00000000",
            INIT_35 => X"0000003a0000000000000032000000000000002c000000000000002600000000",
            INIT_36 => X"0000007b0000000000000073000000000000005a000000000000004600000000",
            INIT_37 => X"000000a0000000000000008b000000000000007b000000000000007300000000",
            INIT_38 => X"000000290000000000000013000000000000001b000000000000002900000000",
            INIT_39 => X"0000001f00000000000000320000000000000046000000000000005100000000",
            INIT_3A => X"0000000000000000000000020000000000000005000000000000000f00000000",
            INIT_3B => X"0000002400000000000000320000000000000040000000000000001100000000",
            INIT_3C => X"00000023000000000000001e000000000000001e000000000000001e00000000",
            INIT_3D => X"0000006100000000000000470000000000000037000000000000002b00000000",
            INIT_3E => X"0000006900000000000000780000000000000083000000000000007c00000000",
            INIT_3F => X"000000b300000000000000980000000000000086000000000000006f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000c000000000000000a000000000000000a000000000000000f00000000",
            INIT_41 => X"00000021000000000000002b0000000000000034000000000000002c00000000",
            INIT_42 => X"0000000100000000000000020000000000000004000000000000001200000000",
            INIT_43 => X"00000080000000000000009e0000000000000075000000000000000800000000",
            INIT_44 => X"0000006900000000000000670000000000000069000000000000007000000000",
            INIT_45 => X"0000007e000000000000007e0000000000000073000000000000006b00000000",
            INIT_46 => X"00000074000000000000005e0000000000000056000000000000006a00000000",
            INIT_47 => X"000000c200000000000000ac0000000000000093000000000000008200000000",
            INIT_48 => X"000000040000000000000003000000000000000a000000000000002800000000",
            INIT_49 => X"0000000a000000000000000c000000000000000c000000000000000600000000",
            INIT_4A => X"0000000200000000000000010000000000000001000000000000000600000000",
            INIT_4B => X"000000820000000000000080000000000000003a000000000000000000000000",
            INIT_4C => X"000000710000000000000077000000000000007b000000000000007f00000000",
            INIT_4D => X"00000042000000000000004b0000000000000060000000000000006e00000000",
            INIT_4E => X"000000840000000000000076000000000000005d000000000000004700000000",
            INIT_4F => X"000000c500000000000000b600000000000000a2000000000000008d00000000",
            INIT_50 => X"000000010000000000000001000000000000001d000000000000004d00000000",
            INIT_51 => X"0000000200000000000000030000000000000002000000000000000100000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_53 => X"0000002f000000000000002d000000000000000c000000000000000100000000",
            INIT_54 => X"0000003100000000000000320000000000000030000000000000002e00000000",
            INIT_55 => X"0000004d00000000000000300000000000000026000000000000002a00000000",
            INIT_56 => X"000000870000000000000080000000000000007e000000000000006e00000000",
            INIT_57 => X"000000c600000000000000bb00000000000000b0000000000000009900000000",
            INIT_58 => X"0000000100000000000000010000000000000034000000000000005e00000000",
            INIT_59 => X"0000000000000000000000010000000000000001000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000002000000000000000190000000000000003000000000000000200000000",
            INIT_5C => X"0000001d00000000000000190000000000000019000000000000001900000000",
            INIT_5D => X"00000071000000000000005c0000000000000042000000000000002900000000",
            INIT_5E => X"0000008b000000000000007f000000000000007e000000000000007c00000000",
            INIT_5F => X"000000c900000000000000bf00000000000000b3000000000000009d00000000",
            INIT_60 => X"000000020000000000000007000000000000003c000000000000006600000000",
            INIT_61 => X"0000000200000000000000030000000000000003000000000000000200000000",
            INIT_62 => X"0000000100000000000000000000000000000000000000000000000100000000",
            INIT_63 => X"0000001f00000000000000130000000000000001000000000000000300000000",
            INIT_64 => X"0000003a000000000000001b000000000000000d000000000000001100000000",
            INIT_65 => X"0000007c000000000000007e0000000000000073000000000000005a00000000",
            INIT_66 => X"0000009100000000000000870000000000000082000000000000007b00000000",
            INIT_67 => X"000000ca00000000000000c000000000000000b0000000000000009f00000000",
            INIT_68 => X"0000000c00000000000000170000000000000033000000000000006300000000",
            INIT_69 => X"00000007000000000000000a000000000000000b000000000000000a00000000",
            INIT_6A => X"0000000300000000000000040000000000000004000000000000000400000000",
            INIT_6B => X"00000015000000000000000d0000000000000005000000000000000600000000",
            INIT_6C => X"00000062000000000000004d0000000000000032000000000000001b00000000",
            INIT_6D => X"0000007d000000000000007e000000000000007e000000000000007100000000",
            INIT_6E => X"0000009a0000000000000094000000000000008a000000000000008000000000",
            INIT_6F => X"000000ca00000000000000c500000000000000b800000000000000a800000000",
            INIT_70 => X"00000023000000000000002c0000000000000039000000000000006000000000",
            INIT_71 => X"00000017000000000000001a000000000000001c000000000000001e00000000",
            INIT_72 => X"0000001700000000000000160000000000000015000000000000001500000000",
            INIT_73 => X"000000370000000000000028000000000000001f000000000000001b00000000",
            INIT_74 => X"0000007000000000000000660000000000000058000000000000004600000000",
            INIT_75 => X"0000007f000000000000007a000000000000007a000000000000007900000000",
            INIT_76 => X"000000a00000000000000095000000000000008b000000000000008500000000",
            INIT_77 => X"000000ca00000000000000c800000000000000bd00000000000000ac00000000",
            INIT_78 => X"0000003d0000000000000043000000000000004b000000000000006500000000",
            INIT_79 => X"0000003700000000000000350000000000000035000000000000003800000000",
            INIT_7A => X"0000003e000000000000003a0000000000000038000000000000003700000000",
            INIT_7B => X"0000006000000000000000540000000000000047000000000000004300000000",
            INIT_7C => X"000000790000000000000074000000000000006d000000000000006700000000",
            INIT_7D => X"00000083000000000000007d000000000000007c000000000000007f00000000",
            INIT_7E => X"000000a200000000000000980000000000000091000000000000008800000000",
            INIT_7F => X"000000c800000000000000c300000000000000b700000000000000ab00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE9;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE10 : if BRAM_NAME = "sampleifmap_layersamples_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e800000000000000e800000000000000e700000000000000eb00000000",
            INIT_01 => X"000000e800000000000000e800000000000000e800000000000000e800000000",
            INIT_02 => X"000000e900000000000000e900000000000000e800000000000000e800000000",
            INIT_03 => X"000000e900000000000000e900000000000000e900000000000000e900000000",
            INIT_04 => X"000000e800000000000000e900000000000000e900000000000000e900000000",
            INIT_05 => X"000000e600000000000000e800000000000000ea00000000000000ea00000000",
            INIT_06 => X"000000e800000000000000e800000000000000e900000000000000e700000000",
            INIT_07 => X"000000e800000000000000e900000000000000e900000000000000e800000000",
            INIT_08 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_09 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_0A => X"000000ec00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_0B => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_0C => X"000000ea00000000000000ea00000000000000e900000000000000e900000000",
            INIT_0D => X"000000eb00000000000000ed00000000000000ee00000000000000ed00000000",
            INIT_0E => X"000000eb00000000000000eb00000000000000ec00000000000000ea00000000",
            INIT_0F => X"000000eb00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_10 => X"000000ea00000000000000ea00000000000000ea00000000000000ed00000000",
            INIT_11 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_12 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_13 => X"000000ea00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_14 => X"000000ec00000000000000ea00000000000000e700000000000000e700000000",
            INIT_15 => X"000000ea00000000000000eb00000000000000ee00000000000000e900000000",
            INIT_16 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_17 => X"000000ea00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_18 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_19 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_1A => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_1B => X"000000ea00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_1C => X"000000e700000000000000e800000000000000e700000000000000e600000000",
            INIT_1D => X"000000e600000000000000d500000000000000db00000000000000c500000000",
            INIT_1E => X"000000ea00000000000000ea00000000000000ea00000000000000eb00000000",
            INIT_1F => X"000000eb00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_20 => X"000000eb00000000000000eb00000000000000ea00000000000000ed00000000",
            INIT_21 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_22 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_23 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_24 => X"000000db00000000000000e600000000000000ed00000000000000ec00000000",
            INIT_25 => X"000000e800000000000000dd00000000000000d000000000000000b300000000",
            INIT_26 => X"000000eb00000000000000eb00000000000000eb00000000000000ed00000000",
            INIT_27 => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_28 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_29 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_2A => X"000000ec00000000000000ec00000000000000eb00000000000000ea00000000",
            INIT_2B => X"000000e800000000000000ed00000000000000ea00000000000000ec00000000",
            INIT_2C => X"000000c800000000000000cf00000000000000d200000000000000da00000000",
            INIT_2D => X"000000e800000000000000dc00000000000000ca00000000000000bd00000000",
            INIT_2E => X"000000eb00000000000000eb00000000000000eb00000000000000ed00000000",
            INIT_2F => X"000000ed00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_30 => X"000000e600000000000000e700000000000000e400000000000000e500000000",
            INIT_31 => X"000000eb00000000000000eb00000000000000ec00000000000000e900000000",
            INIT_32 => X"000000ee00000000000000ed00000000000000ec00000000000000ec00000000",
            INIT_33 => X"000000e400000000000000ee00000000000000e500000000000000e600000000",
            INIT_34 => X"000000be00000000000000bf00000000000000be00000000000000cc00000000",
            INIT_35 => X"000000d300000000000000b100000000000000ab00000000000000b100000000",
            INIT_36 => X"000000eb00000000000000e900000000000000ea00000000000000ef00000000",
            INIT_37 => X"000000ee00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_38 => X"000000ea00000000000000ee00000000000000e900000000000000de00000000",
            INIT_39 => X"000000ec00000000000000eb00000000000000ec00000000000000ea00000000",
            INIT_3A => X"000000ef00000000000000ed00000000000000ee00000000000000ee00000000",
            INIT_3B => X"000000da00000000000000eb00000000000000dd00000000000000cb00000000",
            INIT_3C => X"000000cb00000000000000d300000000000000d200000000000000d200000000",
            INIT_3D => X"000000cc00000000000000b900000000000000bb00000000000000c400000000",
            INIT_3E => X"000000ee00000000000000ed00000000000000ee00000000000000f000000000",
            INIT_3F => X"000000ee00000000000000ee00000000000000ee00000000000000ee00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f300000000000000f600000000000000f300000000000000f100000000",
            INIT_41 => X"000000eb00000000000000eb00000000000000ed00000000000000f000000000",
            INIT_42 => X"000000ef00000000000000ed00000000000000ed00000000000000ed00000000",
            INIT_43 => X"000000e500000000000000e700000000000000da00000000000000c400000000",
            INIT_44 => X"000000e300000000000000eb00000000000000de00000000000000d900000000",
            INIT_45 => X"000000f100000000000000f000000000000000eb00000000000000ea00000000",
            INIT_46 => X"000000f000000000000000f000000000000000f000000000000000f300000000",
            INIT_47 => X"000000ee00000000000000ef00000000000000ef00000000000000ef00000000",
            INIT_48 => X"000000a100000000000000990000000000000094000000000000009500000000",
            INIT_49 => X"000000e800000000000000e900000000000000e900000000000000bf00000000",
            INIT_4A => X"000000eb00000000000000ec00000000000000eb00000000000000ea00000000",
            INIT_4B => X"000000ec00000000000000e800000000000000e200000000000000d600000000",
            INIT_4C => X"000000ef00000000000000f100000000000000eb00000000000000e800000000",
            INIT_4D => X"000000d300000000000000e200000000000000f300000000000000f700000000",
            INIT_4E => X"000000c900000000000000b900000000000000ba00000000000000c300000000",
            INIT_4F => X"000000ef00000000000000ef00000000000000ef00000000000000eb00000000",
            INIT_50 => X"0000008900000000000000890000000000000085000000000000008d00000000",
            INIT_51 => X"000000e000000000000000e100000000000000e700000000000000a500000000",
            INIT_52 => X"000000eb00000000000000ea00000000000000ea00000000000000e900000000",
            INIT_53 => X"000000ec00000000000000ee00000000000000ec00000000000000eb00000000",
            INIT_54 => X"000000ee00000000000000f100000000000000f000000000000000ee00000000",
            INIT_55 => X"000000a300000000000000ac00000000000000bf00000000000000d500000000",
            INIT_56 => X"000000a6000000000000008f0000000000000099000000000000009f00000000",
            INIT_57 => X"000000ef00000000000000ee00000000000000ef00000000000000e500000000",
            INIT_58 => X"000000df00000000000000e000000000000000d700000000000000e000000000",
            INIT_59 => X"000000ce00000000000000d300000000000000e700000000000000e300000000",
            INIT_5A => X"000000db00000000000000e100000000000000de00000000000000d600000000",
            INIT_5B => X"000000e900000000000000e600000000000000e100000000000000df00000000",
            INIT_5C => X"000000ed00000000000000f100000000000000ef00000000000000ed00000000",
            INIT_5D => X"000000ca00000000000000cf00000000000000cb00000000000000d000000000",
            INIT_5E => X"000000ca00000000000000a400000000000000c400000000000000d300000000",
            INIT_5F => X"000000ef00000000000000ef00000000000000ee00000000000000e900000000",
            INIT_60 => X"000000ea00000000000000e000000000000000d900000000000000de00000000",
            INIT_61 => X"000000ae00000000000000d000000000000000e300000000000000f100000000",
            INIT_62 => X"0000007900000000000000bc00000000000000d600000000000000b700000000",
            INIT_63 => X"00000093000000000000008b0000000000000084000000000000007e00000000",
            INIT_64 => X"000000ed00000000000000dc00000000000000ae00000000000000a100000000",
            INIT_65 => X"000000e900000000000000f000000000000000ee00000000000000eb00000000",
            INIT_66 => X"000000ed00000000000000d400000000000000e500000000000000ed00000000",
            INIT_67 => X"000000f200000000000000f200000000000000e900000000000000ea00000000",
            INIT_68 => X"00000097000000000000008d0000000000000093000000000000009800000000",
            INIT_69 => X"000000cc00000000000000cd00000000000000c100000000000000a500000000",
            INIT_6A => X"0000005c00000000000000b700000000000000ea00000000000000e200000000",
            INIT_6B => X"00000062000000000000005a000000000000005b000000000000005b00000000",
            INIT_6C => X"000000f100000000000000e900000000000000b3000000000000008100000000",
            INIT_6D => X"000000d900000000000000e900000000000000ed00000000000000f100000000",
            INIT_6E => X"000000d600000000000000df00000000000000dc00000000000000d400000000",
            INIT_6F => X"000000ea00000000000000e300000000000000cd00000000000000c400000000",
            INIT_70 => X"0000006600000000000000640000000000000072000000000000006c00000000",
            INIT_71 => X"000000cf00000000000000a400000000000000a4000000000000009b00000000",
            INIT_72 => X"0000008a00000000000000be00000000000000e400000000000000ea00000000",
            INIT_73 => X"000000cf00000000000000a80000000000000087000000000000008300000000",
            INIT_74 => X"000000d400000000000000e300000000000000e800000000000000df00000000",
            INIT_75 => X"0000009300000000000000a300000000000000ae00000000000000c300000000",
            INIT_76 => X"0000009700000000000000980000000000000090000000000000008c00000000",
            INIT_77 => X"000000d800000000000000cb00000000000000a0000000000000009300000000",
            INIT_78 => X"000000990000000000000074000000000000005e000000000000004d00000000",
            INIT_79 => X"000000a10000000000000076000000000000006e000000000000009c00000000",
            INIT_7A => X"000000c800000000000000c600000000000000c500000000000000b600000000",
            INIT_7B => X"000000d900000000000000ec00000000000000d900000000000000ca00000000",
            INIT_7C => X"00000095000000000000009f00000000000000ac00000000000000ba00000000",
            INIT_7D => X"0000007b0000000000000076000000000000007b000000000000008a00000000",
            INIT_7E => X"000000a100000000000000910000000000000082000000000000008000000000",
            INIT_7F => X"000000d000000000000000d500000000000000b800000000000000ae00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE10;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE11 : if BRAM_NAME = "sampleifmap_layersamples_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000dc0000000000000097000000000000002f000000000000002300000000",
            INIT_01 => X"000000a20000000000000086000000000000007b000000000000009600000000",
            INIT_02 => X"000000e900000000000000e100000000000000d300000000000000b400000000",
            INIT_03 => X"000000be00000000000000ee00000000000000f000000000000000e800000000",
            INIT_04 => X"000000b100000000000000aa00000000000000a200000000000000a300000000",
            INIT_05 => X"000000bb00000000000000b600000000000000b600000000000000bb00000000",
            INIT_06 => X"000000d900000000000000cc00000000000000bf00000000000000bd00000000",
            INIT_07 => X"000000b700000000000000c100000000000000d000000000000000da00000000",
            INIT_08 => X"000000ef00000000000000d9000000000000004f000000000000001800000000",
            INIT_09 => X"000000e500000000000000da00000000000000d300000000000000d400000000",
            INIT_0A => X"000000ef00000000000000f500000000000000f600000000000000ed00000000",
            INIT_0B => X"000000ea00000000000000f100000000000000ef00000000000000dc00000000",
            INIT_0C => X"000000e500000000000000e600000000000000d600000000000000e400000000",
            INIT_0D => X"000000e000000000000000e800000000000000ea00000000000000e700000000",
            INIT_0E => X"000000b300000000000000c500000000000000d100000000000000d400000000",
            INIT_0F => X"000000a5000000000000009e00000000000000a100000000000000a900000000",
            INIT_10 => X"000000d800000000000000de00000000000000b3000000000000004700000000",
            INIT_11 => X"000000e300000000000000e600000000000000e500000000000000d900000000",
            INIT_12 => X"000000dd00000000000000e400000000000000e400000000000000e300000000",
            INIT_13 => X"000000bc00000000000000c100000000000000d700000000000000cf00000000",
            INIT_14 => X"0000009c00000000000000ba00000000000000c300000000000000b800000000",
            INIT_15 => X"0000009e00000000000000ad00000000000000b400000000000000a100000000",
            INIT_16 => X"0000008300000000000000850000000000000087000000000000008a00000000",
            INIT_17 => X"0000009c000000000000009e0000000000000097000000000000008c00000000",
            INIT_18 => X"000000bd00000000000000c200000000000000cf00000000000000a100000000",
            INIT_19 => X"000000c100000000000000c000000000000000be00000000000000bb00000000",
            INIT_1A => X"000000bd00000000000000bd00000000000000be00000000000000c000000000",
            INIT_1B => X"0000009a00000000000000a300000000000000ba00000000000000bc00000000",
            INIT_1C => X"0000009100000000000000a300000000000000aa000000000000009a00000000",
            INIT_1D => X"0000008800000000000000900000000000000099000000000000009400000000",
            INIT_1E => X"0000008d000000000000008b0000000000000086000000000000008200000000",
            INIT_1F => X"0000009c00000000000000940000000000000092000000000000009000000000",
            INIT_20 => X"0000007f000000000000007a0000000000000071000000000000006d00000000",
            INIT_21 => X"000000960000000000000093000000000000008e000000000000008600000000",
            INIT_22 => X"000000ac00000000000000a500000000000000a0000000000000009800000000",
            INIT_23 => X"000000af00000000000000b400000000000000ba00000000000000b500000000",
            INIT_24 => X"0000009b00000000000000a300000000000000a800000000000000ac00000000",
            INIT_25 => X"0000007f0000000000000084000000000000008b000000000000009400000000",
            INIT_26 => X"0000007a00000000000000810000000000000085000000000000008100000000",
            INIT_27 => X"0000009c0000000000000092000000000000008a000000000000007e00000000",
            INIT_28 => X"0000003000000000000000230000000000000019000000000000002900000000",
            INIT_29 => X"0000003d000000000000003a0000000000000038000000000000003400000000",
            INIT_2A => X"00000057000000000000004d0000000000000046000000000000003e00000000",
            INIT_2B => X"0000007e000000000000007e0000000000000079000000000000006a00000000",
            INIT_2C => X"000000700000000000000078000000000000007e000000000000007f00000000",
            INIT_2D => X"0000006600000000000000670000000000000068000000000000006a00000000",
            INIT_2E => X"000000770000000000000073000000000000006e000000000000006900000000",
            INIT_2F => X"00000095000000000000008d0000000000000088000000000000008000000000",
            INIT_30 => X"0000003500000000000000130000000000000014000000000000003700000000",
            INIT_31 => X"00000018000000000000001e0000000000000029000000000000003a00000000",
            INIT_32 => X"00000014000000000000000f000000000000000f000000000000001100000000",
            INIT_33 => X"0000003e000000000000003c0000000000000038000000000000002a00000000",
            INIT_34 => X"0000004c000000000000004d0000000000000051000000000000004700000000",
            INIT_35 => X"0000005a0000000000000053000000000000004f000000000000004e00000000",
            INIT_36 => X"0000008a000000000000008a0000000000000076000000000000006500000000",
            INIT_37 => X"0000009e00000000000000890000000000000080000000000000007d00000000",
            INIT_38 => X"000000290000000000000012000000000000001a000000000000002d00000000",
            INIT_39 => X"000000250000000000000039000000000000004c000000000000005400000000",
            INIT_3A => X"000000070000000000000007000000000000000b000000000000001500000000",
            INIT_3B => X"0000003e000000000000004e000000000000005b000000000000002300000000",
            INIT_3C => X"00000045000000000000003f000000000000003e000000000000003c00000000",
            INIT_3D => X"0000007b00000000000000630000000000000053000000000000004a00000000",
            INIT_3E => X"0000007200000000000000870000000000000095000000000000009200000000",
            INIT_3F => X"000000af00000000000000920000000000000085000000000000007400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000b00000000000000080000000000000009000000000000001100000000",
            INIT_41 => X"00000023000000000000002f0000000000000039000000000000002e00000000",
            INIT_42 => X"0000000300000000000000040000000000000007000000000000001400000000",
            INIT_43 => X"0000009400000000000000b30000000000000086000000000000000f00000000",
            INIT_44 => X"0000007f000000000000007c000000000000007d000000000000008300000000",
            INIT_45 => X"0000008d00000000000000900000000000000085000000000000007e00000000",
            INIT_46 => X"000000740000000000000061000000000000005b000000000000007400000000",
            INIT_47 => X"000000be00000000000000a50000000000000090000000000000008100000000",
            INIT_48 => X"0000000400000000000000030000000000000007000000000000002300000000",
            INIT_49 => X"0000000c00000000000000110000000000000011000000000000000700000000",
            INIT_4A => X"0000000300000000000000020000000000000003000000000000000700000000",
            INIT_4B => X"0000009400000000000000920000000000000040000000000000000200000000",
            INIT_4C => X"000000810000000000000089000000000000008d000000000000009000000000",
            INIT_4D => X"000000450000000000000053000000000000006a000000000000007a00000000",
            INIT_4E => X"0000007e00000000000000710000000000000058000000000000004600000000",
            INIT_4F => X"000000c200000000000000b0000000000000009e000000000000008700000000",
            INIT_50 => X"0000000200000000000000010000000000000015000000000000004000000000",
            INIT_51 => X"0000000500000000000000090000000000000005000000000000000000000000",
            INIT_52 => X"0000000100000000000000000000000000000000000000000000000200000000",
            INIT_53 => X"00000044000000000000003b000000000000000b000000000000000100000000",
            INIT_54 => X"0000003b00000000000000430000000000000045000000000000004300000000",
            INIT_55 => X"00000047000000000000002e000000000000002a000000000000003100000000",
            INIT_56 => X"0000008000000000000000780000000000000074000000000000006600000000",
            INIT_57 => X"000000c400000000000000b700000000000000ab000000000000009300000000",
            INIT_58 => X"000000020000000000000001000000000000002b000000000000005200000000",
            INIT_59 => X"0000000200000000000000050000000000000002000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000003600000000000000260000000000000002000000000000000000000000",
            INIT_5C => X"000000220000000000000024000000000000002b000000000000002e00000000",
            INIT_5D => X"0000006900000000000000520000000000000038000000000000002700000000",
            INIT_5E => X"0000008300000000000000760000000000000073000000000000007300000000",
            INIT_5F => X"000000c700000000000000bb00000000000000ae000000000000009600000000",
            INIT_60 => X"0000000100000000000000030000000000000032000000000000005d00000000",
            INIT_61 => X"0000000200000000000000030000000000000001000000000000000000000000",
            INIT_62 => X"0000000100000000000000000000000000000000000000000000000100000000",
            INIT_63 => X"0000002f000000000000001c0000000000000000000000000000000200000000",
            INIT_64 => X"000000370000000000000016000000000000000c000000000000001700000000",
            INIT_65 => X"00000070000000000000006f0000000000000063000000000000005100000000",
            INIT_66 => X"00000089000000000000007e0000000000000077000000000000007100000000",
            INIT_67 => X"000000c900000000000000bc00000000000000ab000000000000009700000000",
            INIT_68 => X"00000004000000000000000b0000000000000025000000000000005900000000",
            INIT_69 => X"0000000200000000000000040000000000000004000000000000000200000000",
            INIT_6A => X"0000000200000000000000010000000000000001000000000000000100000000",
            INIT_6B => X"00000018000000000000000d0000000000000002000000000000000600000000",
            INIT_6C => X"00000052000000000000003e0000000000000029000000000000001900000000",
            INIT_6D => X"0000006f00000000000000700000000000000071000000000000006500000000",
            INIT_6E => X"000000910000000000000089000000000000007e000000000000007300000000",
            INIT_6F => X"000000c900000000000000c100000000000000b300000000000000a100000000",
            INIT_70 => X"0000001100000000000000160000000000000024000000000000005200000000",
            INIT_71 => X"0000000c000000000000000d000000000000000f000000000000000f00000000",
            INIT_72 => X"0000000f000000000000000e000000000000000d000000000000000c00000000",
            INIT_73 => X"0000002d000000000000001b0000000000000015000000000000001400000000",
            INIT_74 => X"0000005800000000000000550000000000000051000000000000004300000000",
            INIT_75 => X"00000070000000000000006b000000000000006e000000000000006900000000",
            INIT_76 => X"00000097000000000000008a000000000000007f000000000000007700000000",
            INIT_77 => X"000000c800000000000000c400000000000000b700000000000000a400000000",
            INIT_78 => X"0000002500000000000000260000000000000030000000000000005300000000",
            INIT_79 => X"0000002600000000000000220000000000000021000000000000002300000000",
            INIT_7A => X"0000002e000000000000002c0000000000000029000000000000002800000000",
            INIT_7B => X"0000004a000000000000003b0000000000000030000000000000002d00000000",
            INIT_7C => X"000000610000000000000061000000000000005c000000000000005300000000",
            INIT_7D => X"00000075000000000000006c000000000000006a000000000000006b00000000",
            INIT_7E => X"00000099000000000000008d0000000000000085000000000000007b00000000",
            INIT_7F => X"000000c700000000000000bf00000000000000b200000000000000a300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE11;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE12 : if BRAM_NAME = "sampleifmap_layersamples_instance12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000084000000000000008b000000000000009e000000000000009e00000000",
            INIT_01 => X"000000c100000000000000bb00000000000000b600000000000000a600000000",
            INIT_02 => X"000000ce00000000000000d100000000000000cd00000000000000c700000000",
            INIT_03 => X"000000e600000000000000e300000000000000df00000000000000da00000000",
            INIT_04 => X"000000eb00000000000000e700000000000000e200000000000000d500000000",
            INIT_05 => X"000000ea00000000000000ea00000000000000e800000000000000ec00000000",
            INIT_06 => X"000000ee00000000000000e600000000000000e200000000000000ec00000000",
            INIT_07 => X"000000ee00000000000000ed00000000000000e400000000000000e800000000",
            INIT_08 => X"00000089000000000000009700000000000000ac00000000000000aa00000000",
            INIT_09 => X"000000c700000000000000c500000000000000c100000000000000ae00000000",
            INIT_0A => X"000000d200000000000000d900000000000000d700000000000000ce00000000",
            INIT_0B => X"000000ed00000000000000e900000000000000e700000000000000e100000000",
            INIT_0C => X"000000f200000000000000e800000000000000e400000000000000db00000000",
            INIT_0D => X"000000f200000000000000ec00000000000000ea00000000000000f500000000",
            INIT_0E => X"000000f300000000000000eb00000000000000e400000000000000f100000000",
            INIT_0F => X"000000f600000000000000f600000000000000e800000000000000e900000000",
            INIT_10 => X"0000008e000000000000009d00000000000000b000000000000000ae00000000",
            INIT_11 => X"000000c700000000000000ce00000000000000c900000000000000b500000000",
            INIT_12 => X"000000d400000000000000da00000000000000df00000000000000d100000000",
            INIT_13 => X"000000ef00000000000000e600000000000000e600000000000000e000000000",
            INIT_14 => X"000000ef00000000000000e900000000000000e400000000000000dd00000000",
            INIT_15 => X"000000f300000000000000ec00000000000000d500000000000000e800000000",
            INIT_16 => X"000000f800000000000000ee00000000000000e700000000000000f500000000",
            INIT_17 => X"000000f500000000000000fa00000000000000e600000000000000ed00000000",
            INIT_18 => X"0000009300000000000000a000000000000000b200000000000000b400000000",
            INIT_19 => X"000000cf00000000000000d400000000000000cb00000000000000ba00000000",
            INIT_1A => X"000000d600000000000000dd00000000000000e400000000000000d600000000",
            INIT_1B => X"000000f000000000000000df00000000000000e700000000000000dc00000000",
            INIT_1C => X"000000e400000000000000e900000000000000e400000000000000e000000000",
            INIT_1D => X"000000f300000000000000e600000000000000ac00000000000000b100000000",
            INIT_1E => X"000000fa00000000000000ee00000000000000e800000000000000f800000000",
            INIT_1F => X"000000f400000000000000f900000000000000e400000000000000ee00000000",
            INIT_20 => X"0000009300000000000000a500000000000000b900000000000000ba00000000",
            INIT_21 => X"000000cf00000000000000d900000000000000cc00000000000000bd00000000",
            INIT_22 => X"000000d600000000000000de00000000000000e700000000000000d300000000",
            INIT_23 => X"000000eb00000000000000d300000000000000e700000000000000da00000000",
            INIT_24 => X"000000d400000000000000e800000000000000e000000000000000e200000000",
            INIT_25 => X"000000ed00000000000000e000000000000000a8000000000000009f00000000",
            INIT_26 => X"000000f600000000000000eb00000000000000e700000000000000f700000000",
            INIT_27 => X"000000f200000000000000f800000000000000ea00000000000000e800000000",
            INIT_28 => X"0000008e00000000000000aa00000000000000be00000000000000c100000000",
            INIT_29 => X"000000d300000000000000db00000000000000cb00000000000000bf00000000",
            INIT_2A => X"000000d600000000000000dd00000000000000ea00000000000000d700000000",
            INIT_2B => X"000000cd00000000000000c700000000000000e400000000000000d600000000",
            INIT_2C => X"000000c100000000000000eb00000000000000ce00000000000000cf00000000",
            INIT_2D => X"000000e600000000000000de000000000000009e000000000000007000000000",
            INIT_2E => X"000000f100000000000000e200000000000000e500000000000000f500000000",
            INIT_2F => X"000000eb00000000000000f300000000000000e700000000000000e400000000",
            INIT_30 => X"0000008500000000000000ac00000000000000bf00000000000000c400000000",
            INIT_31 => X"000000d900000000000000de00000000000000ca00000000000000bf00000000",
            INIT_32 => X"000000d600000000000000da00000000000000eb00000000000000df00000000",
            INIT_33 => X"000000b000000000000000bc00000000000000e300000000000000d700000000",
            INIT_34 => X"000000bb00000000000000cd00000000000000ba00000000000000bb00000000",
            INIT_35 => X"000000b700000000000000ac0000000000000089000000000000007800000000",
            INIT_36 => X"000000eb00000000000000d800000000000000df00000000000000db00000000",
            INIT_37 => X"000000eb00000000000000f000000000000000e100000000000000e200000000",
            INIT_38 => X"0000008c00000000000000ae00000000000000c500000000000000cc00000000",
            INIT_39 => X"000000e000000000000000e000000000000000da00000000000000cb00000000",
            INIT_3A => X"000000dc00000000000000dc00000000000000ed00000000000000e800000000",
            INIT_3B => X"000000cd00000000000000c900000000000000dd00000000000000dc00000000",
            INIT_3C => X"000000530000000000000064000000000000008a00000000000000ac00000000",
            INIT_3D => X"0000003c0000000000000041000000000000003e000000000000004700000000",
            INIT_3E => X"000000e400000000000000d100000000000000b6000000000000006800000000",
            INIT_3F => X"000000ec00000000000000ef00000000000000d400000000000000da00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000089000000000000009d00000000000000aa00000000000000af00000000",
            INIT_41 => X"000000c500000000000000af00000000000000ba00000000000000b000000000",
            INIT_42 => X"000000d200000000000000ce00000000000000d400000000000000d100000000",
            INIT_43 => X"000000c100000000000000c100000000000000c900000000000000d400000000",
            INIT_44 => X"0000005b00000000000000590000000000000069000000000000008e00000000",
            INIT_45 => X"00000045000000000000005e0000000000000053000000000000005400000000",
            INIT_46 => X"000000b700000000000000a20000000000000079000000000000004e00000000",
            INIT_47 => X"000000c300000000000000cf00000000000000a300000000000000ae00000000",
            INIT_48 => X"0000006800000000000000710000000000000073000000000000007200000000",
            INIT_49 => X"00000080000000000000006f000000000000006b000000000000006900000000",
            INIT_4A => X"0000009b00000000000000970000000000000092000000000000008b00000000",
            INIT_4B => X"0000009600000000000000970000000000000093000000000000009d00000000",
            INIT_4C => X"0000006300000000000000630000000000000064000000000000007600000000",
            INIT_4D => X"0000005300000000000000560000000000000056000000000000005500000000",
            INIT_4E => X"00000099000000000000009a0000000000000080000000000000008b00000000",
            INIT_4F => X"0000007b0000000000000084000000000000006d000000000000007600000000",
            INIT_50 => X"00000044000000000000004b000000000000004c000000000000004200000000",
            INIT_51 => X"0000005a0000000000000054000000000000005a000000000000005300000000",
            INIT_52 => X"000000670000000000000066000000000000006a000000000000005d00000000",
            INIT_53 => X"0000006c0000000000000072000000000000006b000000000000006a00000000",
            INIT_54 => X"00000055000000000000005b000000000000005a000000000000005a00000000",
            INIT_55 => X"00000072000000000000005f0000000000000042000000000000004800000000",
            INIT_56 => X"000000c70000000000000093000000000000006e000000000000008000000000",
            INIT_57 => X"0000005e000000000000005c0000000000000067000000000000007d00000000",
            INIT_58 => X"0000004d000000000000004b0000000000000041000000000000003500000000",
            INIT_59 => X"000000460000000000000055000000000000006a000000000000006f00000000",
            INIT_5A => X"0000005d000000000000005f0000000000000071000000000000005d00000000",
            INIT_5B => X"00000061000000000000006b0000000000000073000000000000006c00000000",
            INIT_5C => X"000000610000000000000062000000000000005f000000000000006200000000",
            INIT_5D => X"000000bb00000000000000950000000000000055000000000000005a00000000",
            INIT_5E => X"000000cc0000000000000070000000000000009200000000000000b300000000",
            INIT_5F => X"000000550000000000000057000000000000005f000000000000009a00000000",
            INIT_60 => X"0000004a000000000000005e0000000000000056000000000000003a00000000",
            INIT_61 => X"00000055000000000000004d0000000000000064000000000000006400000000",
            INIT_62 => X"0000006c000000000000007f0000000000000085000000000000007800000000",
            INIT_63 => X"000000570000000000000062000000000000006e000000000000006900000000",
            INIT_64 => X"0000005f00000000000000570000000000000051000000000000005100000000",
            INIT_65 => X"000000c300000000000000aa0000000000000070000000000000005f00000000",
            INIT_66 => X"000000ad000000000000007f00000000000000c100000000000000d000000000",
            INIT_67 => X"0000004f0000000000000055000000000000005000000000000000b200000000",
            INIT_68 => X"0000004b00000000000000570000000000000059000000000000004a00000000",
            INIT_69 => X"0000005000000000000000470000000000000044000000000000005200000000",
            INIT_6A => X"0000006f00000000000000760000000000000067000000000000005900000000",
            INIT_6B => X"000000620000000000000069000000000000006a000000000000006500000000",
            INIT_6C => X"0000006d00000000000000620000000000000062000000000000006000000000",
            INIT_6D => X"000000b800000000000000b4000000000000008e000000000000007200000000",
            INIT_6E => X"0000008400000000000000a000000000000000c000000000000000bf00000000",
            INIT_6F => X"00000043000000000000003c000000000000005000000000000000aa00000000",
            INIT_70 => X"0000004e0000000000000052000000000000004f000000000000004d00000000",
            INIT_71 => X"0000005600000000000000460000000000000048000000000000004f00000000",
            INIT_72 => X"0000008500000000000000810000000000000079000000000000006d00000000",
            INIT_73 => X"0000008300000000000000870000000000000088000000000000008900000000",
            INIT_74 => X"0000009600000000000000920000000000000094000000000000009200000000",
            INIT_75 => X"000000b500000000000000b300000000000000a3000000000000009400000000",
            INIT_76 => X"0000006500000000000000aa00000000000000b000000000000000b900000000",
            INIT_77 => X"0000003b00000000000000370000000000000049000000000000005a00000000",
            INIT_78 => X"00000068000000000000006a000000000000005e000000000000006000000000",
            INIT_79 => X"0000008a00000000000000840000000000000083000000000000006d00000000",
            INIT_7A => X"0000009a000000000000009b0000000000000098000000000000009000000000",
            INIT_7B => X"00000094000000000000009e000000000000009b000000000000009b00000000",
            INIT_7C => X"00000092000000000000009c000000000000009d000000000000009600000000",
            INIT_7D => X"000000a900000000000000920000000000000082000000000000007700000000",
            INIT_7E => X"0000006900000000000000a700000000000000a800000000000000b100000000",
            INIT_7F => X"0000004800000000000000560000000000000062000000000000004500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE12;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE13 : if BRAM_NAME = "sampleifmap_layersamples_instance13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000008300000000000000730000000000000065000000000000006a00000000",
            INIT_01 => X"0000008f00000000000000900000000000000087000000000000008100000000",
            INIT_02 => X"0000009a000000000000009a0000000000000096000000000000009200000000",
            INIT_03 => X"0000009000000000000000970000000000000099000000000000009a00000000",
            INIT_04 => X"0000007f000000000000008b0000000000000086000000000000008200000000",
            INIT_05 => X"0000009f00000000000000920000000000000075000000000000005e00000000",
            INIT_06 => X"0000008400000000000000a200000000000000a300000000000000a700000000",
            INIT_07 => X"00000069000000000000009a00000000000000c0000000000000009000000000",
            INIT_08 => X"0000006d0000000000000076000000000000006c000000000000005f00000000",
            INIT_09 => X"000000910000000000000081000000000000005d000000000000005f00000000",
            INIT_0A => X"0000009000000000000000960000000000000097000000000000009500000000",
            INIT_0B => X"0000007b000000000000007a000000000000007e000000000000008600000000",
            INIT_0C => X"00000094000000000000009b0000000000000085000000000000007a00000000",
            INIT_0D => X"0000009c00000000000000a20000000000000093000000000000008300000000",
            INIT_0E => X"0000009500000000000000990000000000000097000000000000009d00000000",
            INIT_0F => X"00000094000000000000009d00000000000000a4000000000000009f00000000",
            INIT_10 => X"0000004600000000000000490000000000000059000000000000006600000000",
            INIT_11 => X"0000008c000000000000007b000000000000006f000000000000005600000000",
            INIT_12 => X"0000007500000000000000780000000000000081000000000000008f00000000",
            INIT_13 => X"0000008d0000000000000085000000000000007e000000000000007800000000",
            INIT_14 => X"0000009f0000000000000099000000000000008e000000000000009600000000",
            INIT_15 => X"000000a100000000000000a5000000000000009d000000000000009700000000",
            INIT_16 => X"00000090000000000000009a0000000000000098000000000000009900000000",
            INIT_17 => X"00000095000000000000007d0000000000000079000000000000008300000000",
            INIT_18 => X"0000006e0000000000000047000000000000003d000000000000005600000000",
            INIT_19 => X"0000007b0000000000000082000000000000008a000000000000008000000000",
            INIT_1A => X"000000840000000000000076000000000000006c000000000000007600000000",
            INIT_1B => X"00000099000000000000009c0000000000000098000000000000008f00000000",
            INIT_1C => X"0000009a00000000000000910000000000000089000000000000009500000000",
            INIT_1D => X"000000a400000000000000a0000000000000009a000000000000009900000000",
            INIT_1E => X"00000069000000000000007d0000000000000090000000000000009800000000",
            INIT_1F => X"000000840000000000000056000000000000004b000000000000005c00000000",
            INIT_20 => X"00000072000000000000006b0000000000000067000000000000006800000000",
            INIT_21 => X"00000076000000000000007b0000000000000074000000000000007300000000",
            INIT_22 => X"00000090000000000000008d0000000000000086000000000000007400000000",
            INIT_23 => X"000000750000000000000085000000000000008d000000000000008f00000000",
            INIT_24 => X"0000009600000000000000820000000000000059000000000000006200000000",
            INIT_25 => X"000000910000000000000098000000000000009a000000000000009700000000",
            INIT_26 => X"00000050000000000000005a0000000000000060000000000000007500000000",
            INIT_27 => X"0000004100000000000000490000000000000047000000000000004100000000",
            INIT_28 => X"0000006f000000000000006f000000000000006b000000000000006300000000",
            INIT_29 => X"0000007e000000000000007d0000000000000077000000000000007200000000",
            INIT_2A => X"00000081000000000000007d000000000000007d000000000000007500000000",
            INIT_2B => X"0000003d000000000000005b0000000000000082000000000000008300000000",
            INIT_2C => X"0000009400000000000000730000000000000038000000000000003900000000",
            INIT_2D => X"0000005f00000000000000720000000000000082000000000000008b00000000",
            INIT_2E => X"0000003a00000000000000490000000000000053000000000000005600000000",
            INIT_2F => X"0000001b0000000000000033000000000000004b000000000000003c00000000",
            INIT_30 => X"0000007200000000000000740000000000000068000000000000003e00000000",
            INIT_31 => X"0000005b00000000000000660000000000000075000000000000007400000000",
            INIT_32 => X"00000070000000000000004e0000000000000051000000000000005400000000",
            INIT_33 => X"0000004c00000000000000600000000000000082000000000000008500000000",
            INIT_34 => X"0000006c000000000000006b0000000000000056000000000000005300000000",
            INIT_35 => X"0000005100000000000000530000000000000058000000000000006000000000",
            INIT_36 => X"0000002d0000000000000033000000000000003d000000000000004600000000",
            INIT_37 => X"00000018000000000000001e000000000000002e000000000000003400000000",
            INIT_38 => X"00000069000000000000006a0000000000000060000000000000003900000000",
            INIT_39 => X"0000003500000000000000410000000000000068000000000000006b00000000",
            INIT_3A => X"0000006e00000000000000440000000000000040000000000000003b00000000",
            INIT_3B => X"0000006200000000000000730000000000000085000000000000008700000000",
            INIT_3C => X"00000050000000000000004e000000000000004f000000000000005800000000",
            INIT_3D => X"0000003700000000000000460000000000000050000000000000005100000000",
            INIT_3E => X"00000029000000000000002d0000000000000031000000000000002c00000000",
            INIT_3F => X"00000018000000000000001b000000000000001e000000000000002200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000690000000000000068000000000000005a000000000000004100000000",
            INIT_41 => X"00000049000000000000004f000000000000006d000000000000006d00000000",
            INIT_42 => X"0000006a00000000000000620000000000000058000000000000005500000000",
            INIT_43 => X"0000004100000000000000440000000000000053000000000000006200000000",
            INIT_44 => X"000000520000000000000051000000000000004a000000000000004600000000",
            INIT_45 => X"0000002c00000000000000290000000000000033000000000000004800000000",
            INIT_46 => X"0000002300000000000000270000000000000037000000000000003d00000000",
            INIT_47 => X"00000019000000000000001b000000000000001e000000000000002000000000",
            INIT_48 => X"0000006700000000000000690000000000000057000000000000004300000000",
            INIT_49 => X"0000005100000000000000580000000000000063000000000000006600000000",
            INIT_4A => X"00000039000000000000003b0000000000000045000000000000004c00000000",
            INIT_4B => X"000000460000000000000042000000000000003f000000000000003a00000000",
            INIT_4C => X"00000036000000000000003e0000000000000044000000000000004800000000",
            INIT_4D => X"0000002c0000000000000031000000000000002f000000000000002e00000000",
            INIT_4E => X"0000001c000000000000001e000000000000002e000000000000003800000000",
            INIT_4F => X"0000001e00000000000000180000000000000019000000000000001d00000000",
            INIT_50 => X"0000003a0000000000000041000000000000003a000000000000003600000000",
            INIT_51 => X"0000002c000000000000002d0000000000000032000000000000003700000000",
            INIT_52 => X"0000003a00000000000000370000000000000033000000000000002e00000000",
            INIT_53 => X"0000003a000000000000003e0000000000000040000000000000003e00000000",
            INIT_54 => X"0000003000000000000000250000000000000026000000000000003300000000",
            INIT_55 => X"00000026000000000000002a0000000000000030000000000000003100000000",
            INIT_56 => X"0000001c000000000000001b0000000000000020000000000000002900000000",
            INIT_57 => X"0000001f000000000000001c0000000000000019000000000000001b00000000",
            INIT_58 => X"0000001b000000000000001a000000000000001d000000000000001e00000000",
            INIT_59 => X"0000002700000000000000210000000000000020000000000000001f00000000",
            INIT_5A => X"0000003300000000000000350000000000000034000000000000003100000000",
            INIT_5B => X"0000002800000000000000260000000000000028000000000000002e00000000",
            INIT_5C => X"000000370000000000000042000000000000002c000000000000002600000000",
            INIT_5D => X"0000002500000000000000240000000000000025000000000000002900000000",
            INIT_5E => X"0000001b000000000000001a000000000000001b000000000000001f00000000",
            INIT_5F => X"000000170000000000000021000000000000001e000000000000001c00000000",
            INIT_60 => X"0000001c000000000000001b000000000000001f000000000000002100000000",
            INIT_61 => X"00000020000000000000001f000000000000001e000000000000001c00000000",
            INIT_62 => X"0000001e000000000000001e0000000000000021000000000000002300000000",
            INIT_63 => X"0000002d00000000000000290000000000000027000000000000002200000000",
            INIT_64 => X"0000003100000000000000490000000000000034000000000000002a00000000",
            INIT_65 => X"0000002000000000000000260000000000000023000000000000001e00000000",
            INIT_66 => X"0000001d000000000000001b000000000000001a000000000000001b00000000",
            INIT_67 => X"0000000d000000000000001a0000000000000026000000000000001e00000000",
            INIT_68 => X"0000001a000000000000001a000000000000001e000000000000001f00000000",
            INIT_69 => X"0000001b000000000000001a0000000000000019000000000000001900000000",
            INIT_6A => X"0000002800000000000000250000000000000020000000000000001d00000000",
            INIT_6B => X"0000002a00000000000000280000000000000029000000000000002a00000000",
            INIT_6C => X"000000260000000000000040000000000000002e000000000000002700000000",
            INIT_6D => X"0000001d000000000000001e0000000000000024000000000000001c00000000",
            INIT_6E => X"0000001c000000000000001b0000000000000019000000000000001a00000000",
            INIT_6F => X"0000000400000000000000090000000000000025000000000000002100000000",
            INIT_70 => X"0000001c0000000000000019000000000000001b000000000000001700000000",
            INIT_71 => X"0000002500000000000000220000000000000020000000000000001e00000000",
            INIT_72 => X"0000002700000000000000280000000000000027000000000000002700000000",
            INIT_73 => X"00000021000000000000001e0000000000000023000000000000002600000000",
            INIT_74 => X"0000002400000000000000390000000000000024000000000000001c00000000",
            INIT_75 => X"0000001d000000000000001d000000000000001d000000000000001e00000000",
            INIT_76 => X"0000001b00000000000000170000000000000018000000000000001800000000",
            INIT_77 => X"0000000500000000000000040000000000000013000000000000002400000000",
            INIT_78 => X"000000220000000000000020000000000000001e000000000000001c00000000",
            INIT_79 => X"0000002500000000000000230000000000000022000000000000002100000000",
            INIT_7A => X"0000002200000000000000240000000000000026000000000000002600000000",
            INIT_7B => X"0000000c000000000000000f0000000000000018000000000000001e00000000",
            INIT_7C => X"00000020000000000000002d0000000000000013000000000000000800000000",
            INIT_7D => X"0000001c000000000000001b000000000000001b000000000000001900000000",
            INIT_7E => X"0000002200000000000000140000000000000015000000000000001800000000",
            INIT_7F => X"0000000700000000000000040000000000000005000000000000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE13;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE14 : if BRAM_NAME = "sampleifmap_layersamples_instance14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009e00000000000000a600000000000000bb00000000000000be00000000",
            INIT_01 => X"000000d800000000000000d300000000000000d000000000000000c100000000",
            INIT_02 => X"000000da00000000000000de00000000000000dd00000000000000db00000000",
            INIT_03 => X"000000ed00000000000000eb00000000000000e800000000000000e500000000",
            INIT_04 => X"000000ef00000000000000ee00000000000000e900000000000000dc00000000",
            INIT_05 => X"000000f100000000000000f100000000000000ef00000000000000f100000000",
            INIT_06 => X"000000f300000000000000eb00000000000000e700000000000000f200000000",
            INIT_07 => X"000000f100000000000000ef00000000000000e700000000000000ed00000000",
            INIT_08 => X"000000a000000000000000b000000000000000c700000000000000c800000000",
            INIT_09 => X"000000da00000000000000da00000000000000d900000000000000c700000000",
            INIT_0A => X"000000db00000000000000e500000000000000e500000000000000df00000000",
            INIT_0B => X"000000f300000000000000ef00000000000000ee00000000000000e900000000",
            INIT_0C => X"000000f500000000000000ee00000000000000ea00000000000000e100000000",
            INIT_0D => X"000000f500000000000000ef00000000000000ed00000000000000f700000000",
            INIT_0E => X"000000f800000000000000ef00000000000000e900000000000000f500000000",
            INIT_0F => X"000000f700000000000000f600000000000000e800000000000000ec00000000",
            INIT_10 => X"000000a200000000000000b300000000000000c800000000000000c900000000",
            INIT_11 => X"000000d600000000000000df00000000000000dc00000000000000c900000000",
            INIT_12 => X"000000db00000000000000e200000000000000e900000000000000dd00000000",
            INIT_13 => X"000000f400000000000000ea00000000000000ea00000000000000e500000000",
            INIT_14 => X"000000f300000000000000ee00000000000000e900000000000000e200000000",
            INIT_15 => X"000000f100000000000000ea00000000000000d600000000000000eb00000000",
            INIT_16 => X"000000fa00000000000000f000000000000000e900000000000000f700000000",
            INIT_17 => X"000000f400000000000000f900000000000000e500000000000000ee00000000",
            INIT_18 => X"000000a400000000000000b300000000000000c700000000000000cb00000000",
            INIT_19 => X"000000d900000000000000e100000000000000d900000000000000c900000000",
            INIT_1A => X"000000d900000000000000e300000000000000eb00000000000000df00000000",
            INIT_1B => X"000000f400000000000000e200000000000000e800000000000000dd00000000",
            INIT_1C => X"000000eb00000000000000ed00000000000000e700000000000000e400000000",
            INIT_1D => X"000000f100000000000000e400000000000000af00000000000000b800000000",
            INIT_1E => X"000000fa00000000000000ee00000000000000e800000000000000f800000000",
            INIT_1F => X"000000f200000000000000f700000000000000e300000000000000ed00000000",
            INIT_20 => X"000000a100000000000000b500000000000000cc00000000000000cf00000000",
            INIT_21 => X"000000d500000000000000e100000000000000d600000000000000c900000000",
            INIT_22 => X"000000d700000000000000e200000000000000ed00000000000000d700000000",
            INIT_23 => X"000000ec00000000000000d400000000000000e500000000000000d900000000",
            INIT_24 => X"000000e100000000000000ec00000000000000e100000000000000e300000000",
            INIT_25 => X"000000ec00000000000000e000000000000000ae00000000000000aa00000000",
            INIT_26 => X"000000f600000000000000eb00000000000000e700000000000000f700000000",
            INIT_27 => X"000000ef00000000000000f500000000000000e700000000000000e700000000",
            INIT_28 => X"0000009a00000000000000b700000000000000cd00000000000000d000000000",
            INIT_29 => X"000000d700000000000000e200000000000000d400000000000000c900000000",
            INIT_2A => X"000000d700000000000000df00000000000000ee00000000000000da00000000",
            INIT_2B => X"000000cd00000000000000c700000000000000e500000000000000d700000000",
            INIT_2C => X"000000cc00000000000000ef00000000000000d000000000000000d100000000",
            INIT_2D => X"000000e900000000000000e300000000000000a7000000000000007c00000000",
            INIT_2E => X"000000ef00000000000000e100000000000000e500000000000000f600000000",
            INIT_2F => X"000000e800000000000000f100000000000000e600000000000000e200000000",
            INIT_30 => X"0000008b00000000000000b300000000000000c700000000000000cc00000000",
            INIT_31 => X"000000d500000000000000dd00000000000000cb00000000000000c200000000",
            INIT_32 => X"000000d400000000000000d800000000000000e900000000000000db00000000",
            INIT_33 => X"000000b000000000000000bc00000000000000e600000000000000d800000000",
            INIT_34 => X"000000c000000000000000d400000000000000c000000000000000be00000000",
            INIT_35 => X"000000be00000000000000b70000000000000097000000000000008100000000",
            INIT_36 => X"000000e500000000000000d600000000000000e000000000000000e000000000",
            INIT_37 => X"000000e000000000000000eb00000000000000de00000000000000db00000000",
            INIT_38 => X"0000008a00000000000000af00000000000000c600000000000000cd00000000",
            INIT_39 => X"000000cc00000000000000ce00000000000000cb00000000000000c000000000",
            INIT_3A => X"000000d200000000000000d000000000000000df00000000000000d400000000",
            INIT_3B => X"000000ce00000000000000c700000000000000d800000000000000d500000000",
            INIT_3C => X"0000005d0000000000000071000000000000009500000000000000b200000000",
            INIT_3D => X"0000004500000000000000500000000000000050000000000000005500000000",
            INIT_3E => X"000000de00000000000000ce00000000000000b7000000000000006c00000000",
            INIT_3F => X"000000d400000000000000dd00000000000000c500000000000000d000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000085000000000000009a00000000000000a800000000000000ad00000000",
            INIT_41 => X"000000b300000000000000a000000000000000ac00000000000000a500000000",
            INIT_42 => X"000000c300000000000000bd00000000000000c200000000000000be00000000",
            INIT_43 => X"000000c600000000000000c100000000000000bf00000000000000c700000000",
            INIT_44 => X"0000006c000000000000006b0000000000000079000000000000009800000000",
            INIT_45 => X"0000004f000000000000006e0000000000000068000000000000006800000000",
            INIT_46 => X"000000af000000000000009f000000000000007a000000000000005200000000",
            INIT_47 => X"000000af00000000000000be000000000000009500000000000000a300000000",
            INIT_48 => X"0000006900000000000000720000000000000074000000000000007300000000",
            INIT_49 => X"0000007f0000000000000070000000000000006e000000000000006d00000000",
            INIT_4A => X"00000093000000000000008c0000000000000088000000000000008700000000",
            INIT_4B => X"000000a1000000000000009e000000000000008f000000000000009700000000",
            INIT_4C => X"0000007800000000000000780000000000000077000000000000008600000000",
            INIT_4D => X"0000005c0000000000000066000000000000006c000000000000006c00000000",
            INIT_4E => X"0000009100000000000000970000000000000080000000000000008f00000000",
            INIT_4F => X"000000780000000000000082000000000000006a000000000000006e00000000",
            INIT_50 => X"0000005200000000000000560000000000000057000000000000004e00000000",
            INIT_51 => X"0000006400000000000000610000000000000069000000000000006300000000",
            INIT_52 => X"0000006f000000000000006a000000000000006d000000000000006500000000",
            INIT_53 => X"0000007f00000000000000840000000000000076000000000000007200000000",
            INIT_54 => X"0000006b000000000000006e000000000000006d000000000000006d00000000",
            INIT_55 => X"00000077000000000000006c0000000000000057000000000000006000000000",
            INIT_56 => X"000000bf0000000000000090000000000000006f000000000000008400000000",
            INIT_57 => X"000000680000000000000066000000000000006f000000000000007800000000",
            INIT_58 => X"00000062000000000000005f0000000000000055000000000000004a00000000",
            INIT_59 => X"000000510000000000000062000000000000007a000000000000008000000000",
            INIT_5A => X"0000007300000000000000710000000000000081000000000000006800000000",
            INIT_5B => X"0000007b0000000000000086000000000000008b000000000000008400000000",
            INIT_5C => X"0000007700000000000000740000000000000073000000000000007800000000",
            INIT_5D => X"000000bd000000000000009e0000000000000068000000000000007100000000",
            INIT_5E => X"000000c5000000000000006d000000000000009400000000000000b700000000",
            INIT_5F => X"0000006300000000000000630000000000000067000000000000009500000000",
            INIT_60 => X"0000005d0000000000000071000000000000006b000000000000005100000000",
            INIT_61 => X"00000066000000000000005d0000000000000073000000000000007500000000",
            INIT_62 => X"0000008300000000000000950000000000000098000000000000008900000000",
            INIT_63 => X"00000071000000000000007d0000000000000088000000000000008200000000",
            INIT_64 => X"0000007b0000000000000072000000000000006c000000000000006c00000000",
            INIT_65 => X"000000c200000000000000af000000000000007f000000000000007600000000",
            INIT_66 => X"000000a2000000000000007600000000000000bd00000000000000ce00000000",
            INIT_67 => X"000000650000000000000062000000000000005000000000000000a700000000",
            INIT_68 => X"0000005d000000000000006a000000000000006e000000000000006100000000",
            INIT_69 => X"0000006400000000000000590000000000000054000000000000006200000000",
            INIT_6A => X"00000086000000000000008a000000000000007b000000000000006e00000000",
            INIT_6B => X"0000007c00000000000000820000000000000083000000000000007e00000000",
            INIT_6C => X"00000087000000000000007e000000000000007f000000000000007b00000000",
            INIT_6D => X"000000b400000000000000b50000000000000099000000000000008600000000",
            INIT_6E => X"0000007a000000000000009700000000000000b700000000000000b800000000",
            INIT_6F => X"000000590000000000000048000000000000004d00000000000000a000000000",
            INIT_70 => X"0000006100000000000000660000000000000065000000000000006600000000",
            INIT_71 => X"0000006b00000000000000580000000000000058000000000000005f00000000",
            INIT_72 => X"0000009e0000000000000097000000000000008e000000000000008200000000",
            INIT_73 => X"0000009d00000000000000a100000000000000a400000000000000a300000000",
            INIT_74 => X"000000a900000000000000aa00000000000000ad00000000000000ab00000000",
            INIT_75 => X"000000ae00000000000000b100000000000000a900000000000000a200000000",
            INIT_76 => X"0000006200000000000000a400000000000000a800000000000000b000000000",
            INIT_77 => X"0000004b000000000000003f0000000000000046000000000000005700000000",
            INIT_78 => X"0000007c000000000000007f0000000000000076000000000000007b00000000",
            INIT_79 => X"000000a000000000000000980000000000000094000000000000007e00000000",
            INIT_7A => X"000000b400000000000000b300000000000000af00000000000000a700000000",
            INIT_7B => X"000000ae00000000000000b900000000000000b800000000000000b700000000",
            INIT_7C => X"000000a000000000000000af00000000000000b200000000000000ad00000000",
            INIT_7D => X"000000a1000000000000008e0000000000000085000000000000008000000000",
            INIT_7E => X"0000006c00000000000000a600000000000000a200000000000000a900000000",
            INIT_7F => X"000000520000000000000059000000000000005f000000000000004600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE14;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE15 : if BRAM_NAME = "sampleifmap_layersamples_instance15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000098000000000000008a000000000000007d000000000000008500000000",
            INIT_01 => X"000000a700000000000000a6000000000000009a000000000000009400000000",
            INIT_02 => X"000000b600000000000000b300000000000000ae00000000000000aa00000000",
            INIT_03 => X"000000ab00000000000000b500000000000000b900000000000000b900000000",
            INIT_04 => X"0000008b000000000000009a0000000000000098000000000000009800000000",
            INIT_05 => X"0000009b00000000000000900000000000000078000000000000006600000000",
            INIT_06 => X"0000008800000000000000a300000000000000a200000000000000a500000000",
            INIT_07 => X"0000006c000000000000009900000000000000bb000000000000009100000000",
            INIT_08 => X"00000083000000000000008d0000000000000085000000000000007c00000000",
            INIT_09 => X"000000aa00000000000000980000000000000072000000000000007400000000",
            INIT_0A => X"000000ad00000000000000b000000000000000af00000000000000af00000000",
            INIT_0B => X"00000097000000000000009a00000000000000a000000000000000a700000000",
            INIT_0C => X"000000a000000000000000a80000000000000096000000000000009000000000",
            INIT_0D => X"0000009e00000000000000a50000000000000098000000000000008c00000000",
            INIT_0E => X"00000097000000000000009c000000000000009b00000000000000a300000000",
            INIT_0F => X"000000930000000000000098000000000000009e000000000000009e00000000",
            INIT_10 => X"0000005d00000000000000600000000000000071000000000000008100000000",
            INIT_11 => X"000000a400000000000000940000000000000087000000000000006e00000000",
            INIT_12 => X"000000920000000000000096000000000000009f00000000000000a900000000",
            INIT_13 => X"000000a5000000000000009f0000000000000099000000000000009400000000",
            INIT_14 => X"000000ac00000000000000a800000000000000a000000000000000aa00000000",
            INIT_15 => X"000000a400000000000000a800000000000000a400000000000000a100000000",
            INIT_16 => X"00000092000000000000009e000000000000009e00000000000000a000000000",
            INIT_17 => X"00000096000000000000007d0000000000000079000000000000008400000000",
            INIT_18 => X"0000008700000000000000600000000000000055000000000000007000000000",
            INIT_19 => X"00000093000000000000009c00000000000000a5000000000000009b00000000",
            INIT_1A => X"000000a00000000000000097000000000000008d000000000000008e00000000",
            INIT_1B => X"000000ab00000000000000ae00000000000000ad00000000000000a700000000",
            INIT_1C => X"000000a800000000000000a2000000000000009b00000000000000a700000000",
            INIT_1D => X"000000a600000000000000a300000000000000a100000000000000a300000000",
            INIT_1E => X"0000006f00000000000000820000000000000097000000000000009e00000000",
            INIT_1F => X"0000008a000000000000005c0000000000000052000000000000006200000000",
            INIT_20 => X"0000008f00000000000000870000000000000084000000000000008500000000",
            INIT_21 => X"0000008e0000000000000096000000000000008f000000000000008f00000000",
            INIT_22 => X"000000ab00000000000000a900000000000000a1000000000000008a00000000",
            INIT_23 => X"00000086000000000000009700000000000000a500000000000000a900000000",
            INIT_24 => X"000000a40000000000000094000000000000006b000000000000007400000000",
            INIT_25 => X"00000098000000000000009f00000000000000a300000000000000a300000000",
            INIT_26 => X"0000005b0000000000000066000000000000006c000000000000008000000000",
            INIT_27 => X"000000480000000000000050000000000000004e000000000000004b00000000",
            INIT_28 => X"0000008f0000000000000090000000000000008c000000000000008400000000",
            INIT_29 => X"0000009600000000000000970000000000000093000000000000009000000000",
            INIT_2A => X"0000009a00000000000000940000000000000092000000000000008b00000000",
            INIT_2B => X"0000004e000000000000006e000000000000009c000000000000009f00000000",
            INIT_2C => X"000000a30000000000000084000000000000004a000000000000004b00000000",
            INIT_2D => X"0000006d000000000000007e000000000000008f000000000000009900000000",
            INIT_2E => X"0000004c000000000000005a0000000000000064000000000000006700000000",
            INIT_2F => X"0000002100000000000000390000000000000052000000000000004b00000000",
            INIT_30 => X"0000009200000000000000940000000000000089000000000000005e00000000",
            INIT_31 => X"0000007300000000000000810000000000000091000000000000009200000000",
            INIT_32 => X"0000008700000000000000630000000000000066000000000000006a00000000",
            INIT_33 => X"0000005d0000000000000072000000000000009a000000000000009d00000000",
            INIT_34 => X"0000007c000000000000007d0000000000000068000000000000006500000000",
            INIT_35 => X"000000650000000000000066000000000000006a000000000000007100000000",
            INIT_36 => X"0000003f0000000000000045000000000000004f000000000000005800000000",
            INIT_37 => X"0000001f00000000000000250000000000000035000000000000004300000000",
            INIT_38 => X"000000860000000000000086000000000000007d000000000000005600000000",
            INIT_39 => X"0000004d000000000000005c0000000000000085000000000000008900000000",
            INIT_3A => X"00000083000000000000005c0000000000000059000000000000005200000000",
            INIT_3B => X"0000007300000000000000840000000000000096000000000000009900000000",
            INIT_3C => X"0000006100000000000000600000000000000061000000000000006a00000000",
            INIT_3D => X"0000004f000000000000005f0000000000000065000000000000006300000000",
            INIT_3E => X"00000039000000000000003c0000000000000040000000000000003c00000000",
            INIT_3F => X"0000001f00000000000000220000000000000026000000000000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008300000000000000810000000000000074000000000000005a00000000",
            INIT_41 => X"00000061000000000000006a000000000000008a000000000000008900000000",
            INIT_42 => X"0000007e000000000000007c0000000000000074000000000000006c00000000",
            INIT_43 => X"000000530000000000000054000000000000005f000000000000007100000000",
            INIT_44 => X"000000640000000000000062000000000000005c000000000000005900000000",
            INIT_45 => X"000000450000000000000043000000000000004a000000000000005c00000000",
            INIT_46 => X"0000002e00000000000000330000000000000042000000000000004a00000000",
            INIT_47 => X"0000002000000000000000230000000000000026000000000000002b00000000",
            INIT_48 => X"0000007f00000000000000820000000000000070000000000000005c00000000",
            INIT_49 => X"00000066000000000000006e0000000000000078000000000000007c00000000",
            INIT_4A => X"0000004c0000000000000050000000000000005a000000000000006100000000",
            INIT_4B => X"0000005b00000000000000540000000000000050000000000000004b00000000",
            INIT_4C => X"0000004900000000000000510000000000000059000000000000005f00000000",
            INIT_4D => X"0000003d00000000000000430000000000000041000000000000004100000000",
            INIT_4E => X"00000028000000000000002a000000000000003a000000000000004500000000",
            INIT_4F => X"0000002500000000000000230000000000000028000000000000002a00000000",
            INIT_50 => X"0000004e0000000000000056000000000000004f000000000000004c00000000",
            INIT_51 => X"0000003f00000000000000400000000000000045000000000000004a00000000",
            INIT_52 => X"0000004d000000000000004a0000000000000046000000000000004100000000",
            INIT_53 => X"0000005000000000000000510000000000000052000000000000005100000000",
            INIT_54 => X"000000440000000000000037000000000000003b000000000000004900000000",
            INIT_55 => X"000000320000000000000036000000000000003f000000000000004300000000",
            INIT_56 => X"000000280000000000000028000000000000002d000000000000003600000000",
            INIT_57 => X"0000002500000000000000270000000000000028000000000000002900000000",
            INIT_58 => X"0000002a0000000000000028000000000000002b000000000000002d00000000",
            INIT_59 => X"0000003a00000000000000350000000000000034000000000000003100000000",
            INIT_5A => X"0000004600000000000000480000000000000047000000000000004400000000",
            INIT_5B => X"0000003b000000000000003a000000000000003b000000000000004100000000",
            INIT_5C => X"000000490000000000000055000000000000003f000000000000003800000000",
            INIT_5D => X"0000002f000000000000002f0000000000000033000000000000003900000000",
            INIT_5E => X"0000002800000000000000270000000000000028000000000000002c00000000",
            INIT_5F => X"0000001d000000000000002a000000000000002a000000000000002900000000",
            INIT_60 => X"0000002600000000000000240000000000000028000000000000002b00000000",
            INIT_61 => X"0000003200000000000000310000000000000030000000000000002c00000000",
            INIT_62 => X"0000003100000000000000310000000000000034000000000000003500000000",
            INIT_63 => X"0000003d000000000000003e000000000000003b000000000000003500000000",
            INIT_64 => X"00000042000000000000005e0000000000000045000000000000003700000000",
            INIT_65 => X"00000028000000000000002f000000000000002e000000000000002c00000000",
            INIT_66 => X"0000002a00000000000000280000000000000027000000000000002700000000",
            INIT_67 => X"000000120000000000000020000000000000002e000000000000002900000000",
            INIT_68 => X"0000002400000000000000230000000000000027000000000000002800000000",
            INIT_69 => X"0000002b00000000000000290000000000000029000000000000002700000000",
            INIT_6A => X"0000003a00000000000000380000000000000033000000000000002e00000000",
            INIT_6B => X"00000037000000000000003c000000000000003d000000000000003d00000000",
            INIT_6C => X"000000360000000000000055000000000000003c000000000000002e00000000",
            INIT_6D => X"000000240000000000000025000000000000002e000000000000002800000000",
            INIT_6E => X"0000002a00000000000000280000000000000026000000000000002600000000",
            INIT_6F => X"00000007000000000000000d0000000000000028000000000000002b00000000",
            INIT_70 => X"0000002800000000000000240000000000000026000000000000002200000000",
            INIT_71 => X"000000330000000000000031000000000000002f000000000000002c00000000",
            INIT_72 => X"00000039000000000000003b0000000000000039000000000000003600000000",
            INIT_73 => X"0000002b00000000000000330000000000000037000000000000003900000000",
            INIT_74 => X"00000032000000000000004e0000000000000030000000000000001f00000000",
            INIT_75 => X"0000002300000000000000230000000000000025000000000000002900000000",
            INIT_76 => X"0000002900000000000000240000000000000025000000000000002500000000",
            INIT_77 => X"0000000700000000000000060000000000000014000000000000002d00000000",
            INIT_78 => X"0000002f000000000000002d000000000000002b000000000000002900000000",
            INIT_79 => X"0000003100000000000000300000000000000030000000000000003000000000",
            INIT_7A => X"0000002d00000000000000310000000000000033000000000000003200000000",
            INIT_7B => X"00000011000000000000001a0000000000000022000000000000002800000000",
            INIT_7C => X"0000002c000000000000003f000000000000001b000000000000000800000000",
            INIT_7D => X"0000002300000000000000220000000000000022000000000000002100000000",
            INIT_7E => X"0000002c00000000000000220000000000000022000000000000002300000000",
            INIT_7F => X"0000000800000000000000050000000000000006000000000000001f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE15;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE16 : if BRAM_NAME = "sampleifmap_layersamples_instance16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ba00000000000000c200000000000000da00000000000000de00000000",
            INIT_01 => X"000000f100000000000000ee00000000000000ec00000000000000de00000000",
            INIT_02 => X"000000eb00000000000000f400000000000000f500000000000000f300000000",
            INIT_03 => X"000000f500000000000000f200000000000000f100000000000000f000000000",
            INIT_04 => X"000000f800000000000000f500000000000000f000000000000000e300000000",
            INIT_05 => X"000000f300000000000000f300000000000000f300000000000000f900000000",
            INIT_06 => X"000000f700000000000000ef00000000000000eb00000000000000f500000000",
            INIT_07 => X"000000f600000000000000f300000000000000ea00000000000000f100000000",
            INIT_08 => X"000000b800000000000000c900000000000000e200000000000000e500000000",
            INIT_09 => X"000000ee00000000000000f000000000000000f000000000000000df00000000",
            INIT_0A => X"000000e800000000000000f500000000000000f700000000000000f300000000",
            INIT_0B => X"000000f800000000000000f500000000000000f500000000000000f300000000",
            INIT_0C => X"000000fb00000000000000f300000000000000ef00000000000000e600000000",
            INIT_0D => X"000000f400000000000000ee00000000000000ee00000000000000fb00000000",
            INIT_0E => X"000000fc00000000000000f300000000000000ec00000000000000f800000000",
            INIT_0F => X"000000fb00000000000000fa00000000000000ec00000000000000f000000000",
            INIT_10 => X"000000b500000000000000c700000000000000de00000000000000e100000000",
            INIT_11 => X"000000e400000000000000ef00000000000000ee00000000000000db00000000",
            INIT_12 => X"000000e400000000000000ec00000000000000f400000000000000eb00000000",
            INIT_13 => X"000000f700000000000000ee00000000000000ef00000000000000eb00000000",
            INIT_14 => X"000000f600000000000000f100000000000000ec00000000000000e500000000",
            INIT_15 => X"000000ef00000000000000e800000000000000d700000000000000ec00000000",
            INIT_16 => X"000000fc00000000000000f200000000000000eb00000000000000f800000000",
            INIT_17 => X"000000f700000000000000fb00000000000000e800000000000000f100000000",
            INIT_18 => X"000000b300000000000000c200000000000000d800000000000000de00000000",
            INIT_19 => X"000000e100000000000000eb00000000000000e400000000000000d600000000",
            INIT_1A => X"000000dd00000000000000e600000000000000ef00000000000000e500000000",
            INIT_1B => X"000000f700000000000000e600000000000000ec00000000000000e100000000",
            INIT_1C => X"000000ee00000000000000f000000000000000ea00000000000000e600000000",
            INIT_1D => X"000000f100000000000000e500000000000000b000000000000000ba00000000",
            INIT_1E => X"000000fb00000000000000ef00000000000000e900000000000000f800000000",
            INIT_1F => X"000000f300000000000000f800000000000000e400000000000000ee00000000",
            INIT_20 => X"000000ac00000000000000c100000000000000d900000000000000df00000000",
            INIT_21 => X"000000d900000000000000e700000000000000dd00000000000000d200000000",
            INIT_22 => X"000000d700000000000000e100000000000000eb00000000000000da00000000",
            INIT_23 => X"000000ee00000000000000d600000000000000e800000000000000db00000000",
            INIT_24 => X"000000e400000000000000ee00000000000000e300000000000000e500000000",
            INIT_25 => X"000000ef00000000000000e500000000000000b200000000000000b000000000",
            INIT_26 => X"000000f500000000000000ea00000000000000e700000000000000f700000000",
            INIT_27 => X"000000f000000000000000f600000000000000e800000000000000e700000000",
            INIT_28 => X"000000a400000000000000bf00000000000000d500000000000000dc00000000",
            INIT_29 => X"000000d500000000000000e100000000000000d500000000000000ce00000000",
            INIT_2A => X"000000d600000000000000da00000000000000e600000000000000d600000000",
            INIT_2B => X"000000ce00000000000000c800000000000000e300000000000000d600000000",
            INIT_2C => X"000000cf00000000000000ed00000000000000ce00000000000000d000000000",
            INIT_2D => X"000000e900000000000000e600000000000000ad000000000000008200000000",
            INIT_2E => X"000000e800000000000000db00000000000000e100000000000000f400000000",
            INIT_2F => X"000000e600000000000000f200000000000000e700000000000000dd00000000",
            INIT_30 => X"0000009600000000000000b900000000000000ca00000000000000d400000000",
            INIT_31 => X"000000d000000000000000d900000000000000c900000000000000c400000000",
            INIT_32 => X"000000d300000000000000d000000000000000db00000000000000d300000000",
            INIT_33 => X"000000af00000000000000b900000000000000dd00000000000000d400000000",
            INIT_34 => X"000000c500000000000000d200000000000000bd00000000000000bb00000000",
            INIT_35 => X"000000bb00000000000000b8000000000000009d000000000000008900000000",
            INIT_36 => X"000000da00000000000000ce00000000000000dc00000000000000dd00000000",
            INIT_37 => X"000000d800000000000000e700000000000000db00000000000000d100000000",
            INIT_38 => X"0000009300000000000000b300000000000000c900000000000000d300000000",
            INIT_39 => X"000000cb00000000000000ce00000000000000cc00000000000000c500000000",
            INIT_3A => X"000000cd00000000000000c600000000000000d200000000000000d000000000",
            INIT_3B => X"000000cb00000000000000c000000000000000ce00000000000000ce00000000",
            INIT_3C => X"0000006a000000000000007a000000000000009b00000000000000b300000000",
            INIT_3D => X"000000490000000000000058000000000000005e000000000000006400000000",
            INIT_3E => X"000000d700000000000000ca00000000000000b7000000000000006f00000000",
            INIT_3F => X"000000c100000000000000ce00000000000000b900000000000000c600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008c00000000000000a000000000000000ad00000000000000b300000000",
            INIT_41 => X"000000b300000000000000a100000000000000af00000000000000aa00000000",
            INIT_42 => X"000000bd00000000000000b400000000000000b800000000000000bb00000000",
            INIT_43 => X"000000c400000000000000ba00000000000000b900000000000000c300000000",
            INIT_44 => X"0000008000000000000000800000000000000089000000000000009f00000000",
            INIT_45 => X"0000005a0000000000000080000000000000007e000000000000007e00000000",
            INIT_46 => X"000000ac000000000000009e000000000000007c000000000000005800000000",
            INIT_47 => X"0000009f00000000000000b00000000000000089000000000000009c00000000",
            INIT_48 => X"00000070000000000000007b000000000000007e000000000000007b00000000",
            INIT_49 => X"0000008000000000000000720000000000000072000000000000007200000000",
            INIT_4A => X"0000009000000000000000890000000000000086000000000000008600000000",
            INIT_4B => X"000000a700000000000000a00000000000000092000000000000009800000000",
            INIT_4C => X"0000008c0000000000000090000000000000008b000000000000009300000000",
            INIT_4D => X"0000006800000000000000780000000000000083000000000000008200000000",
            INIT_4E => X"0000008d00000000000000960000000000000083000000000000009500000000",
            INIT_4F => X"0000007500000000000000800000000000000069000000000000006a00000000",
            INIT_50 => X"0000005800000000000000620000000000000066000000000000005900000000",
            INIT_51 => X"0000006a00000000000000680000000000000073000000000000006b00000000",
            INIT_52 => X"0000007300000000000000710000000000000076000000000000006b00000000",
            INIT_53 => X"0000009200000000000000970000000000000086000000000000007b00000000",
            INIT_54 => X"00000078000000000000007f000000000000007f000000000000008000000000",
            INIT_55 => X"00000080000000000000007a0000000000000068000000000000006f00000000",
            INIT_56 => X"000000b6000000000000008b000000000000006e000000000000008600000000",
            INIT_57 => X"00000070000000000000006d0000000000000075000000000000007200000000",
            INIT_58 => X"0000006a000000000000006e0000000000000068000000000000005800000000",
            INIT_59 => X"0000005e00000000000000710000000000000089000000000000008e00000000",
            INIT_5A => X"0000007d000000000000007f0000000000000092000000000000007400000000",
            INIT_5B => X"0000009700000000000000a500000000000000a5000000000000009400000000",
            INIT_5C => X"0000007f000000000000007f0000000000000082000000000000008e00000000",
            INIT_5D => X"000000bf00000000000000a50000000000000072000000000000007b00000000",
            INIT_5E => X"000000b80000000000000064000000000000008e00000000000000b400000000",
            INIT_5F => X"0000006c000000000000006c000000000000006d000000000000008c00000000",
            INIT_60 => X"0000006800000000000000840000000000000082000000000000006400000000",
            INIT_61 => X"00000076000000000000006d0000000000000082000000000000008100000000",
            INIT_62 => X"0000009700000000000000a800000000000000ab000000000000009a00000000",
            INIT_63 => X"0000008b000000000000009a00000000000000a5000000000000009b00000000",
            INIT_64 => X"0000008c0000000000000081000000000000007d000000000000008200000000",
            INIT_65 => X"000000c100000000000000b30000000000000089000000000000008600000000",
            INIT_66 => X"00000098000000000000007000000000000000b900000000000000cb00000000",
            INIT_67 => X"0000006d0000000000000069000000000000005400000000000000a000000000",
            INIT_68 => X"0000006a000000000000007e0000000000000086000000000000007800000000",
            INIT_69 => X"00000079000000000000006c0000000000000065000000000000007100000000",
            INIT_6A => X"0000009f00000000000000a10000000000000091000000000000008300000000",
            INIT_6B => X"00000095000000000000009e00000000000000a1000000000000009900000000",
            INIT_6C => X"0000009b00000000000000910000000000000093000000000000009200000000",
            INIT_6D => X"000000b100000000000000b600000000000000a1000000000000009600000000",
            INIT_6E => X"00000076000000000000009400000000000000b500000000000000b500000000",
            INIT_6F => X"00000060000000000000004e0000000000000050000000000000009d00000000",
            INIT_70 => X"00000072000000000000007d0000000000000080000000000000007f00000000",
            INIT_71 => X"0000008600000000000000730000000000000071000000000000007400000000",
            INIT_72 => X"000000b800000000000000b000000000000000a8000000000000009f00000000",
            INIT_73 => X"000000b900000000000000be00000000000000bf00000000000000be00000000",
            INIT_74 => X"000000b800000000000000be00000000000000c400000000000000c500000000",
            INIT_75 => X"000000a800000000000000af00000000000000ad00000000000000ac00000000",
            INIT_76 => X"0000006300000000000000a300000000000000a500000000000000ab00000000",
            INIT_77 => X"0000005100000000000000430000000000000047000000000000005700000000",
            INIT_78 => X"00000091000000000000009a0000000000000095000000000000009700000000",
            INIT_79 => X"000000c100000000000000b800000000000000b3000000000000009900000000",
            INIT_7A => X"000000d000000000000000cf00000000000000cd00000000000000c900000000",
            INIT_7B => X"000000c800000000000000d400000000000000d200000000000000d100000000",
            INIT_7C => X"000000ab00000000000000c300000000000000c900000000000000c600000000",
            INIT_7D => X"0000009b000000000000008b0000000000000087000000000000008600000000",
            INIT_7E => X"0000007100000000000000a800000000000000a100000000000000a500000000",
            INIT_7F => X"00000056000000000000005a000000000000005c000000000000004900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE16;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE17 : if BRAM_NAME = "sampleifmap_layersamples_instance17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b000000000000000a7000000000000009f00000000000000a500000000",
            INIT_01 => X"000000c900000000000000c600000000000000b900000000000000af00000000",
            INIT_02 => X"000000d200000000000000d200000000000000d000000000000000cd00000000",
            INIT_03 => X"000000be00000000000000c900000000000000d000000000000000d200000000",
            INIT_04 => X"0000009400000000000000a900000000000000aa00000000000000aa00000000",
            INIT_05 => X"00000099000000000000008e000000000000007a000000000000006c00000000",
            INIT_06 => X"0000008e00000000000000a700000000000000a500000000000000a700000000",
            INIT_07 => X"0000006f000000000000009800000000000000b5000000000000009300000000",
            INIT_08 => X"0000009d00000000000000ae00000000000000aa000000000000009d00000000",
            INIT_09 => X"000000ca00000000000000b6000000000000008f000000000000008d00000000",
            INIT_0A => X"000000ca00000000000000d100000000000000d300000000000000d000000000",
            INIT_0B => X"000000a200000000000000a700000000000000b500000000000000bf00000000",
            INIT_0C => X"000000a900000000000000b200000000000000a0000000000000009b00000000",
            INIT_0D => X"000000a000000000000000a7000000000000009d000000000000009300000000",
            INIT_0E => X"0000009c00000000000000a100000000000000a200000000000000a900000000",
            INIT_0F => X"0000009400000000000000960000000000000096000000000000009e00000000",
            INIT_10 => X"000000790000000000000080000000000000009400000000000000a200000000",
            INIT_11 => X"000000c200000000000000b100000000000000a4000000000000008a00000000",
            INIT_12 => X"000000ab00000000000000b200000000000000bc00000000000000c700000000",
            INIT_13 => X"000000b000000000000000ac00000000000000ac00000000000000aa00000000",
            INIT_14 => X"000000b500000000000000b000000000000000a800000000000000b400000000",
            INIT_15 => X"000000ac00000000000000af00000000000000ad00000000000000aa00000000",
            INIT_16 => X"0000009600000000000000a300000000000000a500000000000000a800000000",
            INIT_17 => X"00000099000000000000007d0000000000000076000000000000008500000000",
            INIT_18 => X"000000a6000000000000007f0000000000000075000000000000008f00000000",
            INIT_19 => X"000000b000000000000000ba00000000000000c500000000000000bc00000000",
            INIT_1A => X"000000b200000000000000ab00000000000000a300000000000000a900000000",
            INIT_1B => X"000000ba00000000000000bf00000000000000be00000000000000b900000000",
            INIT_1C => X"000000b100000000000000ac00000000000000a500000000000000b400000000",
            INIT_1D => X"000000b200000000000000af00000000000000ac00000000000000ad00000000",
            INIT_1E => X"000000740000000000000088000000000000009c00000000000000a400000000",
            INIT_1F => X"0000009000000000000000620000000000000057000000000000006700000000",
            INIT_20 => X"000000b000000000000000a800000000000000a500000000000000a600000000",
            INIT_21 => X"000000aa00000000000000b300000000000000ae00000000000000b000000000",
            INIT_22 => X"000000bd00000000000000be00000000000000b800000000000000a400000000",
            INIT_23 => X"0000009600000000000000a800000000000000b500000000000000b900000000",
            INIT_24 => X"000000ad000000000000009d0000000000000076000000000000008100000000",
            INIT_25 => X"000000a200000000000000ab00000000000000ad00000000000000ad00000000",
            INIT_26 => X"0000005f000000000000006a0000000000000070000000000000008500000000",
            INIT_27 => X"0000004e00000000000000560000000000000054000000000000005000000000",
            INIT_28 => X"000000af00000000000000b100000000000000ac00000000000000a500000000",
            INIT_29 => X"000000b000000000000000b300000000000000b000000000000000ae00000000",
            INIT_2A => X"000000ad00000000000000ab00000000000000ab00000000000000a400000000",
            INIT_2B => X"0000005e000000000000007e00000000000000ab00000000000000af00000000",
            INIT_2C => X"000000ac000000000000008e0000000000000055000000000000005800000000",
            INIT_2D => X"000000750000000000000088000000000000009800000000000000a200000000",
            INIT_2E => X"00000050000000000000005e0000000000000068000000000000006c00000000",
            INIT_2F => X"00000027000000000000003f0000000000000058000000000000004f00000000",
            INIT_30 => X"000000af00000000000000b200000000000000a6000000000000007c00000000",
            INIT_31 => X"0000008b000000000000009a00000000000000ad00000000000000af00000000",
            INIT_32 => X"0000009a000000000000007a000000000000007e000000000000008200000000",
            INIT_33 => X"0000006c000000000000008300000000000000a900000000000000ae00000000",
            INIT_34 => X"0000008500000000000000860000000000000072000000000000007200000000",
            INIT_35 => X"0000006c000000000000006d0000000000000071000000000000007900000000",
            INIT_36 => X"00000045000000000000004b0000000000000056000000000000005f00000000",
            INIT_37 => X"00000026000000000000002b000000000000003b000000000000004900000000",
            INIT_38 => X"0000009f00000000000000a00000000000000096000000000000006f00000000",
            INIT_39 => X"000000640000000000000074000000000000009e00000000000000a300000000",
            INIT_3A => X"0000009700000000000000730000000000000070000000000000006800000000",
            INIT_3B => X"00000083000000000000009500000000000000a800000000000000ac00000000",
            INIT_3C => X"0000006a000000000000006a000000000000006b000000000000007700000000",
            INIT_3D => X"000000540000000000000064000000000000006c000000000000006a00000000",
            INIT_3E => X"0000004100000000000000440000000000000049000000000000004500000000",
            INIT_3F => X"000000250000000000000028000000000000002c000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009a0000000000000097000000000000008a000000000000007100000000",
            INIT_41 => X"00000077000000000000008000000000000000a200000000000000a100000000",
            INIT_42 => X"0000009200000000000000900000000000000088000000000000008100000000",
            INIT_43 => X"0000006200000000000000650000000000000072000000000000008400000000",
            INIT_44 => X"0000006c000000000000006d0000000000000067000000000000006500000000",
            INIT_45 => X"0000004b00000000000000480000000000000050000000000000006300000000",
            INIT_46 => X"0000003a000000000000003d000000000000004d000000000000005500000000",
            INIT_47 => X"000000270000000000000029000000000000002d000000000000003400000000",
            INIT_48 => X"00000097000000000000009a0000000000000088000000000000007400000000",
            INIT_49 => X"0000007c0000000000000084000000000000008f000000000000009400000000",
            INIT_4A => X"00000057000000000000005b0000000000000067000000000000007600000000",
            INIT_4B => X"000000650000000000000063000000000000005b000000000000005600000000",
            INIT_4C => X"00000052000000000000005e0000000000000063000000000000006500000000",
            INIT_4D => X"00000045000000000000004a0000000000000048000000000000004800000000",
            INIT_4E => X"0000003200000000000000340000000000000044000000000000004e00000000",
            INIT_4F => X"00000030000000000000002f0000000000000030000000000000003300000000",
            INIT_50 => X"00000063000000000000006a0000000000000064000000000000006000000000",
            INIT_51 => X"0000005100000000000000520000000000000056000000000000005c00000000",
            INIT_52 => X"000000540000000000000051000000000000004f000000000000005200000000",
            INIT_53 => X"00000058000000000000005e000000000000005b000000000000005700000000",
            INIT_54 => X"0000004c00000000000000440000000000000044000000000000004d00000000",
            INIT_55 => X"0000003b00000000000000400000000000000048000000000000004a00000000",
            INIT_56 => X"0000003200000000000000310000000000000036000000000000003f00000000",
            INIT_57 => X"0000003000000000000000340000000000000030000000000000003100000000",
            INIT_58 => X"0000003700000000000000360000000000000039000000000000003b00000000",
            INIT_59 => X"00000044000000000000003e000000000000003d000000000000003c00000000",
            INIT_5A => X"0000004d000000000000004f000000000000004f000000000000004e00000000",
            INIT_5B => X"0000004200000000000000450000000000000044000000000000004800000000",
            INIT_5C => X"0000005200000000000000610000000000000047000000000000003d00000000",
            INIT_5D => X"000000390000000000000038000000000000003c000000000000004100000000",
            INIT_5E => X"0000003100000000000000300000000000000031000000000000003500000000",
            INIT_5F => X"0000002300000000000000320000000000000032000000000000003200000000",
            INIT_60 => X"0000002d000000000000002c0000000000000030000000000000003200000000",
            INIT_61 => X"0000003700000000000000350000000000000035000000000000003100000000",
            INIT_62 => X"000000380000000000000038000000000000003b000000000000003a00000000",
            INIT_63 => X"0000004400000000000000470000000000000042000000000000003c00000000",
            INIT_64 => X"0000004b0000000000000068000000000000004b000000000000003b00000000",
            INIT_65 => X"00000033000000000000003a0000000000000038000000000000003500000000",
            INIT_66 => X"0000003300000000000000310000000000000030000000000000003100000000",
            INIT_67 => X"0000001400000000000000250000000000000035000000000000003200000000",
            INIT_68 => X"000000290000000000000028000000000000002c000000000000002d00000000",
            INIT_69 => X"00000030000000000000002e000000000000002e000000000000002c00000000",
            INIT_6A => X"00000041000000000000003f0000000000000039000000000000003300000000",
            INIT_6B => X"0000003d00000000000000440000000000000044000000000000004400000000",
            INIT_6C => X"0000003f000000000000005d0000000000000042000000000000003200000000",
            INIT_6D => X"0000002f00000000000000300000000000000038000000000000003100000000",
            INIT_6E => X"000000330000000000000031000000000000002f000000000000002f00000000",
            INIT_6F => X"00000005000000000000000e000000000000002e000000000000003400000000",
            INIT_70 => X"0000002d0000000000000029000000000000002b000000000000002700000000",
            INIT_71 => X"0000003b00000000000000380000000000000036000000000000003200000000",
            INIT_72 => X"0000004000000000000000420000000000000040000000000000003e00000000",
            INIT_73 => X"00000031000000000000003a000000000000003d000000000000004000000000",
            INIT_74 => X"0000003b00000000000000550000000000000035000000000000002400000000",
            INIT_75 => X"0000002f000000000000002f0000000000000030000000000000003200000000",
            INIT_76 => X"00000032000000000000002d000000000000002e000000000000002e00000000",
            INIT_77 => X"0000000300000000000000030000000000000018000000000000003600000000",
            INIT_78 => X"0000003600000000000000340000000000000032000000000000002f00000000",
            INIT_79 => X"0000003a00000000000000380000000000000038000000000000003800000000",
            INIT_7A => X"0000003200000000000000350000000000000037000000000000003a00000000",
            INIT_7B => X"00000014000000000000001e0000000000000027000000000000002d00000000",
            INIT_7C => X"0000003600000000000000480000000000000021000000000000000b00000000",
            INIT_7D => X"0000002e000000000000002d000000000000002d000000000000002c00000000",
            INIT_7E => X"00000034000000000000002b000000000000002c000000000000002c00000000",
            INIT_7F => X"0000000700000000000000030000000000000008000000000000002500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE17;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE18 : if BRAM_NAME = "sampleifmap_layersamples_instance18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000be00000000000000b000000000000000a7000000000000009b00000000",
            INIT_01 => X"000000a600000000000000a800000000000000a600000000000000b100000000",
            INIT_02 => X"000000bb00000000000000bb00000000000000b300000000000000aa00000000",
            INIT_03 => X"000000b800000000000000b800000000000000bb00000000000000bb00000000",
            INIT_04 => X"000000ba00000000000000b800000000000000b400000000000000b600000000",
            INIT_05 => X"000000bd00000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_06 => X"000000c300000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_07 => X"000000c000000000000000ca00000000000000c900000000000000c900000000",
            INIT_08 => X"000000bb00000000000000ab00000000000000a3000000000000009900000000",
            INIT_09 => X"0000009f000000000000009a000000000000009b00000000000000b300000000",
            INIT_0A => X"000000af00000000000000ab00000000000000a5000000000000009f00000000",
            INIT_0B => X"000000a500000000000000a200000000000000ab00000000000000a900000000",
            INIT_0C => X"000000a500000000000000a600000000000000a400000000000000aa00000000",
            INIT_0D => X"000000a800000000000000a900000000000000ad00000000000000a700000000",
            INIT_0E => X"000000ca00000000000000be00000000000000ad00000000000000a900000000",
            INIT_0F => X"000000bd00000000000000cb00000000000000ca00000000000000cc00000000",
            INIT_10 => X"000000b800000000000000a800000000000000a0000000000000009b00000000",
            INIT_11 => X"000000bc00000000000000b000000000000000ae00000000000000bb00000000",
            INIT_12 => X"000000be00000000000000b100000000000000b300000000000000b600000000",
            INIT_13 => X"000000b900000000000000bc00000000000000c200000000000000c000000000",
            INIT_14 => X"000000c200000000000000c100000000000000c200000000000000c100000000",
            INIT_15 => X"000000bf00000000000000c100000000000000c500000000000000c300000000",
            INIT_16 => X"000000cf00000000000000ce00000000000000c500000000000000bf00000000",
            INIT_17 => X"000000bd00000000000000cc00000000000000ce00000000000000d000000000",
            INIT_18 => X"000000b100000000000000a6000000000000009d000000000000009700000000",
            INIT_19 => X"000000c500000000000000c700000000000000b900000000000000b400000000",
            INIT_1A => X"000000c600000000000000cd00000000000000cc00000000000000b600000000",
            INIT_1B => X"000000cb00000000000000c400000000000000c500000000000000d200000000",
            INIT_1C => X"000000cb00000000000000d200000000000000cf00000000000000cd00000000",
            INIT_1D => X"000000cc00000000000000c500000000000000d200000000000000cf00000000",
            INIT_1E => X"000000c900000000000000cc00000000000000c600000000000000d000000000",
            INIT_1F => X"000000c000000000000000ce00000000000000cf00000000000000d100000000",
            INIT_20 => X"000000ae00000000000000a8000000000000009e000000000000009700000000",
            INIT_21 => X"000000c400000000000000bf00000000000000b500000000000000b100000000",
            INIT_22 => X"000000b900000000000000bd00000000000000c200000000000000b700000000",
            INIT_23 => X"000000ca00000000000000b900000000000000b900000000000000c400000000",
            INIT_24 => X"000000c000000000000000c800000000000000c700000000000000c700000000",
            INIT_25 => X"000000bc00000000000000be00000000000000c700000000000000c300000000",
            INIT_26 => X"000000c400000000000000c900000000000000c700000000000000c900000000",
            INIT_27 => X"000000c400000000000000cf00000000000000cc00000000000000ce00000000",
            INIT_28 => X"000000ae00000000000000a7000000000000009c000000000000009400000000",
            INIT_29 => X"000000c300000000000000c400000000000000ae00000000000000ab00000000",
            INIT_2A => X"000000b800000000000000bd00000000000000be00000000000000c000000000",
            INIT_2B => X"000000bf00000000000000bd00000000000000bd00000000000000bb00000000",
            INIT_2C => X"000000c600000000000000bb00000000000000c300000000000000be00000000",
            INIT_2D => X"000000c100000000000000c000000000000000bc00000000000000c000000000",
            INIT_2E => X"000000d100000000000000cb00000000000000ce00000000000000cd00000000",
            INIT_2F => X"000000c400000000000000d100000000000000d000000000000000d400000000",
            INIT_30 => X"000000ae00000000000000a50000000000000099000000000000009400000000",
            INIT_31 => X"000000c300000000000000cb00000000000000b000000000000000a800000000",
            INIT_32 => X"000000be00000000000000bb00000000000000bc00000000000000bc00000000",
            INIT_33 => X"000000c300000000000000c500000000000000c200000000000000b600000000",
            INIT_34 => X"000000cd00000000000000c800000000000000c100000000000000c400000000",
            INIT_35 => X"000000c900000000000000c500000000000000c500000000000000c600000000",
            INIT_36 => X"000000c300000000000000c600000000000000c800000000000000c500000000",
            INIT_37 => X"000000c300000000000000cf00000000000000cb00000000000000c500000000",
            INIT_38 => X"000000ac00000000000000a3000000000000009b000000000000009900000000",
            INIT_39 => X"000000d100000000000000c700000000000000bc00000000000000ac00000000",
            INIT_3A => X"000000bf00000000000000bd00000000000000be00000000000000c400000000",
            INIT_3B => X"000000c400000000000000bb00000000000000bc00000000000000c100000000",
            INIT_3C => X"000000ce00000000000000c400000000000000c200000000000000ca00000000",
            INIT_3D => X"000000c800000000000000c400000000000000c900000000000000c200000000",
            INIT_3E => X"000000c900000000000000c800000000000000bb00000000000000b500000000",
            INIT_3F => X"000000bd00000000000000c700000000000000c400000000000000c800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ac00000000000000a3000000000000009f00000000000000a000000000",
            INIT_41 => X"000000be00000000000000b000000000000000b000000000000000ae00000000",
            INIT_42 => X"000000b000000000000000b000000000000000af00000000000000b400000000",
            INIT_43 => X"000000b600000000000000ac00000000000000aa00000000000000b500000000",
            INIT_44 => X"000000bb00000000000000b500000000000000b200000000000000bb00000000",
            INIT_45 => X"000000bb00000000000000b400000000000000bc00000000000000b100000000",
            INIT_46 => X"000000bc00000000000000bc00000000000000c400000000000000c700000000",
            INIT_47 => X"000000b800000000000000c200000000000000c000000000000000c500000000",
            INIT_48 => X"000000ac00000000000000a200000000000000a700000000000000ab00000000",
            INIT_49 => X"000000b000000000000000b400000000000000ab00000000000000aa00000000",
            INIT_4A => X"0000009c0000000000000096000000000000009c000000000000009b00000000",
            INIT_4B => X"0000009e00000000000000990000000000000092000000000000009600000000",
            INIT_4C => X"0000009d00000000000000a400000000000000a600000000000000a600000000",
            INIT_4D => X"000000a6000000000000009c00000000000000a2000000000000009d00000000",
            INIT_4E => X"000000bd00000000000000bc00000000000000c700000000000000c800000000",
            INIT_4F => X"000000b600000000000000c200000000000000c100000000000000c500000000",
            INIT_50 => X"000000b000000000000000a800000000000000b400000000000000af00000000",
            INIT_51 => X"000000ae00000000000000b600000000000000b100000000000000ad00000000",
            INIT_52 => X"0000009a000000000000009f00000000000000a0000000000000009c00000000",
            INIT_53 => X"000000ad00000000000000a800000000000000a3000000000000009f00000000",
            INIT_54 => X"000000a200000000000000a000000000000000a400000000000000aa00000000",
            INIT_55 => X"000000ac00000000000000a700000000000000a800000000000000a000000000",
            INIT_56 => X"000000c400000000000000c400000000000000c300000000000000c200000000",
            INIT_57 => X"000000b700000000000000c100000000000000bf00000000000000c500000000",
            INIT_58 => X"000000bb00000000000000b200000000000000bb00000000000000b500000000",
            INIT_59 => X"000000b600000000000000ae00000000000000aa00000000000000b700000000",
            INIT_5A => X"000000b500000000000000b400000000000000b300000000000000b300000000",
            INIT_5B => X"000000c100000000000000c100000000000000bb00000000000000b800000000",
            INIT_5C => X"000000b900000000000000bc00000000000000c000000000000000c100000000",
            INIT_5D => X"000000c000000000000000c000000000000000ba00000000000000b800000000",
            INIT_5E => X"000000bd00000000000000c000000000000000bc00000000000000bb00000000",
            INIT_5F => X"000000ba00000000000000c400000000000000bf00000000000000be00000000",
            INIT_60 => X"000000ab00000000000000ba00000000000000be00000000000000b900000000",
            INIT_61 => X"000000c100000000000000950000000000000084000000000000009900000000",
            INIT_62 => X"000000bc00000000000000ba00000000000000bf00000000000000c600000000",
            INIT_63 => X"000000c400000000000000c300000000000000c100000000000000bf00000000",
            INIT_64 => X"000000bc00000000000000be00000000000000c000000000000000c300000000",
            INIT_65 => X"000000bf00000000000000c000000000000000be00000000000000bc00000000",
            INIT_66 => X"000000c500000000000000c300000000000000c100000000000000bf00000000",
            INIT_67 => X"000000c100000000000000cc00000000000000ca00000000000000ca00000000",
            INIT_68 => X"0000009e00000000000000bc00000000000000c200000000000000ba00000000",
            INIT_69 => X"0000006d000000000000005e0000000000000074000000000000008400000000",
            INIT_6A => X"000000c200000000000000c200000000000000b1000000000000009100000000",
            INIT_6B => X"000000c700000000000000c400000000000000c100000000000000bf00000000",
            INIT_6C => X"000000c600000000000000c800000000000000c700000000000000c700000000",
            INIT_6D => X"000000c600000000000000c700000000000000c400000000000000c400000000",
            INIT_6E => X"000000c400000000000000c400000000000000c400000000000000c500000000",
            INIT_6F => X"000000b900000000000000c600000000000000c500000000000000c600000000",
            INIT_70 => X"000000c600000000000000c400000000000000c500000000000000ba00000000",
            INIT_71 => X"0000005c000000000000008d00000000000000b800000000000000c200000000",
            INIT_72 => X"000000b3000000000000008e0000000000000068000000000000005400000000",
            INIT_73 => X"000000cc00000000000000cc00000000000000c900000000000000c300000000",
            INIT_74 => X"000000c700000000000000cc00000000000000cc00000000000000cc00000000",
            INIT_75 => X"000000bf00000000000000c200000000000000c200000000000000c200000000",
            INIT_76 => X"000000be00000000000000be00000000000000be00000000000000bd00000000",
            INIT_77 => X"000000b500000000000000c000000000000000be00000000000000bf00000000",
            INIT_78 => X"000000c800000000000000c600000000000000c700000000000000b800000000",
            INIT_79 => X"000000b100000000000000c900000000000000c800000000000000c500000000",
            INIT_7A => X"00000080000000000000005d0000000000000054000000000000007500000000",
            INIT_7B => X"000000cd00000000000000d000000000000000ca00000000000000ad00000000",
            INIT_7C => X"000000c700000000000000c700000000000000c800000000000000ca00000000",
            INIT_7D => X"000000c300000000000000c500000000000000c400000000000000c300000000",
            INIT_7E => X"000000bf00000000000000c200000000000000c300000000000000c100000000",
            INIT_7F => X"000000b200000000000000be00000000000000bd00000000000000bf00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE18;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE19 : if BRAM_NAME = "sampleifmap_layersamples_instance19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d000000000000000cb00000000000000c900000000000000b900000000",
            INIT_01 => X"000000d600000000000000d000000000000000ce00000000000000cd00000000",
            INIT_02 => X"0000005b000000000000004c000000000000005c00000000000000af00000000",
            INIT_03 => X"000000cb00000000000000b5000000000000008c000000000000006900000000",
            INIT_04 => X"000000c200000000000000c500000000000000ca00000000000000ce00000000",
            INIT_05 => X"000000c200000000000000c200000000000000c200000000000000c100000000",
            INIT_06 => X"000000bf00000000000000c100000000000000c300000000000000c200000000",
            INIT_07 => X"000000b400000000000000be00000000000000be00000000000000c100000000",
            INIT_08 => X"000000d600000000000000cf00000000000000cc00000000000000bb00000000",
            INIT_09 => X"000000d000000000000000d300000000000000d400000000000000d400000000",
            INIT_0A => X"000000570000000000000047000000000000007c00000000000000cb00000000",
            INIT_0B => X"0000008400000000000000630000000000000054000000000000005400000000",
            INIT_0C => X"000000cb00000000000000cb00000000000000be00000000000000a700000000",
            INIT_0D => X"000000c400000000000000c500000000000000c000000000000000c300000000",
            INIT_0E => X"000000bf00000000000000c000000000000000c200000000000000c200000000",
            INIT_0F => X"000000b700000000000000c000000000000000bf00000000000000c100000000",
            INIT_10 => X"000000d600000000000000cf00000000000000cf00000000000000be00000000",
            INIT_11 => X"000000d000000000000000d300000000000000d300000000000000d400000000",
            INIT_12 => X"000000570000000000000048000000000000008900000000000000d300000000",
            INIT_13 => X"0000005300000000000000560000000000000054000000000000005300000000",
            INIT_14 => X"0000009b0000000000000083000000000000006b000000000000005900000000",
            INIT_15 => X"000000cc00000000000000cb00000000000000b600000000000000a300000000",
            INIT_16 => X"000000bf00000000000000c200000000000000c600000000000000ca00000000",
            INIT_17 => X"000000b600000000000000bf00000000000000c000000000000000c100000000",
            INIT_18 => X"000000d700000000000000d100000000000000d200000000000000bf00000000",
            INIT_19 => X"000000d500000000000000d400000000000000d400000000000000d500000000",
            INIT_1A => X"0000003a000000000000002f000000000000007100000000000000cc00000000",
            INIT_1B => X"0000005d0000000000000057000000000000004c000000000000003f00000000",
            INIT_1C => X"0000003e00000000000000460000000000000050000000000000005a00000000",
            INIT_1D => X"0000009f000000000000007a000000000000004d000000000000003a00000000",
            INIT_1E => X"000000c800000000000000c900000000000000c200000000000000b400000000",
            INIT_1F => X"000000b900000000000000c400000000000000c400000000000000c800000000",
            INIT_20 => X"000000d300000000000000cf00000000000000d000000000000000bf00000000",
            INIT_21 => X"000000d400000000000000d100000000000000d200000000000000d100000000",
            INIT_22 => X"0000002500000000000000410000000000000065000000000000009d00000000",
            INIT_23 => X"00000058000000000000004a0000000000000044000000000000003300000000",
            INIT_24 => X"0000004900000000000000550000000000000056000000000000005b00000000",
            INIT_25 => X"00000048000000000000003e000000000000002e000000000000003700000000",
            INIT_26 => X"0000009e0000000000000085000000000000006b000000000000004e00000000",
            INIT_27 => X"000000ba00000000000000c400000000000000c300000000000000b800000000",
            INIT_28 => X"000000d100000000000000cb00000000000000ca00000000000000ba00000000",
            INIT_29 => X"000000c800000000000000d100000000000000ce00000000000000cf00000000",
            INIT_2A => X"000000640000000000000097000000000000008c000000000000009500000000",
            INIT_2B => X"0000006000000000000000320000000000000035000000000000002d00000000",
            INIT_2C => X"00000048000000000000008000000000000000a0000000000000009c00000000",
            INIT_2D => X"0000004200000000000000590000000000000070000000000000006200000000",
            INIT_2E => X"000000a300000000000000a60000000000000083000000000000004300000000",
            INIT_2F => X"000000b200000000000000bc00000000000000b700000000000000ad00000000",
            INIT_30 => X"000000d200000000000000ca00000000000000c900000000000000b900000000",
            INIT_31 => X"000000d100000000000000d100000000000000d000000000000000d200000000",
            INIT_32 => X"000000bd00000000000000d700000000000000d300000000000000d200000000",
            INIT_33 => X"000000a800000000000000940000000000000092000000000000009000000000",
            INIT_34 => X"0000009a00000000000000c000000000000000ce00000000000000ca00000000",
            INIT_35 => X"0000009f00000000000000b100000000000000b200000000000000a300000000",
            INIT_36 => X"000000c200000000000000bf00000000000000b2000000000000009c00000000",
            INIT_37 => X"000000b000000000000000bc00000000000000c100000000000000c400000000",
            INIT_38 => X"000000c400000000000000c000000000000000bc00000000000000b000000000",
            INIT_39 => X"000000b700000000000000b900000000000000bc00000000000000c000000000",
            INIT_3A => X"000000ad00000000000000b300000000000000b200000000000000b600000000",
            INIT_3B => X"000000ad00000000000000ab00000000000000aa00000000000000aa00000000",
            INIT_3C => X"000000a700000000000000a100000000000000a000000000000000a900000000",
            INIT_3D => X"000000aa00000000000000a500000000000000a100000000000000a500000000",
            INIT_3E => X"00000096000000000000009800000000000000a000000000000000aa00000000",
            INIT_3F => X"0000009c00000000000000a400000000000000a3000000000000009d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006b000000000000006e0000000000000063000000000000007200000000",
            INIT_41 => X"0000005d000000000000005e0000000000000061000000000000006600000000",
            INIT_42 => X"0000005000000000000000580000000000000055000000000000005800000000",
            INIT_43 => X"000000650000000000000053000000000000004e000000000000004d00000000",
            INIT_44 => X"0000006b000000000000006a000000000000006c000000000000007100000000",
            INIT_45 => X"00000071000000000000006f000000000000006e000000000000006c00000000",
            INIT_46 => X"0000007700000000000000780000000000000077000000000000007500000000",
            INIT_47 => X"0000007c000000000000007a0000000000000079000000000000007800000000",
            INIT_48 => X"000000750000000000000071000000000000006d000000000000007a00000000",
            INIT_49 => X"0000007100000000000000720000000000000070000000000000007300000000",
            INIT_4A => X"0000006d000000000000006f0000000000000070000000000000006f00000000",
            INIT_4B => X"0000006c000000000000006e000000000000006d000000000000006e00000000",
            INIT_4C => X"0000006b00000000000000690000000000000070000000000000007300000000",
            INIT_4D => X"000000680000000000000065000000000000006a000000000000006c00000000",
            INIT_4E => X"0000006d000000000000006d000000000000006b000000000000006a00000000",
            INIT_4F => X"00000065000000000000005e0000000000000066000000000000006700000000",
            INIT_50 => X"00000070000000000000006b0000000000000061000000000000007800000000",
            INIT_51 => X"0000005e00000000000000620000000000000068000000000000006d00000000",
            INIT_52 => X"000000560000000000000058000000000000005d000000000000005e00000000",
            INIT_53 => X"0000004e0000000000000050000000000000004f000000000000005200000000",
            INIT_54 => X"000000450000000000000048000000000000004f000000000000005000000000",
            INIT_55 => X"0000004100000000000000410000000000000042000000000000004300000000",
            INIT_56 => X"0000004000000000000000420000000000000041000000000000004000000000",
            INIT_57 => X"0000004d0000000000000035000000000000003f000000000000004300000000",
            INIT_58 => X"0000004500000000000000410000000000000037000000000000005b00000000",
            INIT_59 => X"0000003d000000000000003f0000000000000042000000000000004200000000",
            INIT_5A => X"00000039000000000000003c0000000000000040000000000000004200000000",
            INIT_5B => X"0000003f000000000000003d000000000000003c000000000000003900000000",
            INIT_5C => X"0000003a00000000000000400000000000000042000000000000003f00000000",
            INIT_5D => X"0000003c000000000000003b0000000000000039000000000000003800000000",
            INIT_5E => X"0000003900000000000000380000000000000039000000000000003a00000000",
            INIT_5F => X"0000005c000000000000004b0000000000000031000000000000003400000000",
            INIT_60 => X"000000440000000000000042000000000000003c000000000000005d00000000",
            INIT_61 => X"0000004100000000000000400000000000000043000000000000004300000000",
            INIT_62 => X"0000003b000000000000003e0000000000000041000000000000004500000000",
            INIT_63 => X"0000003d000000000000003c000000000000003b000000000000003b00000000",
            INIT_64 => X"00000038000000000000003a000000000000003f000000000000004000000000",
            INIT_65 => X"0000003800000000000000380000000000000037000000000000003700000000",
            INIT_66 => X"000000350000000000000038000000000000003a000000000000003900000000",
            INIT_67 => X"000000510000000000000061000000000000005d000000000000004100000000",
            INIT_68 => X"00000039000000000000003d0000000000000039000000000000005900000000",
            INIT_69 => X"0000003b0000000000000039000000000000003b000000000000003900000000",
            INIT_6A => X"000000360000000000000038000000000000003a000000000000003c00000000",
            INIT_6B => X"0000003d000000000000003b000000000000003d000000000000003c00000000",
            INIT_6C => X"00000039000000000000003a000000000000003d000000000000004100000000",
            INIT_6D => X"0000003d000000000000003d000000000000003c000000000000003c00000000",
            INIT_6E => X"000000460000000000000039000000000000003e000000000000004200000000",
            INIT_6F => X"00000043000000000000003b0000000000000059000000000000006100000000",
            INIT_70 => X"0000003e000000000000003f000000000000003c000000000000005900000000",
            INIT_71 => X"0000003f000000000000003e000000000000003e000000000000003e00000000",
            INIT_72 => X"000000520000000000000041000000000000003d000000000000003e00000000",
            INIT_73 => X"00000051000000000000004e0000000000000051000000000000005400000000",
            INIT_74 => X"0000005300000000000000550000000000000054000000000000005800000000",
            INIT_75 => X"0000004000000000000000420000000000000043000000000000005000000000",
            INIT_76 => X"0000006700000000000000560000000000000038000000000000003400000000",
            INIT_77 => X"0000004b000000000000003d0000000000000039000000000000004c00000000",
            INIT_78 => X"0000003c000000000000003d000000000000003c000000000000005c00000000",
            INIT_79 => X"0000004100000000000000430000000000000042000000000000003f00000000",
            INIT_7A => X"0000004800000000000000410000000000000043000000000000004200000000",
            INIT_7B => X"0000004600000000000000480000000000000049000000000000004900000000",
            INIT_7C => X"0000004b000000000000004b000000000000004a000000000000004900000000",
            INIT_7D => X"0000003e00000000000000400000000000000040000000000000004b00000000",
            INIT_7E => X"0000004000000000000000580000000000000056000000000000004100000000",
            INIT_7F => X"000000490000000000000040000000000000003c000000000000003900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE19;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE20 : if BRAM_NAME = "sampleifmap_layersamples_instance20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000c000000000000000b300000000000000b0000000000000009c00000000",
            INIT_01 => X"000000ad00000000000000ad00000000000000ab00000000000000b900000000",
            INIT_02 => X"000000b800000000000000b600000000000000b300000000000000af00000000",
            INIT_03 => X"000000b500000000000000b600000000000000b800000000000000b900000000",
            INIT_04 => X"000000b900000000000000b700000000000000b300000000000000b300000000",
            INIT_05 => X"000000bd00000000000000bb00000000000000ba00000000000000ba00000000",
            INIT_06 => X"000000c300000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_07 => X"000000b700000000000000ca00000000000000c400000000000000c500000000",
            INIT_08 => X"000000c300000000000000b800000000000000b3000000000000009b00000000",
            INIT_09 => X"000000a4000000000000009f00000000000000a200000000000000be00000000",
            INIT_0A => X"000000b000000000000000a900000000000000a500000000000000a300000000",
            INIT_0B => X"000000a700000000000000a400000000000000ae00000000000000ab00000000",
            INIT_0C => X"000000a600000000000000a800000000000000a600000000000000ac00000000",
            INIT_0D => X"000000a900000000000000ab00000000000000af00000000000000a900000000",
            INIT_0E => X"000000cc00000000000000bf00000000000000ae00000000000000aa00000000",
            INIT_0F => X"000000be00000000000000d700000000000000d000000000000000ce00000000",
            INIT_10 => X"000000c400000000000000b900000000000000b2000000000000009a00000000",
            INIT_11 => X"000000a800000000000000b200000000000000c100000000000000cb00000000",
            INIT_12 => X"000000c400000000000000be00000000000000af00000000000000a000000000",
            INIT_13 => X"000000bc00000000000000be00000000000000c500000000000000c300000000",
            INIT_14 => X"000000c300000000000000c200000000000000c300000000000000c400000000",
            INIT_15 => X"000000bf00000000000000c100000000000000c600000000000000c400000000",
            INIT_16 => X"000000cd00000000000000cd00000000000000c400000000000000c000000000",
            INIT_17 => X"000000bf00000000000000d700000000000000d000000000000000ce00000000",
            INIT_18 => X"000000c300000000000000bc00000000000000b2000000000000009a00000000",
            INIT_19 => X"0000008000000000000000bc00000000000000c500000000000000ca00000000",
            INIT_1A => X"0000009b000000000000009a0000000000000098000000000000006c00000000",
            INIT_1B => X"0000009400000000000000950000000000000095000000000000009e00000000",
            INIT_1C => X"000000ad00000000000000a300000000000000a100000000000000a700000000",
            INIT_1D => X"0000009f00000000000000ae00000000000000a300000000000000a800000000",
            INIT_1E => X"000000ce00000000000000cc00000000000000d000000000000000bc00000000",
            INIT_1F => X"000000bc00000000000000d400000000000000cd00000000000000cc00000000",
            INIT_20 => X"000000bf00000000000000bb00000000000000b1000000000000009a00000000",
            INIT_21 => X"0000007e00000000000000bd00000000000000c400000000000000c600000000",
            INIT_22 => X"0000006b000000000000006a000000000000008b000000000000008000000000",
            INIT_23 => X"0000007100000000000000760000000000000078000000000000007300000000",
            INIT_24 => X"0000007e00000000000000720000000000000072000000000000007700000000",
            INIT_25 => X"0000007000000000000000880000000000000070000000000000007600000000",
            INIT_26 => X"000000ce00000000000000c900000000000000cb00000000000000a000000000",
            INIT_27 => X"000000be00000000000000d600000000000000cd00000000000000ce00000000",
            INIT_28 => X"000000bd00000000000000bb00000000000000ae000000000000009700000000",
            INIT_29 => X"0000009300000000000000b700000000000000c800000000000000c500000000",
            INIT_2A => X"000000a5000000000000009100000000000000a800000000000000a900000000",
            INIT_2B => X"0000009d0000000000000095000000000000009200000000000000aa00000000",
            INIT_2C => X"000000bd00000000000000b000000000000000b200000000000000b400000000",
            INIT_2D => X"000000b100000000000000bc00000000000000b300000000000000b000000000",
            INIT_2E => X"000000d000000000000000cf00000000000000d000000000000000c400000000",
            INIT_2F => X"000000be00000000000000d800000000000000d100000000000000d000000000",
            INIT_30 => X"000000bd00000000000000b900000000000000ac000000000000009800000000",
            INIT_31 => X"00000060000000000000009300000000000000c600000000000000c200000000",
            INIT_32 => X"0000009800000000000000900000000000000097000000000000009500000000",
            INIT_33 => X"0000008b00000000000000800000000000000079000000000000009800000000",
            INIT_34 => X"000000a200000000000000aa0000000000000097000000000000009c00000000",
            INIT_35 => X"000000a4000000000000009600000000000000ad000000000000009600000000",
            INIT_36 => X"000000d200000000000000cc00000000000000a6000000000000009c00000000",
            INIT_37 => X"000000bc00000000000000d400000000000000cf00000000000000d300000000",
            INIT_38 => X"000000bb00000000000000b600000000000000ac000000000000009b00000000",
            INIT_39 => X"00000065000000000000007700000000000000b500000000000000c200000000",
            INIT_3A => X"0000007800000000000000830000000000000083000000000000007b00000000",
            INIT_3B => X"0000007f00000000000000870000000000000087000000000000009200000000",
            INIT_3C => X"0000007b0000000000000083000000000000007b000000000000007b00000000",
            INIT_3D => X"0000009f000000000000007b0000000000000084000000000000006d00000000",
            INIT_3E => X"000000c700000000000000bf0000000000000084000000000000007b00000000",
            INIT_3F => X"000000ba00000000000000d000000000000000c900000000000000c900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b900000000000000b400000000000000af00000000000000a100000000",
            INIT_41 => X"000000af00000000000000ab00000000000000ba00000000000000c000000000",
            INIT_42 => X"000000a600000000000000ac00000000000000a500000000000000a200000000",
            INIT_43 => X"000000aa00000000000000ad00000000000000ac00000000000000af00000000",
            INIT_44 => X"000000af00000000000000b200000000000000b200000000000000ac00000000",
            INIT_45 => X"000000be00000000000000b200000000000000ac00000000000000a300000000",
            INIT_46 => X"000000cd00000000000000c800000000000000b000000000000000ac00000000",
            INIT_47 => X"000000b900000000000000d100000000000000c900000000000000c800000000",
            INIT_48 => X"000000ba00000000000000b400000000000000b700000000000000ac00000000",
            INIT_49 => X"000000b700000000000000c200000000000000c000000000000000be00000000",
            INIT_4A => X"000000a300000000000000a200000000000000a500000000000000a000000000",
            INIT_4B => X"000000a200000000000000a4000000000000009e000000000000009f00000000",
            INIT_4C => X"000000a200000000000000ac00000000000000ae00000000000000a700000000",
            INIT_4D => X"000000b600000000000000a500000000000000a300000000000000a000000000",
            INIT_4E => X"000000cd00000000000000ca00000000000000c600000000000000c800000000",
            INIT_4F => X"000000b800000000000000d000000000000000ca00000000000000ca00000000",
            INIT_50 => X"000000be00000000000000ba00000000000000c400000000000000b100000000",
            INIT_51 => X"000000b700000000000000c100000000000000c100000000000000c000000000",
            INIT_52 => X"0000009f00000000000000a500000000000000a700000000000000a300000000",
            INIT_53 => X"000000ac00000000000000aa00000000000000a600000000000000a400000000",
            INIT_54 => X"000000ab00000000000000a600000000000000a600000000000000a800000000",
            INIT_55 => X"000000b200000000000000ab00000000000000ad00000000000000a800000000",
            INIT_56 => X"000000c700000000000000c700000000000000c600000000000000c700000000",
            INIT_57 => X"000000b800000000000000d000000000000000c800000000000000c800000000",
            INIT_58 => X"000000c800000000000000c300000000000000cc00000000000000b700000000",
            INIT_59 => X"000000c600000000000000be00000000000000bb00000000000000c900000000",
            INIT_5A => X"000000c100000000000000c100000000000000c100000000000000c200000000",
            INIT_5B => X"000000c600000000000000c600000000000000c200000000000000c100000000",
            INIT_5C => X"000000c600000000000000c300000000000000c300000000000000c600000000",
            INIT_5D => X"000000c500000000000000c400000000000000c400000000000000c500000000",
            INIT_5E => X"000000c900000000000000c900000000000000cb00000000000000c900000000",
            INIT_5F => X"000000bb00000000000000d100000000000000c800000000000000ca00000000",
            INIT_60 => X"000000b200000000000000c600000000000000cd00000000000000b900000000",
            INIT_61 => X"000000c4000000000000009a000000000000008d00000000000000a600000000",
            INIT_62 => X"000000c500000000000000c700000000000000ca00000000000000ca00000000",
            INIT_63 => X"000000ca00000000000000c900000000000000c700000000000000c500000000",
            INIT_64 => X"000000c400000000000000c600000000000000c700000000000000c900000000",
            INIT_65 => X"000000c600000000000000c700000000000000c600000000000000c400000000",
            INIT_66 => X"000000ce00000000000000cb00000000000000ca00000000000000c700000000",
            INIT_67 => X"000000bd00000000000000d400000000000000ce00000000000000cf00000000",
            INIT_68 => X"000000a500000000000000c800000000000000d000000000000000ba00000000",
            INIT_69 => X"0000006b000000000000005f000000000000007c000000000000009000000000",
            INIT_6A => X"000000c700000000000000c700000000000000b3000000000000008f00000000",
            INIT_6B => X"000000cc00000000000000c900000000000000c600000000000000c500000000",
            INIT_6C => X"000000cc00000000000000ce00000000000000cd00000000000000cc00000000",
            INIT_6D => X"000000cd00000000000000cd00000000000000c900000000000000c900000000",
            INIT_6E => X"000000cb00000000000000cb00000000000000cb00000000000000cc00000000",
            INIT_6F => X"000000b700000000000000cf00000000000000ca00000000000000ca00000000",
            INIT_70 => X"000000cc00000000000000d000000000000000d400000000000000ba00000000",
            INIT_71 => X"0000005b000000000000008f00000000000000c100000000000000ce00000000",
            INIT_72 => X"000000b5000000000000008e0000000000000065000000000000005100000000",
            INIT_73 => X"000000cf00000000000000cf00000000000000cc00000000000000c600000000",
            INIT_74 => X"000000ca00000000000000cf00000000000000cf00000000000000cf00000000",
            INIT_75 => X"000000c500000000000000c600000000000000c500000000000000c500000000",
            INIT_76 => X"000000c500000000000000c500000000000000c500000000000000c500000000",
            INIT_77 => X"000000b500000000000000cc00000000000000c500000000000000c400000000",
            INIT_78 => X"000000ce00000000000000d200000000000000d600000000000000b800000000",
            INIT_79 => X"000000b300000000000000cf00000000000000d400000000000000d100000000",
            INIT_7A => X"00000080000000000000005d0000000000000053000000000000007400000000",
            INIT_7B => X"000000ce00000000000000d200000000000000cb00000000000000ae00000000",
            INIT_7C => X"000000c900000000000000ca00000000000000ca00000000000000cc00000000",
            INIT_7D => X"000000c900000000000000c900000000000000c700000000000000c600000000",
            INIT_7E => X"000000c700000000000000c900000000000000ca00000000000000c800000000",
            INIT_7F => X"000000b400000000000000cb00000000000000c600000000000000c600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE20;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE21 : if BRAM_NAME = "sampleifmap_layersamples_instance21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d500000000000000d600000000000000d700000000000000ba00000000",
            INIT_01 => X"000000d900000000000000d400000000000000d600000000000000d600000000",
            INIT_02 => X"000000560000000000000049000000000000005b00000000000000af00000000",
            INIT_03 => X"000000cc00000000000000b5000000000000008a000000000000006500000000",
            INIT_04 => X"000000c600000000000000c700000000000000cb00000000000000d000000000",
            INIT_05 => X"000000c800000000000000c900000000000000c900000000000000c700000000",
            INIT_06 => X"000000c900000000000000c900000000000000ca00000000000000c800000000",
            INIT_07 => X"000000b600000000000000cc00000000000000c800000000000000ca00000000",
            INIT_08 => X"000000d900000000000000d800000000000000d800000000000000bb00000000",
            INIT_09 => X"000000d300000000000000d600000000000000d900000000000000db00000000",
            INIT_0A => X"000000520000000000000044000000000000007b00000000000000cc00000000",
            INIT_0B => X"0000008200000000000000610000000000000051000000000000004f00000000",
            INIT_0C => X"000000ca00000000000000c900000000000000bc00000000000000a500000000",
            INIT_0D => X"000000c600000000000000c700000000000000c100000000000000c400000000",
            INIT_0E => X"000000c800000000000000c800000000000000c700000000000000c600000000",
            INIT_0F => X"000000b600000000000000cc00000000000000c700000000000000c900000000",
            INIT_10 => X"000000d600000000000000d500000000000000d900000000000000bc00000000",
            INIT_11 => X"000000d200000000000000d600000000000000d800000000000000d800000000",
            INIT_12 => X"000000530000000000000046000000000000008800000000000000d400000000",
            INIT_13 => X"0000004d00000000000000500000000000000050000000000000004e00000000",
            INIT_14 => X"00000097000000000000007e0000000000000066000000000000005300000000",
            INIT_15 => X"000000cc00000000000000c900000000000000b2000000000000009f00000000",
            INIT_16 => X"000000c600000000000000c800000000000000c900000000000000cb00000000",
            INIT_17 => X"000000b400000000000000c900000000000000c500000000000000c700000000",
            INIT_18 => X"000000d500000000000000d600000000000000da00000000000000bb00000000",
            INIT_19 => X"000000d800000000000000d700000000000000d800000000000000d700000000",
            INIT_1A => X"00000037000000000000002d000000000000007000000000000000cc00000000",
            INIT_1B => X"00000051000000000000004d0000000000000045000000000000003a00000000",
            INIT_1C => X"0000003e0000000000000046000000000000004d000000000000005000000000",
            INIT_1D => X"000000a0000000000000007c000000000000004f000000000000003b00000000",
            INIT_1E => X"000000cd00000000000000cd00000000000000c400000000000000b500000000",
            INIT_1F => X"000000b400000000000000ca00000000000000c800000000000000cb00000000",
            INIT_20 => X"000000d100000000000000d200000000000000d800000000000000bc00000000",
            INIT_21 => X"000000d400000000000000d400000000000000d600000000000000d300000000",
            INIT_22 => X"00000021000000000000003a000000000000005f000000000000009a00000000",
            INIT_23 => X"0000004d0000000000000041000000000000003e000000000000003000000000",
            INIT_24 => X"0000004800000000000000540000000000000054000000000000005200000000",
            INIT_25 => X"00000048000000000000003f000000000000002f000000000000003800000000",
            INIT_26 => X"0000009e0000000000000084000000000000006b000000000000004e00000000",
            INIT_27 => X"000000b600000000000000ca00000000000000c100000000000000b500000000",
            INIT_28 => X"000000cf00000000000000ce00000000000000d200000000000000b800000000",
            INIT_29 => X"000000c800000000000000d400000000000000d300000000000000d100000000",
            INIT_2A => X"00000061000000000000008f0000000000000085000000000000009100000000",
            INIT_2B => X"0000005a000000000000002e0000000000000032000000000000002d00000000",
            INIT_2C => X"00000047000000000000007f000000000000009e000000000000009600000000",
            INIT_2D => X"0000004100000000000000580000000000000070000000000000006100000000",
            INIT_2E => X"000000a200000000000000a50000000000000082000000000000004300000000",
            INIT_2F => X"000000b000000000000000c500000000000000b500000000000000a800000000",
            INIT_30 => X"000000d000000000000000cd00000000000000d200000000000000b700000000",
            INIT_31 => X"000000d200000000000000d500000000000000d400000000000000d300000000",
            INIT_32 => X"000000bf00000000000000d400000000000000d100000000000000d100000000",
            INIT_33 => X"000000a600000000000000930000000000000093000000000000009400000000",
            INIT_34 => X"0000009d00000000000000c300000000000000d000000000000000c800000000",
            INIT_35 => X"000000a200000000000000b400000000000000b500000000000000a600000000",
            INIT_36 => X"000000c500000000000000c100000000000000b4000000000000009f00000000",
            INIT_37 => X"000000b100000000000000c700000000000000c100000000000000c300000000",
            INIT_38 => X"000000c200000000000000c300000000000000c400000000000000ae00000000",
            INIT_39 => X"000000b900000000000000bb00000000000000be00000000000000c200000000",
            INIT_3A => X"000000b500000000000000b700000000000000b500000000000000b800000000",
            INIT_3B => X"000000ad00000000000000ae00000000000000b000000000000000b200000000",
            INIT_3C => X"000000ac00000000000000a600000000000000a400000000000000aa00000000",
            INIT_3D => X"000000b000000000000000aa00000000000000a600000000000000aa00000000",
            INIT_3E => X"0000009b000000000000009d00000000000000a500000000000000af00000000",
            INIT_3F => X"0000009e00000000000000af00000000000000a3000000000000009d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000690000000000000070000000000000006c000000000000007000000000",
            INIT_41 => X"0000006000000000000000610000000000000064000000000000006700000000",
            INIT_42 => X"00000057000000000000005e000000000000005a000000000000005c00000000",
            INIT_43 => X"0000006700000000000000570000000000000053000000000000005400000000",
            INIT_44 => X"00000070000000000000006f0000000000000070000000000000007300000000",
            INIT_45 => X"0000007600000000000000740000000000000073000000000000007100000000",
            INIT_46 => X"0000007b000000000000007c000000000000007b000000000000007a00000000",
            INIT_47 => X"0000007c0000000000000084000000000000007a000000000000007900000000",
            INIT_48 => X"0000007000000000000000710000000000000073000000000000007500000000",
            INIT_49 => X"000000710000000000000071000000000000006f000000000000007100000000",
            INIT_4A => X"0000006e000000000000006f0000000000000070000000000000006f00000000",
            INIT_4B => X"0000006b000000000000006e000000000000006d000000000000006e00000000",
            INIT_4C => X"0000006e000000000000006c0000000000000073000000000000007300000000",
            INIT_4D => X"0000006b0000000000000068000000000000006d000000000000006f00000000",
            INIT_4E => X"000000700000000000000070000000000000006e000000000000006d00000000",
            INIT_4F => X"000000650000000000000062000000000000005f000000000000006400000000",
            INIT_50 => X"0000006a00000000000000690000000000000066000000000000007100000000",
            INIT_51 => X"0000005d00000000000000610000000000000066000000000000006a00000000",
            INIT_52 => X"000000550000000000000059000000000000005e000000000000005f00000000",
            INIT_53 => X"0000004e000000000000004f000000000000004e000000000000005200000000",
            INIT_54 => X"000000440000000000000047000000000000004f000000000000005000000000",
            INIT_55 => X"0000004100000000000000410000000000000041000000000000004300000000",
            INIT_56 => X"0000004100000000000000420000000000000042000000000000004100000000",
            INIT_57 => X"0000006400000000000000470000000000000037000000000000003c00000000",
            INIT_58 => X"000000400000000000000041000000000000003c000000000000005400000000",
            INIT_59 => X"0000003c000000000000003e0000000000000040000000000000004000000000",
            INIT_5A => X"00000038000000000000003d0000000000000040000000000000004200000000",
            INIT_5B => X"0000003f000000000000003d000000000000003c000000000000003900000000",
            INIT_5C => X"0000003b00000000000000410000000000000043000000000000004000000000",
            INIT_5D => X"0000003c000000000000003b000000000000003a000000000000003800000000",
            INIT_5E => X"0000003800000000000000380000000000000039000000000000003a00000000",
            INIT_5F => X"0000008000000000000000750000000000000048000000000000003800000000",
            INIT_60 => X"0000003e000000000000003f000000000000003b000000000000005300000000",
            INIT_61 => X"0000003f000000000000003d0000000000000041000000000000003f00000000",
            INIT_62 => X"00000039000000000000003c000000000000003e000000000000004300000000",
            INIT_63 => X"0000003d000000000000003c000000000000003a000000000000003a00000000",
            INIT_64 => X"0000003e00000000000000400000000000000044000000000000004100000000",
            INIT_65 => X"0000003d000000000000003e000000000000003c000000000000003d00000000",
            INIT_66 => X"00000041000000000000003d000000000000003a000000000000003a00000000",
            INIT_67 => X"0000006300000000000000890000000000000088000000000000005b00000000",
            INIT_68 => X"00000039000000000000003d0000000000000035000000000000004f00000000",
            INIT_69 => X"0000003c000000000000003a000000000000003b000000000000003700000000",
            INIT_6A => X"000000370000000000000039000000000000003c000000000000003d00000000",
            INIT_6B => X"0000003f000000000000003d000000000000003e000000000000003c00000000",
            INIT_6C => X"0000003b000000000000003c000000000000003f000000000000004300000000",
            INIT_6D => X"0000003f0000000000000040000000000000003e000000000000003e00000000",
            INIT_6E => X"0000006e0000000000000047000000000000003c000000000000003e00000000",
            INIT_6F => X"0000004a000000000000004f0000000000000077000000000000008e00000000",
            INIT_70 => X"000000410000000000000042000000000000003a000000000000005200000000",
            INIT_71 => X"0000003e000000000000003e000000000000003e000000000000003f00000000",
            INIT_72 => X"0000004f0000000000000041000000000000003e000000000000003f00000000",
            INIT_73 => X"0000004d000000000000004a000000000000004c000000000000004f00000000",
            INIT_74 => X"0000004e00000000000000500000000000000050000000000000005400000000",
            INIT_75 => X"00000041000000000000003e000000000000003f000000000000004c00000000",
            INIT_76 => X"0000008d000000000000007c0000000000000056000000000000004200000000",
            INIT_77 => X"0000004500000000000000400000000000000042000000000000006600000000",
            INIT_78 => X"0000003a000000000000003a0000000000000034000000000000004e00000000",
            INIT_79 => X"00000039000000000000003b000000000000003a000000000000003a00000000",
            INIT_7A => X"00000045000000000000003a000000000000003b000000000000003a00000000",
            INIT_7B => X"0000004500000000000000460000000000000047000000000000004700000000",
            INIT_7C => X"0000004a00000000000000490000000000000048000000000000004800000000",
            INIT_7D => X"00000044000000000000003f000000000000003f000000000000004900000000",
            INIT_7E => X"0000005800000000000000800000000000000080000000000000005a00000000",
            INIT_7F => X"000000440000000000000041000000000000003f000000000000004200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE21;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE22 : if BRAM_NAME = "sampleifmap_layersamples_instance22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000cd00000000000000c100000000000000bb000000000000009500000000",
            INIT_01 => X"000000b400000000000000b500000000000000b700000000000000ca00000000",
            INIT_02 => X"000000c000000000000000c100000000000000bd00000000000000b600000000",
            INIT_03 => X"000000bd00000000000000bd00000000000000c000000000000000c000000000",
            INIT_04 => X"000000c000000000000000bd00000000000000b900000000000000ba00000000",
            INIT_05 => X"000000be00000000000000c000000000000000c100000000000000c100000000",
            INIT_06 => X"000000c300000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_07 => X"000000ab00000000000000d400000000000000d100000000000000ca00000000",
            INIT_08 => X"000000e300000000000000d700000000000000cc000000000000009d00000000",
            INIT_09 => X"000000b300000000000000b300000000000000be00000000000000e000000000",
            INIT_0A => X"000000c300000000000000c300000000000000bb00000000000000b300000000",
            INIT_0B => X"000000b700000000000000b400000000000000be00000000000000bb00000000",
            INIT_0C => X"000000b700000000000000b800000000000000b700000000000000bc00000000",
            INIT_0D => X"000000bc00000000000000bc00000000000000bf00000000000000b900000000",
            INIT_0E => X"000000e000000000000000d300000000000000c200000000000000be00000000",
            INIT_0F => X"000000b700000000000000e300000000000000de00000000000000df00000000",
            INIT_10 => X"000000db00000000000000d500000000000000c9000000000000009900000000",
            INIT_11 => X"000000b800000000000000c400000000000000d500000000000000df00000000",
            INIT_12 => X"000000d400000000000000d300000000000000c300000000000000b100000000",
            INIT_13 => X"000000ca00000000000000cc00000000000000d200000000000000d000000000",
            INIT_14 => X"000000d100000000000000d000000000000000d100000000000000d100000000",
            INIT_15 => X"000000d000000000000000d000000000000000d400000000000000d200000000",
            INIT_16 => X"000000df00000000000000de00000000000000d500000000000000d000000000",
            INIT_17 => X"000000b800000000000000e000000000000000d700000000000000da00000000",
            INIT_18 => X"000000de00000000000000d300000000000000cf00000000000000a600000000",
            INIT_19 => X"0000008300000000000000c900000000000000dc00000000000000e200000000",
            INIT_1A => X"000000b100000000000000a6000000000000009e000000000000007700000000",
            INIT_1B => X"000000ab00000000000000a600000000000000a700000000000000b200000000",
            INIT_1C => X"000000ba00000000000000b200000000000000b200000000000000b700000000",
            INIT_1D => X"000000a500000000000000b400000000000000ba00000000000000b900000000",
            INIT_1E => X"000000dd00000000000000dc00000000000000e400000000000000cf00000000",
            INIT_1F => X"000000ba00000000000000e600000000000000df00000000000000e000000000",
            INIT_20 => X"000000da00000000000000ca00000000000000cb00000000000000a700000000",
            INIT_21 => X"0000008e00000000000000d600000000000000e100000000000000e000000000",
            INIT_22 => X"0000008100000000000000780000000000000098000000000000009900000000",
            INIT_23 => X"00000083000000000000007c000000000000007e000000000000008100000000",
            INIT_24 => X"0000008a00000000000000820000000000000084000000000000008600000000",
            INIT_25 => X"0000007b000000000000008d0000000000000088000000000000008800000000",
            INIT_26 => X"000000d900000000000000da00000000000000e300000000000000ba00000000",
            INIT_27 => X"000000b900000000000000e300000000000000dc00000000000000de00000000",
            INIT_28 => X"000000d900000000000000cb00000000000000c900000000000000a400000000",
            INIT_29 => X"000000a500000000000000d100000000000000da00000000000000dc00000000",
            INIT_2A => X"000000b4000000000000009c00000000000000b500000000000000c400000000",
            INIT_2B => X"000000ac00000000000000a300000000000000a000000000000000b300000000",
            INIT_2C => X"000000c900000000000000be00000000000000c100000000000000bf00000000",
            INIT_2D => X"000000be00000000000000c600000000000000c000000000000000bf00000000",
            INIT_2E => X"000000e100000000000000e100000000000000e100000000000000d400000000",
            INIT_2F => X"000000bc00000000000000e800000000000000e100000000000000df00000000",
            INIT_30 => X"000000d900000000000000c800000000000000c600000000000000a400000000",
            INIT_31 => X"0000006800000000000000ac00000000000000d600000000000000d900000000",
            INIT_32 => X"000000af00000000000000a600000000000000a5000000000000009e00000000",
            INIT_33 => X"000000a00000000000000097000000000000009000000000000000a500000000",
            INIT_34 => X"000000b600000000000000bd00000000000000ad00000000000000b200000000",
            INIT_35 => X"000000b900000000000000ad00000000000000b700000000000000aa00000000",
            INIT_36 => X"000000e200000000000000dc00000000000000b200000000000000a600000000",
            INIT_37 => X"000000bc00000000000000e700000000000000e000000000000000dd00000000",
            INIT_38 => X"000000d800000000000000c700000000000000c900000000000000a900000000",
            INIT_39 => X"0000006f000000000000009200000000000000cb00000000000000da00000000",
            INIT_3A => X"00000090000000000000009d0000000000000095000000000000008600000000",
            INIT_3B => X"00000090000000000000008f000000000000008f000000000000009b00000000",
            INIT_3C => X"0000008e0000000000000094000000000000008e000000000000009300000000",
            INIT_3D => X"000000b0000000000000008e000000000000008d000000000000007f00000000",
            INIT_3E => X"000000dc00000000000000d10000000000000095000000000000008900000000",
            INIT_3F => X"000000ba00000000000000e400000000000000dc00000000000000d900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d900000000000000c700000000000000ce00000000000000b100000000",
            INIT_41 => X"000000c500000000000000c100000000000000cd00000000000000db00000000",
            INIT_42 => X"000000b800000000000000bb00000000000000b700000000000000b800000000",
            INIT_43 => X"000000bd00000000000000bb00000000000000ba00000000000000c000000000",
            INIT_44 => X"000000bf00000000000000c200000000000000c200000000000000c000000000",
            INIT_45 => X"000000c800000000000000bc00000000000000ba00000000000000b200000000",
            INIT_46 => X"000000db00000000000000d600000000000000c600000000000000c100000000",
            INIT_47 => X"000000b900000000000000e400000000000000dd00000000000000db00000000",
            INIT_48 => X"000000d600000000000000c500000000000000d400000000000000ba00000000",
            INIT_49 => X"000000d200000000000000dc00000000000000d600000000000000d700000000",
            INIT_4A => X"000000ba00000000000000b600000000000000bb00000000000000b900000000",
            INIT_4B => X"000000ba00000000000000b900000000000000b400000000000000b600000000",
            INIT_4C => X"000000b800000000000000c300000000000000c600000000000000c100000000",
            INIT_4D => X"000000c600000000000000b600000000000000b600000000000000b500000000",
            INIT_4E => X"000000df00000000000000dd00000000000000de00000000000000de00000000",
            INIT_4F => X"000000b700000000000000e300000000000000de00000000000000df00000000",
            INIT_50 => X"000000d800000000000000c800000000000000de00000000000000bc00000000",
            INIT_51 => X"000000cc00000000000000d600000000000000d400000000000000d700000000",
            INIT_52 => X"000000b000000000000000b600000000000000b800000000000000b500000000",
            INIT_53 => X"000000bf00000000000000bc00000000000000b800000000000000b500000000",
            INIT_54 => X"000000b900000000000000b800000000000000ba00000000000000bd00000000",
            INIT_55 => X"000000c900000000000000ba00000000000000b800000000000000b600000000",
            INIT_56 => X"000000db00000000000000dc00000000000000dd00000000000000df00000000",
            INIT_57 => X"000000b800000000000000e300000000000000dc00000000000000db00000000",
            INIT_58 => X"000000e000000000000000cf00000000000000e200000000000000bf00000000",
            INIT_59 => X"000000de00000000000000d700000000000000d100000000000000dc00000000",
            INIT_5A => X"000000d700000000000000d600000000000000d700000000000000d900000000",
            INIT_5B => X"000000df00000000000000df00000000000000db00000000000000d900000000",
            INIT_5C => X"000000da00000000000000db00000000000000dd00000000000000df00000000",
            INIT_5D => X"000000db00000000000000d900000000000000d600000000000000d800000000",
            INIT_5E => X"000000d600000000000000d900000000000000db00000000000000db00000000",
            INIT_5F => X"000000ba00000000000000e300000000000000db00000000000000d700000000",
            INIT_60 => X"000000ce00000000000000d400000000000000dc00000000000000bc00000000",
            INIT_61 => X"000000d900000000000000ac000000000000009900000000000000b500000000",
            INIT_62 => X"000000dc00000000000000dd00000000000000e100000000000000e200000000",
            INIT_63 => X"000000e200000000000000e100000000000000df00000000000000de00000000",
            INIT_64 => X"000000da00000000000000dc00000000000000dd00000000000000e100000000",
            INIT_65 => X"000000da00000000000000dc00000000000000db00000000000000d900000000",
            INIT_66 => X"000000e000000000000000de00000000000000dc00000000000000d900000000",
            INIT_67 => X"000000bb00000000000000e600000000000000e000000000000000e000000000",
            INIT_68 => X"000000c100000000000000d600000000000000df00000000000000bd00000000",
            INIT_69 => X"000000730000000000000063000000000000007e000000000000009d00000000",
            INIT_6A => X"000000dd00000000000000dd00000000000000c6000000000000009d00000000",
            INIT_6B => X"000000e200000000000000df00000000000000dc00000000000000da00000000",
            INIT_6C => X"000000df00000000000000e100000000000000e000000000000000e200000000",
            INIT_6D => X"000000e000000000000000e000000000000000dd00000000000000dc00000000",
            INIT_6E => X"000000de00000000000000de00000000000000de00000000000000df00000000",
            INIT_6F => X"000000b700000000000000e200000000000000dd00000000000000dd00000000",
            INIT_70 => X"000000e900000000000000de00000000000000e200000000000000bd00000000",
            INIT_71 => X"0000005a000000000000009200000000000000c400000000000000dc00000000",
            INIT_72 => X"000000ca00000000000000a10000000000000071000000000000005400000000",
            INIT_73 => X"000000e400000000000000e300000000000000e000000000000000da00000000",
            INIT_74 => X"000000dc00000000000000e000000000000000e100000000000000e200000000",
            INIT_75 => X"000000d900000000000000d800000000000000d700000000000000d700000000",
            INIT_76 => X"000000d800000000000000d800000000000000d800000000000000d800000000",
            INIT_77 => X"000000b600000000000000e100000000000000da00000000000000d700000000",
            INIT_78 => X"000000ea00000000000000e000000000000000e500000000000000bb00000000",
            INIT_79 => X"000000b300000000000000da00000000000000e100000000000000e100000000",
            INIT_7A => X"00000091000000000000006a0000000000000058000000000000007300000000",
            INIT_7B => X"000000e100000000000000e400000000000000dd00000000000000c000000000",
            INIT_7C => X"000000d900000000000000da00000000000000db00000000000000df00000000",
            INIT_7D => X"000000db00000000000000d900000000000000d600000000000000d600000000",
            INIT_7E => X"000000da00000000000000dc00000000000000dd00000000000000db00000000",
            INIT_7F => X"000000b700000000000000e200000000000000dc00000000000000d900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE22;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE23 : if BRAM_NAME = "sampleifmap_layersamples_instance23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e900000000000000de00000000000000e900000000000000be00000000",
            INIT_01 => X"000000e100000000000000e000000000000000e200000000000000e400000000",
            INIT_02 => X"0000005b0000000000000050000000000000006200000000000000b500000000",
            INIT_03 => X"000000d900000000000000c00000000000000092000000000000006a00000000",
            INIT_04 => X"000000da00000000000000dd00000000000000e100000000000000e000000000",
            INIT_05 => X"000000d900000000000000da00000000000000da00000000000000d900000000",
            INIT_06 => X"000000dd00000000000000dd00000000000000dd00000000000000da00000000",
            INIT_07 => X"000000bc00000000000000e300000000000000dc00000000000000dd00000000",
            INIT_08 => X"000000e900000000000000dd00000000000000ea00000000000000bf00000000",
            INIT_09 => X"000000dd00000000000000e200000000000000e300000000000000e700000000",
            INIT_0A => X"0000004f0000000000000049000000000000008200000000000000d500000000",
            INIT_0B => X"0000008800000000000000640000000000000050000000000000004b00000000",
            INIT_0C => X"000000dc00000000000000d700000000000000c800000000000000ad00000000",
            INIT_0D => X"000000de00000000000000df00000000000000d900000000000000d900000000",
            INIT_0E => X"000000db00000000000000db00000000000000dd00000000000000dd00000000",
            INIT_0F => X"000000bd00000000000000e300000000000000db00000000000000da00000000",
            INIT_10 => X"000000e400000000000000d900000000000000e800000000000000bd00000000",
            INIT_11 => X"000000dc00000000000000e200000000000000e100000000000000e300000000",
            INIT_12 => X"00000050000000000000004a000000000000009000000000000000dd00000000",
            INIT_13 => X"0000004c000000000000004e000000000000004c000000000000004a00000000",
            INIT_14 => X"000000a100000000000000810000000000000064000000000000005300000000",
            INIT_15 => X"000000e200000000000000e100000000000000c900000000000000b000000000",
            INIT_16 => X"000000d700000000000000d900000000000000dc00000000000000df00000000",
            INIT_17 => X"000000bb00000000000000e100000000000000d900000000000000d700000000",
            INIT_18 => X"000000e100000000000000d700000000000000e800000000000000bb00000000",
            INIT_19 => X"000000e200000000000000e300000000000000e100000000000000e000000000",
            INIT_1A => X"000000380000000000000032000000000000007700000000000000d500000000",
            INIT_1B => X"00000052000000000000004d0000000000000045000000000000003b00000000",
            INIT_1C => X"0000003f00000000000000420000000000000048000000000000005000000000",
            INIT_1D => X"000000a20000000000000085000000000000005b000000000000004100000000",
            INIT_1E => X"000000df00000000000000da00000000000000cc00000000000000b800000000",
            INIT_1F => X"000000bc00000000000000e300000000000000dd00000000000000dd00000000",
            INIT_20 => X"000000df00000000000000de00000000000000e700000000000000b700000000",
            INIT_21 => X"000000e100000000000000e400000000000000e600000000000000df00000000",
            INIT_22 => X"00000027000000000000003c000000000000006200000000000000a200000000",
            INIT_23 => X"0000004e00000000000000440000000000000043000000000000003500000000",
            INIT_24 => X"0000004800000000000000530000000000000052000000000000005100000000",
            INIT_25 => X"00000043000000000000003f0000000000000031000000000000003900000000",
            INIT_26 => X"000000a8000000000000008b000000000000006d000000000000004b00000000",
            INIT_27 => X"000000c300000000000000df00000000000000d700000000000000c600000000",
            INIT_28 => X"000000de00000000000000e200000000000000e200000000000000b000000000",
            INIT_29 => X"000000d400000000000000e200000000000000e200000000000000de00000000",
            INIT_2A => X"0000006a0000000000000096000000000000008b000000000000009b00000000",
            INIT_2B => X"0000005e00000000000000330000000000000039000000000000003500000000",
            INIT_2C => X"00000049000000000000008200000000000000a1000000000000009a00000000",
            INIT_2D => X"00000043000000000000005a0000000000000072000000000000006300000000",
            INIT_2E => X"000000a900000000000000ab0000000000000086000000000000004500000000",
            INIT_2F => X"000000be00000000000000d000000000000000c500000000000000b700000000",
            INIT_30 => X"000000df00000000000000e100000000000000e100000000000000af00000000",
            INIT_31 => X"000000de00000000000000de00000000000000de00000000000000df00000000",
            INIT_32 => X"000000cc00000000000000e400000000000000e000000000000000de00000000",
            INIT_33 => X"000000b300000000000000a0000000000000009f000000000000009f00000000",
            INIT_34 => X"000000a900000000000000cf00000000000000dc00000000000000d600000000",
            INIT_35 => X"000000ad00000000000000c000000000000000c100000000000000b200000000",
            INIT_36 => X"000000d600000000000000d200000000000000c300000000000000ab00000000",
            INIT_37 => X"000000bd00000000000000d200000000000000d100000000000000d800000000",
            INIT_38 => X"000000d100000000000000d700000000000000d400000000000000a600000000",
            INIT_39 => X"000000c700000000000000c900000000000000cc00000000000000ce00000000",
            INIT_3A => X"000000c200000000000000c500000000000000c300000000000000c700000000",
            INIT_3B => X"000000c400000000000000c200000000000000c100000000000000c000000000",
            INIT_3C => X"000000ca00000000000000c400000000000000c200000000000000c400000000",
            INIT_3D => X"000000cd00000000000000c800000000000000c400000000000000c800000000",
            INIT_3E => X"000000bf00000000000000c000000000000000c500000000000000ce00000000",
            INIT_3F => X"000000b500000000000000c900000000000000c500000000000000c500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007800000000000000820000000000000078000000000000006500000000",
            INIT_41 => X"0000006a000000000000006b0000000000000070000000000000007600000000",
            INIT_42 => X"0000006300000000000000660000000000000062000000000000006500000000",
            INIT_43 => X"00000080000000000000006c0000000000000065000000000000006200000000",
            INIT_44 => X"0000009300000000000000920000000000000092000000000000009000000000",
            INIT_45 => X"0000009e00000000000000980000000000000096000000000000009400000000",
            INIT_46 => X"000000a800000000000000a800000000000000a600000000000000a400000000",
            INIT_47 => X"0000009200000000000000a700000000000000a500000000000000a800000000",
            INIT_48 => X"0000008600000000000000860000000000000082000000000000006f00000000",
            INIT_49 => X"0000008800000000000000890000000000000088000000000000008a00000000",
            INIT_4A => X"0000007e00000000000000830000000000000086000000000000008400000000",
            INIT_4B => X"0000008300000000000000830000000000000080000000000000007f00000000",
            INIT_4C => X"00000081000000000000007f0000000000000086000000000000008a00000000",
            INIT_4D => X"0000007e000000000000007c0000000000000080000000000000008100000000",
            INIT_4E => X"0000008400000000000000840000000000000082000000000000008100000000",
            INIT_4F => X"0000006000000000000000730000000000000073000000000000007700000000",
            INIT_50 => X"0000007800000000000000780000000000000071000000000000006800000000",
            INIT_51 => X"00000064000000000000006c0000000000000076000000000000007a00000000",
            INIT_52 => X"000000590000000000000055000000000000005b000000000000006000000000",
            INIT_53 => X"0000005600000000000000570000000000000055000000000000005800000000",
            INIT_54 => X"000000430000000000000046000000000000004f000000000000005600000000",
            INIT_55 => X"0000003c000000000000003f0000000000000041000000000000004200000000",
            INIT_56 => X"0000003b000000000000003c000000000000003c000000000000003b00000000",
            INIT_57 => X"0000004b000000000000003f0000000000000032000000000000003600000000",
            INIT_58 => X"00000039000000000000003d0000000000000037000000000000003d00000000",
            INIT_59 => X"00000036000000000000003b000000000000003f000000000000003a00000000",
            INIT_5A => X"0000002f000000000000002f0000000000000033000000000000003800000000",
            INIT_5B => X"0000003200000000000000310000000000000032000000000000003000000000",
            INIT_5C => X"0000002f00000000000000350000000000000037000000000000003300000000",
            INIT_5D => X"000000370000000000000032000000000000002e000000000000002d00000000",
            INIT_5E => X"0000003400000000000000340000000000000034000000000000003600000000",
            INIT_5F => X"000000680000000000000068000000000000003a000000000000003000000000",
            INIT_60 => X"0000003c0000000000000041000000000000003d000000000000004400000000",
            INIT_61 => X"000000390000000000000037000000000000003d000000000000003e00000000",
            INIT_62 => X"0000003a00000000000000370000000000000038000000000000003d00000000",
            INIT_63 => X"0000003600000000000000380000000000000038000000000000003b00000000",
            INIT_64 => X"000000340000000000000037000000000000003b000000000000003900000000",
            INIT_65 => X"0000003400000000000000340000000000000033000000000000003300000000",
            INIT_66 => X"0000003900000000000000370000000000000035000000000000003300000000",
            INIT_67 => X"0000004b00000000000000780000000000000071000000000000004b00000000",
            INIT_68 => X"00000035000000000000003b0000000000000034000000000000003e00000000",
            INIT_69 => X"0000003600000000000000340000000000000039000000000000003900000000",
            INIT_6A => X"0000003200000000000000300000000000000032000000000000003600000000",
            INIT_6B => X"0000003500000000000000340000000000000038000000000000003900000000",
            INIT_6C => X"0000003300000000000000340000000000000036000000000000003900000000",
            INIT_6D => X"0000003000000000000000350000000000000037000000000000003600000000",
            INIT_6E => X"0000005f000000000000003d0000000000000034000000000000003200000000",
            INIT_6F => X"00000032000000000000003e0000000000000065000000000000007c00000000",
            INIT_70 => X"00000037000000000000003a0000000000000035000000000000003e00000000",
            INIT_71 => X"0000003c000000000000003c000000000000003d000000000000003b00000000",
            INIT_72 => X"0000004b000000000000003a0000000000000037000000000000003900000000",
            INIT_73 => X"0000004500000000000000440000000000000048000000000000004c00000000",
            INIT_74 => X"00000049000000000000004b000000000000004a000000000000004b00000000",
            INIT_75 => X"000000350000000000000037000000000000003a000000000000004600000000",
            INIT_76 => X"0000007f000000000000006b0000000000000045000000000000003300000000",
            INIT_77 => X"000000330000000000000036000000000000003a000000000000005b00000000",
            INIT_78 => X"0000002e00000000000000330000000000000033000000000000004000000000",
            INIT_79 => X"0000003500000000000000390000000000000038000000000000003300000000",
            INIT_7A => X"0000003e00000000000000320000000000000033000000000000003400000000",
            INIT_7B => X"00000039000000000000003c000000000000003e000000000000004000000000",
            INIT_7C => X"000000400000000000000040000000000000003e000000000000003c00000000",
            INIT_7D => X"0000003700000000000000340000000000000035000000000000004000000000",
            INIT_7E => X"0000004800000000000000690000000000000067000000000000004600000000",
            INIT_7F => X"0000003200000000000000340000000000000032000000000000003500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE23;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE24 : if BRAM_NAME = "sampleifmap_layersamples_instance24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001e00000000000000300000000000000046000000000000004100000000",
            INIT_01 => X"0000002d000000000000002c0000000000000028000000000000001700000000",
            INIT_02 => X"0000000f000000000000000a0000000000000028000000000000002d00000000",
            INIT_03 => X"0000003000000000000000330000000000000035000000000000002c00000000",
            INIT_04 => X"0000005b000000000000005d000000000000005a000000000000004100000000",
            INIT_05 => X"00000037000000000000003c0000000000000051000000000000005f00000000",
            INIT_06 => X"000000440000000000000029000000000000006f000000000000007000000000",
            INIT_07 => X"0000004300000000000000360000000000000033000000000000004d00000000",
            INIT_08 => X"0000001e000000000000003c000000000000004f000000000000004500000000",
            INIT_09 => X"0000003100000000000000310000000000000041000000000000002900000000",
            INIT_0A => X"0000001900000000000000070000000000000023000000000000003100000000",
            INIT_0B => X"0000003100000000000000370000000000000045000000000000004100000000",
            INIT_0C => X"0000005000000000000000530000000000000055000000000000004d00000000",
            INIT_0D => X"0000003b00000000000000370000000000000051000000000000005700000000",
            INIT_0E => X"0000002f000000000000001f0000000000000079000000000000008300000000",
            INIT_0F => X"0000003d00000000000000410000000000000036000000000000003800000000",
            INIT_10 => X"0000002900000000000000480000000000000054000000000000004900000000",
            INIT_11 => X"000000360000000000000032000000000000004a000000000000004000000000",
            INIT_12 => X"00000024000000000000000b0000000000000020000000000000003600000000",
            INIT_13 => X"00000027000000000000002f0000000000000043000000000000003c00000000",
            INIT_14 => X"0000003e000000000000003b000000000000004d000000000000004b00000000",
            INIT_15 => X"0000003f00000000000000300000000000000055000000000000005300000000",
            INIT_16 => X"0000002900000000000000170000000000000080000000000000008b00000000",
            INIT_17 => X"000000300000000000000049000000000000004e000000000000004600000000",
            INIT_18 => X"000000360000000000000050000000000000004b000000000000005800000000",
            INIT_19 => X"0000003f00000000000000370000000000000044000000000000005000000000",
            INIT_1A => X"000000250000000000000011000000000000001c000000000000003a00000000",
            INIT_1B => X"0000002700000000000000280000000000000033000000000000002b00000000",
            INIT_1C => X"00000046000000000000004b0000000000000062000000000000005500000000",
            INIT_1D => X"0000004400000000000000320000000000000054000000000000005600000000",
            INIT_1E => X"0000004b000000000000002f0000000000000089000000000000008e00000000",
            INIT_1F => X"000000260000000000000041000000000000005d000000000000006400000000",
            INIT_20 => X"00000042000000000000006f0000000000000059000000000000005f00000000",
            INIT_21 => X"00000044000000000000003d000000000000003d000000000000005100000000",
            INIT_22 => X"00000016000000000000000f0000000000000016000000000000003e00000000",
            INIT_23 => X"0000003f00000000000000330000000000000023000000000000001f00000000",
            INIT_24 => X"000000470000000000000048000000000000004b000000000000004800000000",
            INIT_25 => X"0000004e00000000000000330000000000000053000000000000004d00000000",
            INIT_26 => X"000000570000000000000057000000000000009c000000000000009500000000",
            INIT_27 => X"00000058000000000000004b000000000000005f000000000000006300000000",
            INIT_28 => X"0000004d00000000000000520000000000000053000000000000005200000000",
            INIT_29 => X"000000390000000000000040000000000000003a000000000000004700000000",
            INIT_2A => X"0000001c00000000000000110000000000000014000000000000003b00000000",
            INIT_2B => X"000000470000000000000047000000000000003d000000000000003200000000",
            INIT_2C => X"0000003800000000000000440000000000000043000000000000004500000000",
            INIT_2D => X"0000004e00000000000000460000000000000053000000000000002900000000",
            INIT_2E => X"00000059000000000000006200000000000000ac000000000000009c00000000",
            INIT_2F => X"000000630000000000000070000000000000006f000000000000005e00000000",
            INIT_30 => X"0000003b00000000000000200000000000000040000000000000004500000000",
            INIT_31 => X"000000310000000000000049000000000000004a000000000000004800000000",
            INIT_32 => X"0000003e000000000000001d0000000000000012000000000000003100000000",
            INIT_33 => X"0000003f00000000000000560000000000000055000000000000005200000000",
            INIT_34 => X"0000002b000000000000005f0000000000000034000000000000002200000000",
            INIT_35 => X"0000004e0000000000000055000000000000005e000000000000001900000000",
            INIT_36 => X"0000006b000000000000006d00000000000000b400000000000000a600000000",
            INIT_37 => X"0000002f00000000000000560000000000000083000000000000006c00000000",
            INIT_38 => X"0000004600000000000000190000000000000035000000000000003b00000000",
            INIT_39 => X"0000003d0000000000000050000000000000004e000000000000005100000000",
            INIT_3A => X"0000005e0000000000000035000000000000000a000000000000002800000000",
            INIT_3B => X"00000019000000000000004b0000000000000058000000000000005700000000",
            INIT_3C => X"00000039000000000000005c000000000000002d000000000000000d00000000",
            INIT_3D => X"0000006200000000000000590000000000000065000000000000003200000000",
            INIT_3E => X"0000007c000000000000007800000000000000b3000000000000009000000000",
            INIT_3F => X"0000001800000000000000340000000000000080000000000000007c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000660000000000000031000000000000002f000000000000004400000000",
            INIT_41 => X"0000004f000000000000003f0000000000000059000000000000007700000000",
            INIT_42 => X"0000006000000000000000510000000000000022000000000000004200000000",
            INIT_43 => X"0000000e0000000000000029000000000000005a000000000000005900000000",
            INIT_44 => X"000000470000000000000043000000000000005c000000000000003400000000",
            INIT_45 => X"00000073000000000000006e0000000000000071000000000000006f00000000",
            INIT_46 => X"0000007f0000000000000079000000000000009c000000000000008800000000",
            INIT_47 => X"00000016000000000000001f0000000000000073000000000000007c00000000",
            INIT_48 => X"0000007200000000000000370000000000000035000000000000004d00000000",
            INIT_49 => X"000000370000000000000041000000000000007b000000000000008000000000",
            INIT_4A => X"0000006e000000000000006f0000000000000052000000000000004f00000000",
            INIT_4B => X"0000002500000000000000140000000000000045000000000000006a00000000",
            INIT_4C => X"0000006100000000000000530000000000000069000000000000005c00000000",
            INIT_4D => X"0000005c00000000000000730000000000000078000000000000007600000000",
            INIT_4E => X"0000007f000000000000007d0000000000000093000000000000009000000000",
            INIT_4F => X"00000017000000000000000e000000000000005f000000000000007700000000",
            INIT_50 => X"000000700000000000000036000000000000003a000000000000005500000000",
            INIT_51 => X"0000003100000000000000640000000000000084000000000000008100000000",
            INIT_52 => X"0000006d00000000000000680000000000000054000000000000002700000000",
            INIT_53 => X"00000053000000000000003f000000000000005d000000000000007d00000000",
            INIT_54 => X"0000006e0000000000000068000000000000005e000000000000006100000000",
            INIT_55 => X"000000390000000000000055000000000000007f000000000000006d00000000",
            INIT_56 => X"0000007c000000000000007b0000000000000096000000000000009800000000",
            INIT_57 => X"00000015000000000000000c000000000000005d000000000000007200000000",
            INIT_58 => X"0000006b00000000000000320000000000000035000000000000006c00000000",
            INIT_59 => X"0000004b00000000000000800000000000000083000000000000007e00000000",
            INIT_5A => X"0000006b0000000000000055000000000000005b000000000000003300000000",
            INIT_5B => X"000000930000000000000081000000000000006e000000000000008a00000000",
            INIT_5C => X"0000007700000000000000710000000000000078000000000000008400000000",
            INIT_5D => X"0000005d000000000000005a0000000000000073000000000000007500000000",
            INIT_5E => X"0000007d0000000000000071000000000000008d00000000000000a000000000",
            INIT_5F => X"00000009000000000000000e0000000000000065000000000000007900000000",
            INIT_60 => X"0000005c000000000000002b000000000000002a000000000000006000000000",
            INIT_61 => X"0000007700000000000000820000000000000080000000000000006a00000000",
            INIT_62 => X"000000890000000000000072000000000000007b000000000000007800000000",
            INIT_63 => X"000000840000000000000069000000000000006e000000000000009400000000",
            INIT_64 => X"0000008600000000000000800000000000000087000000000000009200000000",
            INIT_65 => X"00000077000000000000007e0000000000000078000000000000008c00000000",
            INIT_66 => X"0000006a00000000000000630000000000000091000000000000009800000000",
            INIT_67 => X"0000002800000000000000120000000000000063000000000000008200000000",
            INIT_68 => X"00000059000000000000003b0000000000000042000000000000006100000000",
            INIT_69 => X"000000880000000000000085000000000000006f000000000000006400000000",
            INIT_6A => X"000000910000000000000096000000000000008c000000000000009300000000",
            INIT_6B => X"0000007f00000000000000830000000000000088000000000000008e00000000",
            INIT_6C => X"000000930000000000000088000000000000007b000000000000007d00000000",
            INIT_6D => X"00000088000000000000009c000000000000008e000000000000009700000000",
            INIT_6E => X"00000070000000000000006d0000000000000090000000000000009200000000",
            INIT_6F => X"000000530000000000000032000000000000005c000000000000008200000000",
            INIT_70 => X"0000005f000000000000004b0000000000000048000000000000006900000000",
            INIT_71 => X"000000850000000000000085000000000000005e000000000000006800000000",
            INIT_72 => X"0000008500000000000000800000000000000087000000000000008f00000000",
            INIT_73 => X"0000009800000000000000a00000000000000096000000000000009300000000",
            INIT_74 => X"0000008700000000000000840000000000000090000000000000009100000000",
            INIT_75 => X"000000a500000000000000a2000000000000008a000000000000008a00000000",
            INIT_76 => X"00000077000000000000007e000000000000007f00000000000000a300000000",
            INIT_77 => X"0000004d000000000000003b000000000000005f000000000000007600000000",
            INIT_78 => X"0000005b00000000000000440000000000000044000000000000005e00000000",
            INIT_79 => X"00000083000000000000007b0000000000000062000000000000006500000000",
            INIT_7A => X"0000004f000000000000008a00000000000000c1000000000000009300000000",
            INIT_7B => X"000000a200000000000000930000000000000093000000000000007c00000000",
            INIT_7C => X"00000090000000000000009800000000000000ab00000000000000b400000000",
            INIT_7D => X"000000b300000000000000940000000000000079000000000000009000000000",
            INIT_7E => X"0000007b000000000000008000000000000000a000000000000000b400000000",
            INIT_7F => X"00000054000000000000001a000000000000003f000000000000007000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE24;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE25 : if BRAM_NAME = "sampleifmap_layersamples_instance25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000059000000000000004a000000000000004f000000000000005800000000",
            INIT_01 => X"0000008100000000000000780000000000000078000000000000006e00000000",
            INIT_02 => X"0000005700000000000000c000000000000000b8000000000000007800000000",
            INIT_03 => X"000000a600000000000000a4000000000000009c000000000000007200000000",
            INIT_04 => X"000000b600000000000000b700000000000000a1000000000000009a00000000",
            INIT_05 => X"0000008f000000000000009400000000000000ad00000000000000bb00000000",
            INIT_06 => X"0000007c000000000000008e00000000000000c300000000000000b500000000",
            INIT_07 => X"000000760000000000000029000000000000002c000000000000006b00000000",
            INIT_08 => X"0000006000000000000000670000000000000059000000000000005b00000000",
            INIT_09 => X"0000006a000000000000006f0000000000000064000000000000007400000000",
            INIT_0A => X"000000a800000000000000bb0000000000000080000000000000007200000000",
            INIT_0B => X"000000ac00000000000000ac0000000000000099000000000000008c00000000",
            INIT_0C => X"000000a3000000000000009d00000000000000a400000000000000a700000000",
            INIT_0D => X"0000009c00000000000000ab00000000000000a500000000000000a100000000",
            INIT_0E => X"0000007200000000000000a7000000000000009100000000000000a100000000",
            INIT_0F => X"0000005e000000000000002a000000000000004a000000000000006a00000000",
            INIT_10 => X"0000007a00000000000000780000000000000061000000000000006500000000",
            INIT_11 => X"0000005b000000000000005f000000000000004e000000000000007200000000",
            INIT_12 => X"000000cc0000000000000081000000000000006e000000000000007300000000",
            INIT_13 => X"0000009900000000000000a0000000000000008900000000000000a700000000",
            INIT_14 => X"000000b200000000000000aa00000000000000ba00000000000000b300000000",
            INIT_15 => X"000000a500000000000000a2000000000000009c00000000000000b300000000",
            INIT_16 => X"000000480000000000000068000000000000008c000000000000009c00000000",
            INIT_17 => X"0000007200000000000000460000000000000059000000000000005400000000",
            INIT_18 => X"00000060000000000000007a000000000000006b000000000000006e00000000",
            INIT_19 => X"000000640000000000000048000000000000004c000000000000005a00000000",
            INIT_1A => X"0000008c0000000000000057000000000000007f000000000000006d00000000",
            INIT_1B => X"000000b400000000000000a6000000000000009f00000000000000bd00000000",
            INIT_1C => X"000000bc00000000000000be00000000000000ad00000000000000ae00000000",
            INIT_1D => X"000000a100000000000000a2000000000000009900000000000000a200000000",
            INIT_1E => X"0000004a000000000000004b0000000000000095000000000000009900000000",
            INIT_1F => X"0000008a0000000000000070000000000000003e000000000000004200000000",
            INIT_20 => X"0000004e0000000000000059000000000000006a000000000000007700000000",
            INIT_21 => X"00000067000000000000003c0000000000000047000000000000005900000000",
            INIT_22 => X"000000420000000000000072000000000000005f000000000000004b00000000",
            INIT_23 => X"000000be00000000000000ae00000000000000b5000000000000007f00000000",
            INIT_24 => X"000000c100000000000000b800000000000000ab00000000000000ba00000000",
            INIT_25 => X"000000a500000000000000ab00000000000000a000000000000000a400000000",
            INIT_26 => X"0000005c0000000000000068000000000000008b000000000000009200000000",
            INIT_27 => X"000000730000000000000070000000000000005e000000000000004d00000000",
            INIT_28 => X"00000067000000000000003a000000000000005e000000000000007e00000000",
            INIT_29 => X"0000005f0000000000000048000000000000004c000000000000006a00000000",
            INIT_2A => X"0000006300000000000000780000000000000041000000000000005e00000000",
            INIT_2B => X"000000bc00000000000000c400000000000000a1000000000000005b00000000",
            INIT_2C => X"000000a700000000000000a700000000000000c100000000000000b600000000",
            INIT_2D => X"000000a1000000000000009a00000000000000a000000000000000aa00000000",
            INIT_2E => X"00000051000000000000006e000000000000008a000000000000009100000000",
            INIT_2F => X"00000064000000000000006d0000000000000088000000000000006900000000",
            INIT_30 => X"0000006800000000000000460000000000000052000000000000006f00000000",
            INIT_31 => X"000000540000000000000045000000000000005e000000000000007100000000",
            INIT_32 => X"0000007d0000000000000055000000000000006d000000000000007400000000",
            INIT_33 => X"000000c800000000000000ba000000000000009b000000000000007f00000000",
            INIT_34 => X"0000009d00000000000000b100000000000000bb00000000000000bb00000000",
            INIT_35 => X"000000a600000000000000a400000000000000a2000000000000009400000000",
            INIT_36 => X"000000610000000000000079000000000000009500000000000000a200000000",
            INIT_37 => X"0000006100000000000000610000000000000073000000000000007800000000",
            INIT_38 => X"000000b4000000000000008c000000000000005c000000000000006500000000",
            INIT_39 => X"0000004c0000000000000055000000000000007b000000000000009700000000",
            INIT_3A => X"00000054000000000000005a000000000000007c000000000000006700000000",
            INIT_3B => X"000000c800000000000000ad00000000000000af000000000000009200000000",
            INIT_3C => X"0000009f00000000000000ad00000000000000ad00000000000000bc00000000",
            INIT_3D => X"000000ad00000000000000a300000000000000ac000000000000009f00000000",
            INIT_3E => X"000000830000000000000083000000000000008b00000000000000a400000000",
            INIT_3F => X"000000600000000000000064000000000000005f000000000000007000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d100000000000000c00000000000000090000000000000007700000000",
            INIT_41 => X"0000006c000000000000007f000000000000009d00000000000000c200000000",
            INIT_42 => X"0000006f000000000000006a000000000000005e000000000000006a00000000",
            INIT_43 => X"000000c500000000000000b000000000000000af000000000000007c00000000",
            INIT_44 => X"000000a500000000000000b000000000000000aa00000000000000b800000000",
            INIT_45 => X"000000a300000000000000af00000000000000c5000000000000009c00000000",
            INIT_46 => X"00000065000000000000007a0000000000000083000000000000009300000000",
            INIT_47 => X"00000066000000000000006b0000000000000060000000000000006400000000",
            INIT_48 => X"000000a9000000000000008a0000000000000074000000000000006e00000000",
            INIT_49 => X"0000008800000000000000a000000000000000c400000000000000c500000000",
            INIT_4A => X"0000008a000000000000005c0000000000000063000000000000008100000000",
            INIT_4B => X"000000a900000000000000b4000000000000009f000000000000009200000000",
            INIT_4C => X"000000b200000000000000af000000000000008d000000000000008e00000000",
            INIT_4D => X"0000009700000000000000b300000000000000bc00000000000000a600000000",
            INIT_4E => X"0000003a0000000000000070000000000000009a000000000000008f00000000",
            INIT_4F => X"0000004900000000000000660000000000000065000000000000005b00000000",
            INIT_50 => X"0000006b000000000000004a0000000000000057000000000000005b00000000",
            INIT_51 => X"000000a300000000000000bf00000000000000b900000000000000a500000000",
            INIT_52 => X"00000066000000000000006a0000000000000080000000000000008600000000",
            INIT_53 => X"0000007400000000000000920000000000000084000000000000007600000000",
            INIT_54 => X"000000b600000000000000a10000000000000063000000000000004d00000000",
            INIT_55 => X"000000a700000000000000ad000000000000009f00000000000000b700000000",
            INIT_56 => X"0000002b000000000000005e0000000000000087000000000000009c00000000",
            INIT_57 => X"0000004d0000000000000044000000000000005c000000000000005b00000000",
            INIT_58 => X"0000002c0000000000000032000000000000005f000000000000005100000000",
            INIT_59 => X"000000bb00000000000000a60000000000000094000000000000005f00000000",
            INIT_5A => X"00000072000000000000007e000000000000009000000000000000ae00000000",
            INIT_5B => X"0000006b00000000000000770000000000000072000000000000006800000000",
            INIT_5C => X"000000b6000000000000009d0000000000000052000000000000005100000000",
            INIT_5D => X"0000009600000000000000a900000000000000b200000000000000a900000000",
            INIT_5E => X"0000003f000000000000002c000000000000006c000000000000009800000000",
            INIT_5F => X"0000005600000000000000500000000000000045000000000000006100000000",
            INIT_60 => X"000000150000000000000034000000000000005f000000000000005a00000000",
            INIT_61 => X"000000b00000000000000092000000000000006d000000000000001c00000000",
            INIT_62 => X"0000007f000000000000008e00000000000000b500000000000000ca00000000",
            INIT_63 => X"0000008200000000000000720000000000000077000000000000007800000000",
            INIT_64 => X"000000a900000000000000900000000000000076000000000000008100000000",
            INIT_65 => X"0000009800000000000000b400000000000000ad000000000000009f00000000",
            INIT_66 => X"00000055000000000000002c0000000000000044000000000000007700000000",
            INIT_67 => X"0000006a00000000000000a70000000000000072000000000000003300000000",
            INIT_68 => X"000000340000000000000039000000000000005b000000000000005f00000000",
            INIT_69 => X"0000009c00000000000000770000000000000031000000000000001800000000",
            INIT_6A => X"0000009b00000000000000ba00000000000000cb00000000000000bb00000000",
            INIT_6B => X"0000007500000000000000740000000000000085000000000000008d00000000",
            INIT_6C => X"00000099000000000000008b0000000000000077000000000000006d00000000",
            INIT_6D => X"0000007d000000000000009c00000000000000a7000000000000009f00000000",
            INIT_6E => X"0000004000000000000000440000000000000041000000000000006500000000",
            INIT_6F => X"0000007a00000000000000aa0000000000000090000000000000003700000000",
            INIT_70 => X"000000490000000000000020000000000000004b000000000000005e00000000",
            INIT_71 => X"0000007300000000000000360000000000000021000000000000002e00000000",
            INIT_72 => X"000000c200000000000000c300000000000000b0000000000000009600000000",
            INIT_73 => X"000000920000000000000088000000000000009b00000000000000b100000000",
            INIT_74 => X"00000077000000000000005e0000000000000065000000000000008b00000000",
            INIT_75 => X"000000690000000000000060000000000000005f000000000000006500000000",
            INIT_76 => X"0000006d000000000000006b0000000000000076000000000000008300000000",
            INIT_77 => X"0000006a000000000000009a000000000000008f000000000000008000000000",
            INIT_78 => X"0000004c00000000000000180000000000000023000000000000004e00000000",
            INIT_79 => X"0000003b000000000000001b0000000000000028000000000000004100000000",
            INIT_7A => X"000000b000000000000000960000000000000088000000000000007800000000",
            INIT_7B => X"000000ba00000000000000a500000000000000b700000000000000c000000000",
            INIT_7C => X"00000056000000000000006b00000000000000aa00000000000000cf00000000",
            INIT_7D => X"0000008c00000000000000700000000000000055000000000000004200000000",
            INIT_7E => X"000000890000000000000089000000000000009500000000000000a900000000",
            INIT_7F => X"00000080000000000000009a000000000000008f000000000000009600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE25;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE26 : if BRAM_NAME = "sampleifmap_layersamples_instance26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002e00000000000000400000000000000051000000000000004400000000",
            INIT_01 => X"00000050000000000000004b0000000000000039000000000000002100000000",
            INIT_02 => X"0000002200000000000000140000000000000046000000000000005300000000",
            INIT_03 => X"000000420000000000000046000000000000004b000000000000004700000000",
            INIT_04 => X"00000079000000000000007c0000000000000078000000000000005700000000",
            INIT_05 => X"000000520000000000000054000000000000006c000000000000007e00000000",
            INIT_06 => X"0000005b000000000000003b0000000000000081000000000000008800000000",
            INIT_07 => X"00000057000000000000004c0000000000000043000000000000006000000000",
            INIT_08 => X"0000002f000000000000004a0000000000000066000000000000005000000000",
            INIT_09 => X"000000540000000000000054000000000000005c000000000000003800000000",
            INIT_0A => X"000000300000000000000012000000000000003e000000000000005800000000",
            INIT_0B => X"00000049000000000000004d000000000000005c000000000000005d00000000",
            INIT_0C => X"0000006a000000000000006f0000000000000075000000000000006b00000000",
            INIT_0D => X"00000053000000000000004d000000000000006c000000000000007500000000",
            INIT_0E => X"00000041000000000000002d000000000000008b000000000000009700000000",
            INIT_0F => X"00000051000000000000005a0000000000000042000000000000004700000000",
            INIT_10 => X"000000380000000000000058000000000000006d000000000000005f00000000",
            INIT_11 => X"0000005a00000000000000560000000000000069000000000000005400000000",
            INIT_12 => X"0000003c00000000000000140000000000000035000000000000005c00000000",
            INIT_13 => X"0000003c00000000000000420000000000000058000000000000005900000000",
            INIT_14 => X"00000054000000000000004e0000000000000066000000000000006700000000",
            INIT_15 => X"0000005600000000000000420000000000000072000000000000007200000000",
            INIT_16 => X"000000370000000000000023000000000000008f000000000000009e00000000",
            INIT_17 => X"0000003b00000000000000620000000000000062000000000000005400000000",
            INIT_18 => X"0000004900000000000000640000000000000064000000000000007400000000",
            INIT_19 => X"0000006000000000000000580000000000000066000000000000006d00000000",
            INIT_1A => X"00000038000000000000001a000000000000002d000000000000005e00000000",
            INIT_1B => X"0000003700000000000000360000000000000043000000000000004100000000",
            INIT_1C => X"0000006200000000000000610000000000000075000000000000006a00000000",
            INIT_1D => X"0000005b00000000000000450000000000000072000000000000007600000000",
            INIT_1E => X"0000005d0000000000000040000000000000009600000000000000a000000000",
            INIT_1F => X"00000032000000000000005e000000000000007e000000000000007800000000",
            INIT_20 => X"0000005d00000000000000800000000000000068000000000000007800000000",
            INIT_21 => X"0000005e000000000000005a000000000000005e000000000000007200000000",
            INIT_22 => X"00000024000000000000001a0000000000000027000000000000005d00000000",
            INIT_23 => X"0000005600000000000000490000000000000037000000000000002f00000000",
            INIT_24 => X"00000065000000000000006b0000000000000071000000000000006900000000",
            INIT_25 => X"00000067000000000000004a000000000000006d000000000000006700000000",
            INIT_26 => X"00000074000000000000007000000000000000ac00000000000000a200000000",
            INIT_27 => X"0000006c00000000000000670000000000000084000000000000008100000000",
            INIT_28 => X"0000006200000000000000620000000000000066000000000000006900000000",
            INIT_29 => X"0000004e000000000000005b0000000000000059000000000000005f00000000",
            INIT_2A => X"0000002b000000000000001b0000000000000023000000000000005800000000",
            INIT_2B => X"0000006c000000000000006a000000000000005d000000000000004d00000000",
            INIT_2C => X"0000004e00000000000000640000000000000065000000000000006700000000",
            INIT_2D => X"000000660000000000000062000000000000006e000000000000003900000000",
            INIT_2E => X"0000007f000000000000008200000000000000ba00000000000000a700000000",
            INIT_2F => X"0000007800000000000000840000000000000090000000000000008100000000",
            INIT_30 => X"0000004f00000000000000300000000000000060000000000000005e00000000",
            INIT_31 => X"0000003f000000000000005d0000000000000064000000000000005a00000000",
            INIT_32 => X"0000005a0000000000000026000000000000001d000000000000004a00000000",
            INIT_33 => X"0000006300000000000000820000000000000081000000000000007e00000000",
            INIT_34 => X"0000003900000000000000730000000000000047000000000000003a00000000",
            INIT_35 => X"0000006a0000000000000071000000000000007b000000000000002500000000",
            INIT_36 => X"0000008c000000000000008d00000000000000c100000000000000b700000000",
            INIT_37 => X"0000003b000000000000006500000000000000a0000000000000008900000000",
            INIT_38 => X"00000069000000000000002f0000000000000054000000000000005600000000",
            INIT_39 => X"00000047000000000000005e0000000000000061000000000000006700000000",
            INIT_3A => X"0000008b00000000000000490000000000000014000000000000003800000000",
            INIT_3B => X"000000290000000000000072000000000000008c000000000000008a00000000",
            INIT_3C => X"0000004f00000000000000730000000000000041000000000000001a00000000",
            INIT_3D => X"0000008c0000000000000078000000000000007d000000000000003b00000000",
            INIT_3E => X"00000094000000000000009600000000000000c300000000000000b000000000",
            INIT_3F => X"00000018000000000000003f000000000000009b000000000000009000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008c000000000000004a000000000000004e000000000000006200000000",
            INIT_41 => X"0000005c00000000000000500000000000000072000000000000009500000000",
            INIT_42 => X"000000900000000000000071000000000000002c000000000000004700000000",
            INIT_43 => X"00000017000000000000003f0000000000000086000000000000008800000000",
            INIT_44 => X"00000056000000000000005e000000000000007c000000000000004500000000",
            INIT_45 => X"000000a5000000000000009b000000000000008b000000000000007000000000",
            INIT_46 => X"00000096000000000000009600000000000000b100000000000000aa00000000",
            INIT_47 => X"000000160000000000000029000000000000008e000000000000009200000000",
            INIT_48 => X"00000094000000000000004e0000000000000051000000000000007400000000",
            INIT_49 => X"000000450000000000000054000000000000009b00000000000000a300000000",
            INIT_4A => X"0000008e0000000000000089000000000000005a000000000000005100000000",
            INIT_4B => X"000000380000000000000021000000000000005d000000000000008a00000000",
            INIT_4C => X"000000800000000000000073000000000000008f000000000000007c00000000",
            INIT_4D => X"00000081000000000000009c000000000000009c000000000000009700000000",
            INIT_4E => X"0000009a000000000000009800000000000000ad00000000000000a700000000",
            INIT_4F => X"0000001800000000000000160000000000000079000000000000009400000000",
            INIT_50 => X"000000910000000000000049000000000000004f000000000000007800000000",
            INIT_51 => X"00000041000000000000007f00000000000000a600000000000000a500000000",
            INIT_52 => X"0000007f000000000000008e0000000000000072000000000000003600000000",
            INIT_53 => X"0000006c0000000000000047000000000000005d000000000000007e00000000",
            INIT_54 => X"000000a100000000000000920000000000000085000000000000008700000000",
            INIT_55 => X"00000057000000000000007500000000000000a5000000000000009c00000000",
            INIT_56 => X"0000009c000000000000009700000000000000af00000000000000a900000000",
            INIT_57 => X"0000001700000000000000130000000000000074000000000000009100000000",
            INIT_58 => X"0000008a00000000000000420000000000000045000000000000007b00000000",
            INIT_59 => X"0000005f00000000000000a500000000000000a800000000000000a100000000",
            INIT_5A => X"00000070000000000000008a000000000000008c000000000000004b00000000",
            INIT_5B => X"000000a200000000000000880000000000000066000000000000006d00000000",
            INIT_5C => X"000000870000000000000097000000000000009a000000000000009900000000",
            INIT_5D => X"0000008800000000000000760000000000000085000000000000007c00000000",
            INIT_5E => X"0000009d000000000000009200000000000000aa00000000000000bd00000000",
            INIT_5F => X"0000000b00000000000000140000000000000077000000000000009400000000",
            INIT_60 => X"00000079000000000000003c0000000000000039000000000000006a00000000",
            INIT_61 => X"0000009800000000000000ad00000000000000a4000000000000008700000000",
            INIT_62 => X"00000076000000000000007f0000000000000093000000000000009000000000",
            INIT_63 => X"0000008b0000000000000066000000000000005c000000000000007300000000",
            INIT_64 => X"000000740000000000000085000000000000008a000000000000008d00000000",
            INIT_65 => X"000000880000000000000077000000000000006b000000000000007800000000",
            INIT_66 => X"00000091000000000000008700000000000000ae00000000000000b000000000",
            INIT_67 => X"0000002b000000000000001a000000000000007200000000000000a100000000",
            INIT_68 => X"00000074000000000000004e0000000000000055000000000000007400000000",
            INIT_69 => X"000000ab00000000000000ac000000000000008c000000000000007f00000000",
            INIT_6A => X"000000780000000000000082000000000000007c000000000000009900000000",
            INIT_6B => X"0000006e00000000000000710000000000000076000000000000007700000000",
            INIT_6C => X"0000007d0000000000000077000000000000006c000000000000006900000000",
            INIT_6D => X"000000750000000000000081000000000000007a000000000000008300000000",
            INIT_6E => X"0000009a000000000000008d00000000000000a2000000000000009000000000",
            INIT_6F => X"0000005f0000000000000041000000000000007000000000000000a600000000",
            INIT_70 => X"0000007800000000000000630000000000000060000000000000008400000000",
            INIT_71 => X"000000a800000000000000a50000000000000072000000000000008200000000",
            INIT_72 => X"000000700000000000000068000000000000006b000000000000008b00000000",
            INIT_73 => X"00000084000000000000008e0000000000000081000000000000007c00000000",
            INIT_74 => X"0000006f000000000000006b0000000000000077000000000000007a00000000",
            INIT_75 => X"00000090000000000000008d0000000000000076000000000000007300000000",
            INIT_76 => X"0000009f0000000000000092000000000000007b000000000000008e00000000",
            INIT_77 => X"0000005e00000000000000480000000000000070000000000000009d00000000",
            INIT_78 => X"00000076000000000000005d000000000000005a000000000000007900000000",
            INIT_79 => X"000000a60000000000000097000000000000007c000000000000007f00000000",
            INIT_7A => X"00000045000000000000007900000000000000ab000000000000009900000000",
            INIT_7B => X"0000008b000000000000007b000000000000007c000000000000006b00000000",
            INIT_7C => X"0000007700000000000000800000000000000090000000000000009b00000000",
            INIT_7D => X"000000a700000000000000830000000000000067000000000000007a00000000",
            INIT_7E => X"000000a00000000000000080000000000000008c000000000000009f00000000",
            INIT_7F => X"000000680000000000000022000000000000004b000000000000009500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE26;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE27 : if BRAM_NAME = "sampleifmap_layersamples_instance27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007e00000000000000640000000000000064000000000000007000000000",
            INIT_01 => X"000000a300000000000000950000000000000098000000000000008d00000000",
            INIT_02 => X"0000004700000000000000a600000000000000a3000000000000008a00000000",
            INIT_03 => X"0000008d000000000000008b0000000000000085000000000000006400000000",
            INIT_04 => X"0000009e00000000000000a00000000000000088000000000000008100000000",
            INIT_05 => X"0000007e000000000000007d000000000000009700000000000000a300000000",
            INIT_06 => X"0000008f000000000000007a00000000000000b100000000000000a900000000",
            INIT_07 => X"0000008b0000000000000033000000000000003d000000000000008f00000000",
            INIT_08 => X"0000008100000000000000830000000000000070000000000000007000000000",
            INIT_09 => X"000000890000000000000090000000000000007c000000000000009300000000",
            INIT_0A => X"0000009900000000000000a80000000000000079000000000000008f00000000",
            INIT_0B => X"000000930000000000000092000000000000007f000000000000007a00000000",
            INIT_0C => X"0000008a0000000000000084000000000000008b000000000000008d00000000",
            INIT_0D => X"000000860000000000000099000000000000008f000000000000008600000000",
            INIT_0E => X"0000007a00000000000000920000000000000082000000000000009100000000",
            INIT_0F => X"0000006f000000000000003a0000000000000064000000000000008600000000",
            INIT_10 => X"0000008e00000000000000950000000000000076000000000000007900000000",
            INIT_11 => X"00000076000000000000007b0000000000000061000000000000008d00000000",
            INIT_12 => X"000000bb0000000000000079000000000000007e000000000000008f00000000",
            INIT_13 => X"000000820000000000000088000000000000006e000000000000009100000000",
            INIT_14 => X"0000009a000000000000009400000000000000a1000000000000009a00000000",
            INIT_15 => X"0000009100000000000000960000000000000086000000000000009700000000",
            INIT_16 => X"000000570000000000000061000000000000007b000000000000008600000000",
            INIT_17 => X"0000008600000000000000610000000000000077000000000000006700000000",
            INIT_18 => X"0000006f00000000000000970000000000000087000000000000008800000000",
            INIT_19 => X"0000007d000000000000005d0000000000000065000000000000007a00000000",
            INIT_1A => X"0000007d00000000000000600000000000000099000000000000008600000000",
            INIT_1B => X"000000a00000000000000092000000000000008800000000000000a900000000",
            INIT_1C => X"000000a700000000000000a60000000000000094000000000000009600000000",
            INIT_1D => X"0000009100000000000000900000000000000080000000000000008d00000000",
            INIT_1E => X"0000005e000000000000004b0000000000000082000000000000008400000000",
            INIT_1F => X"000000a900000000000000950000000000000057000000000000005300000000",
            INIT_20 => X"0000005e0000000000000070000000000000008c000000000000009400000000",
            INIT_21 => X"0000008200000000000000540000000000000068000000000000007900000000",
            INIT_22 => X"0000004a000000000000008d0000000000000074000000000000006600000000",
            INIT_23 => X"000000aa000000000000009b00000000000000a3000000000000007600000000",
            INIT_24 => X"000000a7000000000000009d000000000000009500000000000000a500000000",
            INIT_25 => X"0000009100000000000000930000000000000089000000000000009200000000",
            INIT_26 => X"00000071000000000000006d000000000000007c000000000000007f00000000",
            INIT_27 => X"000000a1000000000000009c0000000000000077000000000000006000000000",
            INIT_28 => X"0000007d00000000000000480000000000000077000000000000009800000000",
            INIT_29 => X"0000007900000000000000630000000000000065000000000000008100000000",
            INIT_2A => X"0000007d000000000000009a000000000000005b000000000000007800000000",
            INIT_2B => X"000000a900000000000000b50000000000000096000000000000005d00000000",
            INIT_2C => X"0000008f000000000000009100000000000000ad00000000000000a200000000",
            INIT_2D => X"0000008b00000000000000810000000000000087000000000000008f00000000",
            INIT_2E => X"0000006600000000000000750000000000000078000000000000007d00000000",
            INIT_2F => X"00000099000000000000009a00000000000000ab000000000000008100000000",
            INIT_30 => X"0000007b00000000000000520000000000000068000000000000008800000000",
            INIT_31 => X"0000007300000000000000620000000000000076000000000000008800000000",
            INIT_32 => X"000000940000000000000075000000000000008d000000000000009600000000",
            INIT_33 => X"000000b300000000000000ad0000000000000095000000000000008100000000",
            INIT_34 => X"0000008f000000000000009f00000000000000a800000000000000a500000000",
            INIT_35 => X"0000008d000000000000008c000000000000008b000000000000007e00000000",
            INIT_36 => X"0000006d000000000000007a0000000000000085000000000000008800000000",
            INIT_37 => X"00000095000000000000009600000000000000a4000000000000009800000000",
            INIT_38 => X"000000bf0000000000000096000000000000006f000000000000007d00000000",
            INIT_39 => X"0000006f0000000000000079000000000000009e00000000000000ac00000000",
            INIT_3A => X"0000006900000000000000730000000000000099000000000000009100000000",
            INIT_3B => X"000000ac000000000000009a00000000000000a1000000000000009400000000",
            INIT_3C => X"0000008d000000000000009c000000000000009b00000000000000a100000000",
            INIT_3D => X"0000008f00000000000000880000000000000093000000000000008900000000",
            INIT_3E => X"00000086000000000000007b000000000000008c000000000000008900000000",
            INIT_3F => X"00000095000000000000009e0000000000000095000000000000009c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000dc00000000000000c800000000000000a2000000000000009500000000",
            INIT_41 => X"0000009300000000000000aa00000000000000bd00000000000000d100000000",
            INIT_42 => X"00000088000000000000007d000000000000007a000000000000009100000000",
            INIT_43 => X"000000a40000000000000096000000000000009f000000000000008b00000000",
            INIT_44 => X"0000008e000000000000009f000000000000009b000000000000009b00000000",
            INIT_45 => X"00000088000000000000009300000000000000a9000000000000008500000000",
            INIT_46 => X"00000072000000000000006b000000000000007e000000000000007f00000000",
            INIT_47 => X"0000009c00000000000000a0000000000000008f000000000000009a00000000",
            INIT_48 => X"000000be000000000000009d0000000000000089000000000000008b00000000",
            INIT_49 => X"000000b000000000000000bf00000000000000d700000000000000d500000000",
            INIT_4A => X"000000a30000000000000075000000000000008400000000000000a900000000",
            INIT_4B => X"0000008f000000000000009a000000000000009700000000000000ad00000000",
            INIT_4C => X"0000009800000000000000990000000000000081000000000000007c00000000",
            INIT_4D => X"0000007c000000000000009500000000000000a3000000000000009100000000",
            INIT_4E => X"0000004a00000000000000600000000000000083000000000000007700000000",
            INIT_4F => X"0000007800000000000000970000000000000095000000000000009100000000",
            INIT_50 => X"000000860000000000000061000000000000006f000000000000007300000000",
            INIT_51 => X"000000c100000000000000d300000000000000cf00000000000000bf00000000",
            INIT_52 => X"0000007f000000000000009100000000000000ad00000000000000b100000000",
            INIT_53 => X"000000680000000000000086000000000000008f000000000000009000000000",
            INIT_54 => X"0000009b000000000000008b000000000000005c000000000000004900000000",
            INIT_55 => X"0000008e0000000000000094000000000000008a00000000000000a100000000",
            INIT_56 => X"0000003c00000000000000550000000000000075000000000000008300000000",
            INIT_57 => X"0000006d000000000000006f0000000000000091000000000000009200000000",
            INIT_58 => X"0000004000000000000000410000000000000072000000000000006a00000000",
            INIT_59 => X"000000d500000000000000c300000000000000b2000000000000007800000000",
            INIT_5A => X"0000009900000000000000ad00000000000000b900000000000000ca00000000",
            INIT_5B => X"0000007d000000000000008d0000000000000096000000000000008e00000000",
            INIT_5C => X"0000009a000000000000008e0000000000000060000000000000006c00000000",
            INIT_5D => X"0000007f000000000000009500000000000000a1000000000000009000000000",
            INIT_5E => X"0000006100000000000000310000000000000062000000000000008300000000",
            INIT_5F => X"000000750000000000000076000000000000006c000000000000009300000000",
            INIT_60 => X"00000026000000000000003e0000000000000070000000000000007400000000",
            INIT_61 => X"000000c700000000000000b40000000000000087000000000000002900000000",
            INIT_62 => X"000000b200000000000000b700000000000000cc00000000000000d400000000",
            INIT_63 => X"000000a1000000000000009e00000000000000a400000000000000ab00000000",
            INIT_64 => X"0000008d0000000000000087000000000000008b000000000000009d00000000",
            INIT_65 => X"0000007e000000000000009c0000000000000099000000000000008700000000",
            INIT_66 => X"0000007c000000000000003b0000000000000042000000000000006700000000",
            INIT_67 => X"0000008300000000000000c50000000000000088000000000000005400000000",
            INIT_68 => X"0000004e000000000000004f000000000000007b000000000000007f00000000",
            INIT_69 => X"000000bf00000000000000950000000000000042000000000000002500000000",
            INIT_6A => X"000000c200000000000000d600000000000000db00000000000000d000000000",
            INIT_6B => X"0000009f00000000000000a500000000000000b400000000000000b800000000",
            INIT_6C => X"00000083000000000000007b000000000000007d000000000000008700000000",
            INIT_6D => X"0000007200000000000000870000000000000093000000000000008a00000000",
            INIT_6E => X"0000005b0000000000000055000000000000004f000000000000006c00000000",
            INIT_6F => X"0000008f00000000000000c900000000000000ac000000000000004e00000000",
            INIT_70 => X"0000006b00000000000000340000000000000068000000000000007d00000000",
            INIT_71 => X"00000097000000000000004e0000000000000030000000000000004300000000",
            INIT_72 => X"000000da00000000000000d900000000000000cb00000000000000bd00000000",
            INIT_73 => X"000000b600000000000000b400000000000000c300000000000000cd00000000",
            INIT_74 => X"0000007a000000000000005e000000000000007400000000000000a500000000",
            INIT_75 => X"0000006f00000000000000590000000000000059000000000000006100000000",
            INIT_76 => X"000000860000000000000082000000000000008a000000000000009600000000",
            INIT_77 => X"0000008100000000000000bc00000000000000b5000000000000009f00000000",
            INIT_78 => X"0000007300000000000000280000000000000033000000000000006600000000",
            INIT_79 => X"0000004e0000000000000029000000000000003a000000000000006000000000",
            INIT_7A => X"000000cf00000000000000b900000000000000b500000000000000a000000000",
            INIT_7B => X"000000ce00000000000000c400000000000000d200000000000000da00000000",
            INIT_7C => X"00000071000000000000007c00000000000000b400000000000000d600000000",
            INIT_7D => X"000000a000000000000000840000000000000066000000000000005600000000",
            INIT_7E => X"000000a700000000000000a700000000000000a700000000000000ba00000000",
            INIT_7F => X"0000009c00000000000000b900000000000000b300000000000000b400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE27;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE28 : if BRAM_NAME = "sampleifmap_layersamples_instance28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001e000000000000002e0000000000000040000000000000003200000000",
            INIT_01 => X"0000003900000000000000370000000000000024000000000000001600000000",
            INIT_02 => X"00000012000000000000000c0000000000000036000000000000003b00000000",
            INIT_03 => X"000000320000000000000031000000000000002c000000000000002b00000000",
            INIT_04 => X"0000004d0000000000000051000000000000004d000000000000003a00000000",
            INIT_05 => X"000000390000000000000038000000000000004e000000000000005300000000",
            INIT_06 => X"0000003a000000000000001f000000000000005d000000000000006100000000",
            INIT_07 => X"0000004200000000000000350000000000000029000000000000004100000000",
            INIT_08 => X"0000001d00000000000000390000000000000051000000000000003a00000000",
            INIT_09 => X"0000003c000000000000003b000000000000003d000000000000002300000000",
            INIT_0A => X"0000001b0000000000000007000000000000002f000000000000004000000000",
            INIT_0B => X"0000002f000000000000003b000000000000003e000000000000003800000000",
            INIT_0C => X"00000044000000000000004a000000000000004a000000000000004400000000",
            INIT_0D => X"0000003c00000000000000330000000000000051000000000000004e00000000",
            INIT_0E => X"0000002700000000000000150000000000000060000000000000006f00000000",
            INIT_0F => X"000000420000000000000045000000000000002c000000000000002d00000000",
            INIT_10 => X"0000002300000000000000460000000000000057000000000000004800000000",
            INIT_11 => X"00000041000000000000003c0000000000000048000000000000003500000000",
            INIT_12 => X"0000002300000000000000070000000000000026000000000000004500000000",
            INIT_13 => X"0000002100000000000000300000000000000041000000000000003400000000",
            INIT_14 => X"0000003700000000000000320000000000000042000000000000004300000000",
            INIT_15 => X"0000003e000000000000002d0000000000000052000000000000004d00000000",
            INIT_16 => X"0000002600000000000000100000000000000063000000000000007400000000",
            INIT_17 => X"00000033000000000000004d000000000000004b000000000000003f00000000",
            INIT_18 => X"0000002f0000000000000050000000000000004c000000000000005e00000000",
            INIT_19 => X"0000004a00000000000000410000000000000048000000000000004700000000",
            INIT_1A => X"00000022000000000000000c000000000000001e000000000000004800000000",
            INIT_1B => X"0000001e00000000000000230000000000000034000000000000002800000000",
            INIT_1C => X"0000004500000000000000440000000000000057000000000000004b00000000",
            INIT_1D => X"00000043000000000000002e000000000000004d000000000000005100000000",
            INIT_1E => X"00000049000000000000002a000000000000006b000000000000007700000000",
            INIT_1F => X"0000002200000000000000440000000000000060000000000000005f00000000",
            INIT_20 => X"0000003c000000000000006a000000000000004f000000000000006100000000",
            INIT_21 => X"0000004c00000000000000480000000000000044000000000000004b00000000",
            INIT_22 => X"00000011000000000000000c0000000000000018000000000000004900000000",
            INIT_23 => X"0000003b00000000000000330000000000000025000000000000001c00000000",
            INIT_24 => X"00000047000000000000004b000000000000004f000000000000004800000000",
            INIT_25 => X"0000004d000000000000002d0000000000000049000000000000004700000000",
            INIT_26 => X"0000005500000000000000520000000000000081000000000000008000000000",
            INIT_27 => X"0000005000000000000000490000000000000061000000000000005e00000000",
            INIT_28 => X"00000043000000000000004b000000000000004d000000000000005200000000",
            INIT_29 => X"0000003d000000000000004d0000000000000045000000000000003d00000000",
            INIT_2A => X"00000016000000000000000d0000000000000013000000000000004300000000",
            INIT_2B => X"000000490000000000000047000000000000003b000000000000002c00000000",
            INIT_2C => X"0000003500000000000000490000000000000048000000000000004800000000",
            INIT_2D => X"0000004d000000000000003e0000000000000049000000000000002200000000",
            INIT_2E => X"0000005b00000000000000600000000000000093000000000000008800000000",
            INIT_2F => X"0000005c0000000000000068000000000000006e000000000000005c00000000",
            INIT_30 => X"0000003300000000000000190000000000000046000000000000004800000000",
            INIT_31 => X"00000032000000000000004f000000000000004f000000000000003e00000000",
            INIT_32 => X"000000360000000000000018000000000000000f000000000000003800000000",
            INIT_33 => X"0000003e000000000000004d000000000000004b000000000000004900000000",
            INIT_34 => X"0000002a00000000000000600000000000000033000000000000002200000000",
            INIT_35 => X"0000004a00000000000000480000000000000058000000000000001600000000",
            INIT_36 => X"0000006c000000000000006800000000000000a1000000000000009500000000",
            INIT_37 => X"0000002b00000000000000510000000000000083000000000000006b00000000",
            INIT_38 => X"000000460000000000000015000000000000003b000000000000003f00000000",
            INIT_39 => X"0000003a000000000000004b0000000000000048000000000000004d00000000",
            INIT_3A => X"00000051000000000000002f0000000000000008000000000000002900000000",
            INIT_3B => X"00000012000000000000003e000000000000004b000000000000004b00000000",
            INIT_3C => X"0000004000000000000000590000000000000027000000000000000600000000",
            INIT_3D => X"000000530000000000000048000000000000005e000000000000002a00000000",
            INIT_3E => X"00000078000000000000007200000000000000a2000000000000008300000000",
            INIT_3F => X"0000001500000000000000340000000000000085000000000000007600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006800000000000000310000000000000035000000000000004900000000",
            INIT_41 => X"0000004600000000000000390000000000000058000000000000007900000000",
            INIT_42 => X"0000005300000000000000470000000000000017000000000000003300000000",
            INIT_43 => X"000000070000000000000022000000000000004f000000000000004e00000000",
            INIT_44 => X"0000003e000000000000003c0000000000000051000000000000002800000000",
            INIT_45 => X"0000005d000000000000005b0000000000000063000000000000005000000000",
            INIT_46 => X"000000790000000000000078000000000000008d000000000000007300000000",
            INIT_47 => X"000000140000000000000021000000000000007c000000000000007900000000",
            INIT_48 => X"000000760000000000000038000000000000003a000000000000005600000000",
            INIT_49 => X"000000330000000000000040000000000000007f000000000000008300000000",
            INIT_4A => X"0000006300000000000000610000000000000040000000000000003b00000000",
            INIT_4B => X"0000001c000000000000000d000000000000003a000000000000005e00000000",
            INIT_4C => X"000000500000000000000049000000000000005d000000000000005300000000",
            INIT_4D => X"0000004a000000000000005f0000000000000069000000000000006200000000",
            INIT_4E => X"0000007e00000000000000770000000000000084000000000000007400000000",
            INIT_4F => X"00000017000000000000000d0000000000000065000000000000007f00000000",
            INIT_50 => X"000000740000000000000035000000000000003b000000000000005b00000000",
            INIT_51 => X"0000003000000000000000670000000000000087000000000000008400000000",
            INIT_52 => X"000000610000000000000060000000000000004b000000000000002000000000",
            INIT_53 => X"000000490000000000000032000000000000004a000000000000006600000000",
            INIT_54 => X"0000006100000000000000590000000000000052000000000000005a00000000",
            INIT_55 => X"000000310000000000000047000000000000006c000000000000006200000000",
            INIT_56 => X"0000008a0000000000000077000000000000007c000000000000007700000000",
            INIT_57 => X"00000014000000000000000a000000000000005b000000000000007b00000000",
            INIT_58 => X"0000006e000000000000002f0000000000000033000000000000006500000000",
            INIT_59 => X"0000004800000000000000870000000000000087000000000000008100000000",
            INIT_5A => X"0000004f00000000000000520000000000000054000000000000002e00000000",
            INIT_5B => X"0000008700000000000000750000000000000056000000000000005e00000000",
            INIT_5C => X"0000005e000000000000005d0000000000000066000000000000007800000000",
            INIT_5D => X"00000058000000000000004a0000000000000058000000000000005c00000000",
            INIT_5E => X"0000008d00000000000000760000000000000073000000000000008400000000",
            INIT_5F => X"00000007000000000000000b000000000000005b000000000000007700000000",
            INIT_60 => X"0000006000000000000000280000000000000028000000000000005800000000",
            INIT_61 => X"00000077000000000000008b0000000000000083000000000000006b00000000",
            INIT_62 => X"0000005900000000000000570000000000000066000000000000006b00000000",
            INIT_63 => X"0000006c0000000000000051000000000000004a000000000000005f00000000",
            INIT_64 => X"0000005d0000000000000064000000000000006e000000000000007600000000",
            INIT_65 => X"0000005f00000000000000570000000000000055000000000000006600000000",
            INIT_66 => X"0000007100000000000000650000000000000078000000000000007c00000000",
            INIT_67 => X"00000020000000000000000f0000000000000059000000000000007b00000000",
            INIT_68 => X"0000005c0000000000000037000000000000003f000000000000005f00000000",
            INIT_69 => X"00000089000000000000008b000000000000006e000000000000006400000000",
            INIT_6A => X"0000005c00000000000000650000000000000061000000000000007b00000000",
            INIT_6B => X"0000005600000000000000560000000000000058000000000000005a00000000",
            INIT_6C => X"0000006c00000000000000640000000000000058000000000000005500000000",
            INIT_6D => X"0000005f000000000000006e000000000000006c000000000000007200000000",
            INIT_6E => X"00000073000000000000006b0000000000000075000000000000006d00000000",
            INIT_6F => X"0000004c00000000000000310000000000000058000000000000008000000000",
            INIT_70 => X"0000006000000000000000470000000000000045000000000000006a00000000",
            INIT_71 => X"0000008700000000000000860000000000000056000000000000006800000000",
            INIT_72 => X"0000005800000000000000510000000000000057000000000000007400000000",
            INIT_73 => X"0000006a000000000000006e0000000000000060000000000000006000000000",
            INIT_74 => X"0000005c0000000000000057000000000000005f000000000000006200000000",
            INIT_75 => X"00000080000000000000007f000000000000006b000000000000006100000000",
            INIT_76 => X"000000770000000000000074000000000000005e000000000000007a00000000",
            INIT_77 => X"000000460000000000000035000000000000005c000000000000007a00000000",
            INIT_78 => X"0000005c00000000000000400000000000000040000000000000006000000000",
            INIT_79 => X"000000850000000000000079000000000000005f000000000000006700000000",
            INIT_7A => X"0000003300000000000000640000000000000096000000000000008100000000",
            INIT_7B => X"0000007100000000000000620000000000000065000000000000005800000000",
            INIT_7C => X"0000005f00000000000000650000000000000077000000000000008300000000",
            INIT_7D => X"0000009800000000000000710000000000000053000000000000006000000000",
            INIT_7E => X"0000007c00000000000000620000000000000078000000000000009400000000",
            INIT_7F => X"00000048000000000000000d0000000000000039000000000000007600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE28;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE29 : if BRAM_NAME = "sampleifmap_layersamples_instance29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005a0000000000000047000000000000004c000000000000005700000000",
            INIT_01 => X"000000820000000000000078000000000000007c000000000000007300000000",
            INIT_02 => X"0000003a0000000000000096000000000000008e000000000000006e00000000",
            INIT_03 => X"0000007800000000000000770000000000000074000000000000005400000000",
            INIT_04 => X"0000008600000000000000850000000000000071000000000000006c00000000",
            INIT_05 => X"0000006e0000000000000067000000000000007e000000000000008900000000",
            INIT_06 => X"00000072000000000000006300000000000000a3000000000000009f00000000",
            INIT_07 => X"0000006b0000000000000021000000000000002a000000000000007500000000",
            INIT_08 => X"0000005d00000000000000640000000000000058000000000000005600000000",
            INIT_09 => X"0000006900000000000000750000000000000063000000000000007500000000",
            INIT_0A => X"0000008b000000000000009b0000000000000066000000000000006e00000000",
            INIT_0B => X"000000810000000000000081000000000000006f000000000000006b00000000",
            INIT_0C => X"00000076000000000000006d0000000000000077000000000000007c00000000",
            INIT_0D => X"00000071000000000000007c0000000000000076000000000000007100000000",
            INIT_0E => X"0000006300000000000000830000000000000075000000000000008300000000",
            INIT_0F => X"0000005700000000000000270000000000000048000000000000006900000000",
            INIT_10 => X"0000007300000000000000780000000000000060000000000000005f00000000",
            INIT_11 => X"0000005600000000000000630000000000000047000000000000006d00000000",
            INIT_12 => X"000000b0000000000000006a0000000000000063000000000000006c00000000",
            INIT_13 => X"00000075000000000000007b000000000000005e000000000000008200000000",
            INIT_14 => X"000000880000000000000081000000000000008d000000000000008900000000",
            INIT_15 => X"000000790000000000000078000000000000006f000000000000008300000000",
            INIT_16 => X"000000430000000000000050000000000000006b000000000000007500000000",
            INIT_17 => X"0000006e00000000000000430000000000000051000000000000004800000000",
            INIT_18 => X"00000057000000000000007d0000000000000070000000000000006d00000000",
            INIT_19 => X"0000005e00000000000000470000000000000048000000000000005800000000",
            INIT_1A => X"0000007300000000000000490000000000000079000000000000006400000000",
            INIT_1B => X"0000009400000000000000870000000000000076000000000000009800000000",
            INIT_1C => X"0000009500000000000000940000000000000082000000000000008500000000",
            INIT_1D => X"0000007a00000000000000790000000000000071000000000000007d00000000",
            INIT_1E => X"0000004e000000000000003a0000000000000071000000000000007200000000",
            INIT_1F => X"0000008a00000000000000730000000000000038000000000000003d00000000",
            INIT_20 => X"0000004300000000000000590000000000000074000000000000007700000000",
            INIT_21 => X"00000066000000000000003c0000000000000048000000000000005800000000",
            INIT_22 => X"00000037000000000000006d0000000000000057000000000000004800000000",
            INIT_23 => X"0000009c000000000000008d0000000000000092000000000000006500000000",
            INIT_24 => X"00000098000000000000008c0000000000000088000000000000009800000000",
            INIT_25 => X"0000007c000000000000007f000000000000007b000000000000008600000000",
            INIT_26 => X"00000062000000000000005d0000000000000069000000000000006d00000000",
            INIT_27 => X"00000077000000000000007a0000000000000062000000000000004d00000000",
            INIT_28 => X"0000005d00000000000000320000000000000061000000000000007e00000000",
            INIT_29 => X"00000060000000000000004b0000000000000046000000000000006000000000",
            INIT_2A => X"000000610000000000000076000000000000003b000000000000005a00000000",
            INIT_2B => X"0000009700000000000000a20000000000000083000000000000004900000000",
            INIT_2C => X"0000007f000000000000008400000000000000a3000000000000009600000000",
            INIT_2D => X"00000075000000000000006e0000000000000076000000000000007d00000000",
            INIT_2E => X"0000004f000000000000005e0000000000000066000000000000006900000000",
            INIT_2F => X"0000006a0000000000000070000000000000008e000000000000006b00000000",
            INIT_30 => X"0000005900000000000000370000000000000051000000000000007000000000",
            INIT_31 => X"000000590000000000000045000000000000004e000000000000005c00000000",
            INIT_32 => X"000000760000000000000053000000000000006b000000000000007700000000",
            INIT_33 => X"0000009c0000000000000097000000000000007d000000000000006b00000000",
            INIT_34 => X"0000007e0000000000000094000000000000009b000000000000009400000000",
            INIT_35 => X"000000750000000000000078000000000000007b000000000000006c00000000",
            INIT_36 => X"0000005600000000000000540000000000000066000000000000007200000000",
            INIT_37 => X"0000006900000000000000630000000000000079000000000000008100000000",
            INIT_38 => X"0000009a00000000000000780000000000000056000000000000006200000000",
            INIT_39 => X"0000004e0000000000000045000000000000005f000000000000007700000000",
            INIT_3A => X"0000004e0000000000000057000000000000007e000000000000007300000000",
            INIT_3B => X"000000960000000000000084000000000000008b000000000000007d00000000",
            INIT_3C => X"0000007e0000000000000092000000000000008e000000000000008d00000000",
            INIT_3D => X"0000007b00000000000000760000000000000084000000000000007900000000",
            INIT_3E => X"0000006f00000000000000520000000000000058000000000000007300000000",
            INIT_3F => X"00000067000000000000006a0000000000000065000000000000007900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b600000000000000a70000000000000088000000000000007400000000",
            INIT_41 => X"0000005c00000000000000600000000000000077000000000000009f00000000",
            INIT_42 => X"0000006f0000000000000066000000000000005a000000000000006600000000",
            INIT_43 => X"0000008f00000000000000830000000000000088000000000000007000000000",
            INIT_44 => X"000000800000000000000096000000000000008e000000000000008600000000",
            INIT_45 => X"000000770000000000000084000000000000009c000000000000007500000000",
            INIT_46 => X"00000053000000000000004e0000000000000059000000000000006600000000",
            INIT_47 => X"0000006c00000000000000710000000000000060000000000000006a00000000",
            INIT_48 => X"000000920000000000000071000000000000006d000000000000006c00000000",
            INIT_49 => X"00000069000000000000007b000000000000009e00000000000000a600000000",
            INIT_4A => X"0000008c00000000000000550000000000000052000000000000006600000000",
            INIT_4B => X"0000007b0000000000000086000000000000007e000000000000009100000000",
            INIT_4C => X"00000089000000000000008a0000000000000073000000000000006800000000",
            INIT_4D => X"0000006a000000000000008a0000000000000096000000000000008300000000",
            INIT_4E => X"0000002d000000000000004a000000000000006f000000000000006100000000",
            INIT_4F => X"0000004b00000000000000690000000000000065000000000000006000000000",
            INIT_50 => X"0000005600000000000000370000000000000055000000000000005800000000",
            INIT_51 => X"0000007e00000000000000970000000000000097000000000000008b00000000",
            INIT_52 => X"0000005700000000000000570000000000000068000000000000006800000000",
            INIT_53 => X"00000052000000000000006e000000000000006e000000000000006f00000000",
            INIT_54 => X"0000008c0000000000000079000000000000004b000000000000003500000000",
            INIT_55 => X"0000007a00000000000000810000000000000078000000000000009100000000",
            INIT_56 => X"00000020000000000000003e0000000000000062000000000000007400000000",
            INIT_57 => X"0000004000000000000000410000000000000062000000000000006100000000",
            INIT_58 => X"000000200000000000000022000000000000005c000000000000005200000000",
            INIT_59 => X"0000009c00000000000000860000000000000075000000000000004b00000000",
            INIT_5A => X"000000570000000000000062000000000000006d000000000000008d00000000",
            INIT_5B => X"0000005f000000000000005b000000000000005a000000000000005200000000",
            INIT_5C => X"0000008b00000000000000790000000000000046000000000000005200000000",
            INIT_5D => X"0000006b0000000000000080000000000000008f000000000000008100000000",
            INIT_5E => X"0000003f000000000000001d000000000000004e000000000000007100000000",
            INIT_5F => X"0000004200000000000000470000000000000047000000000000006300000000",
            INIT_60 => X"0000000d00000000000000230000000000000056000000000000005a00000000",
            INIT_61 => X"000000940000000000000072000000000000004e000000000000000f00000000",
            INIT_62 => X"00000062000000000000006f000000000000008b00000000000000a200000000",
            INIT_63 => X"000000710000000000000056000000000000005b000000000000006100000000",
            INIT_64 => X"0000007e0000000000000073000000000000006a000000000000007800000000",
            INIT_65 => X"0000006a00000000000000870000000000000087000000000000007600000000",
            INIT_66 => X"0000005b0000000000000026000000000000002a000000000000004f00000000",
            INIT_67 => X"0000005300000000000000990000000000000060000000000000002c00000000",
            INIT_68 => X"00000025000000000000002d0000000000000056000000000000005c00000000",
            INIT_69 => X"0000007a0000000000000057000000000000001f000000000000000d00000000",
            INIT_6A => X"0000007a000000000000009e00000000000000ad000000000000009600000000",
            INIT_6B => X"0000005c000000000000005d0000000000000072000000000000007500000000",
            INIT_6C => X"0000007100000000000000670000000000000055000000000000004d00000000",
            INIT_6D => X"0000005b00000000000000730000000000000085000000000000007e00000000",
            INIT_6E => X"0000003c000000000000003b0000000000000032000000000000004e00000000",
            INIT_6F => X"000000620000000000000086000000000000006c000000000000002a00000000",
            INIT_70 => X"0000003800000000000000180000000000000047000000000000005200000000",
            INIT_71 => X"0000005400000000000000230000000000000017000000000000002400000000",
            INIT_72 => X"000000a500000000000000a50000000000000092000000000000007600000000",
            INIT_73 => X"00000079000000000000006f0000000000000082000000000000009600000000",
            INIT_74 => X"00000062000000000000003f0000000000000042000000000000006c00000000",
            INIT_75 => X"0000005600000000000000460000000000000045000000000000004e00000000",
            INIT_76 => X"000000620000000000000060000000000000006c000000000000007500000000",
            INIT_77 => X"00000059000000000000007b0000000000000074000000000000007800000000",
            INIT_78 => X"000000400000000000000011000000000000001b000000000000004100000000",
            INIT_79 => X"00000025000000000000000f000000000000001d000000000000003400000000",
            INIT_7A => X"0000009600000000000000740000000000000064000000000000005900000000",
            INIT_7B => X"0000009c0000000000000088000000000000009800000000000000aa00000000",
            INIT_7C => X"0000004a0000000000000045000000000000007900000000000000a600000000",
            INIT_7D => X"0000007f00000000000000660000000000000047000000000000002f00000000",
            INIT_7E => X"000000820000000000000083000000000000008b000000000000009c00000000",
            INIT_7F => X"0000007500000000000000920000000000000088000000000000009300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE29;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE30 : if BRAM_NAME = "sampleifmap_layersamples_instance30" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000058000000000000004d000000000000008b00000000000000b300000000",
            INIT_01 => X"00000097000000000000009c000000000000009d000000000000008d00000000",
            INIT_02 => X"000000970000000000000090000000000000009e000000000000009c00000000",
            INIT_03 => X"0000007600000000000000790000000000000088000000000000009700000000",
            INIT_04 => X"000000540000000000000054000000000000006c000000000000007e00000000",
            INIT_05 => X"00000053000000000000005e0000000000000062000000000000006200000000",
            INIT_06 => X"0000006000000000000000540000000000000056000000000000005a00000000",
            INIT_07 => X"0000004d000000000000004c0000000000000057000000000000007500000000",
            INIT_08 => X"000000920000000000000080000000000000008500000000000000b800000000",
            INIT_09 => X"000000a7000000000000009e000000000000009f000000000000009f00000000",
            INIT_0A => X"0000009a000000000000009900000000000000a200000000000000a500000000",
            INIT_0B => X"0000007d00000000000000880000000000000096000000000000009600000000",
            INIT_0C => X"00000052000000000000005a000000000000006d000000000000008100000000",
            INIT_0D => X"00000058000000000000005e0000000000000062000000000000005d00000000",
            INIT_0E => X"0000006a000000000000005b000000000000004c000000000000004e00000000",
            INIT_0F => X"0000005a000000000000005b0000000000000062000000000000007600000000",
            INIT_10 => X"000000aa00000000000000b0000000000000009800000000000000b400000000",
            INIT_11 => X"000000a4000000000000009b000000000000009800000000000000a400000000",
            INIT_12 => X"0000009f00000000000000a200000000000000aa00000000000000a200000000",
            INIT_13 => X"0000008c00000000000000920000000000000097000000000000009c00000000",
            INIT_14 => X"000000470000000000000058000000000000007c000000000000009200000000",
            INIT_15 => X"0000006b00000000000000670000000000000062000000000000005500000000",
            INIT_16 => X"0000006f000000000000006f000000000000006d000000000000006500000000",
            INIT_17 => X"0000005f000000000000005d0000000000000065000000000000006f00000000",
            INIT_18 => X"000000b500000000000000b800000000000000ae00000000000000af00000000",
            INIT_19 => X"000000a300000000000000a4000000000000009800000000000000a800000000",
            INIT_1A => X"000000a800000000000000a700000000000000b300000000000000a600000000",
            INIT_1B => X"000000a4000000000000009f00000000000000a200000000000000ae00000000",
            INIT_1C => X"0000003a00000000000000590000000000000089000000000000009700000000",
            INIT_1D => X"0000006b0000000000000063000000000000005a000000000000004800000000",
            INIT_1E => X"00000079000000000000007d0000000000000080000000000000007500000000",
            INIT_1F => X"0000006f000000000000006d0000000000000061000000000000006900000000",
            INIT_20 => X"000000ac00000000000000a700000000000000ae00000000000000af00000000",
            INIT_21 => X"000000af00000000000000b000000000000000a100000000000000a200000000",
            INIT_22 => X"000000b400000000000000b300000000000000b200000000000000b200000000",
            INIT_23 => X"000000a400000000000000a000000000000000a800000000000000b000000000",
            INIT_24 => X"000000450000000000000078000000000000009c00000000000000ad00000000",
            INIT_25 => X"0000005e0000000000000063000000000000005a000000000000004200000000",
            INIT_26 => X"0000007b000000000000007f000000000000007c000000000000006900000000",
            INIT_27 => X"0000007400000000000000710000000000000068000000000000007000000000",
            INIT_28 => X"000000aa000000000000009000000000000000ae00000000000000b500000000",
            INIT_29 => X"000000b300000000000000b000000000000000a600000000000000a900000000",
            INIT_2A => X"000000b500000000000000b400000000000000b400000000000000b400000000",
            INIT_2B => X"00000096000000000000009f00000000000000ae00000000000000b000000000",
            INIT_2C => X"00000074000000000000009b00000000000000af00000000000000b500000000",
            INIT_2D => X"000000700000000000000083000000000000007d000000000000006000000000",
            INIT_2E => X"00000079000000000000007a0000000000000078000000000000007500000000",
            INIT_2F => X"0000007c00000000000000760000000000000078000000000000007900000000",
            INIT_30 => X"000000b2000000000000008a000000000000009c00000000000000c000000000",
            INIT_31 => X"000000af00000000000000b000000000000000ae00000000000000af00000000",
            INIT_32 => X"000000b800000000000000ba00000000000000b400000000000000b800000000",
            INIT_33 => X"0000009900000000000000ad00000000000000bb00000000000000bb00000000",
            INIT_34 => X"000000a700000000000000ad00000000000000ad00000000000000a600000000",
            INIT_35 => X"0000007900000000000000940000000000000095000000000000009600000000",
            INIT_36 => X"0000006f000000000000006d0000000000000075000000000000007300000000",
            INIT_37 => X"00000080000000000000007b000000000000007a000000000000007800000000",
            INIT_38 => X"000000ab000000000000009c000000000000007d00000000000000b900000000",
            INIT_39 => X"000000b800000000000000af00000000000000af00000000000000ad00000000",
            INIT_3A => X"000000c200000000000000c100000000000000b700000000000000bc00000000",
            INIT_3B => X"000000a600000000000000b800000000000000b900000000000000bd00000000",
            INIT_3C => X"000000b000000000000000b100000000000000ac00000000000000a400000000",
            INIT_3D => X"0000007a000000000000008f000000000000008900000000000000aa00000000",
            INIT_3E => X"000000670000000000000060000000000000006e000000000000006b00000000",
            INIT_3F => X"0000007d000000000000007b0000000000000076000000000000007500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a0000000000000009f0000000000000095000000000000009b00000000",
            INIT_41 => X"000000b400000000000000b200000000000000ad00000000000000ac00000000",
            INIT_42 => X"000000bf00000000000000ba00000000000000ba00000000000000bb00000000",
            INIT_43 => X"000000a000000000000000ac00000000000000af00000000000000bb00000000",
            INIT_44 => X"000000b000000000000000a60000000000000097000000000000009a00000000",
            INIT_45 => X"0000008500000000000000a6000000000000009b00000000000000b700000000",
            INIT_46 => X"0000007700000000000000700000000000000068000000000000006800000000",
            INIT_47 => X"0000007d000000000000007a000000000000007a000000000000007600000000",
            INIT_48 => X"000000a900000000000000930000000000000098000000000000009a00000000",
            INIT_49 => X"000000aa00000000000000b700000000000000b200000000000000b200000000",
            INIT_4A => X"000000c100000000000000c600000000000000bc00000000000000b000000000",
            INIT_4B => X"000000a900000000000000a500000000000000a700000000000000ae00000000",
            INIT_4C => X"000000a90000000000000092000000000000008c000000000000009d00000000",
            INIT_4D => X"0000008d00000000000000ab00000000000000a000000000000000b300000000",
            INIT_4E => X"0000007700000000000000750000000000000068000000000000005f00000000",
            INIT_4F => X"0000007d0000000000000076000000000000007b000000000000007400000000",
            INIT_50 => X"000000b1000000000000009f0000000000000070000000000000008600000000",
            INIT_51 => X"000000ba00000000000000b800000000000000b800000000000000ae00000000",
            INIT_52 => X"000000b000000000000000bf00000000000000c200000000000000ba00000000",
            INIT_53 => X"000000bb00000000000000a7000000000000009e000000000000009b00000000",
            INIT_54 => X"000000970000000000000086000000000000009300000000000000ae00000000",
            INIT_55 => X"0000007c000000000000009b000000000000009c00000000000000a000000000",
            INIT_56 => X"0000006600000000000000690000000000000066000000000000004a00000000",
            INIT_57 => X"0000007f000000000000007b0000000000000075000000000000006b00000000",
            INIT_58 => X"0000009d00000000000000ae000000000000005b000000000000004100000000",
            INIT_59 => X"000000be00000000000000bf00000000000000b1000000000000009300000000",
            INIT_5A => X"000000b000000000000000ac00000000000000b000000000000000bc00000000",
            INIT_5B => X"000000a3000000000000009400000000000000ae00000000000000b800000000",
            INIT_5C => X"000000950000000000000085000000000000009a00000000000000b000000000",
            INIT_5D => X"0000005000000000000000830000000000000095000000000000009800000000",
            INIT_5E => X"0000006600000000000000670000000000000061000000000000004200000000",
            INIT_5F => X"0000007d00000000000000780000000000000071000000000000006700000000",
            INIT_60 => X"000000b100000000000000bf000000000000005c000000000000001500000000",
            INIT_61 => X"000000b600000000000000bd00000000000000ca00000000000000bc00000000",
            INIT_62 => X"000000bc00000000000000a5000000000000009c00000000000000b300000000",
            INIT_63 => X"00000072000000000000009800000000000000ae00000000000000c800000000",
            INIT_64 => X"000000890000000000000078000000000000007f000000000000005f00000000",
            INIT_65 => X"0000004e00000000000000720000000000000088000000000000009700000000",
            INIT_66 => X"0000006200000000000000590000000000000049000000000000004000000000",
            INIT_67 => X"0000007600000000000000750000000000000071000000000000006200000000",
            INIT_68 => X"000000ad00000000000000a80000000000000063000000000000002c00000000",
            INIT_69 => X"000000bb00000000000000bc00000000000000c300000000000000c800000000",
            INIT_6A => X"000000c200000000000000b4000000000000009500000000000000a500000000",
            INIT_6B => X"0000009a00000000000000a800000000000000a800000000000000b900000000",
            INIT_6C => X"0000008a00000000000000910000000000000092000000000000006b00000000",
            INIT_6D => X"000000480000000000000064000000000000007f000000000000009c00000000",
            INIT_6E => X"0000006000000000000000530000000000000040000000000000003900000000",
            INIT_6F => X"0000006f000000000000006c000000000000006a000000000000006200000000",
            INIT_70 => X"0000009f00000000000000750000000000000076000000000000006900000000",
            INIT_71 => X"000000bb00000000000000b400000000000000be00000000000000c400000000",
            INIT_72 => X"000000c100000000000000c600000000000000ad00000000000000ad00000000",
            INIT_73 => X"000000bc00000000000000b400000000000000a500000000000000ab00000000",
            INIT_74 => X"000000b300000000000000ad00000000000000bb00000000000000ae00000000",
            INIT_75 => X"000000480000000000000069000000000000008000000000000000a000000000",
            INIT_76 => X"0000006c00000000000000570000000000000045000000000000004300000000",
            INIT_77 => X"0000006600000000000000610000000000000064000000000000006300000000",
            INIT_78 => X"0000009d00000000000000680000000000000071000000000000008a00000000",
            INIT_79 => X"000000a800000000000000b400000000000000c400000000000000c600000000",
            INIT_7A => X"000000cd00000000000000cb00000000000000bf00000000000000b400000000",
            INIT_7B => X"000000c800000000000000c400000000000000bf00000000000000d200000000",
            INIT_7C => X"000000be00000000000000bc00000000000000bb00000000000000c000000000",
            INIT_7D => X"000000500000000000000071000000000000009900000000000000a800000000",
            INIT_7E => X"0000008700000000000000600000000000000040000000000000004600000000",
            INIT_7F => X"00000062000000000000005a000000000000005a000000000000007800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE30;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE31 : if BRAM_NAME = "sampleifmap_layersamples_instance31" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000930000000000000073000000000000008a000000000000009600000000",
            INIT_01 => X"0000009600000000000000b000000000000000bb00000000000000be00000000",
            INIT_02 => X"000000c600000000000000d300000000000000c700000000000000ab00000000",
            INIT_03 => X"000000cb00000000000000be00000000000000c200000000000000d300000000",
            INIT_04 => X"000000bd00000000000000b800000000000000ba00000000000000bf00000000",
            INIT_05 => X"00000046000000000000006400000000000000a600000000000000be00000000",
            INIT_06 => X"0000008f000000000000006a0000000000000038000000000000002f00000000",
            INIT_07 => X"0000005e000000000000004a000000000000005c000000000000009500000000",
            INIT_08 => X"000000a50000000000000092000000000000009b000000000000009b00000000",
            INIT_09 => X"0000009100000000000000bf00000000000000c000000000000000bd00000000",
            INIT_0A => X"0000009500000000000000a900000000000000d2000000000000009c00000000",
            INIT_0B => X"000000a800000000000000b200000000000000c200000000000000c000000000",
            INIT_0C => X"000000a700000000000000aa00000000000000b500000000000000a900000000",
            INIT_0D => X"0000002b00000000000000430000000000000075000000000000009a00000000",
            INIT_0E => X"0000008f00000000000000680000000000000031000000000000002200000000",
            INIT_0F => X"00000050000000000000003f000000000000006a000000000000009c00000000",
            INIT_10 => X"000000a6000000000000008a00000000000000a200000000000000a500000000",
            INIT_11 => X"0000008900000000000000ba00000000000000be00000000000000c400000000",
            INIT_12 => X"000000a9000000000000009d00000000000000c9000000000000007400000000",
            INIT_13 => X"0000008f000000000000008000000000000000b600000000000000d200000000",
            INIT_14 => X"00000061000000000000007f0000000000000093000000000000007c00000000",
            INIT_15 => X"00000033000000000000002f0000000000000038000000000000005200000000",
            INIT_16 => X"0000009d00000000000000690000000000000040000000000000002b00000000",
            INIT_17 => X"000000410000000000000039000000000000007b000000000000009d00000000",
            INIT_18 => X"0000009e0000000000000078000000000000009600000000000000a900000000",
            INIT_19 => X"0000009800000000000000be00000000000000be00000000000000be00000000",
            INIT_1A => X"000000b900000000000000bc0000000000000099000000000000003c00000000",
            INIT_1B => X"000000ce000000000000009000000000000000a500000000000000c300000000",
            INIT_1C => X"0000003d0000000000000065000000000000008900000000000000b100000000",
            INIT_1D => X"0000005000000000000000470000000000000033000000000000003700000000",
            INIT_1E => X"000000a0000000000000006e000000000000004a000000000000003700000000",
            INIT_1F => X"000000320000000000000036000000000000008e00000000000000b000000000",
            INIT_20 => X"000000a6000000000000009600000000000000a000000000000000aa00000000",
            INIT_21 => X"0000009a00000000000000ba00000000000000bc00000000000000ba00000000",
            INIT_22 => X"00000092000000000000007e0000000000000031000000000000002000000000",
            INIT_23 => X"000000c0000000000000008c000000000000008c000000000000009b00000000",
            INIT_24 => X"0000003e0000000000000061000000000000009c00000000000000cc00000000",
            INIT_25 => X"0000005700000000000000520000000000000049000000000000004900000000",
            INIT_26 => X"000000a6000000000000006b000000000000003e000000000000003a00000000",
            INIT_27 => X"00000033000000000000004800000000000000a700000000000000bc00000000",
            INIT_28 => X"0000009c000000000000009700000000000000ab00000000000000b200000000",
            INIT_29 => X"0000007c00000000000000a300000000000000b200000000000000b500000000",
            INIT_2A => X"000000370000000000000028000000000000001d000000000000002400000000",
            INIT_2B => X"0000008200000000000000650000000000000063000000000000004e00000000",
            INIT_2C => X"00000037000000000000005f000000000000007b000000000000009000000000",
            INIT_2D => X"00000055000000000000003c0000000000000033000000000000003400000000",
            INIT_2E => X"000000990000000000000066000000000000004d000000000000004e00000000",
            INIT_2F => X"00000037000000000000005900000000000000b100000000000000bb00000000",
            INIT_30 => X"00000098000000000000009200000000000000ab00000000000000b500000000",
            INIT_31 => X"00000069000000000000009500000000000000a700000000000000a900000000",
            INIT_32 => X"0000002e0000000000000042000000000000005e000000000000004f00000000",
            INIT_33 => X"00000078000000000000005c0000000000000047000000000000002f00000000",
            INIT_34 => X"0000002900000000000000380000000000000037000000000000005a00000000",
            INIT_35 => X"00000037000000000000001e0000000000000022000000000000002300000000",
            INIT_36 => X"0000007700000000000000610000000000000056000000000000005200000000",
            INIT_37 => X"0000003c000000000000006a00000000000000ae00000000000000ad00000000",
            INIT_38 => X"000000a3000000000000009e000000000000009c00000000000000b100000000",
            INIT_39 => X"00000089000000000000009400000000000000a0000000000000009c00000000",
            INIT_3A => X"0000006b00000000000000660000000000000076000000000000008f00000000",
            INIT_3B => X"00000067000000000000007d000000000000006d000000000000006e00000000",
            INIT_3C => X"0000001300000000000000100000000000000011000000000000002f00000000",
            INIT_3D => X"00000013000000000000000e000000000000001c000000000000001800000000",
            INIT_3E => X"0000006300000000000000600000000000000041000000000000002b00000000",
            INIT_3F => X"00000043000000000000008500000000000000ad000000000000008c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b600000000000000a7000000000000008b000000000000009e00000000",
            INIT_41 => X"000000c000000000000000ab000000000000008c000000000000009700000000",
            INIT_42 => X"000000880000000000000085000000000000007400000000000000ac00000000",
            INIT_43 => X"00000065000000000000007f000000000000008d000000000000009200000000",
            INIT_44 => X"0000001900000000000000200000000000000025000000000000004100000000",
            INIT_45 => X"0000000f000000000000000a0000000000000011000000000000001800000000",
            INIT_46 => X"0000004e00000000000000610000000000000042000000000000001400000000",
            INIT_47 => X"00000069000000000000009c0000000000000094000000000000006200000000",
            INIT_48 => X"000000ab00000000000000ae00000000000000a400000000000000a000000000",
            INIT_49 => X"000000b100000000000000940000000000000088000000000000009e00000000",
            INIT_4A => X"0000009700000000000000a9000000000000009300000000000000b800000000",
            INIT_4B => X"0000007d000000000000008e000000000000008b000000000000007f00000000",
            INIT_4C => X"0000002b000000000000003f000000000000004d000000000000006700000000",
            INIT_4D => X"0000001a00000000000000110000000000000018000000000000002100000000",
            INIT_4E => X"000000320000000000000048000000000000003e000000000000001f00000000",
            INIT_4F => X"000000880000000000000078000000000000005a000000000000004800000000",
            INIT_50 => X"000000a700000000000000a700000000000000a300000000000000a000000000",
            INIT_51 => X"00000078000000000000008c00000000000000a800000000000000b100000000",
            INIT_52 => X"000000820000000000000076000000000000008f00000000000000ab00000000",
            INIT_53 => X"0000009100000000000000a6000000000000009c000000000000007b00000000",
            INIT_54 => X"0000004e000000000000005b0000000000000069000000000000007c00000000",
            INIT_55 => X"0000004300000000000000380000000000000042000000000000004c00000000",
            INIT_56 => X"0000004900000000000000410000000000000041000000000000004600000000",
            INIT_57 => X"0000006a0000000000000051000000000000007b000000000000006400000000",
            INIT_58 => X"00000093000000000000008c000000000000009f000000000000009c00000000",
            INIT_59 => X"0000007b000000000000009900000000000000aa00000000000000b400000000",
            INIT_5A => X"0000007e0000000000000073000000000000009c000000000000008b00000000",
            INIT_5B => X"000000a200000000000000a8000000000000009e000000000000008300000000",
            INIT_5C => X"00000078000000000000007b0000000000000077000000000000007f00000000",
            INIT_5D => X"0000007700000000000000690000000000000068000000000000007000000000",
            INIT_5E => X"0000006d00000000000000680000000000000069000000000000007400000000",
            INIT_5F => X"00000068000000000000005c0000000000000086000000000000007a00000000",
            INIT_60 => X"0000008b000000000000007b000000000000009e00000000000000a400000000",
            INIT_61 => X"0000008c000000000000008d000000000000009c00000000000000ad00000000",
            INIT_62 => X"000000a100000000000000820000000000000079000000000000008d00000000",
            INIT_63 => X"000000a800000000000000a6000000000000009d000000000000009700000000",
            INIT_64 => X"00000084000000000000008f000000000000008a000000000000009000000000",
            INIT_65 => X"00000094000000000000008a0000000000000085000000000000008100000000",
            INIT_66 => X"0000008400000000000000860000000000000089000000000000008f00000000",
            INIT_67 => X"0000009300000000000000730000000000000064000000000000007800000000",
            INIT_68 => X"000000a800000000000000900000000000000095000000000000008e00000000",
            INIT_69 => X"0000009e000000000000009e00000000000000a100000000000000a700000000",
            INIT_6A => X"000000a90000000000000097000000000000009000000000000000a500000000",
            INIT_6B => X"000000a2000000000000009e00000000000000a000000000000000a100000000",
            INIT_6C => X"0000007f00000000000000890000000000000091000000000000009900000000",
            INIT_6D => X"0000009e00000000000000960000000000000095000000000000008d00000000",
            INIT_6E => X"0000008f00000000000000940000000000000096000000000000009f00000000",
            INIT_6F => X"0000009f000000000000008b0000000000000077000000000000007b00000000",
            INIT_70 => X"000000b900000000000000b300000000000000a6000000000000009800000000",
            INIT_71 => X"000000a800000000000000aa00000000000000a700000000000000a700000000",
            INIT_72 => X"000000b200000000000000ad00000000000000a400000000000000a700000000",
            INIT_73 => X"000000850000000000000089000000000000009d00000000000000a900000000",
            INIT_74 => X"00000088000000000000008c000000000000008f000000000000009200000000",
            INIT_75 => X"0000009d00000000000000980000000000000097000000000000008c00000000",
            INIT_76 => X"000000900000000000000099000000000000009c00000000000000a600000000",
            INIT_77 => X"0000009900000000000000900000000000000083000000000000008500000000",
            INIT_78 => X"000000ab00000000000000b700000000000000b2000000000000009f00000000",
            INIT_79 => X"0000009f0000000000000091000000000000007d000000000000008b00000000",
            INIT_7A => X"0000009c0000000000000095000000000000008b00000000000000a200000000",
            INIT_7B => X"0000007300000000000000830000000000000098000000000000009e00000000",
            INIT_7C => X"0000008f0000000000000094000000000000008e000000000000008400000000",
            INIT_7D => X"000000a1000000000000009c000000000000009d000000000000009000000000",
            INIT_7E => X"0000009c0000000000000094000000000000009f00000000000000a700000000",
            INIT_7F => X"0000009800000000000000990000000000000096000000000000009c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE31;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE32 : if BRAM_NAME = "sampleifmap_layersamples_instance32" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003b00000000000000310000000000000060000000000000007600000000",
            INIT_01 => X"000000530000000000000054000000000000005f000000000000006000000000",
            INIT_02 => X"0000005a00000000000000530000000000000061000000000000005f00000000",
            INIT_03 => X"0000004f000000000000004b0000000000000052000000000000005c00000000",
            INIT_04 => X"00000032000000000000003b0000000000000050000000000000005b00000000",
            INIT_05 => X"0000003300000000000000380000000000000038000000000000003700000000",
            INIT_06 => X"0000003a00000000000000330000000000000038000000000000003c00000000",
            INIT_07 => X"0000002f000000000000002f0000000000000035000000000000004c00000000",
            INIT_08 => X"0000006900000000000000590000000000000058000000000000008200000000",
            INIT_09 => X"00000068000000000000005d0000000000000060000000000000006c00000000",
            INIT_0A => X"0000005b000000000000005a0000000000000062000000000000006500000000",
            INIT_0B => X"00000048000000000000004f0000000000000057000000000000005400000000",
            INIT_0C => X"00000032000000000000003d0000000000000048000000000000005200000000",
            INIT_0D => X"0000003300000000000000370000000000000038000000000000003700000000",
            INIT_0E => X"0000004100000000000000350000000000000028000000000000002b00000000",
            INIT_0F => X"00000039000000000000003a000000000000003d000000000000004b00000000",
            INIT_10 => X"0000007a00000000000000810000000000000068000000000000008400000000",
            INIT_11 => X"0000006a000000000000005f0000000000000059000000000000006c00000000",
            INIT_12 => X"0000005e00000000000000620000000000000069000000000000006200000000",
            INIT_13 => X"0000004c000000000000004f0000000000000050000000000000005500000000",
            INIT_14 => X"0000002a0000000000000036000000000000004c000000000000005500000000",
            INIT_15 => X"00000042000000000000003f000000000000003a000000000000003300000000",
            INIT_16 => X"0000004200000000000000430000000000000042000000000000003c00000000",
            INIT_17 => X"000000390000000000000038000000000000003e000000000000004300000000",
            INIT_18 => X"000000840000000000000088000000000000007f000000000000008100000000",
            INIT_19 => X"000000690000000000000068000000000000005a000000000000007000000000",
            INIT_1A => X"0000006600000000000000650000000000000071000000000000006500000000",
            INIT_1B => X"0000005d0000000000000057000000000000005a000000000000006700000000",
            INIT_1C => X"0000001f0000000000000033000000000000004e000000000000004f00000000",
            INIT_1D => X"0000003e00000000000000390000000000000033000000000000002a00000000",
            INIT_1E => X"0000004a000000000000004b000000000000004d000000000000004600000000",
            INIT_1F => X"0000004500000000000000430000000000000037000000000000003c00000000",
            INIT_20 => X"0000007f0000000000000079000000000000007f000000000000008000000000",
            INIT_21 => X"0000007200000000000000720000000000000063000000000000006d00000000",
            INIT_22 => X"000000710000000000000070000000000000006f000000000000006f00000000",
            INIT_23 => X"0000005c00000000000000590000000000000063000000000000006c00000000",
            INIT_24 => X"0000002c000000000000004e0000000000000059000000000000005e00000000",
            INIT_25 => X"0000002e00000000000000380000000000000034000000000000002700000000",
            INIT_26 => X"0000004900000000000000470000000000000043000000000000003500000000",
            INIT_27 => X"000000470000000000000045000000000000003b000000000000004200000000",
            INIT_28 => X"0000007f00000000000000680000000000000083000000000000008900000000",
            INIT_29 => X"000000740000000000000071000000000000006a000000000000007600000000",
            INIT_2A => X"0000007100000000000000740000000000000075000000000000007300000000",
            INIT_2B => X"00000054000000000000005a0000000000000069000000000000006d00000000",
            INIT_2C => X"0000004f00000000000000670000000000000068000000000000006a00000000",
            INIT_2D => X"0000003d0000000000000052000000000000004d000000000000003a00000000",
            INIT_2E => X"000000460000000000000043000000000000003f000000000000003e00000000",
            INIT_2F => X"0000004b00000000000000460000000000000048000000000000004900000000",
            INIT_30 => X"0000008700000000000000660000000000000077000000000000009800000000",
            INIT_31 => X"0000006f00000000000000730000000000000075000000000000007a00000000",
            INIT_32 => X"00000070000000000000007c000000000000007b000000000000007900000000",
            INIT_33 => X"0000005c00000000000000660000000000000071000000000000007300000000",
            INIT_34 => X"0000006e000000000000006d0000000000000065000000000000006400000000",
            INIT_35 => X"00000043000000000000005b0000000000000057000000000000005c00000000",
            INIT_36 => X"0000003b00000000000000380000000000000040000000000000003e00000000",
            INIT_37 => X"0000004e000000000000004a0000000000000048000000000000004500000000",
            INIT_38 => X"0000007e00000000000000780000000000000059000000000000009300000000",
            INIT_39 => X"0000007900000000000000720000000000000076000000000000007800000000",
            INIT_3A => X"00000073000000000000007c000000000000007a000000000000008000000000",
            INIT_3B => X"00000064000000000000006c000000000000006d000000000000007300000000",
            INIT_3C => X"0000006a000000000000006d0000000000000068000000000000006500000000",
            INIT_3D => X"000000480000000000000057000000000000004b000000000000006600000000",
            INIT_3E => X"00000035000000000000002e000000000000003c000000000000003b00000000",
            INIT_3F => X"0000004b00000000000000490000000000000044000000000000004200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000720000000000000078000000000000006f000000000000007600000000",
            INIT_41 => X"0000007700000000000000750000000000000074000000000000007700000000",
            INIT_42 => X"0000006d000000000000006f000000000000007a000000000000008000000000",
            INIT_43 => X"0000005e00000000000000610000000000000067000000000000007300000000",
            INIT_44 => X"0000006400000000000000610000000000000059000000000000005e00000000",
            INIT_45 => X"000000590000000000000072000000000000005f000000000000006d00000000",
            INIT_46 => X"000000470000000000000040000000000000003a000000000000003e00000000",
            INIT_47 => X"0000004b00000000000000480000000000000048000000000000004600000000",
            INIT_48 => X"0000007800000000000000690000000000000071000000000000007700000000",
            INIT_49 => X"0000006f000000000000007b000000000000007a000000000000007c00000000",
            INIT_4A => X"00000079000000000000007d000000000000007b000000000000007600000000",
            INIT_4B => X"0000006f0000000000000065000000000000006d000000000000007600000000",
            INIT_4C => X"0000006000000000000000520000000000000055000000000000006900000000",
            INIT_4D => X"00000067000000000000007a0000000000000064000000000000006a00000000",
            INIT_4E => X"000000490000000000000047000000000000003e000000000000003d00000000",
            INIT_4F => X"0000004b0000000000000044000000000000004b000000000000004700000000",
            INIT_50 => X"0000007e00000000000000720000000000000048000000000000006400000000",
            INIT_51 => X"0000007e000000000000007c000000000000007f000000000000007800000000",
            INIT_52 => X"0000007b00000000000000800000000000000081000000000000007f00000000",
            INIT_53 => X"0000009000000000000000780000000000000077000000000000007900000000",
            INIT_54 => X"00000058000000000000004f0000000000000063000000000000008300000000",
            INIT_55 => X"0000005b000000000000006c0000000000000061000000000000005f00000000",
            INIT_56 => X"0000003b000000000000003d000000000000003e000000000000002e00000000",
            INIT_57 => X"0000004c00000000000000490000000000000046000000000000004000000000",
            INIT_58 => X"00000069000000000000007f0000000000000034000000000000002200000000",
            INIT_59 => X"000000830000000000000084000000000000007a000000000000005d00000000",
            INIT_5A => X"0000008c00000000000000780000000000000073000000000000008100000000",
            INIT_5B => X"000000850000000000000074000000000000009700000000000000a600000000",
            INIT_5C => X"000000610000000000000056000000000000006e000000000000008d00000000",
            INIT_5D => X"000000310000000000000056000000000000005c000000000000006000000000",
            INIT_5E => X"0000003c000000000000003e000000000000003c000000000000002a00000000",
            INIT_5F => X"0000004a00000000000000450000000000000042000000000000003e00000000",
            INIT_60 => X"0000007d000000000000008e0000000000000040000000000000000400000000",
            INIT_61 => X"00000084000000000000008c000000000000009a000000000000008c00000000",
            INIT_62 => X"0000009c000000000000007b000000000000006b000000000000007f00000000",
            INIT_63 => X"000000530000000000000077000000000000009300000000000000b200000000",
            INIT_64 => X"000000640000000000000053000000000000005b000000000000004000000000",
            INIT_65 => X"00000031000000000000004d000000000000005c000000000000006f00000000",
            INIT_66 => X"000000390000000000000037000000000000002f000000000000002900000000",
            INIT_67 => X"0000004400000000000000420000000000000043000000000000003b00000000",
            INIT_68 => X"0000007b000000000000007a0000000000000048000000000000001800000000",
            INIT_69 => X"0000008d000000000000008f0000000000000096000000000000009c00000000",
            INIT_6A => X"000000a0000000000000008f000000000000006a000000000000007700000000",
            INIT_6B => X"0000007700000000000000800000000000000081000000000000009700000000",
            INIT_6C => X"0000006d00000000000000730000000000000074000000000000004d00000000",
            INIT_6D => X"0000002d0000000000000044000000000000005a000000000000007b00000000",
            INIT_6E => X"000000370000000000000033000000000000002b000000000000002300000000",
            INIT_6F => X"0000003e000000000000003a000000000000003e000000000000003b00000000",
            INIT_70 => X"00000070000000000000004a0000000000000052000000000000004500000000",
            INIT_71 => X"0000008f00000000000000860000000000000091000000000000009600000000",
            INIT_72 => X"0000009c00000000000000a10000000000000084000000000000008300000000",
            INIT_73 => X"0000009700000000000000850000000000000072000000000000007d00000000",
            INIT_74 => X"00000098000000000000009200000000000000a0000000000000009100000000",
            INIT_75 => X"0000002f000000000000004b000000000000005d000000000000008100000000",
            INIT_76 => X"0000004400000000000000380000000000000030000000000000002f00000000",
            INIT_77 => X"000000390000000000000036000000000000003c000000000000003c00000000",
            INIT_78 => X"00000070000000000000003b0000000000000041000000000000005700000000",
            INIT_79 => X"0000007d00000000000000860000000000000096000000000000009800000000",
            INIT_7A => X"000000a500000000000000a7000000000000009b000000000000008f00000000",
            INIT_7B => X"000000a0000000000000008f0000000000000084000000000000009b00000000",
            INIT_7C => X"000000a1000000000000009f000000000000009e00000000000000a200000000",
            INIT_7D => X"0000003900000000000000540000000000000078000000000000008900000000",
            INIT_7E => X"0000005f0000000000000040000000000000002b000000000000003300000000",
            INIT_7F => X"0000003900000000000000360000000000000037000000000000005100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE32;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE33 : if BRAM_NAME = "sampleifmap_layersamples_instance33" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000660000000000000040000000000000004e000000000000005800000000",
            INIT_01 => X"0000006c0000000000000081000000000000008d000000000000009000000000",
            INIT_02 => X"0000009d00000000000000af00000000000000a5000000000000008b00000000",
            INIT_03 => X"0000009f00000000000000860000000000000086000000000000009e00000000",
            INIT_04 => X"0000009800000000000000930000000000000094000000000000009a00000000",
            INIT_05 => X"0000003100000000000000490000000000000087000000000000009a00000000",
            INIT_06 => X"00000067000000000000004b0000000000000023000000000000001e00000000",
            INIT_07 => X"00000039000000000000002c000000000000003d000000000000006f00000000",
            INIT_08 => X"0000007400000000000000570000000000000057000000000000005600000000",
            INIT_09 => X"0000006900000000000000910000000000000093000000000000008f00000000",
            INIT_0A => X"0000006c000000000000008500000000000000b3000000000000008000000000",
            INIT_0B => X"00000079000000000000007a000000000000008b000000000000009100000000",
            INIT_0C => X"00000079000000000000007c0000000000000087000000000000007d00000000",
            INIT_0D => X"00000018000000000000002a0000000000000058000000000000007200000000",
            INIT_0E => X"000000660000000000000049000000000000001d000000000000001300000000",
            INIT_0F => X"0000002e00000000000000270000000000000050000000000000007500000000",
            INIT_10 => X"00000076000000000000004d000000000000005c000000000000005c00000000",
            INIT_11 => X"0000006200000000000000910000000000000099000000000000009c00000000",
            INIT_12 => X"0000007a000000000000007400000000000000aa000000000000005c00000000",
            INIT_13 => X"00000062000000000000004b000000000000008300000000000000a500000000",
            INIT_14 => X"0000004000000000000000550000000000000061000000000000004c00000000",
            INIT_15 => X"0000001b0000000000000011000000000000001b000000000000003600000000",
            INIT_16 => X"0000007500000000000000450000000000000028000000000000001a00000000",
            INIT_17 => X"0000002800000000000000240000000000000064000000000000007f00000000",
            INIT_18 => X"0000006e000000000000003c0000000000000054000000000000005e00000000",
            INIT_19 => X"00000073000000000000009b00000000000000a3000000000000009c00000000",
            INIT_1A => X"000000890000000000000094000000000000007c000000000000002700000000",
            INIT_1B => X"0000009c00000000000000570000000000000071000000000000009500000000",
            INIT_1C => X"00000027000000000000003d0000000000000050000000000000007800000000",
            INIT_1D => X"0000002e00000000000000220000000000000018000000000000002700000000",
            INIT_1E => X"000000780000000000000045000000000000002d000000000000001f00000000",
            INIT_1F => X"000000200000000000000022000000000000007b000000000000009900000000",
            INIT_20 => X"000000720000000000000059000000000000005d000000000000006100000000",
            INIT_21 => X"00000075000000000000009800000000000000a2000000000000009600000000",
            INIT_22 => X"000000740000000000000064000000000000001d000000000000000d00000000",
            INIT_23 => X"0000007c00000000000000490000000000000056000000000000007300000000",
            INIT_24 => X"0000001b000000000000002f000000000000005b000000000000008600000000",
            INIT_25 => X"0000003200000000000000310000000000000032000000000000003100000000",
            INIT_26 => X"0000007d0000000000000042000000000000001e000000000000001900000000",
            INIT_27 => X"000000200000000000000038000000000000009600000000000000a200000000",
            INIT_28 => X"0000006300000000000000570000000000000068000000000000006a00000000",
            INIT_29 => X"0000005700000000000000810000000000000096000000000000008d00000000",
            INIT_2A => X"000000250000000000000016000000000000000b000000000000000f00000000",
            INIT_2B => X"0000003e00000000000000290000000000000039000000000000003600000000",
            INIT_2C => X"0000001a00000000000000360000000000000048000000000000005300000000",
            INIT_2D => X"0000003300000000000000220000000000000023000000000000002000000000",
            INIT_2E => X"00000070000000000000003e000000000000002b000000000000002800000000",
            INIT_2F => X"0000001f000000000000004a000000000000009e000000000000009b00000000",
            INIT_30 => X"0000005a000000000000004f0000000000000068000000000000007000000000",
            INIT_31 => X"0000004200000000000000730000000000000089000000000000007b00000000",
            INIT_32 => X"0000001700000000000000280000000000000042000000000000002f00000000",
            INIT_33 => X"00000045000000000000002c0000000000000026000000000000001b00000000",
            INIT_34 => X"0000001d0000000000000026000000000000001f000000000000003600000000",
            INIT_35 => X"0000001f000000000000000f0000000000000016000000000000001900000000",
            INIT_36 => X"0000004e000000000000003a0000000000000033000000000000003100000000",
            INIT_37 => X"0000001f00000000000000570000000000000094000000000000008600000000",
            INIT_38 => X"0000006000000000000000590000000000000058000000000000006d00000000",
            INIT_39 => X"0000005e00000000000000730000000000000081000000000000006900000000",
            INIT_3A => X"0000003c00000000000000360000000000000047000000000000006100000000",
            INIT_3B => X"0000003c000000000000004b000000000000003e000000000000004200000000",
            INIT_3C => X"0000000e0000000000000009000000000000000a000000000000001a00000000",
            INIT_3D => X"0000000c000000000000000b0000000000000013000000000000001100000000",
            INIT_3E => X"0000003b000000000000003a000000000000001f000000000000001700000000",
            INIT_3F => X"0000002300000000000000690000000000000088000000000000005e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007000000000000000600000000000000046000000000000005b00000000",
            INIT_41 => X"0000009300000000000000890000000000000068000000000000006000000000",
            INIT_42 => X"000000430000000000000045000000000000003a000000000000007500000000",
            INIT_43 => X"00000035000000000000003f0000000000000045000000000000004a00000000",
            INIT_44 => X"0000000d00000000000000130000000000000019000000000000002900000000",
            INIT_45 => X"00000012000000000000000d0000000000000009000000000000000c00000000",
            INIT_46 => X"00000027000000000000003e0000000000000024000000000000000c00000000",
            INIT_47 => X"0000004700000000000000790000000000000068000000000000003400000000",
            INIT_48 => X"000000620000000000000062000000000000005c000000000000005b00000000",
            INIT_49 => X"0000008600000000000000690000000000000056000000000000006100000000",
            INIT_4A => X"00000061000000000000007c000000000000006b000000000000008e00000000",
            INIT_4B => X"00000049000000000000004e0000000000000049000000000000004400000000",
            INIT_4C => X"0000001c0000000000000026000000000000002b000000000000003e00000000",
            INIT_4D => X"00000014000000000000000b000000000000000e000000000000001600000000",
            INIT_4E => X"000000140000000000000030000000000000002a000000000000001400000000",
            INIT_4F => X"0000006400000000000000580000000000000038000000000000002500000000",
            INIT_50 => X"000000620000000000000061000000000000005e000000000000005b00000000",
            INIT_51 => X"0000004c000000000000005b000000000000006f000000000000007100000000",
            INIT_52 => X"000000510000000000000050000000000000006e000000000000008400000000",
            INIT_53 => X"000000540000000000000063000000000000005f000000000000004700000000",
            INIT_54 => X"000000330000000000000038000000000000003d000000000000004800000000",
            INIT_55 => X"0000002b0000000000000020000000000000002b000000000000003500000000",
            INIT_56 => X"0000002800000000000000250000000000000028000000000000002e00000000",
            INIT_57 => X"000000420000000000000030000000000000005a000000000000004000000000",
            INIT_58 => X"0000005200000000000000500000000000000060000000000000005700000000",
            INIT_59 => X"000000480000000000000062000000000000006d000000000000007100000000",
            INIT_5A => X"0000004600000000000000450000000000000073000000000000005c00000000",
            INIT_5B => X"000000580000000000000060000000000000005e000000000000004a00000000",
            INIT_5C => X"0000004a000000000000004c0000000000000047000000000000004500000000",
            INIT_5D => X"0000004b000000000000003d000000000000003c000000000000004200000000",
            INIT_5E => X"00000041000000000000003f0000000000000040000000000000004900000000",
            INIT_5F => X"0000003a0000000000000036000000000000005e000000000000004c00000000",
            INIT_60 => X"0000004c00000000000000430000000000000061000000000000006000000000",
            INIT_61 => X"00000050000000000000004e000000000000005a000000000000006900000000",
            INIT_62 => X"00000062000000000000004c0000000000000048000000000000005700000000",
            INIT_63 => X"0000005a000000000000005d000000000000005c000000000000005700000000",
            INIT_64 => X"0000004600000000000000550000000000000054000000000000004f00000000",
            INIT_65 => X"00000057000000000000004d0000000000000048000000000000004200000000",
            INIT_66 => X"0000004f00000000000000500000000000000052000000000000005300000000",
            INIT_67 => X"0000005e00000000000000460000000000000035000000000000004300000000",
            INIT_68 => X"0000006500000000000000510000000000000054000000000000004900000000",
            INIT_69 => X"0000005b0000000000000058000000000000005b000000000000006100000000",
            INIT_6A => X"00000063000000000000005b0000000000000059000000000000006900000000",
            INIT_6B => X"0000005a000000000000005d000000000000005d000000000000005900000000",
            INIT_6C => X"0000003c00000000000000490000000000000055000000000000005800000000",
            INIT_6D => X"0000005b00000000000000540000000000000052000000000000004900000000",
            INIT_6E => X"0000005500000000000000570000000000000056000000000000005d00000000",
            INIT_6F => X"0000006400000000000000570000000000000044000000000000004300000000",
            INIT_70 => X"00000071000000000000006a0000000000000060000000000000005300000000",
            INIT_71 => X"0000005f0000000000000060000000000000005f000000000000006000000000",
            INIT_72 => X"00000068000000000000006d0000000000000069000000000000006600000000",
            INIT_73 => X"0000004a0000000000000052000000000000005a000000000000005b00000000",
            INIT_74 => X"0000004a000000000000004d000000000000004e000000000000005200000000",
            INIT_75 => X"0000005c00000000000000570000000000000055000000000000004d00000000",
            INIT_76 => X"00000054000000000000005a0000000000000059000000000000006400000000",
            INIT_77 => X"0000005a0000000000000057000000000000004d000000000000004e00000000",
            INIT_78 => X"000000680000000000000071000000000000006b000000000000005c00000000",
            INIT_79 => X"0000005c000000000000004d0000000000000042000000000000005200000000",
            INIT_7A => X"0000005a000000000000005b0000000000000051000000000000005f00000000",
            INIT_7B => X"0000003d000000000000004d000000000000005b000000000000005800000000",
            INIT_7C => X"000000520000000000000056000000000000004d000000000000004600000000",
            INIT_7D => X"00000060000000000000005b000000000000005c000000000000005300000000",
            INIT_7E => X"0000005b0000000000000057000000000000005c000000000000006500000000",
            INIT_7F => X"00000057000000000000005b000000000000005a000000000000005c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE33;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE34 : if BRAM_NAME = "sampleifmap_layersamples_instance34" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000024000000000000001a000000000000003d000000000000005300000000",
            INIT_01 => X"00000036000000000000003a0000000000000043000000000000004100000000",
            INIT_02 => X"0000003b00000000000000340000000000000041000000000000003f00000000",
            INIT_03 => X"00000034000000000000002e0000000000000035000000000000003e00000000",
            INIT_04 => X"00000027000000000000002b0000000000000041000000000000004700000000",
            INIT_05 => X"00000026000000000000002d000000000000002f000000000000002f00000000",
            INIT_06 => X"00000032000000000000002a000000000000002d000000000000002f00000000",
            INIT_07 => X"000000290000000000000029000000000000002e000000000000004500000000",
            INIT_08 => X"00000046000000000000003a0000000000000035000000000000006100000000",
            INIT_09 => X"0000004d00000000000000440000000000000043000000000000004600000000",
            INIT_0A => X"0000003900000000000000380000000000000041000000000000004400000000",
            INIT_0B => X"0000002e00000000000000320000000000000039000000000000003400000000",
            INIT_0C => X"00000026000000000000002b0000000000000034000000000000003c00000000",
            INIT_0D => X"00000028000000000000002c000000000000002f000000000000002f00000000",
            INIT_0E => X"00000038000000000000002b000000000000001e000000000000002000000000",
            INIT_0F => X"0000003100000000000000330000000000000035000000000000004300000000",
            INIT_10 => X"00000051000000000000005c0000000000000047000000000000006400000000",
            INIT_11 => X"0000004e00000000000000440000000000000039000000000000004400000000",
            INIT_12 => X"0000003b000000000000003f0000000000000047000000000000004000000000",
            INIT_13 => X"0000003000000000000000310000000000000030000000000000003400000000",
            INIT_14 => X"0000001e00000000000000210000000000000032000000000000003b00000000",
            INIT_15 => X"0000003800000000000000350000000000000030000000000000002b00000000",
            INIT_16 => X"0000003800000000000000390000000000000038000000000000003300000000",
            INIT_17 => X"00000031000000000000002f0000000000000035000000000000003900000000",
            INIT_18 => X"000000590000000000000061000000000000005f000000000000006000000000",
            INIT_19 => X"0000004800000000000000490000000000000037000000000000004900000000",
            INIT_1A => X"000000420000000000000042000000000000004e000000000000004100000000",
            INIT_1B => X"0000003f00000000000000360000000000000037000000000000004300000000",
            INIT_1C => X"00000012000000000000001a000000000000002e000000000000002f00000000",
            INIT_1D => X"00000035000000000000002f0000000000000029000000000000002200000000",
            INIT_1E => X"0000003e00000000000000400000000000000044000000000000003d00000000",
            INIT_1F => X"0000003c000000000000003a000000000000002d000000000000003000000000",
            INIT_20 => X"0000005700000000000000540000000000000061000000000000005c00000000",
            INIT_21 => X"0000004b000000000000004c000000000000003f000000000000004900000000",
            INIT_22 => X"0000004b000000000000004b000000000000004a000000000000004a00000000",
            INIT_23 => X"0000003b0000000000000035000000000000003b000000000000004300000000",
            INIT_24 => X"0000001e00000000000000330000000000000034000000000000003b00000000",
            INIT_25 => X"00000027000000000000002e0000000000000029000000000000001f00000000",
            INIT_26 => X"0000003d000000000000003d000000000000003b000000000000002e00000000",
            INIT_27 => X"0000003c000000000000003a0000000000000030000000000000003400000000",
            INIT_28 => X"0000005900000000000000470000000000000066000000000000006500000000",
            INIT_29 => X"0000004c000000000000004c0000000000000046000000000000005100000000",
            INIT_2A => X"00000047000000000000004e0000000000000051000000000000004c00000000",
            INIT_2B => X"0000003100000000000000350000000000000043000000000000004400000000",
            INIT_2C => X"0000003900000000000000480000000000000041000000000000004300000000",
            INIT_2D => X"000000320000000000000042000000000000003e000000000000002b00000000",
            INIT_2E => X"0000003a00000000000000380000000000000036000000000000003800000000",
            INIT_2F => X"00000041000000000000003c000000000000003d000000000000003c00000000",
            INIT_30 => X"0000006300000000000000490000000000000059000000000000007800000000",
            INIT_31 => X"0000004b00000000000000510000000000000050000000000000005300000000",
            INIT_32 => X"0000004200000000000000550000000000000057000000000000005100000000",
            INIT_33 => X"000000350000000000000043000000000000004f000000000000004c00000000",
            INIT_34 => X"0000004d000000000000004a0000000000000040000000000000003c00000000",
            INIT_35 => X"0000002f00000000000000410000000000000040000000000000004100000000",
            INIT_36 => X"00000030000000000000002d0000000000000036000000000000003500000000",
            INIT_37 => X"00000042000000000000003f000000000000003d000000000000003a00000000",
            INIT_38 => X"0000005b000000000000005b000000000000003b000000000000007500000000",
            INIT_39 => X"00000054000000000000004f0000000000000051000000000000005100000000",
            INIT_3A => X"0000004800000000000000560000000000000056000000000000005700000000",
            INIT_3B => X"0000003f000000000000004a000000000000004c000000000000004d00000000",
            INIT_3C => X"00000049000000000000004c0000000000000049000000000000004200000000",
            INIT_3D => X"0000002f0000000000000038000000000000002f000000000000004700000000",
            INIT_3E => X"0000002a00000000000000230000000000000031000000000000002c00000000",
            INIT_3F => X"00000040000000000000003e0000000000000039000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000051000000000000005b0000000000000054000000000000005c00000000",
            INIT_41 => X"000000500000000000000050000000000000004f000000000000005300000000",
            INIT_42 => X"0000004600000000000000490000000000000053000000000000005800000000",
            INIT_43 => X"0000003d00000000000000430000000000000048000000000000005100000000",
            INIT_44 => X"0000004600000000000000460000000000000041000000000000004300000000",
            INIT_45 => X"0000003c000000000000004f0000000000000040000000000000004f00000000",
            INIT_46 => X"0000003b0000000000000034000000000000002d000000000000002c00000000",
            INIT_47 => X"00000040000000000000003d000000000000003d000000000000003a00000000",
            INIT_48 => X"0000005a000000000000004c0000000000000058000000000000006100000000",
            INIT_49 => X"0000004700000000000000530000000000000056000000000000005b00000000",
            INIT_4A => X"0000005300000000000000540000000000000052000000000000004f00000000",
            INIT_4B => X"00000055000000000000004d0000000000000053000000000000005800000000",
            INIT_4C => X"000000460000000000000039000000000000003e000000000000005100000000",
            INIT_4D => X"0000004b00000000000000590000000000000048000000000000005000000000",
            INIT_4E => X"0000003c000000000000003a0000000000000031000000000000002b00000000",
            INIT_4F => X"000000400000000000000039000000000000003f000000000000003a00000000",
            INIT_50 => X"0000006200000000000000560000000000000030000000000000005100000000",
            INIT_51 => X"000000540000000000000052000000000000005b000000000000005900000000",
            INIT_52 => X"0000005000000000000000500000000000000054000000000000005b00000000",
            INIT_53 => X"0000007e00000000000000670000000000000065000000000000005e00000000",
            INIT_54 => X"0000004300000000000000370000000000000049000000000000006b00000000",
            INIT_55 => X"000000440000000000000051000000000000004c000000000000004b00000000",
            INIT_56 => X"0000002d000000000000002f0000000000000031000000000000002000000000",
            INIT_57 => X"00000041000000000000003e000000000000003a000000000000003300000000",
            INIT_58 => X"0000004d0000000000000063000000000000001f000000000000001400000000",
            INIT_59 => X"0000005a000000000000005a0000000000000056000000000000004000000000",
            INIT_5A => X"0000005f00000000000000450000000000000045000000000000005f00000000",
            INIT_5B => X"0000007900000000000000670000000000000088000000000000008f00000000",
            INIT_5C => X"00000050000000000000003f0000000000000052000000000000007600000000",
            INIT_5D => X"000000210000000000000042000000000000004d000000000000005200000000",
            INIT_5E => X"0000002e00000000000000300000000000000030000000000000002100000000",
            INIT_5F => X"0000003f000000000000003b0000000000000036000000000000003000000000",
            INIT_60 => X"0000005c00000000000000700000000000000032000000000000000000000000",
            INIT_61 => X"000000620000000000000069000000000000007a000000000000006e00000000",
            INIT_62 => X"0000007700000000000000540000000000000048000000000000006000000000",
            INIT_63 => X"00000049000000000000005f000000000000007d000000000000009d00000000",
            INIT_64 => X"0000005400000000000000410000000000000047000000000000003400000000",
            INIT_65 => X"0000002a0000000000000041000000000000004f000000000000006000000000",
            INIT_66 => X"0000002900000000000000290000000000000025000000000000002500000000",
            INIT_67 => X"0000003a00000000000000390000000000000038000000000000002d00000000",
            INIT_68 => X"0000005c0000000000000061000000000000003c000000000000001400000000",
            INIT_69 => X"0000006f00000000000000700000000000000078000000000000007d00000000",
            INIT_6A => X"00000080000000000000006e000000000000004c000000000000005900000000",
            INIT_6B => X"0000006c00000000000000620000000000000064000000000000007f00000000",
            INIT_6C => X"0000005b00000000000000620000000000000063000000000000004400000000",
            INIT_6D => X"00000029000000000000003a000000000000004c000000000000006a00000000",
            INIT_6E => X"0000002600000000000000250000000000000023000000000000002100000000",
            INIT_6F => X"0000003500000000000000320000000000000034000000000000002e00000000",
            INIT_70 => X"00000058000000000000003a0000000000000046000000000000003b00000000",
            INIT_71 => X"00000073000000000000006a0000000000000075000000000000007b00000000",
            INIT_72 => X"0000007d00000000000000820000000000000067000000000000006600000000",
            INIT_73 => X"0000008900000000000000660000000000000050000000000000005f00000000",
            INIT_74 => X"00000084000000000000007e000000000000008c000000000000008300000000",
            INIT_75 => X"0000002a0000000000000040000000000000004e000000000000006f00000000",
            INIT_76 => X"00000032000000000000002a0000000000000028000000000000002b00000000",
            INIT_77 => X"00000031000000000000002e0000000000000032000000000000002f00000000",
            INIT_78 => X"0000005e00000000000000320000000000000035000000000000004900000000",
            INIT_79 => X"00000062000000000000006c000000000000007c000000000000007e00000000",
            INIT_7A => X"00000088000000000000008a000000000000007d000000000000007200000000",
            INIT_7B => X"0000008c00000000000000710000000000000062000000000000007b00000000",
            INIT_7C => X"0000008c000000000000008a0000000000000089000000000000008f00000000",
            INIT_7D => X"0000003300000000000000490000000000000069000000000000007500000000",
            INIT_7E => X"0000004d00000000000000320000000000000023000000000000002f00000000",
            INIT_7F => X"00000032000000000000002d000000000000002d000000000000004300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE34;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE35 : if BRAM_NAME = "sampleifmap_layersamples_instance35" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000056000000000000003a0000000000000041000000000000004800000000",
            INIT_01 => X"0000005300000000000000690000000000000075000000000000007700000000",
            INIT_02 => X"0000008200000000000000930000000000000089000000000000006e00000000",
            INIT_03 => X"00000087000000000000006d000000000000006b000000000000008200000000",
            INIT_04 => X"00000083000000000000007e000000000000007f000000000000008400000000",
            INIT_05 => X"0000002a000000000000003d0000000000000077000000000000008700000000",
            INIT_06 => X"00000055000000000000003c000000000000001b000000000000001a00000000",
            INIT_07 => X"0000003300000000000000240000000000000033000000000000006100000000",
            INIT_08 => X"0000006600000000000000510000000000000048000000000000004700000000",
            INIT_09 => X"00000050000000000000007a000000000000007c000000000000007800000000",
            INIT_0A => X"00000054000000000000006a0000000000000097000000000000006300000000",
            INIT_0B => X"0000005c00000000000000650000000000000079000000000000007c00000000",
            INIT_0C => X"0000006500000000000000680000000000000073000000000000006300000000",
            INIT_0D => X"00000011000000000000001f0000000000000048000000000000005e00000000",
            INIT_0E => X"00000055000000000000003a0000000000000015000000000000000e00000000",
            INIT_0F => X"00000029000000000000001f0000000000000046000000000000006800000000",
            INIT_10 => X"000000640000000000000044000000000000004e000000000000004f00000000",
            INIT_11 => X"0000004b000000000000007d0000000000000088000000000000008600000000",
            INIT_12 => X"00000061000000000000005b0000000000000093000000000000004700000000",
            INIT_13 => X"0000004800000000000000370000000000000071000000000000008e00000000",
            INIT_14 => X"000000320000000000000045000000000000004f000000000000003500000000",
            INIT_15 => X"00000016000000000000000d0000000000000014000000000000002a00000000",
            INIT_16 => X"0000006000000000000000370000000000000023000000000000001400000000",
            INIT_17 => X"00000023000000000000001e000000000000005b000000000000006f00000000",
            INIT_18 => X"0000005800000000000000320000000000000048000000000000005100000000",
            INIT_19 => X"0000005d000000000000008a0000000000000099000000000000008700000000",
            INIT_1A => X"00000071000000000000007f000000000000006f000000000000001f00000000",
            INIT_1B => X"0000008d0000000000000047000000000000005c000000000000007c00000000",
            INIT_1C => X"0000002100000000000000330000000000000041000000000000006700000000",
            INIT_1D => X"0000002c00000000000000240000000000000019000000000000002400000000",
            INIT_1E => X"000000600000000000000036000000000000002b000000000000001a00000000",
            INIT_1F => X"0000001a000000000000001e0000000000000073000000000000008900000000",
            INIT_20 => X"0000005f000000000000004f0000000000000052000000000000005300000000",
            INIT_21 => X"0000006200000000000000860000000000000096000000000000008200000000",
            INIT_22 => X"0000006300000000000000560000000000000017000000000000000a00000000",
            INIT_23 => X"000000740000000000000042000000000000004c000000000000006500000000",
            INIT_24 => X"000000170000000000000027000000000000004e000000000000007a00000000",
            INIT_25 => X"0000002e000000000000002f000000000000002f000000000000002e00000000",
            INIT_26 => X"000000670000000000000034000000000000001b000000000000001400000000",
            INIT_27 => X"00000019000000000000002f0000000000000089000000000000009200000000",
            INIT_28 => X"00000053000000000000004e000000000000005c000000000000005c00000000",
            INIT_29 => X"00000046000000000000006e0000000000000087000000000000007b00000000",
            INIT_2A => X"0000001d00000000000000100000000000000008000000000000000c00000000",
            INIT_2B => X"0000003800000000000000250000000000000034000000000000002f00000000",
            INIT_2C => X"00000012000000000000002b0000000000000039000000000000004600000000",
            INIT_2D => X"0000002c000000000000001d000000000000001c000000000000001900000000",
            INIT_2E => X"0000005e00000000000000310000000000000026000000000000002100000000",
            INIT_2F => X"00000018000000000000003d000000000000008d000000000000008c00000000",
            INIT_30 => X"0000004e0000000000000046000000000000005d000000000000006100000000",
            INIT_31 => X"0000003000000000000000600000000000000076000000000000006b00000000",
            INIT_32 => X"000000130000000000000022000000000000003a000000000000002500000000",
            INIT_33 => X"0000003b0000000000000026000000000000001f000000000000001300000000",
            INIT_34 => X"00000012000000000000001b0000000000000013000000000000002700000000",
            INIT_35 => X"00000018000000000000000a0000000000000011000000000000001100000000",
            INIT_36 => X"000000400000000000000030000000000000002c000000000000002a00000000",
            INIT_37 => X"0000001800000000000000460000000000000080000000000000007800000000",
            INIT_38 => X"000000580000000000000052000000000000004d000000000000005e00000000",
            INIT_39 => X"0000004b000000000000005f000000000000006b000000000000005b00000000",
            INIT_3A => X"0000003900000000000000300000000000000037000000000000004a00000000",
            INIT_3B => X"0000003300000000000000430000000000000035000000000000003a00000000",
            INIT_3C => X"0000000800000000000000030000000000000004000000000000001000000000",
            INIT_3D => X"0000000600000000000000070000000000000013000000000000000e00000000",
            INIT_3E => X"0000002f00000000000000300000000000000017000000000000001100000000",
            INIT_3F => X"0000001b00000000000000570000000000000073000000000000005100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000690000000000000057000000000000003b000000000000004b00000000",
            INIT_41 => X"0000007e00000000000000750000000000000052000000000000005300000000",
            INIT_42 => X"0000003e00000000000000390000000000000022000000000000005500000000",
            INIT_43 => X"0000002e0000000000000039000000000000003d000000000000004200000000",
            INIT_44 => X"0000000d00000000000000120000000000000017000000000000002400000000",
            INIT_45 => X"0000000e000000000000000c000000000000000e000000000000000f00000000",
            INIT_46 => X"0000001e0000000000000036000000000000001c000000000000000700000000",
            INIT_47 => X"0000003e00000000000000680000000000000055000000000000002800000000",
            INIT_48 => X"000000560000000000000051000000000000004d000000000000004d00000000",
            INIT_49 => X"0000007000000000000000570000000000000045000000000000005500000000",
            INIT_4A => X"0000004f0000000000000064000000000000004f000000000000006f00000000",
            INIT_4B => X"0000003a00000000000000450000000000000043000000000000003b00000000",
            INIT_4C => X"0000001500000000000000200000000000000026000000000000003300000000",
            INIT_4D => X"0000000e0000000000000006000000000000000c000000000000001100000000",
            INIT_4E => X"0000000f00000000000000290000000000000022000000000000000f00000000",
            INIT_4F => X"0000005a000000000000004c000000000000002e000000000000001f00000000",
            INIT_50 => X"0000005500000000000000520000000000000051000000000000004f00000000",
            INIT_51 => X"00000039000000000000004a0000000000000060000000000000006500000000",
            INIT_52 => X"0000003e000000000000003a0000000000000057000000000000006d00000000",
            INIT_53 => X"00000044000000000000005a0000000000000058000000000000003d00000000",
            INIT_54 => X"0000002a000000000000002f0000000000000035000000000000003b00000000",
            INIT_55 => X"0000002300000000000000180000000000000023000000000000002c00000000",
            INIT_56 => X"0000001f000000000000001b000000000000001d000000000000002600000000",
            INIT_57 => X"0000003800000000000000270000000000000052000000000000003900000000",
            INIT_58 => X"0000004a000000000000004a0000000000000057000000000000004c00000000",
            INIT_59 => X"000000390000000000000053000000000000005f000000000000006600000000",
            INIT_5A => X"0000003a00000000000000370000000000000063000000000000004d00000000",
            INIT_5B => X"0000004d00000000000000570000000000000054000000000000003f00000000",
            INIT_5C => X"000000440000000000000043000000000000003c000000000000003900000000",
            INIT_5D => X"0000003f00000000000000310000000000000031000000000000003b00000000",
            INIT_5E => X"0000003300000000000000300000000000000031000000000000003c00000000",
            INIT_5F => X"0000002f000000000000002d0000000000000054000000000000003f00000000",
            INIT_60 => X"000000450000000000000040000000000000005a000000000000005500000000",
            INIT_61 => X"000000440000000000000041000000000000004e000000000000005e00000000",
            INIT_62 => X"0000005a0000000000000042000000000000003c000000000000004c00000000",
            INIT_63 => X"000000510000000000000053000000000000004e000000000000004a00000000",
            INIT_64 => X"00000040000000000000004c0000000000000047000000000000004300000000",
            INIT_65 => X"00000048000000000000003e0000000000000039000000000000003b00000000",
            INIT_66 => X"0000003e00000000000000400000000000000042000000000000004400000000",
            INIT_67 => X"00000053000000000000003d0000000000000029000000000000003200000000",
            INIT_68 => X"0000005c0000000000000049000000000000004b000000000000003d00000000",
            INIT_69 => X"00000050000000000000004e0000000000000051000000000000005700000000",
            INIT_6A => X"000000590000000000000050000000000000004c000000000000005d00000000",
            INIT_6B => X"00000050000000000000004e000000000000004c000000000000004a00000000",
            INIT_6C => X"00000035000000000000003e0000000000000045000000000000004a00000000",
            INIT_6D => X"0000004b00000000000000440000000000000042000000000000004000000000",
            INIT_6E => X"0000004400000000000000480000000000000048000000000000004d00000000",
            INIT_6F => X"00000059000000000000004e0000000000000038000000000000003200000000",
            INIT_70 => X"00000064000000000000005a0000000000000051000000000000004600000000",
            INIT_71 => X"0000005500000000000000570000000000000055000000000000005600000000",
            INIT_72 => X"0000005a000000000000005d0000000000000057000000000000005600000000",
            INIT_73 => X"0000003c000000000000003f0000000000000046000000000000004a00000000",
            INIT_74 => X"0000003e000000000000003e000000000000003c000000000000004200000000",
            INIT_75 => X"0000004c00000000000000470000000000000046000000000000004100000000",
            INIT_76 => X"00000047000000000000004e000000000000004d000000000000005500000000",
            INIT_77 => X"0000004f000000000000004d0000000000000041000000000000003e00000000",
            INIT_78 => X"00000059000000000000005f000000000000005d000000000000004f00000000",
            INIT_79 => X"0000005100000000000000460000000000000039000000000000004600000000",
            INIT_7A => X"0000004700000000000000470000000000000040000000000000005300000000",
            INIT_7B => X"0000002f000000000000003d000000000000004c000000000000004a00000000",
            INIT_7C => X"000000460000000000000048000000000000003f000000000000003800000000",
            INIT_7D => X"00000050000000000000004b000000000000004c000000000000004500000000",
            INIT_7E => X"0000004e0000000000000049000000000000004f000000000000005600000000",
            INIT_7F => X"00000049000000000000004f000000000000004c000000000000004f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE35;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE36 : if BRAM_NAME = "sampleifmap_layersamples_instance36" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d900000000000000d100000000000000b900000000000000a000000000",
            INIT_01 => X"000000f600000000000000f900000000000000f600000000000000e600000000",
            INIT_02 => X"000000dd00000000000000e600000000000000f300000000000000f800000000",
            INIT_03 => X"000000c700000000000000d800000000000000dd00000000000000da00000000",
            INIT_04 => X"000000b400000000000000b800000000000000bb00000000000000bc00000000",
            INIT_05 => X"0000008b0000000000000079000000000000009000000000000000a600000000",
            INIT_06 => X"0000004f00000000000000660000000000000066000000000000006a00000000",
            INIT_07 => X"0000005e000000000000005b0000000000000065000000000000005e00000000",
            INIT_08 => X"000000e600000000000000f200000000000000ef00000000000000e100000000",
            INIT_09 => X"000000eb00000000000000f300000000000000f500000000000000e800000000",
            INIT_0A => X"000000cd00000000000000d800000000000000e600000000000000ed00000000",
            INIT_0B => X"000000ba00000000000000c800000000000000cb00000000000000c900000000",
            INIT_0C => X"0000007f00000000000000a100000000000000ab00000000000000af00000000",
            INIT_0D => X"00000087000000000000007a000000000000008d000000000000008e00000000",
            INIT_0E => X"0000003400000000000000250000000000000052000000000000007600000000",
            INIT_0F => X"000000640000000000000061000000000000006b000000000000005f00000000",
            INIT_10 => X"000000dc00000000000000f100000000000000f900000000000000fc00000000",
            INIT_11 => X"000000d600000000000000df00000000000000e200000000000000d900000000",
            INIT_12 => X"000000b800000000000000c300000000000000cf00000000000000d500000000",
            INIT_13 => X"000000a700000000000000b300000000000000b600000000000000b300000000",
            INIT_14 => X"0000008100000000000000940000000000000098000000000000009f00000000",
            INIT_15 => X"000000720000000000000080000000000000008c000000000000008000000000",
            INIT_16 => X"0000002600000000000000040000000000000028000000000000005700000000",
            INIT_17 => X"0000006900000000000000690000000000000073000000000000006300000000",
            INIT_18 => X"000000d300000000000000de00000000000000e100000000000000e900000000",
            INIT_19 => X"000000c000000000000000c800000000000000cb00000000000000d300000000",
            INIT_1A => X"000000a400000000000000ae00000000000000b700000000000000bb00000000",
            INIT_1B => X"0000009900000000000000a000000000000000a500000000000000a000000000",
            INIT_1C => X"0000008a000000000000008c000000000000008d000000000000009100000000",
            INIT_1D => X"00000069000000000000007f000000000000007d000000000000007d00000000",
            INIT_1E => X"00000037000000000000001a0000000000000025000000000000003b00000000",
            INIT_1F => X"0000006d00000000000000700000000000000078000000000000007000000000",
            INIT_20 => X"000000c900000000000000cf00000000000000c300000000000000cf00000000",
            INIT_21 => X"000000ab00000000000000b300000000000000b400000000000000be00000000",
            INIT_22 => X"000000920000000000000099000000000000009f00000000000000a300000000",
            INIT_23 => X"0000008d00000000000000930000000000000097000000000000009100000000",
            INIT_24 => X"0000008700000000000000830000000000000088000000000000008700000000",
            INIT_25 => X"0000005a0000000000000084000000000000007a000000000000008100000000",
            INIT_26 => X"000000560000000000000030000000000000003d000000000000003a00000000",
            INIT_27 => X"0000006d00000000000000720000000000000078000000000000007500000000",
            INIT_28 => X"000000a200000000000000aa00000000000000ab00000000000000b600000000",
            INIT_29 => X"00000097000000000000009f000000000000009c000000000000009900000000",
            INIT_2A => X"0000008a000000000000008c000000000000008d000000000000009000000000",
            INIT_2B => X"0000008a000000000000008a000000000000008d000000000000008b00000000",
            INIT_2C => X"0000008a0000000000000086000000000000008c000000000000008700000000",
            INIT_2D => X"0000004500000000000000660000000000000089000000000000008c00000000",
            INIT_2E => X"000000740000000000000043000000000000003e000000000000004b00000000",
            INIT_2F => X"0000006e00000000000000700000000000000080000000000000008100000000",
            INIT_30 => X"0000008600000000000000880000000000000088000000000000008d00000000",
            INIT_31 => X"00000085000000000000008c0000000000000086000000000000008800000000",
            INIT_32 => X"0000008d000000000000008b0000000000000089000000000000008700000000",
            INIT_33 => X"00000091000000000000008e0000000000000092000000000000008f00000000",
            INIT_34 => X"0000008f000000000000008a0000000000000091000000000000009100000000",
            INIT_35 => X"00000021000000000000002f000000000000006b000000000000008e00000000",
            INIT_36 => X"0000007f000000000000006c000000000000004b000000000000004800000000",
            INIT_37 => X"00000070000000000000006f0000000000000084000000000000008400000000",
            INIT_38 => X"000000810000000000000080000000000000007d000000000000007600000000",
            INIT_39 => X"00000084000000000000008a0000000000000083000000000000008800000000",
            INIT_3A => X"000000930000000000000090000000000000008c000000000000008800000000",
            INIT_3B => X"00000099000000000000009a000000000000009e000000000000009600000000",
            INIT_3C => X"0000009400000000000000930000000000000095000000000000009200000000",
            INIT_3D => X"00000011000000000000000d0000000000000042000000000000008000000000",
            INIT_3E => X"0000007a00000000000000800000000000000075000000000000005000000000",
            INIT_3F => X"0000007000000000000000720000000000000080000000000000007b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000850000000000000084000000000000007e000000000000007300000000",
            INIT_41 => X"00000089000000000000008f0000000000000087000000000000008b00000000",
            INIT_42 => X"0000009800000000000000950000000000000091000000000000008b00000000",
            INIT_43 => X"000000aa00000000000000a3000000000000009a000000000000009400000000",
            INIT_44 => X"00000094000000000000009d00000000000000a2000000000000009e00000000",
            INIT_45 => X"0000001e000000000000000e000000000000002c000000000000007300000000",
            INIT_46 => X"0000007e0000000000000088000000000000008b000000000000006900000000",
            INIT_47 => X"0000006f0000000000000074000000000000007a000000000000007700000000",
            INIT_48 => X"0000008800000000000000880000000000000080000000000000007600000000",
            INIT_49 => X"0000008d00000000000000910000000000000088000000000000008d00000000",
            INIT_4A => X"000000a5000000000000009a0000000000000093000000000000008d00000000",
            INIT_4B => X"000000a700000000000000a2000000000000009a000000000000009d00000000",
            INIT_4C => X"0000008a00000000000000910000000000000093000000000000009b00000000",
            INIT_4D => X"00000037000000000000002e0000000000000038000000000000006300000000",
            INIT_4E => X"0000007e000000000000007a000000000000007c000000000000006d00000000",
            INIT_4F => X"0000006e00000000000000750000000000000074000000000000007300000000",
            INIT_50 => X"00000089000000000000008b0000000000000084000000000000007d00000000",
            INIT_51 => X"0000008c00000000000000900000000000000088000000000000008e00000000",
            INIT_52 => X"0000009900000000000000960000000000000090000000000000008b00000000",
            INIT_53 => X"000000980000000000000090000000000000008b000000000000008300000000",
            INIT_54 => X"000000d600000000000000d300000000000000ba00000000000000a600000000",
            INIT_55 => X"0000002a0000000000000045000000000000005c000000000000008000000000",
            INIT_56 => X"000000730000000000000063000000000000005f000000000000005500000000",
            INIT_57 => X"0000006b0000000000000071000000000000006f000000000000007000000000",
            INIT_58 => X"0000008a000000000000008e0000000000000089000000000000008500000000",
            INIT_59 => X"0000008a000000000000008e0000000000000088000000000000008d00000000",
            INIT_5A => X"000000840000000000000088000000000000008f000000000000008900000000",
            INIT_5B => X"000000cb00000000000000c900000000000000b6000000000000008e00000000",
            INIT_5C => X"000000c000000000000000cf00000000000000ce00000000000000d200000000",
            INIT_5D => X"0000002a000000000000009200000000000000bd00000000000000a200000000",
            INIT_5E => X"0000007200000000000000670000000000000028000000000000001b00000000",
            INIT_5F => X"00000068000000000000006c000000000000006a000000000000006d00000000",
            INIT_60 => X"0000008b000000000000008f000000000000008b000000000000008c00000000",
            INIT_61 => X"00000089000000000000008a000000000000008c000000000000008f00000000",
            INIT_62 => X"000000a400000000000000900000000000000085000000000000008700000000",
            INIT_63 => X"00000073000000000000008900000000000000a000000000000000ab00000000",
            INIT_64 => X"0000003b000000000000004b000000000000005d000000000000006a00000000",
            INIT_65 => X"0000005f00000000000000c900000000000000dc000000000000006f00000000",
            INIT_66 => X"00000074000000000000003e0000000000000007000000000000000d00000000",
            INIT_67 => X"0000006400000000000000690000000000000065000000000000006300000000",
            INIT_68 => X"0000008c000000000000008f000000000000008a000000000000009000000000",
            INIT_69 => X"0000008700000000000000820000000000000092000000000000009200000000",
            INIT_6A => X"0000006e000000000000008c0000000000000091000000000000008200000000",
            INIT_6B => X"000000130000000000000031000000000000005c000000000000005e00000000",
            INIT_6C => X"0000001200000000000000190000000000000032000000000000001d00000000",
            INIT_6D => X"0000009d00000000000000d200000000000000d1000000000000007800000000",
            INIT_6E => X"0000004400000000000000130000000000000006000000000000002600000000",
            INIT_6F => X"0000005f00000000000000630000000000000052000000000000004500000000",
            INIT_70 => X"0000008e0000000000000092000000000000008b000000000000009100000000",
            INIT_71 => X"000000800000000000000079000000000000008e000000000000009000000000",
            INIT_72 => X"000000440000000000000054000000000000007f000000000000008500000000",
            INIT_73 => X"00000016000000000000002e0000000000000052000000000000005600000000",
            INIT_74 => X"00000041000000000000001e0000000000000032000000000000001300000000",
            INIT_75 => X"000000cb00000000000000cd00000000000000c900000000000000af00000000",
            INIT_76 => X"0000001600000000000000120000000000000010000000000000006600000000",
            INIT_77 => X"00000058000000000000004f0000000000000038000000000000002300000000",
            INIT_78 => X"000000900000000000000094000000000000008b000000000000008f00000000",
            INIT_79 => X"00000083000000000000008b0000000000000084000000000000008a00000000",
            INIT_7A => X"0000005600000000000000480000000000000042000000000000007500000000",
            INIT_7B => X"000000220000000000000028000000000000004e000000000000006a00000000",
            INIT_7C => X"000000b600000000000000730000000000000046000000000000002400000000",
            INIT_7D => X"000000c300000000000000cd00000000000000c500000000000000cb00000000",
            INIT_7E => X"000000120000000000000025000000000000003d000000000000006c00000000",
            INIT_7F => X"000000530000000000000064000000000000004f000000000000001800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE36;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE37 : if BRAM_NAME = "sampleifmap_layersamples_instance37" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000900000000000000093000000000000008b000000000000008e00000000",
            INIT_01 => X"0000007900000000000000840000000000000072000000000000008500000000",
            INIT_02 => X"00000045000000000000003c0000000000000059000000000000005100000000",
            INIT_03 => X"0000009b00000000000000530000000000000044000000000000005500000000",
            INIT_04 => X"000000eb00000000000000ed00000000000000db00000000000000c000000000",
            INIT_05 => X"0000007200000000000000d300000000000000d700000000000000d700000000",
            INIT_06 => X"000000140000000000000035000000000000005d000000000000003000000000",
            INIT_07 => X"00000054000000000000008f000000000000008b000000000000004100000000",
            INIT_08 => X"00000089000000000000008e000000000000008d000000000000008f00000000",
            INIT_09 => X"00000043000000000000003a0000000000000045000000000000007400000000",
            INIT_0A => X"0000001c000000000000001d000000000000004b000000000000005100000000",
            INIT_0B => X"000000f2000000000000008c0000000000000019000000000000002400000000",
            INIT_0C => X"000000dc00000000000000e300000000000000eb00000000000000ec00000000",
            INIT_0D => X"0000003a000000000000009500000000000000df00000000000000db00000000",
            INIT_0E => X"0000004e000000000000004e0000000000000054000000000000003900000000",
            INIT_0F => X"0000005b00000000000000a700000000000000a1000000000000008500000000",
            INIT_10 => X"000000860000000000000088000000000000008c000000000000008f00000000",
            INIT_11 => X"00000034000000000000002d0000000000000047000000000000008d00000000",
            INIT_12 => X"0000001600000000000000170000000000000021000000000000004300000000",
            INIT_13 => X"000000d9000000000000009b0000000000000029000000000000002f00000000",
            INIT_14 => X"000000d000000000000000bf00000000000000be00000000000000c700000000",
            INIT_15 => X"0000006700000000000000ad00000000000000df00000000000000dc00000000",
            INIT_16 => X"0000009500000000000000870000000000000073000000000000005d00000000",
            INIT_17 => X"0000005900000000000000a50000000000000094000000000000009800000000",
            INIT_18 => X"000000b5000000000000007e000000000000008c000000000000008f00000000",
            INIT_19 => X"0000002b0000000000000021000000000000004c00000000000000bd00000000",
            INIT_1A => X"0000001700000000000000100000000000000015000000000000003900000000",
            INIT_1B => X"000000c2000000000000009e0000000000000042000000000000003900000000",
            INIT_1C => X"000000c900000000000000c400000000000000b300000000000000b600000000",
            INIT_1D => X"000000b300000000000000de00000000000000ce00000000000000c200000000",
            INIT_1E => X"000000970000000000000095000000000000009c000000000000009700000000",
            INIT_1F => X"0000004200000000000000880000000000000092000000000000009600000000",
            INIT_20 => X"000000ea000000000000009a0000000000000085000000000000008c00000000",
            INIT_21 => X"0000002a0000000000000026000000000000005a00000000000000b500000000",
            INIT_22 => X"0000000b000000000000000b000000000000000b000000000000003400000000",
            INIT_23 => X"000000ba00000000000000a00000000000000031000000000000001400000000",
            INIT_24 => X"0000007300000000000000b900000000000000b900000000000000b000000000",
            INIT_25 => X"000000c400000000000000a1000000000000005a000000000000004500000000",
            INIT_26 => X"0000009900000000000000a000000000000000aa00000000000000b700000000",
            INIT_27 => X"00000026000000000000004d0000000000000088000000000000009300000000",
            INIT_28 => X"000000a300000000000000a30000000000000080000000000000008200000000",
            INIT_29 => X"0000002e000000000000002d000000000000006a000000000000008b00000000",
            INIT_2A => X"0000000f00000000000000090000000000000003000000000000001c00000000",
            INIT_2B => X"000000b400000000000000a20000000000000036000000000000001e00000000",
            INIT_2C => X"00000015000000000000007100000000000000be00000000000000ac00000000",
            INIT_2D => X"0000009500000000000000300000000000000015000000000000001400000000",
            INIT_2E => X"00000085000000000000008e00000000000000ab00000000000000bb00000000",
            INIT_2F => X"0000002700000000000000150000000000000043000000000000008000000000",
            INIT_30 => X"0000001a00000000000000670000000000000084000000000000007c00000000",
            INIT_31 => X"000000300000000000000034000000000000006c000000000000004800000000",
            INIT_32 => X"0000003b000000000000000b0000000000000007000000000000001200000000",
            INIT_33 => X"000000b000000000000000a50000000000000063000000000000005a00000000",
            INIT_34 => X"0000001d000000000000002a00000000000000a900000000000000b100000000",
            INIT_35 => X"00000046000000000000000e0000000000000026000000000000002f00000000",
            INIT_36 => X"0000007500000000000000750000000000000088000000000000009500000000",
            INIT_37 => X"000000300000000000000015000000000000000e000000000000003c00000000",
            INIT_38 => X"0000001e0000000000000049000000000000007c000000000000007900000000",
            INIT_39 => X"0000001f00000000000000440000000000000072000000000000003b00000000",
            INIT_3A => X"000000480000000000000018000000000000000e000000000000000d00000000",
            INIT_3B => X"000000bb00000000000000bb000000000000006c000000000000004f00000000",
            INIT_3C => X"0000002b000000000000001b000000000000008b00000000000000bf00000000",
            INIT_3D => X"0000001b000000000000001c000000000000001b000000000000001e00000000",
            INIT_3E => X"00000059000000000000007b0000000000000084000000000000006c00000000",
            INIT_3F => X"0000003b000000000000002a0000000000000015000000000000001600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003f00000000000000470000000000000066000000000000006d00000000",
            INIT_41 => X"0000001c000000000000004d0000000000000071000000000000003c00000000",
            INIT_42 => X"000000470000000000000030000000000000001f000000000000001000000000",
            INIT_43 => X"000000b300000000000000bd0000000000000088000000000000004600000000",
            INIT_44 => X"00000036000000000000001f000000000000007400000000000000b400000000",
            INIT_45 => X"0000000e000000000000001b0000000000000029000000000000003500000000",
            INIT_46 => X"0000003c000000000000007c0000000000000085000000000000004800000000",
            INIT_47 => X"0000003b00000000000000320000000000000022000000000000001200000000",
            INIT_48 => X"0000003c000000000000003d0000000000000051000000000000005700000000",
            INIT_49 => X"00000015000000000000004b0000000000000069000000000000003a00000000",
            INIT_4A => X"00000060000000000000004c000000000000002e000000000000001400000000",
            INIT_4B => X"000000a300000000000000a40000000000000091000000000000006100000000",
            INIT_4C => X"000000390000000000000020000000000000007100000000000000aa00000000",
            INIT_4D => X"0000001100000000000000250000000000000031000000000000004700000000",
            INIT_4E => X"000000210000000000000060000000000000006c000000000000002900000000",
            INIT_4F => X"000000320000000000000028000000000000001d000000000000000c00000000",
            INIT_50 => X"0000003c00000000000000400000000000000049000000000000004900000000",
            INIT_51 => X"0000002f0000000000000057000000000000005f000000000000003900000000",
            INIT_52 => X"000000a500000000000000890000000000000062000000000000003d00000000",
            INIT_53 => X"000000b600000000000000b700000000000000b000000000000000a900000000",
            INIT_54 => X"000000360000000000000022000000000000007c00000000000000b600000000",
            INIT_55 => X"0000001b0000000000000033000000000000005c000000000000006000000000",
            INIT_56 => X"0000000c000000000000003b0000000000000046000000000000001100000000",
            INIT_57 => X"00000028000000000000001d0000000000000012000000000000000600000000",
            INIT_58 => X"0000004e00000000000000450000000000000049000000000000004900000000",
            INIT_59 => X"0000002f00000000000000450000000000000059000000000000004100000000",
            INIT_5A => X"00000056000000000000004a000000000000003c000000000000003400000000",
            INIT_5B => X"0000006000000000000000620000000000000060000000000000005b00000000",
            INIT_5C => X"0000003c00000000000000200000000000000053000000000000006200000000",
            INIT_5D => X"00000014000000000000001d000000000000003e000000000000003b00000000",
            INIT_5E => X"00000003000000000000000a0000000000000011000000000000000400000000",
            INIT_5F => X"000000210000000000000011000000000000000a000000000000000700000000",
            INIT_60 => X"0000003600000000000000480000000000000053000000000000004b00000000",
            INIT_61 => X"00000004000000000000000f0000000000000027000000000000002d00000000",
            INIT_62 => X"0000000700000000000000050000000000000002000000000000000300000000",
            INIT_63 => X"0000000b000000000000000a0000000000000008000000000000000700000000",
            INIT_64 => X"000000420000000000000008000000000000000d000000000000000b00000000",
            INIT_65 => X"0000000f0000000000000038000000000000002f000000000000004300000000",
            INIT_66 => X"0000000300000000000000010000000000000002000000000000000200000000",
            INIT_67 => X"00000020000000000000000f000000000000000a000000000000000600000000",
            INIT_68 => X"0000002f00000000000000510000000000000059000000000000005000000000",
            INIT_69 => X"000000190000000000000010000000000000000a000000000000001500000000",
            INIT_6A => X"0000000e000000000000000e000000000000000a000000000000000e00000000",
            INIT_6B => X"0000000c000000000000000e000000000000000e000000000000000e00000000",
            INIT_6C => X"0000001700000000000000060000000000000009000000000000000a00000000",
            INIT_6D => X"00000007000000000000002a0000000000000048000000000000003e00000000",
            INIT_6E => X"0000000500000000000000050000000000000004000000000000000300000000",
            INIT_6F => X"000000210000000000000015000000000000000b000000000000000700000000",
            INIT_70 => X"000000370000000000000049000000000000004f000000000000004900000000",
            INIT_71 => X"0000003a000000000000003b000000000000002f000000000000002e00000000",
            INIT_72 => X"0000001c00000000000000190000000000000011000000000000001a00000000",
            INIT_73 => X"0000001c000000000000001d0000000000000020000000000000001f00000000",
            INIT_74 => X"0000000c00000000000000100000000000000015000000000000001800000000",
            INIT_75 => X"0000000600000000000000080000000000000016000000000000001400000000",
            INIT_76 => X"0000000800000000000000080000000000000007000000000000000800000000",
            INIT_77 => X"0000001f000000000000001b000000000000000f000000000000000b00000000",
            INIT_78 => X"0000004e000000000000004c0000000000000048000000000000004500000000",
            INIT_79 => X"0000003800000000000000480000000000000053000000000000005800000000",
            INIT_7A => X"0000002a000000000000002b0000000000000026000000000000002000000000",
            INIT_7B => X"0000003100000000000000320000000000000033000000000000002f00000000",
            INIT_7C => X"0000001c000000000000001e0000000000000026000000000000002c00000000",
            INIT_7D => X"0000000c00000000000000130000000000000022000000000000002200000000",
            INIT_7E => X"0000000d000000000000000f0000000000000010000000000000000e00000000",
            INIT_7F => X"0000001d000000000000001e000000000000001a000000000000001200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE37;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE38 : if BRAM_NAME = "sampleifmap_layersamples_instance38" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003a00000000000000390000000000000031000000000000002500000000",
            INIT_01 => X"000000510000000000000050000000000000004e000000000000004200000000",
            INIT_02 => X"0000004200000000000000490000000000000052000000000000005600000000",
            INIT_03 => X"0000003800000000000000430000000000000043000000000000004100000000",
            INIT_04 => X"0000007300000000000000400000000000000032000000000000003200000000",
            INIT_05 => X"0000002700000000000000320000000000000038000000000000003400000000",
            INIT_06 => X"00000024000000000000002e0000000000000022000000000000001600000000",
            INIT_07 => X"0000001300000000000000150000000000000012000000000000001d00000000",
            INIT_08 => X"00000044000000000000004d0000000000000048000000000000004300000000",
            INIT_09 => X"000000420000000000000048000000000000004a000000000000004300000000",
            INIT_0A => X"0000003400000000000000390000000000000040000000000000004400000000",
            INIT_0B => X"0000002e00000000000000370000000000000036000000000000003200000000",
            INIT_0C => X"000000290000000000000027000000000000002a000000000000002900000000",
            INIT_0D => X"00000021000000000000001e0000000000000023000000000000002800000000",
            INIT_0E => X"0000001b000000000000001e000000000000002e000000000000002200000000",
            INIT_0F => X"0000001200000000000000160000000000000015000000000000001c00000000",
            INIT_10 => X"0000003e00000000000000480000000000000044000000000000004800000000",
            INIT_11 => X"000000310000000000000038000000000000003d000000000000003a00000000",
            INIT_12 => X"00000028000000000000002b000000000000002d000000000000003000000000",
            INIT_13 => X"00000026000000000000002b000000000000002a000000000000002600000000",
            INIT_14 => X"0000001c000000000000001e0000000000000023000000000000002200000000",
            INIT_15 => X"00000022000000000000001f0000000000000021000000000000002300000000",
            INIT_16 => X"0000000e000000000000000d0000000000000022000000000000003000000000",
            INIT_17 => X"0000001100000000000000130000000000000014000000000000001500000000",
            INIT_18 => X"0000003c000000000000003d0000000000000036000000000000003800000000",
            INIT_19 => X"00000024000000000000002b0000000000000030000000000000003e00000000",
            INIT_1A => X"0000002000000000000000220000000000000023000000000000002300000000",
            INIT_1B => X"0000002000000000000000220000000000000021000000000000001f00000000",
            INIT_1C => X"0000001d000000000000001b000000000000001e000000000000001d00000000",
            INIT_1D => X"00000025000000000000001d000000000000001c000000000000002000000000",
            INIT_1E => X"0000000f000000000000000b0000000000000012000000000000002a00000000",
            INIT_1F => X"0000001100000000000000100000000000000013000000000000001600000000",
            INIT_20 => X"0000003b00000000000000420000000000000039000000000000003900000000",
            INIT_21 => X"0000001b00000000000000200000000000000024000000000000003400000000",
            INIT_22 => X"0000001a000000000000001c000000000000001d000000000000001c00000000",
            INIT_23 => X"0000001e000000000000001c000000000000001a000000000000001a00000000",
            INIT_24 => X"0000001c000000000000001c000000000000001c000000000000001c00000000",
            INIT_25 => X"0000002a00000000000000430000000000000030000000000000001c00000000",
            INIT_26 => X"00000019000000000000000d0000000000000012000000000000001900000000",
            INIT_27 => X"000000110000000000000013000000000000001f000000000000001b00000000",
            INIT_28 => X"00000021000000000000002f000000000000003a000000000000003b00000000",
            INIT_29 => X"000000160000000000000019000000000000001a000000000000001a00000000",
            INIT_2A => X"00000019000000000000001a0000000000000019000000000000001700000000",
            INIT_2B => X"0000001f000000000000001b0000000000000018000000000000001800000000",
            INIT_2C => X"0000001e0000000000000021000000000000001e000000000000001d00000000",
            INIT_2D => X"0000003c000000000000005e000000000000005d000000000000002100000000",
            INIT_2E => X"0000002c000000000000001e000000000000001b000000000000002900000000",
            INIT_2F => X"000000130000000000000018000000000000002d000000000000002b00000000",
            INIT_30 => X"000000140000000000000017000000000000001c000000000000002200000000",
            INIT_31 => X"0000001500000000000000160000000000000017000000000000001600000000",
            INIT_32 => X"0000001a00000000000000190000000000000016000000000000001600000000",
            INIT_33 => X"00000023000000000000001d0000000000000019000000000000001800000000",
            INIT_34 => X"0000001e0000000000000023000000000000001f000000000000002000000000",
            INIT_35 => X"0000002500000000000000370000000000000059000000000000003300000000",
            INIT_36 => X"0000002d000000000000002b0000000000000028000000000000003800000000",
            INIT_37 => X"000000150000000000000017000000000000001e000000000000002400000000",
            INIT_38 => X"0000001200000000000000100000000000000011000000000000001100000000",
            INIT_39 => X"0000001600000000000000160000000000000017000000000000001600000000",
            INIT_3A => X"0000001b000000000000001a0000000000000017000000000000001800000000",
            INIT_3B => X"00000027000000000000001d000000000000001b000000000000001900000000",
            INIT_3C => X"000000300000000000000033000000000000002d000000000000002800000000",
            INIT_3D => X"0000000b00000000000000120000000000000040000000000000004100000000",
            INIT_3E => X"00000020000000000000001f0000000000000025000000000000002200000000",
            INIT_3F => X"0000001500000000000000160000000000000016000000000000001900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001200000000000000120000000000000012000000000000001100000000",
            INIT_41 => X"0000001700000000000000170000000000000016000000000000001500000000",
            INIT_42 => X"0000001e000000000000001c0000000000000018000000000000001900000000",
            INIT_43 => X"0000003b00000000000000330000000000000038000000000000002500000000",
            INIT_44 => X"000000360000000000000037000000000000003a000000000000003b00000000",
            INIT_45 => X"0000001000000000000000110000000000000028000000000000003d00000000",
            INIT_46 => X"0000001b00000000000000180000000000000019000000000000001a00000000",
            INIT_47 => X"0000001400000000000000150000000000000017000000000000001a00000000",
            INIT_48 => X"0000001200000000000000120000000000000012000000000000001300000000",
            INIT_49 => X"0000001800000000000000160000000000000014000000000000001500000000",
            INIT_4A => X"0000003100000000000000200000000000000019000000000000001800000000",
            INIT_4B => X"000000340000000000000039000000000000004c000000000000003e00000000",
            INIT_4C => X"0000003a0000000000000032000000000000002e000000000000003100000000",
            INIT_4D => X"0000002c00000000000000300000000000000031000000000000003800000000",
            INIT_4E => X"0000001900000000000000190000000000000023000000000000002900000000",
            INIT_4F => X"0000001400000000000000140000000000000018000000000000001900000000",
            INIT_50 => X"0000001200000000000000130000000000000012000000000000001400000000",
            INIT_51 => X"0000001700000000000000150000000000000015000000000000001500000000",
            INIT_52 => X"0000003500000000000000240000000000000019000000000000001900000000",
            INIT_53 => X"0000004a000000000000003e0000000000000042000000000000003100000000",
            INIT_54 => X"000000b800000000000000a60000000000000089000000000000006800000000",
            INIT_55 => X"00000021000000000000004b0000000000000068000000000000007c00000000",
            INIT_56 => X"000000190000000000000026000000000000003d000000000000003800000000",
            INIT_57 => X"0000001300000000000000120000000000000019000000000000001800000000",
            INIT_58 => X"0000001300000000000000140000000000000012000000000000001500000000",
            INIT_59 => X"0000001800000000000000160000000000000018000000000000001800000000",
            INIT_5A => X"00000030000000000000001f000000000000001d000000000000001900000000",
            INIT_5B => X"000000be00000000000000b20000000000000097000000000000005500000000",
            INIT_5C => X"000000c500000000000000ca00000000000000cd00000000000000cd00000000",
            INIT_5D => X"00000016000000000000009800000000000000d000000000000000b200000000",
            INIT_5E => X"0000002800000000000000460000000000000025000000000000001800000000",
            INIT_5F => X"0000001100000000000000110000000000000016000000000000001500000000",
            INIT_60 => X"0000001500000000000000160000000000000014000000000000001400000000",
            INIT_61 => X"0000001a00000000000000190000000000000018000000000000001800000000",
            INIT_62 => X"0000007000000000000000420000000000000020000000000000001900000000",
            INIT_63 => X"00000075000000000000008c000000000000009b000000000000009000000000",
            INIT_64 => X"0000003d00000000000000470000000000000058000000000000006400000000",
            INIT_65 => X"0000004e00000000000000d500000000000000e8000000000000007500000000",
            INIT_66 => X"000000460000000000000032000000000000000a000000000000000f00000000",
            INIT_67 => X"0000001000000000000000110000000000000015000000000000001a00000000",
            INIT_68 => X"0000001600000000000000190000000000000016000000000000001400000000",
            INIT_69 => X"0000001a00000000000000190000000000000017000000000000001700000000",
            INIT_6A => X"0000005b00000000000000670000000000000048000000000000001a00000000",
            INIT_6B => X"0000001200000000000000340000000000000056000000000000005000000000",
            INIT_6C => X"00000010000000000000000f0000000000000022000000000000001100000000",
            INIT_6D => X"0000009b00000000000000e000000000000000dd000000000000007c00000000",
            INIT_6E => X"0000003b00000000000000160000000000000007000000000000002400000000",
            INIT_6F => X"0000001000000000000000120000000000000013000000000000002100000000",
            INIT_70 => X"00000016000000000000001b0000000000000017000000000000001800000000",
            INIT_71 => X"0000001500000000000000130000000000000019000000000000001800000000",
            INIT_72 => X"00000029000000000000003a0000000000000055000000000000003700000000",
            INIT_73 => X"000000180000000000000032000000000000004e000000000000003d00000000",
            INIT_74 => X"00000049000000000000001e000000000000002b000000000000000b00000000",
            INIT_75 => X"000000cd00000000000000d100000000000000d800000000000000bf00000000",
            INIT_76 => X"000000170000000000000010000000000000000e000000000000006700000000",
            INIT_77 => X"0000001200000000000000140000000000000016000000000000001b00000000",
            INIT_78 => X"00000017000000000000001a0000000000000016000000000000001a00000000",
            INIT_79 => X"00000034000000000000003c0000000000000025000000000000001900000000",
            INIT_7A => X"0000003b00000000000000380000000000000034000000000000004c00000000",
            INIT_7B => X"00000026000000000000002e000000000000004d000000000000005000000000",
            INIT_7C => X"000000c4000000000000007c0000000000000049000000000000002300000000",
            INIT_7D => X"000000d200000000000000d900000000000000d800000000000000df00000000",
            INIT_7E => X"0000000e00000000000000150000000000000039000000000000007600000000",
            INIT_7F => X"00000011000000000000003e0000000000000047000000000000001f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE38;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE39 : if BRAM_NAME = "sampleifmap_layersamples_instance39" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001700000000000000190000000000000014000000000000001900000000",
            INIT_01 => X"0000005c00000000000000600000000000000035000000000000002100000000",
            INIT_02 => X"00000042000000000000003e000000000000005d000000000000004900000000",
            INIT_03 => X"000000a2000000000000005a0000000000000047000000000000005100000000",
            INIT_04 => X"000000f500000000000000f500000000000000df00000000000000c400000000",
            INIT_05 => X"0000007900000000000000de00000000000000e400000000000000e300000000",
            INIT_06 => X"000000090000000000000011000000000000003b000000000000002500000000",
            INIT_07 => X"000000130000000000000075000000000000008c000000000000004800000000",
            INIT_08 => X"0000001a00000000000000180000000000000015000000000000001900000000",
            INIT_09 => X"000000450000000000000035000000000000002c000000000000002800000000",
            INIT_0A => X"0000002900000000000000250000000000000052000000000000005800000000",
            INIT_0B => X"000000fb00000000000000940000000000000020000000000000003100000000",
            INIT_0C => X"000000e200000000000000e900000000000000f200000000000000f600000000",
            INIT_0D => X"0000001f000000000000008b00000000000000e200000000000000e100000000",
            INIT_0E => X"0000004300000000000000280000000000000019000000000000000b00000000",
            INIT_0F => X"00000022000000000000009700000000000000a2000000000000008500000000",
            INIT_10 => X"0000002600000000000000160000000000000013000000000000001600000000",
            INIT_11 => X"00000036000000000000002e0000000000000046000000000000005d00000000",
            INIT_12 => X"0000001b00000000000000180000000000000026000000000000004b00000000",
            INIT_13 => X"000000e300000000000000a30000000000000031000000000000003800000000",
            INIT_14 => X"000000da00000000000000cb00000000000000cd00000000000000d600000000",
            INIT_15 => X"0000004a00000000000000a300000000000000e400000000000000e500000000",
            INIT_16 => X"000000950000000000000080000000000000005a000000000000003900000000",
            INIT_17 => X"0000003300000000000000a00000000000000096000000000000009700000000",
            INIT_18 => X"0000007c0000000000000026000000000000000f000000000000001300000000",
            INIT_19 => X"0000002a0000000000000024000000000000005a00000000000000af00000000",
            INIT_1A => X"00000015000000000000000b0000000000000017000000000000003f00000000",
            INIT_1B => X"000000d000000000000000aa000000000000004f000000000000004000000000",
            INIT_1C => X"000000d600000000000000d300000000000000c500000000000000c700000000",
            INIT_1D => X"000000b100000000000000e300000000000000d900000000000000ce00000000",
            INIT_1E => X"000000a200000000000000a700000000000000a8000000000000009800000000",
            INIT_1F => X"0000002a00000000000000880000000000000097000000000000009a00000000",
            INIT_20 => X"000000dc0000000000000065000000000000000a000000000000001200000000",
            INIT_21 => X"0000002e000000000000002f000000000000006f00000000000000be00000000",
            INIT_22 => X"0000000e0000000000000009000000000000000a000000000000003900000000",
            INIT_23 => X"000000cc00000000000000b10000000000000042000000000000001f00000000",
            INIT_24 => X"0000007c00000000000000c600000000000000ca00000000000000c200000000",
            INIT_25 => X"000000d300000000000000ac0000000000000066000000000000004f00000000",
            INIT_26 => X"000000a900000000000000b100000000000000b800000000000000c800000000",
            INIT_27 => X"00000011000000000000004a000000000000008c000000000000009c00000000",
            INIT_28 => X"000000a500000000000000840000000000000014000000000000000e00000000",
            INIT_29 => X"0000003400000000000000370000000000000080000000000000009600000000",
            INIT_2A => X"00000016000000000000000a0000000000000003000000000000001e00000000",
            INIT_2B => X"000000c600000000000000b40000000000000048000000000000002d00000000",
            INIT_2C => X"00000019000000000000007b00000000000000cd00000000000000be00000000",
            INIT_2D => X"000000a30000000000000038000000000000001e000000000000001a00000000",
            INIT_2E => X"00000093000000000000009e00000000000000b800000000000000ca00000000",
            INIT_2F => X"00000011000000000000000d0000000000000044000000000000008800000000",
            INIT_30 => X"0000002100000000000000530000000000000023000000000000000a00000000",
            INIT_31 => X"00000035000000000000003e0000000000000082000000000000005300000000",
            INIT_32 => X"0000004800000000000000100000000000000007000000000000001300000000",
            INIT_33 => X"000000c200000000000000b70000000000000075000000000000006c00000000",
            INIT_34 => X"0000001e000000000000002f00000000000000b700000000000000c300000000",
            INIT_35 => X"0000004f0000000000000014000000000000002b000000000000003100000000",
            INIT_36 => X"000000810000000000000084000000000000009400000000000000a100000000",
            INIT_37 => X"000000180000000000000009000000000000000a000000000000004000000000",
            INIT_38 => X"0000002300000000000000370000000000000021000000000000000a00000000",
            INIT_39 => X"00000024000000000000004e0000000000000088000000000000004600000000",
            INIT_3A => X"0000005800000000000000220000000000000011000000000000000f00000000",
            INIT_3B => X"000000cd00000000000000cd000000000000007e000000000000006100000000",
            INIT_3C => X"0000002b0000000000000020000000000000009800000000000000d000000000",
            INIT_3D => X"0000001f0000000000000020000000000000001f000000000000002000000000",
            INIT_3E => X"00000063000000000000008a0000000000000091000000000000007500000000",
            INIT_3F => X"000000210000000000000019000000000000000c000000000000001700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004100000000000000360000000000000015000000000000000a00000000",
            INIT_41 => X"0000002100000000000000570000000000000088000000000000004700000000",
            INIT_42 => X"00000057000000000000003f0000000000000027000000000000001500000000",
            INIT_43 => X"000000c500000000000000cf000000000000009a000000000000005600000000",
            INIT_44 => X"000000380000000000000025000000000000008100000000000000c600000000",
            INIT_45 => X"0000000f000000000000001c000000000000002c000000000000003700000000",
            INIT_46 => X"00000043000000000000008b0000000000000093000000000000004d00000000",
            INIT_47 => X"0000001f000000000000001c0000000000000014000000000000000e00000000",
            INIT_48 => X"0000003e000000000000002f000000000000000e000000000000000700000000",
            INIT_49 => X"0000001c00000000000000560000000000000080000000000000004500000000",
            INIT_4A => X"0000006f000000000000005e000000000000003c000000000000001e00000000",
            INIT_4B => X"000000b400000000000000b600000000000000a2000000000000006f00000000",
            INIT_4C => X"0000003c0000000000000029000000000000007f00000000000000bc00000000",
            INIT_4D => X"0000000f00000000000000230000000000000035000000000000004b00000000",
            INIT_4E => X"00000026000000000000006f000000000000007a000000000000002c00000000",
            INIT_4F => X"000000160000000000000010000000000000000d000000000000000700000000",
            INIT_50 => X"0000003b00000000000000270000000000000011000000000000000b00000000",
            INIT_51 => X"0000003d00000000000000680000000000000075000000000000004600000000",
            INIT_52 => X"000000b7000000000000009f0000000000000079000000000000005100000000",
            INIT_53 => X"000000c700000000000000c900000000000000c300000000000000b900000000",
            INIT_54 => X"0000003c000000000000002a000000000000008800000000000000c600000000",
            INIT_55 => X"0000001c00000000000000340000000000000062000000000000006600000000",
            INIT_56 => X"000000100000000000000045000000000000004f000000000000001500000000",
            INIT_57 => X"00000016000000000000000c0000000000000007000000000000000300000000",
            INIT_58 => X"00000043000000000000001d0000000000000014000000000000001300000000",
            INIT_59 => X"0000003c00000000000000550000000000000067000000000000004900000000",
            INIT_5A => X"00000064000000000000005b0000000000000050000000000000004500000000",
            INIT_5B => X"0000006d00000000000000710000000000000071000000000000006800000000",
            INIT_5C => X"0000004100000000000000250000000000000059000000000000006d00000000",
            INIT_5D => X"00000017000000000000001f0000000000000042000000000000004000000000",
            INIT_5E => X"00000005000000000000000e0000000000000014000000000000000800000000",
            INIT_5F => X"00000018000000000000000b0000000000000006000000000000000600000000",
            INIT_60 => X"00000025000000000000001d000000000000001c000000000000001700000000",
            INIT_61 => X"000000070000000000000016000000000000002c000000000000002c00000000",
            INIT_62 => X"0000000c000000000000000c000000000000000a000000000000000a00000000",
            INIT_63 => X"0000001000000000000000110000000000000010000000000000000d00000000",
            INIT_64 => X"000000430000000000000009000000000000000f000000000000000f00000000",
            INIT_65 => X"0000001000000000000000380000000000000030000000000000004400000000",
            INIT_66 => X"0000000400000000000000030000000000000003000000000000000400000000",
            INIT_67 => X"00000019000000000000000e0000000000000009000000000000000600000000",
            INIT_68 => X"0000002000000000000000270000000000000025000000000000002100000000",
            INIT_69 => X"0000002000000000000000190000000000000012000000000000001700000000",
            INIT_6A => X"0000001700000000000000170000000000000015000000000000001700000000",
            INIT_6B => X"0000000f00000000000000130000000000000015000000000000001700000000",
            INIT_6C => X"000000180000000000000007000000000000000a000000000000000b00000000",
            INIT_6D => X"0000000800000000000000290000000000000047000000000000003e00000000",
            INIT_6E => X"0000000600000000000000050000000000000005000000000000000400000000",
            INIT_6F => X"0000001d0000000000000018000000000000000e000000000000000900000000",
            INIT_70 => X"0000003200000000000000290000000000000025000000000000002300000000",
            INIT_71 => X"0000004d00000000000000510000000000000043000000000000003c00000000",
            INIT_72 => X"00000030000000000000002d0000000000000024000000000000002c00000000",
            INIT_73 => X"000000230000000000000027000000000000002c000000000000003100000000",
            INIT_74 => X"000000100000000000000015000000000000001b000000000000001d00000000",
            INIT_75 => X"00000009000000000000000a0000000000000019000000000000001700000000",
            INIT_76 => X"0000000b000000000000000a0000000000000009000000000000000b00000000",
            INIT_77 => X"0000001e000000000000001f0000000000000014000000000000000e00000000",
            INIT_78 => X"00000057000000000000003b000000000000002a000000000000002a00000000",
            INIT_79 => X"000000520000000000000066000000000000006f000000000000006d00000000",
            INIT_7A => X"000000470000000000000045000000000000003e000000000000003700000000",
            INIT_7B => X"0000004300000000000000460000000000000048000000000000004a00000000",
            INIT_7C => X"00000029000000000000002b0000000000000033000000000000003b00000000",
            INIT_7D => X"000000120000000000000018000000000000002c000000000000002f00000000",
            INIT_7E => X"0000001300000000000000150000000000000016000000000000001400000000",
            INIT_7F => X"0000001e0000000000000020000000000000001c000000000000001600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE39;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE40 : if BRAM_NAME = "sampleifmap_layersamples_instance40" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000a000000000000000e000000000000000b000000000000000d00000000",
            INIT_01 => X"000000020000000000000005000000000000000a000000000000000900000000",
            INIT_02 => X"0000000200000000000000010000000000000003000000000000000300000000",
            INIT_03 => X"0000000000000000000000050000000000000006000000000000000400000000",
            INIT_04 => X"0000005600000000000000230000000000000000000000000000000100000000",
            INIT_05 => X"00000008000000000000001d0000000000000017000000000000001600000000",
            INIT_06 => X"0000001d0000000000000027000000000000001b000000000000000d00000000",
            INIT_07 => X"0000000500000000000000060000000000000008000000000000001300000000",
            INIT_08 => X"00000004000000000000000a000000000000000c000000000000000d00000000",
            INIT_09 => X"0000000000000000000000030000000000000008000000000000000700000000",
            INIT_0A => X"0000000100000000000000010000000000000002000000000000000400000000",
            INIT_0B => X"0000000100000000000000040000000000000004000000000000000200000000",
            INIT_0C => X"0000001300000000000000100000000000000001000000000000000100000000",
            INIT_0D => X"0000000700000000000000060000000000000006000000000000000700000000",
            INIT_0E => X"000000160000000000000017000000000000002e000000000000002100000000",
            INIT_0F => X"0000000600000000000000040000000000000008000000000000001300000000",
            INIT_10 => X"0000000000000000000000030000000000000004000000000000000700000000",
            INIT_11 => X"0000000000000000000000010000000000000004000000000000000400000000",
            INIT_12 => X"0000000400000000000000040000000000000004000000000000000400000000",
            INIT_13 => X"0000000300000000000000050000000000000006000000000000000400000000",
            INIT_14 => X"00000009000000000000000c0000000000000003000000000000000400000000",
            INIT_15 => X"0000000a00000000000000060000000000000007000000000000000400000000",
            INIT_16 => X"0000000c000000000000000d0000000000000023000000000000002800000000",
            INIT_17 => X"0000000600000000000000030000000000000006000000000000000f00000000",
            INIT_18 => X"0000000b00000000000000080000000000000003000000000000000100000000",
            INIT_19 => X"0000000300000000000000030000000000000004000000000000001200000000",
            INIT_1A => X"0000000700000000000000080000000000000006000000000000000500000000",
            INIT_1B => X"0000000600000000000000060000000000000009000000000000000800000000",
            INIT_1C => X"00000009000000000000000a0000000000000005000000000000000700000000",
            INIT_1D => X"000000170000000000000010000000000000000a000000000000000400000000",
            INIT_1E => X"0000000e00000000000000110000000000000016000000000000001e00000000",
            INIT_1F => X"0000000800000000000000050000000000000006000000000000000f00000000",
            INIT_20 => X"0000001a000000000000001d0000000000000013000000000000000c00000000",
            INIT_21 => X"0000000800000000000000070000000000000006000000000000001700000000",
            INIT_22 => X"0000000800000000000000090000000000000008000000000000000700000000",
            INIT_23 => X"000000080000000000000007000000000000000a000000000000000900000000",
            INIT_24 => X"0000000700000000000000080000000000000007000000000000000900000000",
            INIT_25 => X"0000002700000000000000400000000000000025000000000000000800000000",
            INIT_26 => X"00000015000000000000000e0000000000000010000000000000001000000000",
            INIT_27 => X"00000009000000000000000d000000000000000f000000000000000e00000000",
            INIT_28 => X"0000000c0000000000000016000000000000001e000000000000001800000000",
            INIT_29 => X"0000000800000000000000090000000000000006000000000000000900000000",
            INIT_2A => X"0000000a00000000000000090000000000000005000000000000000500000000",
            INIT_2B => X"000000090000000000000007000000000000000a000000000000000b00000000",
            INIT_2C => X"00000007000000000000000b000000000000000b000000000000000a00000000",
            INIT_2D => X"0000003b000000000000005d0000000000000055000000000000001400000000",
            INIT_2E => X"000000200000000000000013000000000000000e000000000000002200000000",
            INIT_2F => X"000000090000000000000010000000000000001b000000000000001700000000",
            INIT_30 => X"00000007000000000000000a000000000000000b000000000000000c00000000",
            INIT_31 => X"00000007000000000000000a0000000000000008000000000000000800000000",
            INIT_32 => X"0000000e000000000000000a0000000000000005000000000000000600000000",
            INIT_33 => X"0000000c000000000000000a000000000000000c000000000000000d00000000",
            INIT_34 => X"00000007000000000000000e000000000000000e000000000000000900000000",
            INIT_35 => X"00000028000000000000003c0000000000000056000000000000002500000000",
            INIT_36 => X"0000001c000000000000001c000000000000001c000000000000003500000000",
            INIT_37 => X"0000000700000000000000060000000000000010000000000000001400000000",
            INIT_38 => X"0000000700000000000000060000000000000006000000000000000300000000",
            INIT_39 => X"00000009000000000000000c000000000000000a000000000000000b00000000",
            INIT_3A => X"0000000e000000000000000c0000000000000008000000000000000900000000",
            INIT_3B => X"0000001300000000000000100000000000000012000000000000000e00000000",
            INIT_3C => X"00000016000000000000001a0000000000000015000000000000001000000000",
            INIT_3D => X"0000000a0000000000000014000000000000003e000000000000003100000000",
            INIT_3E => X"0000000d0000000000000010000000000000001a000000000000001e00000000",
            INIT_3F => X"0000000700000000000000040000000000000008000000000000000900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000080000000000000009000000000000000a000000000000000700000000",
            INIT_41 => X"0000000b000000000000000e000000000000000a000000000000000b00000000",
            INIT_42 => X"0000000f000000000000000e000000000000000c000000000000000d00000000",
            INIT_43 => X"0000002800000000000000220000000000000024000000000000001300000000",
            INIT_44 => X"0000002200000000000000220000000000000020000000000000002400000000",
            INIT_45 => X"00000009000000000000000f000000000000002b000000000000003300000000",
            INIT_46 => X"0000000a0000000000000009000000000000000c000000000000001400000000",
            INIT_47 => X"0000000800000000000000080000000000000008000000000000000800000000",
            INIT_48 => X"00000008000000000000000b000000000000000c000000000000000c00000000",
            INIT_49 => X"0000000d000000000000000e000000000000000a000000000000000c00000000",
            INIT_4A => X"000000220000000000000014000000000000000e000000000000000e00000000",
            INIT_4B => X"0000002600000000000000280000000000000031000000000000002700000000",
            INIT_4C => X"000000320000000000000027000000000000001b000000000000002000000000",
            INIT_4D => X"000000260000000000000034000000000000003b000000000000003600000000",
            INIT_4E => X"0000000c000000000000000b0000000000000015000000000000002300000000",
            INIT_4F => X"0000000a000000000000000b0000000000000009000000000000000600000000",
            INIT_50 => X"00000009000000000000000b000000000000000b000000000000000c00000000",
            INIT_51 => X"0000000d000000000000000d000000000000000a000000000000000c00000000",
            INIT_52 => X"00000028000000000000001b0000000000000010000000000000000d00000000",
            INIT_53 => X"0000003f00000000000000320000000000000032000000000000002000000000",
            INIT_54 => X"000000b400000000000000a10000000000000077000000000000005800000000",
            INIT_55 => X"0000002200000000000000540000000000000071000000000000007900000000",
            INIT_56 => X"00000011000000000000001d0000000000000031000000000000003200000000",
            INIT_57 => X"0000000a000000000000000c000000000000000a000000000000000900000000",
            INIT_58 => X"0000000b000000000000000e000000000000000a000000000000000900000000",
            INIT_59 => X"0000000c000000000000000d000000000000000c000000000000000e00000000",
            INIT_5A => X"0000002700000000000000180000000000000012000000000000000c00000000",
            INIT_5B => X"000000ba00000000000000af0000000000000093000000000000004d00000000",
            INIT_5C => X"000000ca00000000000000d200000000000000c800000000000000c800000000",
            INIT_5D => X"0000001c000000000000009e00000000000000d500000000000000b100000000",
            INIT_5E => X"0000002500000000000000460000000000000022000000000000001300000000",
            INIT_5F => X"00000009000000000000000b0000000000000009000000000000000a00000000",
            INIT_60 => X"0000000d000000000000000f000000000000000a000000000000000800000000",
            INIT_61 => X"0000000e000000000000000d000000000000000e000000000000001000000000",
            INIT_62 => X"0000006c000000000000003e0000000000000018000000000000000c00000000",
            INIT_63 => X"0000007d000000000000009300000000000000a2000000000000008e00000000",
            INIT_64 => X"0000004a0000000000000054000000000000005e000000000000006e00000000",
            INIT_65 => X"0000005400000000000000d700000000000000f1000000000000007e00000000",
            INIT_66 => X"0000004900000000000000340000000000000009000000000000000c00000000",
            INIT_67 => X"000000080000000000000009000000000000000d000000000000001900000000",
            INIT_68 => X"0000000e000000000000000f000000000000000b000000000000000b00000000",
            INIT_69 => X"0000000e000000000000000c0000000000000010000000000000001100000000",
            INIT_6A => X"0000005d00000000000000670000000000000044000000000000001400000000",
            INIT_6B => X"00000019000000000000003d000000000000005f000000000000005600000000",
            INIT_6C => X"0000001700000000000000110000000000000023000000000000001600000000",
            INIT_6D => X"000000a700000000000000eb00000000000000eb000000000000008900000000",
            INIT_6E => X"0000004200000000000000170000000000000007000000000000002a00000000",
            INIT_6F => X"0000000700000000000000090000000000000011000000000000002800000000",
            INIT_70 => X"0000000e0000000000000012000000000000000d000000000000000f00000000",
            INIT_71 => X"00000012000000000000000b0000000000000012000000000000001000000000",
            INIT_72 => X"0000002e000000000000003b0000000000000053000000000000003600000000",
            INIT_73 => X"0000001b00000000000000370000000000000053000000000000004400000000",
            INIT_74 => X"0000004c000000000000001c0000000000000027000000000000000c00000000",
            INIT_75 => X"000000e000000000000000e700000000000000e800000000000000c800000000",
            INIT_76 => X"0000001a00000000000000130000000000000016000000000000007300000000",
            INIT_77 => X"00000008000000000000000d0000000000000016000000000000001f00000000",
            INIT_78 => X"0000000e0000000000000013000000000000000d000000000000001000000000",
            INIT_79 => X"000000370000000000000039000000000000001e000000000000000e00000000",
            INIT_7A => X"0000003c00000000000000390000000000000035000000000000004f00000000",
            INIT_7B => X"000000290000000000000032000000000000004e000000000000005200000000",
            INIT_7C => X"000000c8000000000000007c0000000000000047000000000000002300000000",
            INIT_7D => X"000000dd00000000000000ec00000000000000e600000000000000e700000000",
            INIT_7E => X"0000000e000000000000001a0000000000000044000000000000007e00000000",
            INIT_7F => X"00000009000000000000003f0000000000000049000000000000002000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE40;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE41 : if BRAM_NAME = "sampleifmap_layersamples_instance41" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000110000000000000013000000000000000e000000000000001100000000",
            INIT_01 => X"0000005c000000000000005d000000000000002f000000000000001800000000",
            INIT_02 => X"0000003d000000000000003c0000000000000062000000000000004f00000000",
            INIT_03 => X"000000a6000000000000005e0000000000000047000000000000004c00000000",
            INIT_04 => X"000000fc00000000000000fa00000000000000e200000000000000c600000000",
            INIT_05 => X"0000007c00000000000000e700000000000000f000000000000000ed00000000",
            INIT_06 => X"0000000c000000000000001c000000000000004a000000000000002a00000000",
            INIT_07 => X"00000011000000000000007e0000000000000095000000000000004c00000000",
            INIT_08 => X"0000001500000000000000120000000000000010000000000000001200000000",
            INIT_09 => X"000000480000000000000038000000000000002a000000000000002400000000",
            INIT_0A => X"0000002400000000000000240000000000000058000000000000006000000000",
            INIT_0B => X"00000100000000000000009a0000000000000022000000000000002d00000000",
            INIT_0C => X"000000ed00000000000000f400000000000000f900000000000000fa00000000",
            INIT_0D => X"00000027000000000000009600000000000000ee00000000000000ed00000000",
            INIT_0E => X"0000004d000000000000003b000000000000002e000000000000001500000000",
            INIT_0F => X"0000002600000000000000a300000000000000ae000000000000008e00000000",
            INIT_10 => X"0000002200000000000000100000000000000010000000000000001100000000",
            INIT_11 => X"00000042000000000000003c0000000000000049000000000000005c00000000",
            INIT_12 => X"00000021000000000000001c000000000000002c000000000000005400000000",
            INIT_13 => X"000000f000000000000000ae0000000000000037000000000000003e00000000",
            INIT_14 => X"000000e700000000000000d900000000000000d900000000000000e100000000",
            INIT_15 => X"0000005600000000000000b100000000000000ee00000000000000ef00000000",
            INIT_16 => X"000000a40000000000000092000000000000006a000000000000004500000000",
            INIT_17 => X"0000003700000000000000a900000000000000a100000000000000a400000000",
            INIT_18 => X"0000007d0000000000000020000000000000000a000000000000000d00000000",
            INIT_19 => X"000000380000000000000035000000000000006200000000000000b400000000",
            INIT_1A => X"0000001b000000000000000e000000000000001c000000000000004800000000",
            INIT_1B => X"000000e000000000000000b90000000000000059000000000000004900000000",
            INIT_1C => X"000000e300000000000000e400000000000000d500000000000000d500000000",
            INIT_1D => X"000000c000000000000000f200000000000000e100000000000000d700000000",
            INIT_1E => X"000000b000000000000000b500000000000000b400000000000000a500000000",
            INIT_1F => X"0000002a000000000000008d000000000000009f00000000000000a600000000",
            INIT_20 => X"000000e500000000000000650000000000000007000000000000000c00000000",
            INIT_21 => X"00000039000000000000003e000000000000007b00000000000000c900000000",
            INIT_22 => X"0000000f0000000000000009000000000000000f000000000000004100000000",
            INIT_23 => X"000000da00000000000000bf000000000000004f000000000000002600000000",
            INIT_24 => X"0000008a00000000000000d800000000000000db00000000000000d000000000",
            INIT_25 => X"000000e400000000000000b8000000000000006d000000000000005800000000",
            INIT_26 => X"000000b500000000000000bf00000000000000c900000000000000da00000000",
            INIT_27 => X"0000000e000000000000004d000000000000009300000000000000a600000000",
            INIT_28 => X"000000b3000000000000008b0000000000000018000000000000000d00000000",
            INIT_29 => X"0000003d0000000000000045000000000000008d00000000000000a200000000",
            INIT_2A => X"0000001b000000000000000b0000000000000004000000000000002300000000",
            INIT_2B => X"000000d400000000000000c20000000000000056000000000000003600000000",
            INIT_2C => X"00000024000000000000008800000000000000db00000000000000cc00000000",
            INIT_2D => X"000000b100000000000000400000000000000022000000000000002000000000",
            INIT_2E => X"0000009f00000000000000ad00000000000000cc00000000000000dd00000000",
            INIT_2F => X"0000000d000000000000000f0000000000000049000000000000009000000000",
            INIT_30 => X"00000031000000000000005b0000000000000027000000000000000900000000",
            INIT_31 => X"0000003e000000000000004c000000000000008f000000000000006000000000",
            INIT_32 => X"0000005100000000000000150000000000000007000000000000001500000000",
            INIT_33 => X"000000d000000000000000c50000000000000083000000000000007900000000",
            INIT_34 => X"00000026000000000000003800000000000000c100000000000000d100000000",
            INIT_35 => X"000000590000000000000019000000000000002e000000000000003700000000",
            INIT_36 => X"0000008d000000000000009500000000000000a900000000000000b200000000",
            INIT_37 => X"000000140000000000000008000000000000000e000000000000004800000000",
            INIT_38 => X"00000030000000000000003b0000000000000022000000000000000500000000",
            INIT_39 => X"0000002d000000000000005c0000000000000095000000000000005300000000",
            INIT_3A => X"00000064000000000000002a0000000000000013000000000000000f00000000",
            INIT_3B => X"000000db00000000000000db000000000000008c000000000000006f00000000",
            INIT_3C => X"00000033000000000000002600000000000000a000000000000000de00000000",
            INIT_3D => X"0000002700000000000000240000000000000023000000000000002500000000",
            INIT_3E => X"0000006e000000000000009b00000000000000a4000000000000008200000000",
            INIT_3F => X"0000001e0000000000000016000000000000000c000000000000001d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004d000000000000003a0000000000000017000000000000000700000000",
            INIT_41 => X"0000002a00000000000000650000000000000094000000000000005400000000",
            INIT_42 => X"00000065000000000000004a000000000000002b000000000000001600000000",
            INIT_43 => X"000000d300000000000000dd00000000000000a8000000000000006400000000",
            INIT_44 => X"00000040000000000000002b000000000000008900000000000000d400000000",
            INIT_45 => X"0000001500000000000000230000000000000034000000000000003f00000000",
            INIT_46 => X"0000004e000000000000009a00000000000000a2000000000000005600000000",
            INIT_47 => X"0000001c00000000000000180000000000000012000000000000001300000000",
            INIT_48 => X"0000004c00000000000000370000000000000015000000000000000900000000",
            INIT_49 => X"000000250000000000000065000000000000008c000000000000005200000000",
            INIT_4A => X"0000007f000000000000006c0000000000000043000000000000002100000000",
            INIT_4B => X"000000c200000000000000c300000000000000b0000000000000007e00000000",
            INIT_4C => X"000000460000000000000030000000000000008700000000000000c900000000",
            INIT_4D => X"00000015000000000000002e0000000000000041000000000000005600000000",
            INIT_4E => X"00000031000000000000007b0000000000000083000000000000003200000000",
            INIT_4F => X"00000014000000000000000b000000000000000a000000000000000b00000000",
            INIT_50 => X"0000004900000000000000310000000000000017000000000000000b00000000",
            INIT_51 => X"0000004b00000000000000780000000000000084000000000000005700000000",
            INIT_52 => X"000000c800000000000000b10000000000000086000000000000005d00000000",
            INIT_53 => X"000000d500000000000000d400000000000000cf00000000000000c800000000",
            INIT_54 => X"000000480000000000000035000000000000009400000000000000d600000000",
            INIT_55 => X"000000220000000000000040000000000000006e000000000000007100000000",
            INIT_56 => X"00000016000000000000004c0000000000000055000000000000001800000000",
            INIT_57 => X"00000016000000000000000d0000000000000009000000000000000700000000",
            INIT_58 => X"0000004e00000000000000250000000000000016000000000000000f00000000",
            INIT_59 => X"0000004800000000000000600000000000000073000000000000005700000000",
            INIT_5A => X"000000720000000000000069000000000000005d000000000000005200000000",
            INIT_5B => X"0000007b000000000000007e000000000000007d000000000000007700000000",
            INIT_5C => X"0000004c00000000000000300000000000000066000000000000007c00000000",
            INIT_5D => X"0000001b0000000000000029000000000000004e000000000000004b00000000",
            INIT_5E => X"0000000600000000000000100000000000000018000000000000000900000000",
            INIT_5F => X"00000019000000000000000f000000000000000a000000000000000800000000",
            INIT_60 => X"0000002b0000000000000023000000000000001f000000000000001500000000",
            INIT_61 => X"0000000c00000000000000190000000000000030000000000000003200000000",
            INIT_62 => X"000000110000000000000011000000000000000e000000000000000e00000000",
            INIT_63 => X"00000019000000000000001a0000000000000018000000000000001400000000",
            INIT_64 => X"0000004a000000000000000d0000000000000014000000000000001800000000",
            INIT_65 => X"000000120000000000000041000000000000003b000000000000004e00000000",
            INIT_66 => X"0000000300000000000000040000000000000005000000000000000300000000",
            INIT_67 => X"0000001a000000000000000d0000000000000009000000000000000500000000",
            INIT_68 => X"00000025000000000000002c0000000000000028000000000000002100000000",
            INIT_69 => X"00000025000000000000001e0000000000000017000000000000001e00000000",
            INIT_6A => X"0000001c000000000000001c0000000000000019000000000000001c00000000",
            INIT_6B => X"0000001300000000000000170000000000000018000000000000001b00000000",
            INIT_6C => X"0000001c00000000000000060000000000000009000000000000000f00000000",
            INIT_6D => X"00000008000000000000002f0000000000000053000000000000004700000000",
            INIT_6E => X"0000000400000000000000050000000000000005000000000000000200000000",
            INIT_6F => X"0000001c0000000000000015000000000000000b000000000000000600000000",
            INIT_70 => X"0000003b00000000000000300000000000000029000000000000002500000000",
            INIT_71 => X"00000059000000000000005c000000000000004f000000000000004900000000",
            INIT_72 => X"0000003b0000000000000038000000000000002f000000000000003800000000",
            INIT_73 => X"00000028000000000000002b0000000000000030000000000000003900000000",
            INIT_74 => X"000000150000000000000015000000000000001b000000000000002300000000",
            INIT_75 => X"0000000800000000000000100000000000000025000000000000002100000000",
            INIT_76 => X"0000000a000000000000000a0000000000000009000000000000000800000000",
            INIT_77 => X"0000001c000000000000001d0000000000000012000000000000000d00000000",
            INIT_78 => X"0000006500000000000000460000000000000031000000000000002c00000000",
            INIT_79 => X"0000006300000000000000760000000000000080000000000000008000000000",
            INIT_7A => X"000000550000000000000054000000000000004e000000000000004700000000",
            INIT_7B => X"0000004f00000000000000510000000000000053000000000000005700000000",
            INIT_7C => X"000000310000000000000031000000000000003c000000000000004700000000",
            INIT_7D => X"0000001300000000000000200000000000000038000000000000003a00000000",
            INIT_7E => X"0000001500000000000000180000000000000018000000000000001300000000",
            INIT_7F => X"0000001c0000000000000022000000000000001f000000000000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE41;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE42 : if BRAM_NAME = "sampleifmap_layersamples_instance42" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004d00000000000000510000000000000052000000000000005300000000",
            INIT_01 => X"0000005c000000000000005b0000000000000055000000000000005100000000",
            INIT_02 => X"0000005c0000000000000065000000000000005f000000000000005c00000000",
            INIT_03 => X"0000004c00000000000000500000000000000052000000000000005700000000",
            INIT_04 => X"0000003e000000000000003f0000000000000041000000000000004400000000",
            INIT_05 => X"0000002f00000000000000340000000000000038000000000000003c00000000",
            INIT_06 => X"0000002200000000000000230000000000000025000000000000002a00000000",
            INIT_07 => X"000000150000000000000019000000000000001d000000000000002400000000",
            INIT_08 => X"0000004d00000000000000530000000000000053000000000000005400000000",
            INIT_09 => X"0000005d000000000000005a0000000000000054000000000000005000000000",
            INIT_0A => X"00000061000000000000005f0000000000000058000000000000005a00000000",
            INIT_0B => X"0000004c000000000000004e0000000000000052000000000000005800000000",
            INIT_0C => X"0000004200000000000000400000000000000044000000000000004700000000",
            INIT_0D => X"0000002e00000000000000340000000000000036000000000000003d00000000",
            INIT_0E => X"0000002300000000000000240000000000000026000000000000002a00000000",
            INIT_0F => X"0000001f000000000000001d000000000000001e000000000000002400000000",
            INIT_10 => X"0000004b00000000000000500000000000000051000000000000005200000000",
            INIT_11 => X"0000004c00000000000000580000000000000054000000000000004b00000000",
            INIT_12 => X"0000006300000000000000570000000000000056000000000000005200000000",
            INIT_13 => X"0000004c000000000000004d0000000000000058000000000000006500000000",
            INIT_14 => X"0000004000000000000000400000000000000044000000000000004900000000",
            INIT_15 => X"0000002d00000000000000340000000000000037000000000000003a00000000",
            INIT_16 => X"0000002c00000000000000290000000000000028000000000000002b00000000",
            INIT_17 => X"0000003500000000000000310000000000000030000000000000003100000000",
            INIT_18 => X"0000004e00000000000000500000000000000051000000000000005300000000",
            INIT_19 => X"0000003200000000000000500000000000000057000000000000004a00000000",
            INIT_1A => X"0000005b00000000000000570000000000000061000000000000005500000000",
            INIT_1B => X"0000005000000000000000580000000000000066000000000000006800000000",
            INIT_1C => X"0000003f000000000000003f0000000000000040000000000000004900000000",
            INIT_1D => X"0000003a00000000000000390000000000000038000000000000003b00000000",
            INIT_1E => X"000000470000000000000044000000000000003f000000000000003d00000000",
            INIT_1F => X"0000004500000000000000450000000000000047000000000000004900000000",
            INIT_20 => X"0000004f000000000000004f000000000000004f000000000000004f00000000",
            INIT_21 => X"00000037000000000000004c0000000000000053000000000000004a00000000",
            INIT_22 => X"0000004b000000000000004b0000000000000054000000000000005300000000",
            INIT_23 => X"00000057000000000000005a0000000000000059000000000000004e00000000",
            INIT_24 => X"0000004600000000000000430000000000000042000000000000005300000000",
            INIT_25 => X"0000005700000000000000540000000000000050000000000000004e00000000",
            INIT_26 => X"0000005900000000000000590000000000000056000000000000005700000000",
            INIT_27 => X"00000049000000000000004f0000000000000054000000000000005800000000",
            INIT_28 => X"0000004d000000000000004b000000000000004a000000000000004c00000000",
            INIT_29 => X"0000004600000000000000460000000000000049000000000000004900000000",
            INIT_2A => X"0000004900000000000000470000000000000045000000000000004600000000",
            INIT_2B => X"00000051000000000000004e000000000000004e000000000000004b00000000",
            INIT_2C => X"0000006200000000000000600000000000000059000000000000005a00000000",
            INIT_2D => X"0000006800000000000000660000000000000068000000000000006400000000",
            INIT_2E => X"0000005e0000000000000061000000000000005f000000000000006300000000",
            INIT_2F => X"0000004200000000000000490000000000000050000000000000005700000000",
            INIT_30 => X"0000004900000000000000470000000000000048000000000000004a00000000",
            INIT_31 => X"00000033000000000000002b000000000000003e000000000000004a00000000",
            INIT_32 => X"0000004700000000000000440000000000000040000000000000004400000000",
            INIT_33 => X"0000005e0000000000000051000000000000004a000000000000004b00000000",
            INIT_34 => X"00000072000000000000006e0000000000000062000000000000006000000000",
            INIT_35 => X"0000006d00000000000000680000000000000064000000000000006600000000",
            INIT_36 => X"000000500000000000000055000000000000005b000000000000006300000000",
            INIT_37 => X"0000004300000000000000460000000000000049000000000000004c00000000",
            INIT_38 => X"0000004800000000000000470000000000000048000000000000004700000000",
            INIT_39 => X"00000029000000000000002a000000000000003a000000000000004700000000",
            INIT_3A => X"0000003f000000000000003a0000000000000036000000000000003900000000",
            INIT_3B => X"0000006000000000000000520000000000000047000000000000004100000000",
            INIT_3C => X"00000067000000000000005d000000000000005e000000000000006900000000",
            INIT_3D => X"00000061000000000000006c000000000000006a000000000000006700000000",
            INIT_3E => X"000000500000000000000054000000000000005b000000000000005d00000000",
            INIT_3F => X"0000004d000000000000004f0000000000000050000000000000005000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000052000000000000004b0000000000000049000000000000004900000000",
            INIT_41 => X"0000002e00000000000000570000000000000067000000000000005800000000",
            INIT_42 => X"0000005200000000000000450000000000000038000000000000003800000000",
            INIT_43 => X"00000057000000000000005a0000000000000057000000000000005100000000",
            INIT_44 => X"0000005b000000000000005e0000000000000063000000000000006200000000",
            INIT_45 => X"00000066000000000000006a0000000000000066000000000000006100000000",
            INIT_46 => X"0000005c00000000000000610000000000000063000000000000005e00000000",
            INIT_47 => X"0000005f000000000000005b0000000000000059000000000000005900000000",
            INIT_48 => X"0000007b000000000000006d000000000000005f000000000000005600000000",
            INIT_49 => X"0000003300000000000000680000000000000099000000000000008800000000",
            INIT_4A => X"000000610000000000000049000000000000003b000000000000003c00000000",
            INIT_4B => X"0000005a0000000000000066000000000000006c000000000000006500000000",
            INIT_4C => X"0000005d00000000000000610000000000000061000000000000005f00000000",
            INIT_4D => X"0000006e00000000000000690000000000000063000000000000005d00000000",
            INIT_4E => X"0000006c000000000000006c0000000000000069000000000000006700000000",
            INIT_4F => X"0000006e000000000000006e000000000000006e000000000000006d00000000",
            INIT_50 => X"0000009d0000000000000096000000000000008b000000000000007f00000000",
            INIT_51 => X"00000032000000000000005700000000000000a200000000000000a000000000",
            INIT_52 => X"0000005800000000000000350000000000000038000000000000004300000000",
            INIT_53 => X"0000005a000000000000006b0000000000000070000000000000006500000000",
            INIT_54 => X"00000060000000000000005e0000000000000060000000000000005e00000000",
            INIT_55 => X"000000650000000000000060000000000000005f000000000000006000000000",
            INIT_56 => X"0000007e000000000000007d0000000000000071000000000000006800000000",
            INIT_57 => X"0000007000000000000000740000000000000077000000000000007b00000000",
            INIT_58 => X"000000a2000000000000009f000000000000009d000000000000009800000000",
            INIT_59 => X"0000002c000000000000005a000000000000009f00000000000000a000000000",
            INIT_5A => X"00000056000000000000003a0000000000000045000000000000004800000000",
            INIT_5B => X"0000005c0000000000000061000000000000005a000000000000006700000000",
            INIT_5C => X"0000005e000000000000005f0000000000000060000000000000005a00000000",
            INIT_5D => X"0000005c00000000000000570000000000000062000000000000006300000000",
            INIT_5E => X"0000008300000000000000830000000000000070000000000000006100000000",
            INIT_5F => X"0000006c00000000000000740000000000000079000000000000007f00000000",
            INIT_60 => X"0000009d00000000000000a0000000000000009e000000000000009b00000000",
            INIT_61 => X"0000003000000000000000720000000000000094000000000000009800000000",
            INIT_62 => X"00000067000000000000005e0000000000000058000000000000004400000000",
            INIT_63 => X"0000005d00000000000000580000000000000060000000000000007300000000",
            INIT_64 => X"0000005e00000000000000620000000000000065000000000000005900000000",
            INIT_65 => X"0000005500000000000000540000000000000065000000000000006300000000",
            INIT_66 => X"00000084000000000000007d000000000000006e000000000000006900000000",
            INIT_67 => X"0000005f000000000000006b0000000000000076000000000000007f00000000",
            INIT_68 => X"0000009200000000000000950000000000000094000000000000009400000000",
            INIT_69 => X"000000500000000000000088000000000000008e000000000000009000000000",
            INIT_6A => X"00000068000000000000005e0000000000000048000000000000002f00000000",
            INIT_6B => X"0000005e000000000000005c0000000000000071000000000000007200000000",
            INIT_6C => X"0000005d00000000000000610000000000000067000000000000005d00000000",
            INIT_6D => X"0000005200000000000000550000000000000061000000000000006000000000",
            INIT_6E => X"00000079000000000000006f000000000000006b000000000000006b00000000",
            INIT_6F => X"0000004d00000000000000570000000000000064000000000000007000000000",
            INIT_70 => X"0000008c000000000000008a0000000000000087000000000000008600000000",
            INIT_71 => X"0000008900000000000000970000000000000093000000000000008e00000000",
            INIT_72 => X"0000003e00000000000000320000000000000049000000000000005d00000000",
            INIT_73 => X"00000062000000000000005a000000000000005e000000000000005900000000",
            INIT_74 => X"0000006100000000000000670000000000000069000000000000006600000000",
            INIT_75 => X"000000530000000000000056000000000000005e000000000000005e00000000",
            INIT_76 => X"00000066000000000000005c0000000000000065000000000000005f00000000",
            INIT_77 => X"0000004b000000000000004a0000000000000052000000000000005f00000000",
            INIT_78 => X"00000090000000000000008b0000000000000086000000000000008300000000",
            INIT_79 => X"00000098000000000000009a000000000000009f000000000000009800000000",
            INIT_7A => X"0000003900000000000000350000000000000076000000000000009e00000000",
            INIT_7B => X"00000066000000000000005f0000000000000064000000000000006700000000",
            INIT_7C => X"0000006a000000000000006f0000000000000074000000000000006e00000000",
            INIT_7D => X"000000550000000000000057000000000000005b000000000000006100000000",
            INIT_7E => X"0000005300000000000000550000000000000062000000000000005400000000",
            INIT_7F => X"0000005f000000000000005a0000000000000055000000000000005300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE42;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE43 : if BRAM_NAME = "sampleifmap_layersamples_instance43" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a000000000000000980000000000000090000000000000008700000000",
            INIT_01 => X"00000073000000000000008900000000000000a100000000000000a400000000",
            INIT_02 => X"0000006e00000000000000800000000000000091000000000000009d00000000",
            INIT_03 => X"000000670000000000000068000000000000007a000000000000007b00000000",
            INIT_04 => X"00000068000000000000006c000000000000006d000000000000006900000000",
            INIT_05 => X"000000570000000000000058000000000000005a000000000000006100000000",
            INIT_06 => X"000000550000000000000057000000000000005c000000000000004f00000000",
            INIT_07 => X"0000005e00000000000000690000000000000069000000000000006500000000",
            INIT_08 => X"000000a4000000000000009f000000000000009a000000000000009400000000",
            INIT_09 => X"0000007f00000000000000b000000000000000b300000000000000aa00000000",
            INIT_0A => X"00000098000000000000009d00000000000000c500000000000000b000000000",
            INIT_0B => X"0000006700000000000000800000000000000091000000000000007100000000",
            INIT_0C => X"0000006600000000000000680000000000000065000000000000006700000000",
            INIT_0D => X"00000059000000000000005b000000000000005f000000000000006100000000",
            INIT_0E => X"0000005b000000000000005b0000000000000056000000000000004f00000000",
            INIT_0F => X"0000004600000000000000560000000000000068000000000000006d00000000",
            INIT_10 => X"000000c500000000000000b200000000000000a4000000000000009b00000000",
            INIT_11 => X"000000c400000000000000f800000000000000ee00000000000000dd00000000",
            INIT_12 => X"000000b800000000000000b000000000000000c8000000000000009c00000000",
            INIT_13 => X"0000006a0000000000000089000000000000008e000000000000006c00000000",
            INIT_14 => X"0000006500000000000000640000000000000063000000000000006400000000",
            INIT_15 => X"00000059000000000000005f0000000000000063000000000000006500000000",
            INIT_16 => X"00000053000000000000005c0000000000000051000000000000005000000000",
            INIT_17 => X"0000004700000000000000490000000000000052000000000000005800000000",
            INIT_18 => X"000000f900000000000000eb00000000000000d600000000000000bf00000000",
            INIT_19 => X"000000f400000000000000fb00000000000000f600000000000000fd00000000",
            INIT_1A => X"000000c300000000000000ac000000000000009e00000000000000a000000000",
            INIT_1B => X"0000006e000000000000008b0000000000000072000000000000007100000000",
            INIT_1C => X"0000006300000000000000610000000000000062000000000000006200000000",
            INIT_1D => X"0000005c00000000000000660000000000000068000000000000006700000000",
            INIT_1E => X"000000490000000000000055000000000000004e000000000000005300000000",
            INIT_1F => X"00000048000000000000004a0000000000000050000000000000004b00000000",
            INIT_20 => X"000000fe00000000000000fd00000000000000fc00000000000000f500000000",
            INIT_21 => X"000000c900000000000000ba00000000000000bb00000000000000f300000000",
            INIT_22 => X"0000009c00000000000000970000000000000080000000000000009100000000",
            INIT_23 => X"000000720000000000000080000000000000006a000000000000007400000000",
            INIT_24 => X"0000006700000000000000650000000000000067000000000000006800000000",
            INIT_25 => X"0000005c0000000000000069000000000000006e000000000000006c00000000",
            INIT_26 => X"000000550000000000000054000000000000004c000000000000005200000000",
            INIT_27 => X"00000049000000000000004d0000000000000053000000000000004e00000000",
            INIT_28 => X"0000010000000000000000fc00000000000000fc00000000000000fb00000000",
            INIT_29 => X"00000072000000000000006b000000000000007e00000000000000e900000000",
            INIT_2A => X"0000006e00000000000000780000000000000073000000000000006900000000",
            INIT_2B => X"0000006700000000000000680000000000000063000000000000006300000000",
            INIT_2C => X"0000006b000000000000006b000000000000006e000000000000006d00000000",
            INIT_2D => X"000000560000000000000060000000000000006e000000000000007000000000",
            INIT_2E => X"00000068000000000000005a000000000000004c000000000000004e00000000",
            INIT_2F => X"0000004f00000000000000520000000000000052000000000000005b00000000",
            INIT_30 => X"000000eb00000000000000f600000000000000f800000000000000f800000000",
            INIT_31 => X"000000760000000000000072000000000000007c00000000000000c800000000",
            INIT_32 => X"0000004f00000000000000530000000000000057000000000000005d00000000",
            INIT_33 => X"00000044000000000000004b0000000000000056000000000000005000000000",
            INIT_34 => X"0000006100000000000000620000000000000064000000000000005f00000000",
            INIT_35 => X"0000006100000000000000610000000000000061000000000000006200000000",
            INIT_36 => X"0000006f000000000000005b0000000000000057000000000000005b00000000",
            INIT_37 => X"0000005200000000000000520000000000000055000000000000006e00000000",
            INIT_38 => X"0000009600000000000000b500000000000000d600000000000000eb00000000",
            INIT_39 => X"0000008400000000000000850000000000000088000000000000008a00000000",
            INIT_3A => X"0000003c0000000000000039000000000000003d000000000000006400000000",
            INIT_3B => X"0000003a00000000000000600000000000000059000000000000004300000000",
            INIT_3C => X"0000005000000000000000470000000000000045000000000000003300000000",
            INIT_3D => X"0000006500000000000000680000000000000065000000000000005e00000000",
            INIT_3E => X"0000006d000000000000005e0000000000000057000000000000005d00000000",
            INIT_3F => X"0000005100000000000000510000000000000062000000000000007700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000078000000000000007a0000000000000082000000000000009900000000",
            INIT_41 => X"00000067000000000000006f000000000000007a000000000000007c00000000",
            INIT_42 => X"000000340000000000000039000000000000005a000000000000006a00000000",
            INIT_43 => X"00000053000000000000006a0000000000000066000000000000004500000000",
            INIT_44 => X"00000055000000000000004d0000000000000047000000000000004000000000",
            INIT_45 => X"0000006d00000000000000660000000000000067000000000000006400000000",
            INIT_46 => X"00000063000000000000005d0000000000000057000000000000006a00000000",
            INIT_47 => X"00000050000000000000005c0000000000000073000000000000007100000000",
            INIT_48 => X"0000006d0000000000000072000000000000006f000000000000006d00000000",
            INIT_49 => X"0000006d00000000000000660000000000000061000000000000006500000000",
            INIT_4A => X"0000005500000000000000670000000000000078000000000000007500000000",
            INIT_4B => X"00000059000000000000005f0000000000000065000000000000005d00000000",
            INIT_4C => X"0000005a0000000000000052000000000000004b000000000000004a00000000",
            INIT_4D => X"0000006600000000000000690000000000000077000000000000007200000000",
            INIT_4E => X"00000062000000000000005e000000000000006b000000000000006f00000000",
            INIT_4F => X"0000004f000000000000006b0000000000000075000000000000006500000000",
            INIT_50 => X"0000005b000000000000005d0000000000000062000000000000006900000000",
            INIT_51 => X"00000071000000000000006f000000000000006a000000000000006300000000",
            INIT_52 => X"0000005f00000000000000610000000000000068000000000000007000000000",
            INIT_53 => X"0000005c0000000000000054000000000000004c000000000000005000000000",
            INIT_54 => X"00000059000000000000004f0000000000000048000000000000005100000000",
            INIT_55 => X"0000005e0000000000000069000000000000007b000000000000007500000000",
            INIT_56 => X"0000006500000000000000670000000000000067000000000000006000000000",
            INIT_57 => X"0000005a000000000000006f0000000000000069000000000000006000000000",
            INIT_58 => X"00000065000000000000005e0000000000000057000000000000005700000000",
            INIT_59 => X"00000064000000000000006b000000000000006e000000000000006c00000000",
            INIT_5A => X"0000006800000000000000560000000000000051000000000000005b00000000",
            INIT_5B => X"0000005c000000000000004c0000000000000049000000000000005d00000000",
            INIT_5C => X"0000004f000000000000004f000000000000004d000000000000005800000000",
            INIT_5D => X"00000056000000000000005d0000000000000064000000000000005b00000000",
            INIT_5E => X"000000600000000000000061000000000000005c000000000000005700000000",
            INIT_5F => X"0000006500000000000000660000000000000060000000000000006000000000",
            INIT_60 => X"0000006900000000000000670000000000000060000000000000005a00000000",
            INIT_61 => X"000000500000000000000056000000000000005f000000000000006500000000",
            INIT_62 => X"0000006a00000000000000600000000000000055000000000000005100000000",
            INIT_63 => X"0000005d00000000000000600000000000000055000000000000006200000000",
            INIT_64 => X"0000004c000000000000004f0000000000000051000000000000005800000000",
            INIT_65 => X"0000005b0000000000000054000000000000004c000000000000004700000000",
            INIT_66 => X"0000005a00000000000000530000000000000056000000000000005c00000000",
            INIT_67 => X"00000060000000000000005b0000000000000060000000000000006200000000",
            INIT_68 => X"00000056000000000000005f0000000000000063000000000000006400000000",
            INIT_69 => X"0000004f000000000000004f000000000000004f000000000000005000000000",
            INIT_6A => X"0000006c00000000000000620000000000000053000000000000005200000000",
            INIT_6B => X"0000005900000000000000610000000000000060000000000000006300000000",
            INIT_6C => X"00000051000000000000004f0000000000000054000000000000005c00000000",
            INIT_6D => X"000000590000000000000052000000000000004a000000000000004c00000000",
            INIT_6E => X"0000005600000000000000520000000000000055000000000000005a00000000",
            INIT_6F => X"000000530000000000000053000000000000005c000000000000005d00000000",
            INIT_70 => X"000000470000000000000049000000000000004e000000000000005700000000",
            INIT_71 => X"0000005300000000000000590000000000000057000000000000004d00000000",
            INIT_72 => X"0000006a0000000000000061000000000000004f000000000000005100000000",
            INIT_73 => X"0000005c00000000000000590000000000000067000000000000006400000000",
            INIT_74 => X"0000005900000000000000580000000000000057000000000000006000000000",
            INIT_75 => X"000000530000000000000054000000000000004f000000000000005200000000",
            INIT_76 => X"000000530000000000000056000000000000005a000000000000005600000000",
            INIT_77 => X"00000049000000000000004f0000000000000056000000000000005600000000",
            INIT_78 => X"000000490000000000000046000000000000003f000000000000003e00000000",
            INIT_79 => X"0000005100000000000000530000000000000056000000000000005400000000",
            INIT_7A => X"0000006b000000000000005e000000000000004a000000000000004e00000000",
            INIT_7B => X"00000058000000000000005b0000000000000068000000000000005f00000000",
            INIT_7C => X"0000005900000000000000580000000000000058000000000000005b00000000",
            INIT_7D => X"0000005300000000000000550000000000000050000000000000005500000000",
            INIT_7E => X"0000005000000000000000560000000000000059000000000000005400000000",
            INIT_7F => X"00000048000000000000004c000000000000004d000000000000004c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE43;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE44 : if BRAM_NAME = "sampleifmap_layersamples_instance44" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000059000000000000005d000000000000005e000000000000005e00000000",
            INIT_01 => X"000000600000000000000060000000000000005a000000000000005a00000000",
            INIT_02 => X"00000065000000000000006e0000000000000066000000000000006100000000",
            INIT_03 => X"0000005200000000000000550000000000000058000000000000005e00000000",
            INIT_04 => X"000000480000000000000049000000000000004b000000000000004e00000000",
            INIT_05 => X"00000038000000000000003d0000000000000041000000000000004500000000",
            INIT_06 => X"000000270000000000000029000000000000002e000000000000003300000000",
            INIT_07 => X"00000019000000000000001d0000000000000022000000000000002800000000",
            INIT_08 => X"00000059000000000000005f000000000000005f000000000000006000000000",
            INIT_09 => X"00000062000000000000005f0000000000000059000000000000005900000000",
            INIT_0A => X"0000006b000000000000006a0000000000000060000000000000006100000000",
            INIT_0B => X"0000005200000000000000550000000000000059000000000000006000000000",
            INIT_0C => X"000000490000000000000047000000000000004b000000000000004f00000000",
            INIT_0D => X"00000035000000000000003b000000000000003d000000000000004400000000",
            INIT_0E => X"000000250000000000000027000000000000002c000000000000003100000000",
            INIT_0F => X"0000001f000000000000001f0000000000000020000000000000002600000000",
            INIT_10 => X"00000057000000000000005c000000000000005c000000000000005e00000000",
            INIT_11 => X"00000051000000000000005d000000000000005a000000000000005400000000",
            INIT_12 => X"0000006e00000000000000630000000000000060000000000000005900000000",
            INIT_13 => X"0000005400000000000000560000000000000062000000000000007000000000",
            INIT_14 => X"0000004600000000000000440000000000000049000000000000004f00000000",
            INIT_15 => X"000000300000000000000036000000000000003a000000000000003f00000000",
            INIT_16 => X"0000002b0000000000000029000000000000002b000000000000002e00000000",
            INIT_17 => X"000000310000000000000030000000000000002e000000000000002f00000000",
            INIT_18 => X"0000005a000000000000005c000000000000005d000000000000005f00000000",
            INIT_19 => X"000000390000000000000056000000000000005d000000000000005300000000",
            INIT_1A => X"000000680000000000000063000000000000006b000000000000005d00000000",
            INIT_1B => X"0000005a00000000000000650000000000000072000000000000007400000000",
            INIT_1C => X"0000004200000000000000420000000000000043000000000000004e00000000",
            INIT_1D => X"0000003900000000000000380000000000000038000000000000003e00000000",
            INIT_1E => X"000000420000000000000041000000000000003e000000000000003c00000000",
            INIT_1F => X"0000003d000000000000003f0000000000000041000000000000004300000000",
            INIT_20 => X"0000005b000000000000005b000000000000005b000000000000005c00000000",
            INIT_21 => X"0000003e00000000000000520000000000000059000000000000005300000000",
            INIT_22 => X"000000580000000000000058000000000000005f000000000000005c00000000",
            INIT_23 => X"0000006400000000000000690000000000000068000000000000005c00000000",
            INIT_24 => X"0000004800000000000000450000000000000046000000000000005b00000000",
            INIT_25 => X"000000530000000000000050000000000000004d000000000000005000000000",
            INIT_26 => X"0000005000000000000000510000000000000051000000000000005300000000",
            INIT_27 => X"0000003f0000000000000046000000000000004b000000000000004f00000000",
            INIT_28 => X"0000005900000000000000570000000000000056000000000000005800000000",
            INIT_29 => X"0000004d000000000000004c000000000000004f000000000000005200000000",
            INIT_2A => X"0000005700000000000000550000000000000052000000000000005000000000",
            INIT_2B => X"0000005f000000000000005e000000000000005e000000000000005a00000000",
            INIT_2C => X"000000630000000000000062000000000000005e000000000000006300000000",
            INIT_2D => X"0000006200000000000000600000000000000064000000000000006400000000",
            INIT_2E => X"0000005300000000000000580000000000000058000000000000005d00000000",
            INIT_2F => X"00000037000000000000003e0000000000000045000000000000004c00000000",
            INIT_30 => X"0000005400000000000000520000000000000054000000000000005500000000",
            INIT_31 => X"00000037000000000000002a000000000000003d000000000000005100000000",
            INIT_32 => X"0000005900000000000000580000000000000057000000000000005300000000",
            INIT_33 => X"00000065000000000000005d0000000000000057000000000000005b00000000",
            INIT_34 => X"0000007300000000000000700000000000000064000000000000006200000000",
            INIT_35 => X"0000006700000000000000670000000000000067000000000000006900000000",
            INIT_36 => X"0000004a000000000000004e0000000000000050000000000000005b00000000",
            INIT_37 => X"000000360000000000000039000000000000003f000000000000004400000000",
            INIT_38 => X"0000005400000000000000520000000000000053000000000000005200000000",
            INIT_39 => X"0000002c00000000000000260000000000000037000000000000004c00000000",
            INIT_3A => X"0000005100000000000000520000000000000055000000000000004c00000000",
            INIT_3B => X"00000063000000000000005b0000000000000053000000000000005000000000",
            INIT_3C => X"0000006c00000000000000610000000000000060000000000000006700000000",
            INIT_3D => X"0000005e00000000000000710000000000000072000000000000006d00000000",
            INIT_3E => X"0000004b000000000000004d000000000000004d000000000000005200000000",
            INIT_3F => X"0000003b00000000000000400000000000000044000000000000004700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005b00000000000000540000000000000052000000000000005100000000",
            INIT_41 => X"0000003100000000000000550000000000000068000000000000005e00000000",
            INIT_42 => X"00000063000000000000005b0000000000000054000000000000004900000000",
            INIT_43 => X"0000005e00000000000000650000000000000064000000000000006100000000",
            INIT_44 => X"0000006200000000000000650000000000000068000000000000006500000000",
            INIT_45 => X"000000670000000000000072000000000000006f000000000000006a00000000",
            INIT_46 => X"0000004e00000000000000520000000000000055000000000000005700000000",
            INIT_47 => X"0000004800000000000000470000000000000046000000000000004a00000000",
            INIT_48 => X"0000008000000000000000730000000000000065000000000000005c00000000",
            INIT_49 => X"000000360000000000000068000000000000009d000000000000008e00000000",
            INIT_4A => X"00000071000000000000005d0000000000000054000000000000004b00000000",
            INIT_4B => X"000000650000000000000075000000000000007c000000000000007500000000",
            INIT_4C => X"00000067000000000000006b000000000000006a000000000000006700000000",
            INIT_4D => X"000000760000000000000074000000000000006e000000000000006800000000",
            INIT_4E => X"000000540000000000000055000000000000005a000000000000006400000000",
            INIT_4F => X"0000005200000000000000550000000000000055000000000000005500000000",
            INIT_50 => X"000000a00000000000000099000000000000008e000000000000008200000000",
            INIT_51 => X"00000035000000000000005900000000000000aa00000000000000a600000000",
            INIT_52 => X"000000680000000000000046000000000000004d000000000000005000000000",
            INIT_53 => X"0000006b000000000000007f0000000000000082000000000000007700000000",
            INIT_54 => X"0000006a0000000000000069000000000000006c000000000000006a00000000",
            INIT_55 => X"00000072000000000000006e0000000000000069000000000000006a00000000",
            INIT_56 => X"0000006000000000000000620000000000000062000000000000006900000000",
            INIT_57 => X"000000550000000000000059000000000000005b000000000000005e00000000",
            INIT_58 => X"000000a400000000000000a2000000000000009f000000000000009a00000000",
            INIT_59 => X"0000002e000000000000005d00000000000000a900000000000000a700000000",
            INIT_5A => X"00000067000000000000004a0000000000000056000000000000005100000000",
            INIT_5B => X"00000072000000000000007a0000000000000070000000000000007b00000000",
            INIT_5C => X"00000067000000000000006a000000000000006d000000000000006a00000000",
            INIT_5D => X"0000006e00000000000000670000000000000069000000000000006b00000000",
            INIT_5E => X"0000006300000000000000650000000000000061000000000000006600000000",
            INIT_5F => X"00000055000000000000005a000000000000005e000000000000006000000000",
            INIT_60 => X"0000009e00000000000000a1000000000000009f000000000000009d00000000",
            INIT_61 => X"000000300000000000000075000000000000009f000000000000009e00000000",
            INIT_62 => X"00000078000000000000006c0000000000000065000000000000004900000000",
            INIT_63 => X"0000007500000000000000740000000000000078000000000000008700000000",
            INIT_64 => X"00000066000000000000006c0000000000000073000000000000006b00000000",
            INIT_65 => X"000000690000000000000064000000000000006a000000000000006900000000",
            INIT_66 => X"0000006500000000000000600000000000000060000000000000007000000000",
            INIT_67 => X"0000004c0000000000000055000000000000005d000000000000006200000000",
            INIT_68 => X"0000009300000000000000970000000000000098000000000000009900000000",
            INIT_69 => X"0000004c00000000000000870000000000000093000000000000009300000000",
            INIT_6A => X"0000007500000000000000670000000000000049000000000000002c00000000",
            INIT_6B => X"0000007100000000000000730000000000000085000000000000008300000000",
            INIT_6C => X"0000006b00000000000000710000000000000077000000000000006c00000000",
            INIT_6D => X"000000640000000000000065000000000000006a000000000000006a00000000",
            INIT_6E => X"00000062000000000000005d0000000000000069000000000000007500000000",
            INIT_6F => X"00000040000000000000004a0000000000000055000000000000005d00000000",
            INIT_70 => X"0000008e000000000000008e000000000000008e000000000000008f00000000",
            INIT_71 => X"0000008300000000000000950000000000000094000000000000008f00000000",
            INIT_72 => X"0000004600000000000000350000000000000041000000000000005400000000",
            INIT_73 => X"0000006d0000000000000068000000000000006b000000000000006300000000",
            INIT_74 => X"00000075000000000000007d000000000000007c000000000000007200000000",
            INIT_75 => X"000000620000000000000065000000000000006c000000000000006e00000000",
            INIT_76 => X"0000005a0000000000000058000000000000006f000000000000006c00000000",
            INIT_77 => X"0000003f00000000000000410000000000000048000000000000005500000000",
            INIT_78 => X"00000091000000000000008e000000000000008d000000000000008c00000000",
            INIT_79 => X"00000093000000000000009900000000000000a0000000000000009900000000",
            INIT_7A => X"0000003a0000000000000034000000000000006f000000000000009700000000",
            INIT_7B => X"0000006e00000000000000650000000000000068000000000000006a00000000",
            INIT_7C => X"0000008000000000000000870000000000000089000000000000007b00000000",
            INIT_7D => X"000000650000000000000068000000000000006c000000000000007300000000",
            INIT_7E => X"0000004e0000000000000059000000000000006f000000000000006300000000",
            INIT_7F => X"0000004d000000000000004a0000000000000048000000000000004a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE44;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE45 : if BRAM_NAME = "sampleifmap_layersamples_instance45" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009f000000000000009b0000000000000095000000000000008f00000000",
            INIT_01 => X"00000072000000000000008800000000000000a000000000000000a400000000",
            INIT_02 => X"00000068000000000000007a000000000000008f000000000000009b00000000",
            INIT_03 => X"0000006c00000000000000660000000000000077000000000000007600000000",
            INIT_04 => X"0000008000000000000000850000000000000084000000000000007800000000",
            INIT_05 => X"0000006a000000000000006b000000000000006d000000000000007500000000",
            INIT_06 => X"000000560000000000000062000000000000006c000000000000006100000000",
            INIT_07 => X"00000044000000000000004f0000000000000054000000000000005a00000000",
            INIT_08 => X"000000a1000000000000009f000000000000009d000000000000009a00000000",
            INIT_09 => X"0000008100000000000000b000000000000000b100000000000000a700000000",
            INIT_0A => X"0000008e000000000000009700000000000000c700000000000000b300000000",
            INIT_0B => X"0000006c000000000000007b0000000000000089000000000000006800000000",
            INIT_0C => X"000000800000000000000083000000000000007e000000000000007900000000",
            INIT_0D => X"0000006e00000000000000700000000000000073000000000000007700000000",
            INIT_0E => X"0000005e000000000000006a0000000000000069000000000000006300000000",
            INIT_0F => X"000000270000000000000034000000000000004a000000000000005c00000000",
            INIT_10 => X"000000c100000000000000b000000000000000a4000000000000009d00000000",
            INIT_11 => X"000000c700000000000000f700000000000000ec00000000000000da00000000",
            INIT_12 => X"000000b100000000000000ad00000000000000ce00000000000000a300000000",
            INIT_13 => X"0000007100000000000000860000000000000088000000000000006500000000",
            INIT_14 => X"000000810000000000000082000000000000007e000000000000007700000000",
            INIT_15 => X"000000710000000000000076000000000000007a000000000000007d00000000",
            INIT_16 => X"00000050000000000000006a0000000000000067000000000000006800000000",
            INIT_17 => X"000000270000000000000025000000000000002c000000000000003e00000000",
            INIT_18 => X"000000f600000000000000e800000000000000d400000000000000c000000000",
            INIT_19 => X"000000f700000000000000fa00000000000000f200000000000000fa00000000",
            INIT_1A => X"000000c100000000000000ae00000000000000aa00000000000000a900000000",
            INIT_1B => X"00000078000000000000008b0000000000000070000000000000006e00000000",
            INIT_1C => X"000000800000000000000080000000000000007e000000000000007600000000",
            INIT_1D => X"00000074000000000000007e000000000000007f000000000000008000000000",
            INIT_1E => X"0000003e00000000000000600000000000000066000000000000006c00000000",
            INIT_1F => X"0000002b00000000000000270000000000000025000000000000002a00000000",
            INIT_20 => X"000000fb00000000000000fa00000000000000fb00000000000000f500000000",
            INIT_21 => X"000000d200000000000000be00000000000000ba00000000000000f100000000",
            INIT_22 => X"000000a0000000000000009c000000000000009200000000000000a100000000",
            INIT_23 => X"0000007a00000000000000870000000000000073000000000000007d00000000",
            INIT_24 => X"000000800000000000000081000000000000007f000000000000007800000000",
            INIT_25 => X"00000074000000000000007d000000000000007f000000000000007f00000000",
            INIT_26 => X"0000004200000000000000570000000000000062000000000000006a00000000",
            INIT_27 => X"000000290000000000000029000000000000002a000000000000002d00000000",
            INIT_28 => X"000000fe00000000000000fb00000000000000fb00000000000000fb00000000",
            INIT_29 => X"000000820000000000000074000000000000008300000000000000ea00000000",
            INIT_2A => X"0000007c0000000000000082000000000000008a000000000000007f00000000",
            INIT_2B => X"0000006b00000000000000720000000000000077000000000000007a00000000",
            INIT_2C => X"0000007f00000000000000820000000000000080000000000000007600000000",
            INIT_2D => X"0000006c000000000000006f0000000000000077000000000000007d00000000",
            INIT_2E => X"000000500000000000000052000000000000005a000000000000006300000000",
            INIT_2F => X"00000029000000000000002c000000000000002f000000000000003d00000000",
            INIT_30 => X"000000ef00000000000000f900000000000000fc00000000000000fc00000000",
            INIT_31 => X"00000083000000000000007b000000000000008000000000000000cb00000000",
            INIT_32 => X"000000670000000000000066000000000000006c000000000000006f00000000",
            INIT_33 => X"0000004400000000000000510000000000000069000000000000006a00000000",
            INIT_34 => X"0000007400000000000000780000000000000075000000000000006600000000",
            INIT_35 => X"000000730000000000000070000000000000006b000000000000006e00000000",
            INIT_36 => X"00000054000000000000004b0000000000000059000000000000006800000000",
            INIT_37 => X"0000002d000000000000002d0000000000000034000000000000005100000000",
            INIT_38 => X"000000a000000000000000bf00000000000000df00000000000000f500000000",
            INIT_39 => X"0000008a00000000000000890000000000000089000000000000009000000000",
            INIT_3A => X"000000570000000000000051000000000000004b000000000000006d00000000",
            INIT_3B => X"0000003a00000000000000630000000000000066000000000000005a00000000",
            INIT_3C => X"00000065000000000000005f0000000000000056000000000000003a00000000",
            INIT_3D => X"00000074000000000000007a0000000000000074000000000000006d00000000",
            INIT_3E => X"000000500000000000000046000000000000004d000000000000006100000000",
            INIT_3F => X"0000002f000000000000002f0000000000000042000000000000005900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000840000000000000086000000000000008d00000000000000a500000000",
            INIT_41 => X"000000690000000000000070000000000000007b000000000000008200000000",
            INIT_42 => X"00000047000000000000004a000000000000005e000000000000006b00000000",
            INIT_43 => X"00000056000000000000006f000000000000006e000000000000005300000000",
            INIT_44 => X"0000006c0000000000000066000000000000005a000000000000004800000000",
            INIT_45 => X"0000007c000000000000007b000000000000007b000000000000007600000000",
            INIT_46 => X"0000004400000000000000420000000000000049000000000000006c00000000",
            INIT_47 => X"00000030000000000000003d0000000000000054000000000000005200000000",
            INIT_48 => X"00000075000000000000007a0000000000000078000000000000007500000000",
            INIT_49 => X"0000006a00000000000000650000000000000061000000000000006a00000000",
            INIT_4A => X"00000057000000000000006a0000000000000073000000000000007000000000",
            INIT_4B => X"0000006100000000000000680000000000000068000000000000005c00000000",
            INIT_4C => X"00000072000000000000006c000000000000005f000000000000005400000000",
            INIT_4D => X"0000007a0000000000000082000000000000008e000000000000008600000000",
            INIT_4E => X"0000004000000000000000450000000000000064000000000000007700000000",
            INIT_4F => X"00000032000000000000004f0000000000000057000000000000004500000000",
            INIT_50 => X"0000005e00000000000000600000000000000066000000000000006c00000000",
            INIT_51 => X"0000006b000000000000006e000000000000006b000000000000006500000000",
            INIT_52 => X"000000510000000000000056000000000000005d000000000000006700000000",
            INIT_53 => X"00000068000000000000005d0000000000000048000000000000004200000000",
            INIT_54 => X"00000071000000000000006b000000000000005f000000000000005e00000000",
            INIT_55 => X"0000007a00000000000000850000000000000094000000000000008900000000",
            INIT_56 => X"000000420000000000000051000000000000006b000000000000007200000000",
            INIT_57 => X"0000003f0000000000000055000000000000004b000000000000004000000000",
            INIT_58 => X"00000063000000000000005d0000000000000057000000000000005800000000",
            INIT_59 => X"000000570000000000000065000000000000006c000000000000006b00000000",
            INIT_5A => X"000000530000000000000041000000000000003c000000000000004900000000",
            INIT_5B => X"0000005e000000000000004e000000000000003f000000000000004a00000000",
            INIT_5C => X"0000005d000000000000005f0000000000000057000000000000005900000000",
            INIT_5D => X"00000072000000000000007a000000000000007b000000000000006900000000",
            INIT_5E => X"0000003b000000000000004e0000000000000068000000000000006d00000000",
            INIT_5F => X"0000004b000000000000004a000000000000003f000000000000003c00000000",
            INIT_60 => X"0000005f0000000000000061000000000000005f000000000000005d00000000",
            INIT_61 => X"0000003800000000000000450000000000000054000000000000005b00000000",
            INIT_62 => X"0000005500000000000000420000000000000031000000000000003200000000",
            INIT_63 => X"0000004800000000000000550000000000000049000000000000005300000000",
            INIT_64 => X"000000440000000000000043000000000000003e000000000000003e00000000",
            INIT_65 => X"0000006800000000000000640000000000000058000000000000004500000000",
            INIT_66 => X"000000330000000000000040000000000000005a000000000000006500000000",
            INIT_67 => X"00000045000000000000003a0000000000000036000000000000003500000000",
            INIT_68 => X"000000440000000000000051000000000000005b000000000000006000000000",
            INIT_69 => X"0000003000000000000000340000000000000037000000000000003b00000000",
            INIT_6A => X"000000520000000000000040000000000000002e000000000000002f00000000",
            INIT_6B => X"00000039000000000000004d000000000000004f000000000000005200000000",
            INIT_6C => X"0000003a00000000000000340000000000000032000000000000003500000000",
            INIT_6D => X"0000004a0000000000000047000000000000003f000000000000003a00000000",
            INIT_6E => X"0000002e00000000000000340000000000000041000000000000004800000000",
            INIT_6F => X"0000003600000000000000300000000000000031000000000000003000000000",
            INIT_70 => X"0000002b0000000000000031000000000000003c000000000000004900000000",
            INIT_71 => X"0000003000000000000000340000000000000030000000000000002c00000000",
            INIT_72 => X"00000049000000000000003a000000000000002c000000000000003000000000",
            INIT_73 => X"00000035000000000000003e000000000000004f000000000000004b00000000",
            INIT_74 => X"000000390000000000000034000000000000002e000000000000003200000000",
            INIT_75 => X"0000002f0000000000000033000000000000002f000000000000003400000000",
            INIT_76 => X"0000002a000000000000002e0000000000000031000000000000002f00000000",
            INIT_77 => X"0000002a000000000000002b000000000000002d000000000000002b00000000",
            INIT_78 => X"0000002500000000000000270000000000000025000000000000002900000000",
            INIT_79 => X"0000002d00000000000000290000000000000029000000000000002a00000000",
            INIT_7A => X"000000470000000000000036000000000000002b000000000000002f00000000",
            INIT_7B => X"0000002e000000000000003b000000000000004c000000000000004300000000",
            INIT_7C => X"00000030000000000000002d000000000000002a000000000000002b00000000",
            INIT_7D => X"0000002d0000000000000031000000000000002d000000000000002f00000000",
            INIT_7E => X"00000027000000000000002a000000000000002d000000000000002b00000000",
            INIT_7F => X"0000002600000000000000280000000000000028000000000000002500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE45;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE46 : if BRAM_NAME = "sampleifmap_layersamples_instance46" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004f00000000000000530000000000000054000000000000005500000000",
            INIT_01 => X"0000005f000000000000005d0000000000000052000000000000005000000000",
            INIT_02 => X"00000048000000000000004f0000000000000055000000000000005a00000000",
            INIT_03 => X"0000004f0000000000000054000000000000004e000000000000004b00000000",
            INIT_04 => X"0000003d000000000000003c000000000000003e000000000000004400000000",
            INIT_05 => X"000000330000000000000038000000000000003b000000000000003c00000000",
            INIT_06 => X"0000002300000000000000250000000000000029000000000000002e00000000",
            INIT_07 => X"000000150000000000000019000000000000001e000000000000002400000000",
            INIT_08 => X"0000004f00000000000000550000000000000055000000000000005600000000",
            INIT_09 => X"0000005d000000000000005a0000000000000050000000000000004e00000000",
            INIT_0A => X"0000004700000000000000460000000000000049000000000000005400000000",
            INIT_0B => X"0000004800000000000000470000000000000045000000000000004400000000",
            INIT_0C => X"0000003e000000000000003e0000000000000043000000000000004600000000",
            INIT_0D => X"0000002e00000000000000340000000000000035000000000000003800000000",
            INIT_0E => X"0000002000000000000000220000000000000025000000000000002900000000",
            INIT_0F => X"0000001b000000000000001a000000000000001b000000000000002100000000",
            INIT_10 => X"0000004e00000000000000520000000000000053000000000000005400000000",
            INIT_11 => X"0000004800000000000000560000000000000050000000000000004900000000",
            INIT_12 => X"0000004300000000000000380000000000000041000000000000004600000000",
            INIT_13 => X"0000003c0000000000000036000000000000003f000000000000004800000000",
            INIT_14 => X"0000003a000000000000003d0000000000000041000000000000004200000000",
            INIT_15 => X"00000026000000000000002d000000000000002f000000000000003000000000",
            INIT_16 => X"0000002500000000000000220000000000000021000000000000002400000000",
            INIT_17 => X"0000002c000000000000002a0000000000000029000000000000002a00000000",
            INIT_18 => X"0000005000000000000000520000000000000053000000000000005500000000",
            INIT_19 => X"0000002b000000000000004d0000000000000052000000000000004800000000",
            INIT_1A => X"0000003400000000000000320000000000000045000000000000004300000000",
            INIT_1B => X"0000002f0000000000000032000000000000003f000000000000004100000000",
            INIT_1C => X"0000003600000000000000390000000000000034000000000000003200000000",
            INIT_1D => X"0000002c000000000000002b000000000000002b000000000000002d00000000",
            INIT_1E => X"0000003b00000000000000380000000000000032000000000000002f00000000",
            INIT_1F => X"000000370000000000000038000000000000003b000000000000003c00000000",
            INIT_20 => X"0000005100000000000000510000000000000051000000000000005200000000",
            INIT_21 => X"0000002c0000000000000046000000000000004c000000000000004800000000",
            INIT_22 => X"0000001d00000000000000220000000000000033000000000000003d00000000",
            INIT_23 => X"0000002300000000000000260000000000000027000000000000001f00000000",
            INIT_24 => X"0000003b0000000000000039000000000000002b000000000000002900000000",
            INIT_25 => X"000000440000000000000041000000000000003d000000000000003d00000000",
            INIT_26 => X"0000004800000000000000470000000000000042000000000000004400000000",
            INIT_27 => X"00000038000000000000003e0000000000000043000000000000004700000000",
            INIT_28 => X"0000004f000000000000004c000000000000004c000000000000004d00000000",
            INIT_29 => X"00000038000000000000003e0000000000000042000000000000004700000000",
            INIT_2A => X"00000017000000000000001a0000000000000021000000000000002c00000000",
            INIT_2B => X"0000000e000000000000000f0000000000000014000000000000001600000000",
            INIT_2C => X"00000054000000000000004f0000000000000035000000000000001f00000000",
            INIT_2D => X"00000050000000000000004e0000000000000052000000000000005300000000",
            INIT_2E => X"0000004b000000000000004d0000000000000048000000000000004c00000000",
            INIT_2F => X"0000002e0000000000000035000000000000003c000000000000004400000000",
            INIT_30 => X"0000004800000000000000460000000000000047000000000000004900000000",
            INIT_31 => X"0000002000000000000000200000000000000037000000000000004700000000",
            INIT_32 => X"0000001300000000000000140000000000000018000000000000002600000000",
            INIT_33 => X"00000015000000000000000e000000000000000b000000000000001200000000",
            INIT_34 => X"0000005900000000000000460000000000000029000000000000001800000000",
            INIT_35 => X"00000052000000000000004f0000000000000050000000000000005600000000",
            INIT_36 => X"0000004300000000000000480000000000000048000000000000004b00000000",
            INIT_37 => X"0000002a000000000000002d0000000000000034000000000000003b00000000",
            INIT_38 => X"0000004500000000000000440000000000000045000000000000004400000000",
            INIT_39 => X"00000011000000000000001c0000000000000033000000000000004300000000",
            INIT_3A => X"0000000b000000000000000a000000000000000c000000000000001700000000",
            INIT_3B => X"000000180000000000000011000000000000000b000000000000000900000000",
            INIT_3C => X"0000003f00000000000000210000000000000016000000000000001c00000000",
            INIT_3D => X"00000040000000000000004d000000000000004f000000000000004d00000000",
            INIT_3E => X"0000004200000000000000480000000000000049000000000000004100000000",
            INIT_3F => X"0000002b000000000000002f0000000000000036000000000000003c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004e00000000000000470000000000000045000000000000004400000000",
            INIT_41 => X"000000130000000000000046000000000000005d000000000000005200000000",
            INIT_42 => X"000000250000000000000019000000000000000c000000000000001200000000",
            INIT_43 => X"0000001400000000000000210000000000000021000000000000002000000000",
            INIT_44 => X"0000002100000000000000190000000000000018000000000000001600000000",
            INIT_45 => X"0000003b000000000000003c0000000000000038000000000000003100000000",
            INIT_46 => X"0000003f0000000000000049000000000000004b000000000000003b00000000",
            INIT_47 => X"0000003500000000000000340000000000000034000000000000003900000000",
            INIT_48 => X"0000007500000000000000670000000000000059000000000000005000000000",
            INIT_49 => X"000000160000000000000055000000000000008d000000000000008000000000",
            INIT_4A => X"000000380000000000000021000000000000000f000000000000001500000000",
            INIT_4B => X"0000001c0000000000000035000000000000003d000000000000003900000000",
            INIT_4C => X"0000001400000000000000160000000000000016000000000000001500000000",
            INIT_4D => X"0000003a000000000000002d0000000000000023000000000000001800000000",
            INIT_4E => X"0000004100000000000000460000000000000048000000000000003d00000000",
            INIT_4F => X"0000003d000000000000003f0000000000000040000000000000004100000000",
            INIT_50 => X"00000095000000000000008e0000000000000083000000000000007700000000",
            INIT_51 => X"0000001800000000000000470000000000000098000000000000009800000000",
            INIT_52 => X"0000003100000000000000150000000000000011000000000000001e00000000",
            INIT_53 => X"00000021000000000000003f0000000000000044000000000000003c00000000",
            INIT_54 => X"000000110000000000000015000000000000001b000000000000001900000000",
            INIT_55 => X"0000002b000000000000001c0000000000000014000000000000000f00000000",
            INIT_56 => X"0000004a000000000000004d0000000000000046000000000000003700000000",
            INIT_57 => X"0000004100000000000000440000000000000047000000000000004900000000",
            INIT_58 => X"0000009900000000000000960000000000000094000000000000008f00000000",
            INIT_59 => X"00000017000000000000004f0000000000000099000000000000009900000000",
            INIT_5A => X"0000002e00000000000000190000000000000022000000000000002800000000",
            INIT_5B => X"0000002700000000000000370000000000000030000000000000003d00000000",
            INIT_5C => X"00000015000000000000001f0000000000000024000000000000001d00000000",
            INIT_5D => X"0000001f00000000000000120000000000000015000000000000001300000000",
            INIT_5E => X"0000004d000000000000004c000000000000003b000000000000002a00000000",
            INIT_5F => X"00000045000000000000004a000000000000004c000000000000004d00000000",
            INIT_60 => X"0000009400000000000000970000000000000095000000000000009200000000",
            INIT_61 => X"00000020000000000000006b0000000000000092000000000000009200000000",
            INIT_62 => X"0000003b00000000000000340000000000000037000000000000002b00000000",
            INIT_63 => X"00000029000000000000002c0000000000000034000000000000004700000000",
            INIT_64 => X"0000001e000000000000002c0000000000000032000000000000002200000000",
            INIT_65 => X"000000190000000000000012000000000000001c000000000000001a00000000",
            INIT_66 => X"0000005100000000000000450000000000000032000000000000002e00000000",
            INIT_67 => X"000000420000000000000049000000000000004f000000000000005100000000",
            INIT_68 => X"0000008b000000000000008f000000000000008f000000000000009000000000",
            INIT_69 => X"00000040000000000000007e0000000000000089000000000000008a00000000",
            INIT_6A => X"00000041000000000000003d000000000000002e000000000000001a00000000",
            INIT_6B => X"0000002400000000000000280000000000000040000000000000004600000000",
            INIT_6C => X"0000002800000000000000330000000000000036000000000000002400000000",
            INIT_6D => X"000000130000000000000012000000000000001d000000000000002100000000",
            INIT_6E => X"0000004e000000000000003c0000000000000033000000000000002f00000000",
            INIT_6F => X"000000370000000000000040000000000000004a000000000000004f00000000",
            INIT_70 => X"0000008600000000000000860000000000000084000000000000008500000000",
            INIT_71 => X"0000007700000000000000890000000000000088000000000000008600000000",
            INIT_72 => X"00000021000000000000001b0000000000000031000000000000004700000000",
            INIT_73 => X"000000220000000000000020000000000000002a000000000000002e00000000",
            INIT_74 => X"00000032000000000000003d0000000000000039000000000000002800000000",
            INIT_75 => X"000000110000000000000011000000000000001c000000000000002700000000",
            INIT_76 => X"0000004100000000000000300000000000000033000000000000002400000000",
            INIT_77 => X"000000320000000000000036000000000000003e000000000000004600000000",
            INIT_78 => X"000000850000000000000081000000000000007f000000000000007d00000000",
            INIT_79 => X"0000008100000000000000880000000000000091000000000000008c00000000",
            INIT_7A => X"0000001e000000000000001e000000000000005a000000000000008400000000",
            INIT_7B => X"0000002700000000000000270000000000000033000000000000004000000000",
            INIT_7C => X"0000003d00000000000000450000000000000045000000000000003100000000",
            INIT_7D => X"000000130000000000000014000000000000001c000000000000002c00000000",
            INIT_7E => X"0000002d00000000000000290000000000000030000000000000001900000000",
            INIT_7F => X"0000003d000000000000003c0000000000000039000000000000003500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE46;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE47 : if BRAM_NAME = "sampleifmap_layersamples_instance47" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000091000000000000008b0000000000000084000000000000007d00000000",
            INIT_01 => X"0000005a00000000000000750000000000000091000000000000009500000000",
            INIT_02 => X"0000005000000000000000620000000000000072000000000000008000000000",
            INIT_03 => X"000000280000000000000031000000000000004d000000000000005700000000",
            INIT_04 => X"0000003c0000000000000044000000000000003f000000000000002e00000000",
            INIT_05 => X"000000170000000000000019000000000000001f000000000000002d00000000",
            INIT_06 => X"0000002d000000000000002b000000000000002a000000000000001500000000",
            INIT_07 => X"00000032000000000000003e0000000000000042000000000000004000000000",
            INIT_08 => X"000000930000000000000090000000000000008c000000000000008800000000",
            INIT_09 => X"00000068000000000000009e00000000000000a4000000000000009a00000000",
            INIT_0A => X"00000077000000000000007a00000000000000a6000000000000009500000000",
            INIT_0B => X"00000029000000000000004b0000000000000067000000000000005000000000",
            INIT_0C => X"0000003c00000000000000410000000000000038000000000000002d00000000",
            INIT_0D => X"0000001b000000000000001f0000000000000028000000000000003000000000",
            INIT_0E => X"00000032000000000000002f0000000000000023000000000000001500000000",
            INIT_0F => X"0000001400000000000000230000000000000039000000000000004100000000",
            INIT_10 => X"000000b600000000000000a40000000000000097000000000000009000000000",
            INIT_11 => X"000000b200000000000000eb00000000000000e600000000000000d200000000",
            INIT_12 => X"00000095000000000000008a00000000000000ab000000000000008500000000",
            INIT_13 => X"0000002d00000000000000550000000000000067000000000000004d00000000",
            INIT_14 => X"0000003c000000000000003f0000000000000038000000000000002b00000000",
            INIT_15 => X"0000001d00000000000000270000000000000030000000000000003500000000",
            INIT_16 => X"00000027000000000000002f000000000000001d000000000000001700000000",
            INIT_17 => X"000000150000000000000016000000000000001f000000000000002700000000",
            INIT_18 => X"000000f000000000000000e100000000000000cd00000000000000b700000000",
            INIT_19 => X"000000e600000000000000f200000000000000f200000000000000f800000000",
            INIT_1A => X"0000009f00000000000000840000000000000084000000000000008d00000000",
            INIT_1B => X"000000310000000000000056000000000000004d000000000000005300000000",
            INIT_1C => X"0000003a000000000000003c0000000000000037000000000000002a00000000",
            INIT_1D => X"00000021000000000000002f0000000000000037000000000000003900000000",
            INIT_1E => X"0000001c0000000000000027000000000000001a000000000000001900000000",
            INIT_1F => X"0000001b000000000000001c000000000000001d000000000000001900000000",
            INIT_20 => X"000000f900000000000000f700000000000000f800000000000000f100000000",
            INIT_21 => X"000000b500000000000000ab00000000000000b000000000000000ec00000000",
            INIT_22 => X"0000007600000000000000720000000000000062000000000000007800000000",
            INIT_23 => X"000000340000000000000047000000000000003c000000000000004d00000000",
            INIT_24 => X"0000003a00000000000000390000000000000036000000000000002e00000000",
            INIT_25 => X"0000002000000000000000300000000000000039000000000000003b00000000",
            INIT_26 => X"0000002500000000000000250000000000000017000000000000001800000000",
            INIT_27 => X"0000001a000000000000001f0000000000000020000000000000001c00000000",
            INIT_28 => X"000000fd00000000000000f900000000000000f900000000000000f800000000",
            INIT_29 => X"000000550000000000000053000000000000006a00000000000000e000000000",
            INIT_2A => X"000000410000000000000051000000000000004e000000000000004700000000",
            INIT_2B => X"000000310000000000000034000000000000002e000000000000003000000000",
            INIT_2C => X"0000003900000000000000360000000000000037000000000000003300000000",
            INIT_2D => X"0000001b00000000000000240000000000000033000000000000003d00000000",
            INIT_2E => X"0000003600000000000000270000000000000016000000000000001500000000",
            INIT_2F => X"0000001c000000000000001f000000000000001f000000000000002800000000",
            INIT_30 => X"000000eb00000000000000f500000000000000f800000000000000f700000000",
            INIT_31 => X"0000005e0000000000000060000000000000006d00000000000000c200000000",
            INIT_32 => X"0000001900000000000000230000000000000035000000000000004100000000",
            INIT_33 => X"00000020000000000000002d000000000000002b000000000000001c00000000",
            INIT_34 => X"0000002f000000000000002f0000000000000033000000000000002e00000000",
            INIT_35 => X"00000029000000000000002b000000000000002d000000000000003000000000",
            INIT_36 => X"0000003a0000000000000024000000000000001e000000000000002200000000",
            INIT_37 => X"0000001e000000000000001d0000000000000021000000000000003900000000",
            INIT_38 => X"0000009800000000000000b600000000000000d700000000000000ec00000000",
            INIT_39 => X"00000074000000000000007a0000000000000081000000000000008800000000",
            INIT_3A => X"00000009000000000000000d0000000000000023000000000000005100000000",
            INIT_3B => X"0000002200000000000000490000000000000034000000000000001400000000",
            INIT_3C => X"00000020000000000000001a000000000000001c000000000000001100000000",
            INIT_3D => X"00000031000000000000003b000000000000003b000000000000002f00000000",
            INIT_3E => X"000000340000000000000022000000000000001a000000000000002300000000",
            INIT_3F => X"0000001d000000000000001c000000000000002c000000000000003f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000078000000000000007a0000000000000082000000000000009a00000000",
            INIT_41 => X"0000005c00000000000000680000000000000076000000000000007b00000000",
            INIT_42 => X"00000012000000000000001f0000000000000046000000000000005a00000000",
            INIT_43 => X"000000340000000000000045000000000000003d000000000000001d00000000",
            INIT_44 => X"0000002800000000000000240000000000000024000000000000002200000000",
            INIT_45 => X"0000003d00000000000000410000000000000047000000000000003a00000000",
            INIT_46 => X"00000028000000000000001f0000000000000017000000000000003000000000",
            INIT_47 => X"0000001c0000000000000027000000000000003c000000000000003800000000",
            INIT_48 => X"00000068000000000000006d000000000000006b000000000000006900000000",
            INIT_49 => X"0000005d000000000000005b0000000000000058000000000000005f00000000",
            INIT_4A => X"0000003e00000000000000560000000000000062000000000000006000000000",
            INIT_4B => X"00000031000000000000002f0000000000000038000000000000003800000000",
            INIT_4C => X"00000030000000000000002a0000000000000025000000000000002800000000",
            INIT_4D => X"000000390000000000000048000000000000005b000000000000004c00000000",
            INIT_4E => X"00000023000000000000001d000000000000002c000000000000003600000000",
            INIT_4F => X"0000001d0000000000000037000000000000003d000000000000002a00000000",
            INIT_50 => X"0000005100000000000000530000000000000059000000000000005f00000000",
            INIT_51 => X"00000058000000000000005b0000000000000058000000000000005600000000",
            INIT_52 => X"0000003e00000000000000440000000000000049000000000000005300000000",
            INIT_53 => X"00000034000000000000002c0000000000000023000000000000002800000000",
            INIT_54 => X"000000310000000000000027000000000000001e000000000000002800000000",
            INIT_55 => X"000000320000000000000047000000000000005f000000000000005100000000",
            INIT_56 => X"000000230000000000000025000000000000002a000000000000002900000000",
            INIT_57 => X"00000028000000000000003a0000000000000030000000000000002200000000",
            INIT_58 => X"00000055000000000000004f0000000000000049000000000000004b00000000",
            INIT_59 => X"00000040000000000000004c0000000000000053000000000000005700000000",
            INIT_5A => X"0000003b000000000000002a0000000000000027000000000000003300000000",
            INIT_5B => X"0000003100000000000000290000000000000022000000000000003200000000",
            INIT_5C => X"000000270000000000000024000000000000001e000000000000002600000000",
            INIT_5D => X"0000002d000000000000003c0000000000000045000000000000003700000000",
            INIT_5E => X"0000001d00000000000000220000000000000026000000000000002600000000",
            INIT_5F => X"0000003300000000000000300000000000000024000000000000002000000000",
            INIT_60 => X"0000004d000000000000004f000000000000004e000000000000004c00000000",
            INIT_61 => X"00000021000000000000002c0000000000000039000000000000004400000000",
            INIT_62 => X"0000003d000000000000002e000000000000001e000000000000001d00000000",
            INIT_63 => X"0000002600000000000000320000000000000029000000000000003700000000",
            INIT_64 => X"0000001e000000000000001d000000000000001a000000000000001d00000000",
            INIT_65 => X"00000030000000000000002e0000000000000025000000000000001d00000000",
            INIT_66 => X"0000001800000000000000190000000000000025000000000000002e00000000",
            INIT_67 => X"0000002f00000000000000240000000000000020000000000000001e00000000",
            INIT_68 => X"000000320000000000000040000000000000004a000000000000005000000000",
            INIT_69 => X"0000001b000000000000001e0000000000000020000000000000002600000000",
            INIT_6A => X"0000003c000000000000002d000000000000001b000000000000001b00000000",
            INIT_6B => X"0000001d000000000000002c000000000000002f000000000000003500000000",
            INIT_6C => X"0000001c00000000000000170000000000000017000000000000001c00000000",
            INIT_6D => X"0000002500000000000000200000000000000018000000000000001900000000",
            INIT_6E => X"000000150000000000000015000000000000001d000000000000002300000000",
            INIT_6F => X"00000022000000000000001c000000000000001e000000000000001a00000000",
            INIT_70 => X"0000001a0000000000000021000000000000002d000000000000003a00000000",
            INIT_71 => X"0000001c0000000000000021000000000000001d000000000000001a00000000",
            INIT_72 => X"0000003300000000000000270000000000000018000000000000001b00000000",
            INIT_73 => X"0000001c00000000000000210000000000000032000000000000003100000000",
            INIT_74 => X"0000001d00000000000000190000000000000015000000000000001b00000000",
            INIT_75 => X"0000001700000000000000190000000000000015000000000000001800000000",
            INIT_76 => X"000000120000000000000016000000000000001a000000000000001700000000",
            INIT_77 => X"000000170000000000000019000000000000001a000000000000001500000000",
            INIT_78 => X"0000001500000000000000180000000000000017000000000000001b00000000",
            INIT_79 => X"0000001900000000000000180000000000000019000000000000001a00000000",
            INIT_7A => X"0000003000000000000000210000000000000016000000000000001a00000000",
            INIT_7B => X"0000001800000000000000230000000000000033000000000000002a00000000",
            INIT_7C => X"0000001800000000000000150000000000000014000000000000001500000000",
            INIT_7D => X"00000019000000000000001d0000000000000017000000000000001700000000",
            INIT_7E => X"000000120000000000000016000000000000001b000000000000001800000000",
            INIT_7F => X"0000001600000000000000180000000000000016000000000000001100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE47;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE48 : if BRAM_NAME = "sampleifmap_layersamples_instance48" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004100000000000000150000000000000013000000000000001700000000",
            INIT_01 => X"000000b200000000000000b700000000000000bc00000000000000a400000000",
            INIT_02 => X"000000ba00000000000000ba00000000000000ac00000000000000aa00000000",
            INIT_03 => X"000000b700000000000000b600000000000000b700000000000000b800000000",
            INIT_04 => X"0000005c000000000000007f00000000000000a400000000000000b400000000",
            INIT_05 => X"000000c20000000000000099000000000000006e000000000000006b00000000",
            INIT_06 => X"000000c600000000000000c500000000000000c900000000000000c300000000",
            INIT_07 => X"000000c500000000000000c700000000000000c800000000000000c900000000",
            INIT_08 => X"0000002e00000000000000150000000000000013000000000000001700000000",
            INIT_09 => X"000000b200000000000000bf00000000000000ca000000000000009900000000",
            INIT_0A => X"000000b700000000000000a9000000000000009e00000000000000a400000000",
            INIT_0B => X"000000b200000000000000b400000000000000b800000000000000ba00000000",
            INIT_0C => X"00000056000000000000008a00000000000000ad00000000000000b400000000",
            INIT_0D => X"000000ce00000000000000b4000000000000006a000000000000004a00000000",
            INIT_0E => X"000000ce00000000000000d000000000000000d500000000000000cf00000000",
            INIT_0F => X"000000ca00000000000000cc00000000000000cd00000000000000cf00000000",
            INIT_10 => X"0000001f00000000000000170000000000000014000000000000001700000000",
            INIT_11 => X"000000a800000000000000b900000000000000c8000000000000007f00000000",
            INIT_12 => X"000000a2000000000000009a000000000000009e000000000000009f00000000",
            INIT_13 => X"000000b200000000000000b300000000000000b200000000000000b200000000",
            INIT_14 => X"0000007d00000000000000b600000000000000be00000000000000b500000000",
            INIT_15 => X"000000d100000000000000c50000000000000072000000000000004700000000",
            INIT_16 => X"000000d300000000000000d500000000000000d800000000000000d500000000",
            INIT_17 => X"000000ce00000000000000d000000000000000d300000000000000d400000000",
            INIT_18 => X"0000001700000000000000180000000000000015000000000000001700000000",
            INIT_19 => X"000000a000000000000000af00000000000000bd000000000000006300000000",
            INIT_1A => X"0000009500000000000000a600000000000000a800000000000000a800000000",
            INIT_1B => X"000000c300000000000000bf00000000000000ba00000000000000aa00000000",
            INIT_1C => X"0000008d00000000000000bc00000000000000c800000000000000c300000000",
            INIT_1D => X"000000d600000000000000d20000000000000092000000000000006300000000",
            INIT_1E => X"000000d500000000000000d400000000000000d400000000000000d500000000",
            INIT_1F => X"000000d600000000000000d700000000000000d900000000000000d900000000",
            INIT_20 => X"0000001500000000000000170000000000000017000000000000001900000000",
            INIT_21 => X"0000009700000000000000a500000000000000aa000000000000004800000000",
            INIT_22 => X"0000009b00000000000000b900000000000000b700000000000000af00000000",
            INIT_23 => X"000000bc00000000000000a9000000000000009d000000000000009200000000",
            INIT_24 => X"0000008d00000000000000b200000000000000c400000000000000c500000000",
            INIT_25 => X"000000db00000000000000d300000000000000ac000000000000007900000000",
            INIT_26 => X"000000d900000000000000d900000000000000d900000000000000dd00000000",
            INIT_27 => X"000000ce00000000000000d100000000000000d400000000000000d600000000",
            INIT_28 => X"00000017000000000000001a000000000000001b000000000000001a00000000",
            INIT_29 => X"0000009a00000000000000a4000000000000008f000000000000003100000000",
            INIT_2A => X"000000a600000000000000c800000000000000c200000000000000a900000000",
            INIT_2B => X"000000970000000000000080000000000000007d000000000000008200000000",
            INIT_2C => X"0000008f000000000000009400000000000000a500000000000000a500000000",
            INIT_2D => X"000000c900000000000000bc00000000000000b6000000000000009300000000",
            INIT_2E => X"000000db00000000000000d500000000000000d900000000000000d400000000",
            INIT_2F => X"000000d300000000000000d700000000000000d700000000000000dc00000000",
            INIT_30 => X"00000019000000000000001b000000000000001a000000000000001e00000000",
            INIT_31 => X"000000ab00000000000000b4000000000000007d000000000000002500000000",
            INIT_32 => X"000000b300000000000000ca00000000000000c500000000000000a900000000",
            INIT_33 => X"00000082000000000000007a0000000000000071000000000000008b00000000",
            INIT_34 => X"0000008c000000000000007a0000000000000085000000000000007700000000",
            INIT_35 => X"000000c900000000000000bf00000000000000cb00000000000000b900000000",
            INIT_36 => X"000000db00000000000000d700000000000000da00000000000000d700000000",
            INIT_37 => X"000000e000000000000000dc00000000000000da00000000000000dc00000000",
            INIT_38 => X"00000024000000000000001f0000000000000030000000000000005e00000000",
            INIT_39 => X"000000a800000000000000c100000000000000af000000000000006400000000",
            INIT_3A => X"000000c300000000000000c600000000000000c000000000000000a300000000",
            INIT_3B => X"00000084000000000000008e000000000000009100000000000000ae00000000",
            INIT_3C => X"0000008b000000000000007a0000000000000079000000000000006a00000000",
            INIT_3D => X"000000d500000000000000bd00000000000000d100000000000000c000000000",
            INIT_3E => X"000000e800000000000000ef00000000000000ed00000000000000f200000000",
            INIT_3F => X"000000e500000000000000de00000000000000d500000000000000d000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007a0000000000000072000000000000009e00000000000000b400000000",
            INIT_41 => X"000000a000000000000000be00000000000000be00000000000000b100000000",
            INIT_42 => X"000000c800000000000000c500000000000000ad000000000000008500000000",
            INIT_43 => X"0000009200000000000000a700000000000000b900000000000000c200000000",
            INIT_44 => X"0000008d00000000000000850000000000000081000000000000008100000000",
            INIT_45 => X"000000dc00000000000000bd00000000000000c900000000000000b100000000",
            INIT_46 => X"000000d500000000000000e800000000000000eb00000000000000f100000000",
            INIT_47 => X"000000ea00000000000000e100000000000000c700000000000000bd00000000",
            INIT_48 => X"000000ba00000000000000b200000000000000c000000000000000c500000000",
            INIT_49 => X"0000009d00000000000000c500000000000000c300000000000000c100000000",
            INIT_4A => X"000000bf00000000000000b900000000000000a3000000000000008000000000",
            INIT_4B => X"0000009700000000000000b200000000000000c300000000000000c100000000",
            INIT_4C => X"0000008600000000000000830000000000000081000000000000007200000000",
            INIT_4D => X"000000ea00000000000000d000000000000000c200000000000000aa00000000",
            INIT_4E => X"000000c900000000000000eb00000000000000f000000000000000ec00000000",
            INIT_4F => X"000000eb00000000000000d000000000000000bb00000000000000b900000000",
            INIT_50 => X"000000c000000000000000bb00000000000000c400000000000000ca00000000",
            INIT_51 => X"0000009700000000000000c500000000000000cd00000000000000c800000000",
            INIT_52 => X"000000bd00000000000000b800000000000000af000000000000009500000000",
            INIT_53 => X"0000008800000000000000a800000000000000bb00000000000000c100000000",
            INIT_54 => X"0000008100000000000000800000000000000080000000000000007500000000",
            INIT_55 => X"000000f000000000000000cd00000000000000b500000000000000a700000000",
            INIT_56 => X"000000ce00000000000000ee00000000000000f300000000000000f300000000",
            INIT_57 => X"000000dd00000000000000c100000000000000bb00000000000000ba00000000",
            INIT_58 => X"000000c000000000000000c500000000000000cd00000000000000cd00000000",
            INIT_59 => X"000000a000000000000000c200000000000000d000000000000000cb00000000",
            INIT_5A => X"000000bf00000000000000c100000000000000bf00000000000000a800000000",
            INIT_5B => X"00000077000000000000009200000000000000ac00000000000000c100000000",
            INIT_5C => X"000000870000000000000085000000000000008e000000000000007c00000000",
            INIT_5D => X"000000ea00000000000000bf00000000000000b000000000000000a700000000",
            INIT_5E => X"000000d700000000000000ec00000000000000f100000000000000f300000000",
            INIT_5F => X"000000c400000000000000b900000000000000b800000000000000ba00000000",
            INIT_60 => X"000000c100000000000000c800000000000000cc00000000000000ce00000000",
            INIT_61 => X"000000b400000000000000bf00000000000000c700000000000000c500000000",
            INIT_62 => X"000000ad00000000000000b700000000000000b300000000000000ac00000000",
            INIT_63 => X"00000083000000000000009800000000000000ae00000000000000ae00000000",
            INIT_64 => X"0000009a000000000000008e00000000000000a6000000000000008d00000000",
            INIT_65 => X"000000e600000000000000bf00000000000000ac00000000000000a900000000",
            INIT_66 => X"000000e400000000000000ef00000000000000f100000000000000f000000000",
            INIT_67 => X"000000c000000000000000b800000000000000ba00000000000000c800000000",
            INIT_68 => X"000000bf00000000000000c600000000000000ca00000000000000d200000000",
            INIT_69 => X"000000ca00000000000000b100000000000000b400000000000000c900000000",
            INIT_6A => X"0000008e000000000000008e000000000000009a00000000000000ab00000000",
            INIT_6B => X"0000009c000000000000009300000000000000a800000000000000a800000000",
            INIT_6C => X"000000a4000000000000009600000000000000a900000000000000af00000000",
            INIT_6D => X"000000e600000000000000c500000000000000a0000000000000009e00000000",
            INIT_6E => X"000000f200000000000000f400000000000000f100000000000000f100000000",
            INIT_6F => X"000000d700000000000000c300000000000000bf00000000000000e200000000",
            INIT_70 => X"000000c000000000000000c700000000000000c900000000000000d300000000",
            INIT_71 => X"000000d700000000000000a100000000000000aa00000000000000cf00000000",
            INIT_72 => X"000000ac00000000000000ad00000000000000ba00000000000000bd00000000",
            INIT_73 => X"0000007f000000000000008900000000000000b100000000000000be00000000",
            INIT_74 => X"000000a0000000000000009600000000000000ae00000000000000b400000000",
            INIT_75 => X"000000ec00000000000000c100000000000000b000000000000000af00000000",
            INIT_76 => X"000000fb00000000000000f300000000000000f200000000000000f500000000",
            INIT_77 => X"000000e100000000000000d400000000000000c900000000000000ef00000000",
            INIT_78 => X"000000c100000000000000c500000000000000c400000000000000d300000000",
            INIT_79 => X"000000d9000000000000009a00000000000000b500000000000000d100000000",
            INIT_7A => X"000000b900000000000000c300000000000000c500000000000000ce00000000",
            INIT_7B => X"0000009800000000000000a600000000000000ad00000000000000aa00000000",
            INIT_7C => X"0000009800000000000000a600000000000000b800000000000000a300000000",
            INIT_7D => X"000000cc00000000000000af00000000000000b500000000000000c000000000",
            INIT_7E => X"000000f700000000000000f400000000000000f300000000000000ee00000000",
            INIT_7F => X"000000e200000000000000e200000000000000d500000000000000df00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE48;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE49 : if BRAM_NAME = "sampleifmap_layersamples_instance49" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b500000000000000b400000000000000c200000000000000d600000000",
            INIT_01 => X"000000c6000000000000009b00000000000000c400000000000000c500000000",
            INIT_02 => X"000000b700000000000000ae00000000000000c000000000000000d600000000",
            INIT_03 => X"000000b200000000000000ae00000000000000a100000000000000ad00000000",
            INIT_04 => X"0000009300000000000000bd00000000000000a4000000000000008000000000",
            INIT_05 => X"00000076000000000000009c00000000000000b400000000000000a700000000",
            INIT_06 => X"000000eb00000000000000ef00000000000000d7000000000000009d00000000",
            INIT_07 => X"000000e400000000000000ea00000000000000d600000000000000ce00000000",
            INIT_08 => X"000000a300000000000000a600000000000000c600000000000000d700000000",
            INIT_09 => X"000000b900000000000000be00000000000000ca00000000000000b400000000",
            INIT_0A => X"000000d600000000000000cd00000000000000d200000000000000cf00000000",
            INIT_0B => X"000000ad00000000000000b000000000000000ae00000000000000c100000000",
            INIT_0C => X"0000009900000000000000bf0000000000000089000000000000008100000000",
            INIT_0D => X"0000008700000000000000ab00000000000000c800000000000000a300000000",
            INIT_0E => X"000000c100000000000000b80000000000000090000000000000007400000000",
            INIT_0F => X"000000eb00000000000000ef00000000000000d200000000000000bb00000000",
            INIT_10 => X"000000a400000000000000ae00000000000000cd00000000000000d800000000",
            INIT_11 => X"000000c200000000000000d200000000000000cb00000000000000b900000000",
            INIT_12 => X"000000e200000000000000da00000000000000d300000000000000bf00000000",
            INIT_13 => X"000000b300000000000000be00000000000000cb00000000000000e100000000",
            INIT_14 => X"0000009e00000000000000a80000000000000079000000000000009700000000",
            INIT_15 => X"000000ac00000000000000aa00000000000000c200000000000000a700000000",
            INIT_16 => X"000000a900000000000000990000000000000083000000000000009a00000000",
            INIT_17 => X"000000ec00000000000000de00000000000000b800000000000000a200000000",
            INIT_18 => X"000000b400000000000000c000000000000000d000000000000000d800000000",
            INIT_19 => X"000000d200000000000000d100000000000000ca00000000000000c500000000",
            INIT_1A => X"000000cc00000000000000c500000000000000bd00000000000000ba00000000",
            INIT_1B => X"000000b500000000000000cf00000000000000d500000000000000d100000000",
            INIT_1C => X"000000af0000000000000092000000000000009500000000000000b200000000",
            INIT_1D => X"000000ab000000000000009c00000000000000ae00000000000000b700000000",
            INIT_1E => X"000000b400000000000000a9000000000000009400000000000000a300000000",
            INIT_1F => X"000000cc00000000000000ac00000000000000a000000000000000a600000000",
            INIT_20 => X"000000b600000000000000ca00000000000000d500000000000000da00000000",
            INIT_21 => X"000000ca00000000000000c900000000000000cb00000000000000bf00000000",
            INIT_22 => X"000000c000000000000000c100000000000000c300000000000000ca00000000",
            INIT_23 => X"000000c700000000000000cf00000000000000c600000000000000b200000000",
            INIT_24 => X"000000bb00000000000000a600000000000000cb00000000000000d300000000",
            INIT_25 => X"000000a60000000000000093000000000000009b00000000000000b100000000",
            INIT_26 => X"000000af00000000000000b600000000000000ab00000000000000a700000000",
            INIT_27 => X"000000a7000000000000009f000000000000009c000000000000009c00000000",
            INIT_28 => X"000000ba00000000000000d100000000000000d700000000000000d900000000",
            INIT_29 => X"000000c800000000000000d000000000000000c800000000000000b300000000",
            INIT_2A => X"000000ba00000000000000d200000000000000d700000000000000d100000000",
            INIT_2B => X"000000c200000000000000c400000000000000b600000000000000a100000000",
            INIT_2C => X"000000b900000000000000be00000000000000cf00000000000000cb00000000",
            INIT_2D => X"000000a6000000000000009b000000000000008e000000000000009b00000000",
            INIT_2E => X"0000009f00000000000000ad00000000000000b300000000000000ac00000000",
            INIT_2F => X"0000008f000000000000009e000000000000009e000000000000009600000000",
            INIT_30 => X"000000c000000000000000d600000000000000d500000000000000d600000000",
            INIT_31 => X"000000d900000000000000da00000000000000c500000000000000a900000000",
            INIT_32 => X"000000c300000000000000d400000000000000d900000000000000d700000000",
            INIT_33 => X"000000bf00000000000000c300000000000000b300000000000000aa00000000",
            INIT_34 => X"000000aa00000000000000c000000000000000c000000000000000be00000000",
            INIT_35 => X"000000aa00000000000000a7000000000000008e000000000000008400000000",
            INIT_36 => X"0000009d00000000000000ad00000000000000b300000000000000aa00000000",
            INIT_37 => X"0000007d00000000000000860000000000000093000000000000009d00000000",
            INIT_38 => X"000000ca00000000000000d300000000000000d100000000000000d500000000",
            INIT_39 => X"000000de00000000000000d800000000000000c100000000000000a800000000",
            INIT_3A => X"000000cd00000000000000d300000000000000de00000000000000df00000000",
            INIT_3B => X"000000c600000000000000c900000000000000c200000000000000c200000000",
            INIT_3C => X"0000009900000000000000bc00000000000000c400000000000000c600000000",
            INIT_3D => X"000000a700000000000000ab000000000000009b000000000000008600000000",
            INIT_3E => X"000000a500000000000000b200000000000000bd00000000000000a600000000",
            INIT_3F => X"000000890000000000000085000000000000008e00000000000000a300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ca00000000000000ce00000000000000ce00000000000000d300000000",
            INIT_41 => X"000000d500000000000000d300000000000000bf00000000000000af00000000",
            INIT_42 => X"000000ab00000000000000c600000000000000d800000000000000d600000000",
            INIT_43 => X"000000c900000000000000c900000000000000ce00000000000000c200000000",
            INIT_44 => X"0000009600000000000000b100000000000000c500000000000000c800000000",
            INIT_45 => X"0000009d00000000000000a7000000000000009e000000000000009000000000",
            INIT_46 => X"000000a800000000000000b000000000000000b5000000000000009f00000000",
            INIT_47 => X"0000009000000000000000950000000000000096000000000000009800000000",
            INIT_48 => X"000000c100000000000000c900000000000000cc00000000000000d200000000",
            INIT_49 => X"000000d200000000000000d000000000000000bc00000000000000b500000000",
            INIT_4A => X"0000007a00000000000000a000000000000000ce00000000000000cd00000000",
            INIT_4B => X"000000c200000000000000c600000000000000d000000000000000b100000000",
            INIT_4C => X"0000009600000000000000a600000000000000b800000000000000c100000000",
            INIT_4D => X"0000009900000000000000a0000000000000009c000000000000008b00000000",
            INIT_4E => X"0000009b000000000000009f00000000000000a0000000000000009b00000000",
            INIT_4F => X"00000083000000000000008c0000000000000098000000000000009800000000",
            INIT_50 => X"000000bb00000000000000c600000000000000ca00000000000000d200000000",
            INIT_51 => X"000000d600000000000000cd00000000000000b200000000000000ae00000000",
            INIT_52 => X"0000008300000000000000a400000000000000cb00000000000000d100000000",
            INIT_53 => X"000000b600000000000000bb00000000000000ca00000000000000b400000000",
            INIT_54 => X"0000008b000000000000009d00000000000000a900000000000000b600000000",
            INIT_55 => X"00000090000000000000009a0000000000000099000000000000008600000000",
            INIT_56 => X"0000008d0000000000000083000000000000008d000000000000009700000000",
            INIT_57 => X"000000930000000000000096000000000000009b000000000000009d00000000",
            INIT_58 => X"000000b500000000000000c200000000000000c800000000000000d200000000",
            INIT_59 => X"000000d700000000000000c400000000000000a800000000000000a800000000",
            INIT_5A => X"000000b800000000000000bd00000000000000c700000000000000d400000000",
            INIT_5B => X"000000ac00000000000000ad00000000000000b900000000000000cb00000000",
            INIT_5C => X"000000760000000000000093000000000000009b00000000000000a300000000",
            INIT_5D => X"0000008d00000000000000910000000000000094000000000000008300000000",
            INIT_5E => X"00000085000000000000007f0000000000000084000000000000009000000000",
            INIT_5F => X"0000009c00000000000000a200000000000000a3000000000000009500000000",
            INIT_60 => X"000000b400000000000000bd00000000000000c200000000000000d000000000",
            INIT_61 => X"000000d300000000000000bd000000000000009e00000000000000a200000000",
            INIT_62 => X"000000c700000000000000c200000000000000c500000000000000d300000000",
            INIT_63 => X"000000a400000000000000a300000000000000ac00000000000000bf00000000",
            INIT_64 => X"0000006d00000000000000820000000000000093000000000000009e00000000",
            INIT_65 => X"0000009100000000000000900000000000000090000000000000008900000000",
            INIT_66 => X"00000086000000000000007c0000000000000084000000000000009000000000",
            INIT_67 => X"00000093000000000000009f00000000000000a2000000000000009700000000",
            INIT_68 => X"000000b500000000000000b000000000000000b100000000000000c200000000",
            INIT_69 => X"000000cd00000000000000b3000000000000008f000000000000009f00000000",
            INIT_6A => X"000000be00000000000000c200000000000000c700000000000000d000000000",
            INIT_6B => X"000000a1000000000000009c00000000000000a500000000000000b500000000",
            INIT_6C => X"0000007200000000000000700000000000000088000000000000009500000000",
            INIT_6D => X"00000092000000000000008a0000000000000085000000000000008900000000",
            INIT_6E => X"0000009000000000000000830000000000000083000000000000009200000000",
            INIT_6F => X"0000008d00000000000000940000000000000095000000000000009600000000",
            INIT_70 => X"000000b200000000000000a5000000000000009d00000000000000ac00000000",
            INIT_71 => X"000000c7000000000000009c000000000000008500000000000000a700000000",
            INIT_72 => X"000000c200000000000000c700000000000000c700000000000000ce00000000",
            INIT_73 => X"0000008b0000000000000084000000000000008500000000000000a000000000",
            INIT_74 => X"0000007e000000000000006b000000000000007e000000000000008c00000000",
            INIT_75 => X"00000095000000000000008a0000000000000081000000000000008200000000",
            INIT_76 => X"0000008e0000000000000091000000000000008c000000000000008d00000000",
            INIT_77 => X"000000980000000000000095000000000000008c000000000000008800000000",
            INIT_78 => X"0000009b00000000000000900000000000000086000000000000009700000000",
            INIT_79 => X"000000b70000000000000082000000000000007d000000000000009e00000000",
            INIT_7A => X"000000a500000000000000b700000000000000bf00000000000000c500000000",
            INIT_7B => X"00000069000000000000005e0000000000000067000000000000008000000000",
            INIT_7C => X"0000007c00000000000000750000000000000070000000000000007700000000",
            INIT_7D => X"0000008f000000000000008b000000000000007d000000000000007900000000",
            INIT_7E => X"0000007d0000000000000081000000000000008c000000000000008b00000000",
            INIT_7F => X"00000096000000000000009b0000000000000095000000000000008400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE49;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE50 : if BRAM_NAME = "sampleifmap_layersamples_instance50" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002f00000000000000100000000000000015000000000000001300000000",
            INIT_01 => X"0000008e00000000000000930000000000000093000000000000008300000000",
            INIT_02 => X"0000008e00000000000000900000000000000089000000000000008700000000",
            INIT_03 => X"0000008f000000000000008c000000000000008c000000000000008d00000000",
            INIT_04 => X"000000490000000000000060000000000000007e000000000000008c00000000",
            INIT_05 => X"000000a40000000000000082000000000000005d000000000000005f00000000",
            INIT_06 => X"0000009d000000000000009b000000000000009c000000000000009b00000000",
            INIT_07 => X"000000970000000000000098000000000000009b000000000000009e00000000",
            INIT_08 => X"0000001f00000000000000110000000000000014000000000000001400000000",
            INIT_09 => X"00000092000000000000009b00000000000000a1000000000000007a00000000",
            INIT_0A => X"00000095000000000000008b0000000000000088000000000000008a00000000",
            INIT_0B => X"0000009700000000000000920000000000000096000000000000009800000000",
            INIT_0C => X"0000004900000000000000750000000000000096000000000000009f00000000",
            INIT_0D => X"000000af000000000000009c0000000000000058000000000000004100000000",
            INIT_0E => X"000000ad00000000000000ab00000000000000a900000000000000a800000000",
            INIT_0F => X"000000a300000000000000a400000000000000a800000000000000ac00000000",
            INIT_10 => X"0000001500000000000000140000000000000014000000000000001400000000",
            INIT_11 => X"0000008c000000000000009700000000000000a2000000000000006600000000",
            INIT_12 => X"0000008b00000000000000880000000000000095000000000000008d00000000",
            INIT_13 => X"0000009f00000000000000980000000000000099000000000000009a00000000",
            INIT_14 => X"0000006d00000000000000a100000000000000ab00000000000000a600000000",
            INIT_15 => X"000000b700000000000000b10000000000000061000000000000003a00000000",
            INIT_16 => X"000000b200000000000000b100000000000000b200000000000000b300000000",
            INIT_17 => X"000000a600000000000000a900000000000000ad00000000000000b100000000",
            INIT_18 => X"0000001100000000000000150000000000000014000000000000001400000000",
            INIT_19 => X"00000082000000000000008c0000000000000099000000000000004f00000000",
            INIT_1A => X"00000087000000000000009d00000000000000a4000000000000009700000000",
            INIT_1B => X"000000b000000000000000a900000000000000a6000000000000009900000000",
            INIT_1C => X"0000007600000000000000a100000000000000af00000000000000b000000000",
            INIT_1D => X"000000c300000000000000c40000000000000085000000000000005200000000",
            INIT_1E => X"000000b300000000000000b400000000000000b700000000000000bd00000000",
            INIT_1F => X"000000ab00000000000000ad00000000000000b100000000000000b300000000",
            INIT_20 => X"0000001300000000000000150000000000000014000000000000001500000000",
            INIT_21 => X"0000007700000000000000820000000000000089000000000000003800000000",
            INIT_22 => X"0000009200000000000000b300000000000000b2000000000000009c00000000",
            INIT_23 => X"000000a70000000000000094000000000000008b000000000000008400000000",
            INIT_24 => X"00000078000000000000009800000000000000a900000000000000af00000000",
            INIT_25 => X"000000d200000000000000ce00000000000000a7000000000000006d00000000",
            INIT_26 => X"000000bf00000000000000c300000000000000c900000000000000d100000000",
            INIT_27 => X"000000ac00000000000000b100000000000000b600000000000000ba00000000",
            INIT_28 => X"0000001600000000000000170000000000000016000000000000001600000000",
            INIT_29 => X"0000007800000000000000820000000000000073000000000000002600000000",
            INIT_2A => X"0000009e00000000000000c300000000000000b9000000000000009200000000",
            INIT_2B => X"00000084000000000000006b000000000000006c000000000000007600000000",
            INIT_2C => X"000000840000000000000081000000000000008f000000000000009200000000",
            INIT_2D => X"000000c700000000000000be00000000000000b7000000000000008f00000000",
            INIT_2E => X"000000d100000000000000cc00000000000000d100000000000000cf00000000",
            INIT_2F => X"000000c200000000000000c700000000000000ca00000000000000d100000000",
            INIT_30 => X"0000001400000000000000150000000000000013000000000000001800000000",
            INIT_31 => X"0000009400000000000000a10000000000000071000000000000001e00000000",
            INIT_32 => X"000000aa00000000000000c200000000000000ba000000000000009700000000",
            INIT_33 => X"0000007100000000000000690000000000000062000000000000008000000000",
            INIT_34 => X"00000080000000000000006b0000000000000074000000000000006800000000",
            INIT_35 => X"000000c500000000000000c000000000000000ca00000000000000b200000000",
            INIT_36 => X"000000d700000000000000d100000000000000cf00000000000000ce00000000",
            INIT_37 => X"000000da00000000000000d700000000000000d600000000000000d800000000",
            INIT_38 => X"0000001d00000000000000180000000000000029000000000000005800000000",
            INIT_39 => X"0000009c00000000000000ba00000000000000ae000000000000006000000000",
            INIT_3A => X"000000ba00000000000000bd00000000000000b5000000000000009500000000",
            INIT_3B => X"000000760000000000000081000000000000008400000000000000a400000000",
            INIT_3C => X"0000007c000000000000006c000000000000006b000000000000005c00000000",
            INIT_3D => X"000000ce00000000000000bb00000000000000cc00000000000000b400000000",
            INIT_3E => X"000000e400000000000000e700000000000000e000000000000000e600000000",
            INIT_3F => X"000000e200000000000000dc00000000000000d300000000000000cd00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000075000000000000006d000000000000009900000000000000b100000000",
            INIT_41 => X"0000009300000000000000b700000000000000bd00000000000000af00000000",
            INIT_42 => X"000000c000000000000000bc00000000000000a1000000000000007800000000",
            INIT_43 => X"00000083000000000000009a00000000000000ad00000000000000b800000000",
            INIT_44 => X"0000007f00000000000000770000000000000073000000000000007300000000",
            INIT_45 => X"000000d800000000000000bc00000000000000c500000000000000a600000000",
            INIT_46 => X"000000d300000000000000e300000000000000e200000000000000e900000000",
            INIT_47 => X"000000e800000000000000e000000000000000c600000000000000bc00000000",
            INIT_48 => X"000000b600000000000000af00000000000000bc00000000000000c200000000",
            INIT_49 => X"0000009000000000000000be00000000000000c200000000000000bf00000000",
            INIT_4A => X"000000b600000000000000b10000000000000098000000000000007300000000",
            INIT_4B => X"0000008a00000000000000a400000000000000b600000000000000b700000000",
            INIT_4C => X"0000007b00000000000000770000000000000076000000000000006600000000",
            INIT_4D => X"000000e900000000000000d000000000000000bd00000000000000a000000000",
            INIT_4E => X"000000cb00000000000000ea00000000000000eb00000000000000e800000000",
            INIT_4F => X"000000eb00000000000000d100000000000000bd00000000000000bb00000000",
            INIT_50 => X"000000bb00000000000000b700000000000000c000000000000000c700000000",
            INIT_51 => X"0000008a00000000000000bf00000000000000cd00000000000000c600000000",
            INIT_52 => X"000000b500000000000000b000000000000000a5000000000000008800000000",
            INIT_53 => X"0000007c000000000000009a00000000000000af00000000000000b800000000",
            INIT_54 => X"0000007800000000000000770000000000000076000000000000006b00000000",
            INIT_55 => X"000000f000000000000000cd00000000000000b0000000000000009e00000000",
            INIT_56 => X"000000d400000000000000f200000000000000f400000000000000f300000000",
            INIT_57 => X"000000e000000000000000c600000000000000c000000000000000c000000000",
            INIT_58 => X"000000bb00000000000000c100000000000000c900000000000000c900000000",
            INIT_59 => X"0000009200000000000000bc00000000000000d100000000000000c900000000",
            INIT_5A => X"000000b700000000000000b900000000000000b6000000000000009b00000000",
            INIT_5B => X"0000006b0000000000000084000000000000009f00000000000000b700000000",
            INIT_5C => X"0000007e000000000000007c0000000000000085000000000000007300000000",
            INIT_5D => X"000000eb00000000000000bd00000000000000aa000000000000009e00000000",
            INIT_5E => X"000000de00000000000000f200000000000000f600000000000000f600000000",
            INIT_5F => X"000000ca00000000000000c000000000000000c000000000000000c200000000",
            INIT_60 => X"000000bd00000000000000c500000000000000c900000000000000cb00000000",
            INIT_61 => X"000000a500000000000000b700000000000000c600000000000000c400000000",
            INIT_62 => X"000000a500000000000000b000000000000000aa000000000000009f00000000",
            INIT_63 => X"00000078000000000000008a00000000000000a200000000000000a400000000",
            INIT_64 => X"000000920000000000000087000000000000009f000000000000008500000000",
            INIT_65 => X"000000e700000000000000bd00000000000000a500000000000000a100000000",
            INIT_66 => X"000000ea00000000000000f700000000000000f800000000000000f400000000",
            INIT_67 => X"000000c700000000000000c100000000000000c300000000000000d000000000",
            INIT_68 => X"000000b900000000000000c400000000000000ca00000000000000d000000000",
            INIT_69 => X"000000b9000000000000009c00000000000000a700000000000000c100000000",
            INIT_6A => X"000000870000000000000087000000000000009100000000000000a100000000",
            INIT_6B => X"0000008f0000000000000089000000000000009e00000000000000a100000000",
            INIT_6C => X"000000a2000000000000009500000000000000a400000000000000a400000000",
            INIT_6D => X"000000e400000000000000c3000000000000009d000000000000009900000000",
            INIT_6E => X"000000f500000000000000f900000000000000f700000000000000f200000000",
            INIT_6F => X"000000de00000000000000cc00000000000000c700000000000000e800000000",
            INIT_70 => X"000000b600000000000000c500000000000000cc00000000000000d200000000",
            INIT_71 => X"000000c1000000000000007d000000000000008e00000000000000bf00000000",
            INIT_72 => X"000000a700000000000000a600000000000000b100000000000000b500000000",
            INIT_73 => X"00000072000000000000008200000000000000aa00000000000000b800000000",
            INIT_74 => X"0000009e000000000000009800000000000000aa00000000000000a500000000",
            INIT_75 => X"000000e700000000000000bd00000000000000ae00000000000000ab00000000",
            INIT_76 => X"000000fb00000000000000f500000000000000f400000000000000f200000000",
            INIT_77 => X"000000e900000000000000dd00000000000000cf00000000000000f200000000",
            INIT_78 => X"000000b900000000000000c500000000000000c800000000000000d400000000",
            INIT_79 => X"000000c00000000000000070000000000000009100000000000000bd00000000",
            INIT_7A => X"000000b400000000000000bd00000000000000be00000000000000c700000000",
            INIT_7B => X"0000008900000000000000a000000000000000a700000000000000a400000000",
            INIT_7C => X"0000009100000000000000a200000000000000b0000000000000009200000000",
            INIT_7D => X"000000c300000000000000a800000000000000b100000000000000b800000000",
            INIT_7E => X"000000f900000000000000f500000000000000f100000000000000e800000000",
            INIT_7F => X"000000eb00000000000000ec00000000000000dd00000000000000e400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE50;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE51 : if BRAM_NAME = "sampleifmap_layersamples_instance51" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ae00000000000000b600000000000000c700000000000000d800000000",
            INIT_01 => X"000000ad000000000000006e000000000000009b00000000000000b000000000",
            INIT_02 => X"000000b200000000000000a800000000000000ba00000000000000d000000000",
            INIT_03 => X"000000a400000000000000a7000000000000009b00000000000000a800000000",
            INIT_04 => X"0000008600000000000000b10000000000000096000000000000006e00000000",
            INIT_05 => X"00000068000000000000009000000000000000ab000000000000009a00000000",
            INIT_06 => X"000000ed00000000000000ee00000000000000d1000000000000009100000000",
            INIT_07 => X"000000ed00000000000000f300000000000000dd00000000000000d200000000",
            INIT_08 => X"0000009e00000000000000a900000000000000ce00000000000000db00000000",
            INIT_09 => X"000000a2000000000000009500000000000000a700000000000000a300000000",
            INIT_0A => X"000000d100000000000000c800000000000000cd00000000000000ca00000000",
            INIT_0B => X"000000a100000000000000aa00000000000000a800000000000000bc00000000",
            INIT_0C => X"0000008700000000000000ad0000000000000078000000000000007000000000",
            INIT_0D => X"00000073000000000000009b00000000000000ba000000000000009300000000",
            INIT_0E => X"000000bc00000000000000b20000000000000084000000000000006200000000",
            INIT_0F => X"000000ef00000000000000f300000000000000d400000000000000b900000000",
            INIT_10 => X"000000a100000000000000b300000000000000d600000000000000dd00000000",
            INIT_11 => X"000000b100000000000000b300000000000000b500000000000000af00000000",
            INIT_12 => X"000000dd00000000000000d400000000000000cf00000000000000bd00000000",
            INIT_13 => X"000000ab00000000000000b800000000000000c500000000000000dc00000000",
            INIT_14 => X"0000008c00000000000000950000000000000067000000000000008b00000000",
            INIT_15 => X"00000093000000000000009400000000000000b1000000000000009700000000",
            INIT_16 => X"0000009c000000000000008a0000000000000070000000000000008300000000",
            INIT_17 => X"000000ea00000000000000d900000000000000b1000000000000009700000000",
            INIT_18 => X"000000b200000000000000c600000000000000da00000000000000df00000000",
            INIT_19 => X"000000c800000000000000be00000000000000c200000000000000c200000000",
            INIT_1A => X"000000c700000000000000bf00000000000000b800000000000000ba00000000",
            INIT_1B => X"000000b100000000000000c800000000000000d000000000000000cb00000000",
            INIT_1C => X"0000009e000000000000007f000000000000008700000000000000ab00000000",
            INIT_1D => X"0000008f0000000000000083000000000000009b00000000000000a800000000",
            INIT_1E => X"0000009f0000000000000094000000000000007e000000000000008900000000",
            INIT_1F => X"000000c5000000000000009e0000000000000090000000000000009300000000",
            INIT_20 => X"000000b700000000000000d000000000000000dd00000000000000e100000000",
            INIT_21 => X"000000c200000000000000be00000000000000c700000000000000bf00000000",
            INIT_22 => X"000000ba00000000000000be00000000000000bc00000000000000c600000000",
            INIT_23 => X"000000bf00000000000000c600000000000000c100000000000000ab00000000",
            INIT_24 => X"000000a9000000000000009400000000000000bf00000000000000cf00000000",
            INIT_25 => X"0000008d000000000000007b000000000000008700000000000000a000000000",
            INIT_26 => X"00000098000000000000009f0000000000000095000000000000008e00000000",
            INIT_27 => X"0000009a000000000000008c0000000000000088000000000000008700000000",
            INIT_28 => X"000000be00000000000000d600000000000000dd00000000000000de00000000",
            INIT_29 => X"000000be00000000000000c800000000000000c300000000000000b300000000",
            INIT_2A => X"000000b200000000000000d100000000000000cd00000000000000c600000000",
            INIT_2B => X"000000b500000000000000b600000000000000b3000000000000009700000000",
            INIT_2C => X"000000a500000000000000ae00000000000000c400000000000000c500000000",
            INIT_2D => X"000000930000000000000089000000000000007c000000000000008600000000",
            INIT_2E => X"0000008b000000000000009900000000000000a1000000000000009900000000",
            INIT_2F => X"0000007d000000000000008b000000000000008b000000000000008300000000",
            INIT_30 => X"000000c600000000000000db00000000000000da00000000000000db00000000",
            INIT_31 => X"000000cf00000000000000d200000000000000bf00000000000000aa00000000",
            INIT_32 => X"000000b400000000000000cf00000000000000ce00000000000000cb00000000",
            INIT_33 => X"000000b000000000000000b400000000000000ae000000000000009c00000000",
            INIT_34 => X"0000009600000000000000b000000000000000b500000000000000b600000000",
            INIT_35 => X"000000980000000000000096000000000000007d000000000000006f00000000",
            INIT_36 => X"0000008a000000000000009a00000000000000a1000000000000009800000000",
            INIT_37 => X"0000006a00000000000000730000000000000080000000000000008a00000000",
            INIT_38 => X"000000cf00000000000000d900000000000000d600000000000000da00000000",
            INIT_39 => X"000000d500000000000000d200000000000000bc00000000000000aa00000000",
            INIT_3A => X"000000b600000000000000c700000000000000d300000000000000d400000000",
            INIT_3B => X"000000b500000000000000ba00000000000000ba00000000000000ae00000000",
            INIT_3C => X"0000008500000000000000ab00000000000000b600000000000000ba00000000",
            INIT_3D => X"00000095000000000000009a0000000000000089000000000000007200000000",
            INIT_3E => X"00000092000000000000009f00000000000000ab000000000000009400000000",
            INIT_3F => X"000000760000000000000073000000000000007b000000000000009000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d100000000000000d400000000000000d400000000000000d800000000",
            INIT_41 => X"000000cd00000000000000cf00000000000000bd00000000000000b300000000",
            INIT_42 => X"0000008a00000000000000b100000000000000cd00000000000000cd00000000",
            INIT_43 => X"000000b600000000000000bb00000000000000c300000000000000a700000000",
            INIT_44 => X"00000082000000000000009e00000000000000b500000000000000b900000000",
            INIT_45 => X"0000008c0000000000000096000000000000008d000000000000007d00000000",
            INIT_46 => X"00000095000000000000009d00000000000000a3000000000000008d00000000",
            INIT_47 => X"0000007c00000000000000820000000000000083000000000000008500000000",
            INIT_48 => X"000000c800000000000000d000000000000000d200000000000000d700000000",
            INIT_49 => X"000000cc00000000000000ce00000000000000be00000000000000bb00000000",
            INIT_4A => X"00000050000000000000008300000000000000c400000000000000c600000000",
            INIT_4B => X"000000ae00000000000000b800000000000000c2000000000000009100000000",
            INIT_4C => X"00000083000000000000009300000000000000a500000000000000ae00000000",
            INIT_4D => X"00000088000000000000008f000000000000008b000000000000007800000000",
            INIT_4E => X"00000088000000000000008c000000000000008e000000000000008900000000",
            INIT_4F => X"0000007000000000000000790000000000000085000000000000008500000000",
            INIT_50 => X"000000c200000000000000cd00000000000000d000000000000000d700000000",
            INIT_51 => X"000000d100000000000000cd00000000000000b700000000000000b500000000",
            INIT_52 => X"00000051000000000000008100000000000000c200000000000000cc00000000",
            INIT_53 => X"000000a100000000000000ab00000000000000ba000000000000008e00000000",
            INIT_54 => X"000000780000000000000089000000000000009500000000000000a100000000",
            INIT_55 => X"0000007e00000000000000890000000000000087000000000000007300000000",
            INIT_56 => X"0000007a0000000000000070000000000000007b000000000000008500000000",
            INIT_57 => X"0000008000000000000000830000000000000088000000000000008a00000000",
            INIT_58 => X"000000bc00000000000000c800000000000000cd00000000000000d600000000",
            INIT_59 => X"000000d400000000000000c600000000000000af00000000000000b000000000",
            INIT_5A => X"0000008e00000000000000a000000000000000c000000000000000d000000000",
            INIT_5B => X"00000095000000000000009b00000000000000a800000000000000aa00000000",
            INIT_5C => X"00000064000000000000007f0000000000000085000000000000008d00000000",
            INIT_5D => X"0000007b00000000000000800000000000000083000000000000007100000000",
            INIT_5E => X"00000072000000000000006c0000000000000072000000000000007e00000000",
            INIT_5F => X"0000008900000000000000900000000000000090000000000000008200000000",
            INIT_60 => X"000000b700000000000000c000000000000000c400000000000000d200000000",
            INIT_61 => X"000000d200000000000000c000000000000000a600000000000000a900000000",
            INIT_62 => X"000000b400000000000000b600000000000000c000000000000000d100000000",
            INIT_63 => X"0000008c000000000000008d000000000000009900000000000000ab00000000",
            INIT_64 => X"0000005c000000000000006f000000000000007d000000000000008600000000",
            INIT_65 => X"0000007f000000000000007e000000000000007e000000000000007800000000",
            INIT_66 => X"0000007400000000000000690000000000000072000000000000007e00000000",
            INIT_67 => X"00000081000000000000008d0000000000000090000000000000008500000000",
            INIT_68 => X"000000b900000000000000b300000000000000b300000000000000c400000000",
            INIT_69 => X"000000cc00000000000000b5000000000000009700000000000000a600000000",
            INIT_6A => X"000000b300000000000000ba00000000000000c200000000000000cd00000000",
            INIT_6B => X"000000880000000000000085000000000000009200000000000000a600000000",
            INIT_6C => X"00000061000000000000005d0000000000000072000000000000007e00000000",
            INIT_6D => X"0000008000000000000000780000000000000073000000000000007800000000",
            INIT_6E => X"0000007e00000000000000710000000000000071000000000000008000000000",
            INIT_6F => X"0000007b00000000000000820000000000000083000000000000008400000000",
            INIT_70 => X"000000b800000000000000aa00000000000000a100000000000000b100000000",
            INIT_71 => X"000000c3000000000000009c000000000000008c00000000000000ae00000000",
            INIT_72 => X"000000b600000000000000bf00000000000000c100000000000000c900000000",
            INIT_73 => X"00000073000000000000006c0000000000000071000000000000009100000000",
            INIT_74 => X"0000006e0000000000000059000000000000006a000000000000007600000000",
            INIT_75 => X"0000008300000000000000780000000000000070000000000000007200000000",
            INIT_76 => X"0000007c000000000000007f000000000000007a000000000000007b00000000",
            INIT_77 => X"000000860000000000000082000000000000007a000000000000007500000000",
            INIT_78 => X"000000a10000000000000097000000000000008c000000000000009d00000000",
            INIT_79 => X"000000b10000000000000080000000000000008200000000000000a600000000",
            INIT_7A => X"0000009a00000000000000af00000000000000b700000000000000bf00000000",
            INIT_7B => X"0000005300000000000000470000000000000053000000000000007000000000",
            INIT_7C => X"0000006e0000000000000065000000000000005e000000000000006300000000",
            INIT_7D => X"0000007e0000000000000079000000000000006c000000000000006c00000000",
            INIT_7E => X"0000006b000000000000006f000000000000007a000000000000007900000000",
            INIT_7F => X"0000008400000000000000890000000000000084000000000000007300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE51;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE52 : if BRAM_NAME = "sampleifmap_layersamples_instance52" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000280000000000000013000000000000001c000000000000001700000000",
            INIT_01 => X"00000074000000000000006d0000000000000073000000000000007100000000",
            INIT_02 => X"00000069000000000000006a0000000000000067000000000000007100000000",
            INIT_03 => X"0000006b00000000000000690000000000000069000000000000006900000000",
            INIT_04 => X"0000003a000000000000004c0000000000000063000000000000006a00000000",
            INIT_05 => X"0000008900000000000000720000000000000056000000000000005400000000",
            INIT_06 => X"0000007d000000000000007c000000000000007d000000000000007c00000000",
            INIT_07 => X"00000078000000000000007a000000000000007d000000000000007f00000000",
            INIT_08 => X"0000001a0000000000000014000000000000001b000000000000001800000000",
            INIT_09 => X"0000007c00000000000000760000000000000082000000000000006a00000000",
            INIT_0A => X"00000075000000000000006d0000000000000072000000000000007d00000000",
            INIT_0B => X"0000007900000000000000720000000000000076000000000000007800000000",
            INIT_0C => X"00000044000000000000006a0000000000000083000000000000008500000000",
            INIT_0D => X"00000096000000000000008c0000000000000051000000000000003e00000000",
            INIT_0E => X"000000880000000000000089000000000000008c000000000000008a00000000",
            INIT_0F => X"0000008000000000000000810000000000000085000000000000008800000000",
            INIT_10 => X"000000120000000000000017000000000000001a000000000000001800000000",
            INIT_11 => X"0000007b00000000000000740000000000000083000000000000005800000000",
            INIT_12 => X"000000740000000000000074000000000000008d000000000000008b00000000",
            INIT_13 => X"00000084000000000000007d000000000000007f000000000000008100000000",
            INIT_14 => X"000000690000000000000098000000000000009a000000000000008e00000000",
            INIT_15 => X"0000009e000000000000009f0000000000000059000000000000003700000000",
            INIT_16 => X"0000008e00000000000000920000000000000097000000000000009700000000",
            INIT_17 => X"000000840000000000000088000000000000008b000000000000008e00000000",
            INIT_18 => X"0000001200000000000000190000000000000019000000000000001800000000",
            INIT_19 => X"00000073000000000000006a000000000000007c000000000000004500000000",
            INIT_1A => X"00000078000000000000009200000000000000a6000000000000009c00000000",
            INIT_1B => X"0000009700000000000000950000000000000094000000000000008900000000",
            INIT_1C => X"0000006d0000000000000094000000000000009c000000000000009600000000",
            INIT_1D => X"000000a900000000000000b1000000000000007a000000000000004a00000000",
            INIT_1E => X"000000950000000000000098000000000000009d00000000000000a100000000",
            INIT_1F => X"0000008e00000000000000910000000000000094000000000000009600000000",
            INIT_20 => X"0000001700000000000000190000000000000018000000000000001900000000",
            INIT_21 => X"000000680000000000000060000000000000006d000000000000003300000000",
            INIT_22 => X"0000008d00000000000000b200000000000000b800000000000000a100000000",
            INIT_23 => X"0000009300000000000000860000000000000080000000000000007c00000000",
            INIT_24 => X"0000006c00000000000000890000000000000096000000000000009700000000",
            INIT_25 => X"000000b500000000000000b70000000000000098000000000000006000000000",
            INIT_26 => X"000000a400000000000000a800000000000000ae00000000000000b300000000",
            INIT_27 => X"000000930000000000000098000000000000009c00000000000000a000000000",
            INIT_28 => X"0000001c000000000000001b000000000000001a000000000000001a00000000",
            INIT_29 => X"00000066000000000000005f0000000000000059000000000000002300000000",
            INIT_2A => X"0000009f00000000000000c700000000000000c1000000000000009600000000",
            INIT_2B => X"0000007600000000000000620000000000000066000000000000007400000000",
            INIT_2C => X"0000007a00000000000000770000000000000083000000000000008200000000",
            INIT_2D => X"000000aa00000000000000a600000000000000a7000000000000008400000000",
            INIT_2E => X"000000b700000000000000b300000000000000b700000000000000b200000000",
            INIT_2F => X"000000a900000000000000af00000000000000b100000000000000b700000000",
            INIT_30 => X"0000001a00000000000000190000000000000016000000000000001a00000000",
            INIT_31 => X"0000007b0000000000000080000000000000005c000000000000001d00000000",
            INIT_32 => X"000000ab00000000000000c700000000000000c3000000000000009300000000",
            INIT_33 => X"0000006a0000000000000063000000000000005e000000000000007e00000000",
            INIT_34 => X"0000007a0000000000000065000000000000006d000000000000006000000000",
            INIT_35 => X"000000b000000000000000aa00000000000000c000000000000000ac00000000",
            INIT_36 => X"000000ca00000000000000c500000000000000c400000000000000c300000000",
            INIT_37 => X"000000c200000000000000bf00000000000000bf00000000000000c500000000",
            INIT_38 => X"0000001900000000000000110000000000000021000000000000004d00000000",
            INIT_39 => X"0000007e000000000000009b000000000000009a000000000000005800000000",
            INIT_3A => X"000000b900000000000000c100000000000000be000000000000008c00000000",
            INIT_3B => X"00000071000000000000007b000000000000008100000000000000a300000000",
            INIT_3C => X"0000007900000000000000680000000000000067000000000000005800000000",
            INIT_3D => X"000000bd00000000000000a500000000000000c600000000000000b100000000",
            INIT_3E => X"000000da00000000000000e000000000000000db00000000000000e400000000",
            INIT_3F => X"000000cd00000000000000c400000000000000bb00000000000000ba00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006000000000000000560000000000000080000000000000009500000000",
            INIT_41 => X"00000077000000000000009900000000000000a7000000000000009b00000000",
            INIT_42 => X"000000bf00000000000000bf00000000000000a8000000000000006f00000000",
            INIT_43 => X"0000007f000000000000009400000000000000aa00000000000000b700000000",
            INIT_44 => X"0000007c00000000000000740000000000000070000000000000007000000000",
            INIT_45 => X"000000c100000000000000a200000000000000bb00000000000000a300000000",
            INIT_46 => X"000000bb00000000000000cf00000000000000d500000000000000df00000000",
            INIT_47 => X"000000d200000000000000c400000000000000a6000000000000009d00000000",
            INIT_48 => X"0000009b0000000000000092000000000000009e00000000000000a100000000",
            INIT_49 => X"00000075000000000000009f00000000000000a900000000000000a700000000",
            INIT_4A => X"000000b500000000000000b3000000000000009b000000000000006800000000",
            INIT_4B => X"00000087000000000000009f00000000000000b400000000000000b600000000",
            INIT_4C => X"0000007900000000000000750000000000000074000000000000006400000000",
            INIT_4D => X"000000cc00000000000000b200000000000000b2000000000000009e00000000",
            INIT_4E => X"000000a700000000000000cb00000000000000d600000000000000d800000000",
            INIT_4F => X"000000cf00000000000000b00000000000000096000000000000009300000000",
            INIT_50 => X"000000a5000000000000009e00000000000000a500000000000000aa00000000",
            INIT_51 => X"0000007000000000000000a000000000000000b000000000000000af00000000",
            INIT_52 => X"000000b400000000000000b100000000000000a4000000000000007b00000000",
            INIT_53 => X"00000079000000000000009500000000000000ac00000000000000b600000000",
            INIT_54 => X"0000007600000000000000750000000000000074000000000000006a00000000",
            INIT_55 => X"000000d100000000000000af00000000000000a6000000000000009c00000000",
            INIT_56 => X"000000a900000000000000cd00000000000000d800000000000000de00000000",
            INIT_57 => X"000000ba000000000000009f0000000000000093000000000000009100000000",
            INIT_58 => X"000000a600000000000000a900000000000000ae00000000000000ac00000000",
            INIT_59 => X"0000007a000000000000009d00000000000000b000000000000000b000000000",
            INIT_5A => X"000000b600000000000000b900000000000000b1000000000000008d00000000",
            INIT_5B => X"00000068000000000000007f000000000000009d00000000000000b600000000",
            INIT_5C => X"0000007d000000000000007b0000000000000084000000000000007300000000",
            INIT_5D => X"000000ce00000000000000a300000000000000a4000000000000009f00000000",
            INIT_5E => X"000000b500000000000000cd00000000000000d900000000000000e000000000",
            INIT_5F => X"0000009c0000000000000093000000000000008e000000000000009200000000",
            INIT_60 => X"000000a000000000000000a500000000000000a700000000000000a700000000",
            INIT_61 => X"0000008f000000000000009900000000000000a400000000000000a500000000",
            INIT_62 => X"000000a400000000000000ae00000000000000a3000000000000009100000000",
            INIT_63 => X"000000760000000000000085000000000000009f00000000000000a300000000",
            INIT_64 => X"000000920000000000000087000000000000009f000000000000008600000000",
            INIT_65 => X"000000cd00000000000000a800000000000000a300000000000000a300000000",
            INIT_66 => X"000000c700000000000000d600000000000000dc00000000000000df00000000",
            INIT_67 => X"000000980000000000000090000000000000009000000000000000a300000000",
            INIT_68 => X"0000009b00000000000000a000000000000000a200000000000000a900000000",
            INIT_69 => X"000000a40000000000000083000000000000008800000000000000a300000000",
            INIT_6A => X"0000008500000000000000840000000000000088000000000000009200000000",
            INIT_6B => X"000000920000000000000087000000000000009e000000000000009f00000000",
            INIT_6C => X"0000009e000000000000009000000000000000a200000000000000a700000000",
            INIT_6D => X"000000cb00000000000000b00000000000000098000000000000009800000000",
            INIT_6E => X"000000da00000000000000dd00000000000000d800000000000000d700000000",
            INIT_6F => X"000000b600000000000000a2000000000000009f00000000000000c500000000",
            INIT_70 => X"0000009d00000000000000a200000000000000a400000000000000ae00000000",
            INIT_71 => X"000000b2000000000000006d000000000000007800000000000000a800000000",
            INIT_72 => X"000000a300000000000000a100000000000000a700000000000000a600000000",
            INIT_73 => X"00000078000000000000008400000000000000ab00000000000000b600000000",
            INIT_74 => X"00000095000000000000008c00000000000000a300000000000000a900000000",
            INIT_75 => X"000000cc00000000000000aa00000000000000a400000000000000a600000000",
            INIT_76 => X"000000e400000000000000da00000000000000d500000000000000d300000000",
            INIT_77 => X"000000c700000000000000bb00000000000000b000000000000000d600000000",
            INIT_78 => X"0000009f00000000000000a100000000000000a000000000000000af00000000",
            INIT_79 => X"000000b70000000000000068000000000000008400000000000000aa00000000",
            INIT_7A => X"000000b000000000000000b800000000000000b600000000000000bc00000000",
            INIT_7B => X"0000008d00000000000000a300000000000000a800000000000000a200000000",
            INIT_7C => X"00000085000000000000009200000000000000a5000000000000009100000000",
            INIT_7D => X"000000a9000000000000009600000000000000a500000000000000af00000000",
            INIT_7E => X"000000dd00000000000000d900000000000000d400000000000000ca00000000",
            INIT_7F => X"000000c700000000000000c700000000000000ba00000000000000c400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE52;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE53 : if BRAM_NAME = "sampleifmap_layersamples_instance53" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000940000000000000092000000000000009f00000000000000b300000000",
            INIT_01 => X"000000a8000000000000006d000000000000009700000000000000a100000000",
            INIT_02 => X"000000ae00000000000000a400000000000000b500000000000000c700000000",
            INIT_03 => X"000000a600000000000000aa000000000000009c00000000000000a500000000",
            INIT_04 => X"00000077000000000000009f0000000000000088000000000000006900000000",
            INIT_05 => X"00000050000000000000007e000000000000009e000000000000008f00000000",
            INIT_06 => X"000000cd00000000000000d100000000000000b7000000000000007600000000",
            INIT_07 => X"000000c500000000000000c900000000000000b700000000000000af00000000",
            INIT_08 => X"00000083000000000000008500000000000000a400000000000000b500000000",
            INIT_09 => X"0000009f000000000000009700000000000000a5000000000000009500000000",
            INIT_0A => X"000000cd00000000000000c400000000000000c700000000000000c200000000",
            INIT_0B => X"000000a200000000000000ac00000000000000a800000000000000b900000000",
            INIT_0C => X"00000077000000000000009b0000000000000069000000000000006800000000",
            INIT_0D => X"0000005c000000000000008800000000000000ad000000000000008600000000",
            INIT_0E => X"0000009e0000000000000098000000000000006f000000000000004b00000000",
            INIT_0F => X"000000c800000000000000cb00000000000000b0000000000000009800000000",
            INIT_10 => X"00000085000000000000008e00000000000000ac00000000000000b700000000",
            INIT_11 => X"000000aa00000000000000b100000000000000b0000000000000009f00000000",
            INIT_12 => X"000000d900000000000000cf00000000000000c500000000000000b100000000",
            INIT_13 => X"000000aa00000000000000bb00000000000000c600000000000000d900000000",
            INIT_14 => X"0000007e0000000000000085000000000000005a000000000000008300000000",
            INIT_15 => X"0000007e000000000000008200000000000000a2000000000000008b00000000",
            INIT_16 => X"0000008400000000000000760000000000000060000000000000006f00000000",
            INIT_17 => X"000000c700000000000000b80000000000000092000000000000007c00000000",
            INIT_18 => X"0000009500000000000000a100000000000000b000000000000000b900000000",
            INIT_19 => X"000000bc00000000000000b600000000000000b700000000000000af00000000",
            INIT_1A => X"000000c200000000000000b900000000000000aa00000000000000aa00000000",
            INIT_1B => X"000000af00000000000000ca00000000000000d000000000000000c900000000",
            INIT_1C => X"000000910000000000000071000000000000007b00000000000000a400000000",
            INIT_1D => X"0000007b0000000000000071000000000000008c000000000000009d00000000",
            INIT_1E => X"0000008e00000000000000860000000000000070000000000000007700000000",
            INIT_1F => X"000000a600000000000000840000000000000079000000000000007f00000000",
            INIT_20 => X"0000009b00000000000000ad00000000000000b700000000000000bd00000000",
            INIT_21 => X"000000b200000000000000b100000000000000ba00000000000000ab00000000",
            INIT_22 => X"000000b100000000000000b200000000000000ac00000000000000b400000000",
            INIT_23 => X"000000bd00000000000000c300000000000000bc00000000000000a400000000",
            INIT_24 => X"0000009d000000000000008800000000000000b600000000000000c900000000",
            INIT_25 => X"0000007c000000000000006a0000000000000078000000000000009300000000",
            INIT_26 => X"0000008a0000000000000094000000000000008a000000000000008000000000",
            INIT_27 => X"00000082000000000000007a0000000000000077000000000000007800000000",
            INIT_28 => X"000000a100000000000000b700000000000000bc00000000000000bd00000000",
            INIT_29 => X"000000b000000000000000bb00000000000000b7000000000000009e00000000",
            INIT_2A => X"000000a400000000000000c000000000000000bf00000000000000b800000000",
            INIT_2B => X"000000b100000000000000ad00000000000000a6000000000000008b00000000",
            INIT_2C => X"0000009600000000000000a200000000000000bc00000000000000c000000000",
            INIT_2D => X"000000850000000000000079000000000000006b000000000000007600000000",
            INIT_2E => X"0000007d000000000000008d0000000000000096000000000000008e00000000",
            INIT_2F => X"0000006c000000000000007d000000000000007c000000000000007500000000",
            INIT_30 => X"000000a600000000000000bb00000000000000ba00000000000000ba00000000",
            INIT_31 => X"000000c500000000000000c700000000000000b4000000000000009400000000",
            INIT_32 => X"000000a800000000000000c000000000000000c300000000000000c100000000",
            INIT_33 => X"000000aa00000000000000a9000000000000009f000000000000009100000000",
            INIT_34 => X"0000008600000000000000a300000000000000ac00000000000000af00000000",
            INIT_35 => X"0000008b0000000000000086000000000000006c000000000000005d00000000",
            INIT_36 => X"0000007c000000000000008e0000000000000097000000000000008d00000000",
            INIT_37 => X"0000005b00000000000000650000000000000072000000000000007c00000000",
            INIT_38 => X"000000ac00000000000000b700000000000000b500000000000000ba00000000",
            INIT_39 => X"000000cf00000000000000c900000000000000b0000000000000008f00000000",
            INIT_3A => X"000000af00000000000000bd00000000000000cb00000000000000ce00000000",
            INIT_3B => X"000000ac00000000000000ae00000000000000ab00000000000000a500000000",
            INIT_3C => X"00000075000000000000009e00000000000000ab00000000000000b200000000",
            INIT_3D => X"00000088000000000000008a0000000000000078000000000000006100000000",
            INIT_3E => X"00000084000000000000009200000000000000a1000000000000008a00000000",
            INIT_3F => X"000000680000000000000064000000000000006d000000000000008200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a900000000000000af00000000000000b200000000000000b800000000",
            INIT_41 => X"000000ca00000000000000c600000000000000aa000000000000009200000000",
            INIT_42 => X"0000008800000000000000ab00000000000000c500000000000000c800000000",
            INIT_43 => X"000000aa00000000000000ab00000000000000b400000000000000a100000000",
            INIT_44 => X"00000073000000000000009000000000000000a800000000000000ad00000000",
            INIT_45 => X"0000007e0000000000000086000000000000007c000000000000006c00000000",
            INIT_46 => X"0000008700000000000000910000000000000099000000000000008200000000",
            INIT_47 => X"0000006f00000000000000740000000000000075000000000000007700000000",
            INIT_48 => X"0000009d00000000000000a800000000000000b000000000000000b800000000",
            INIT_49 => X"000000c800000000000000c000000000000000a2000000000000009300000000",
            INIT_4A => X"00000052000000000000008100000000000000b900000000000000bf00000000",
            INIT_4B => X"0000009f00000000000000a600000000000000b3000000000000008d00000000",
            INIT_4C => X"0000007400000000000000840000000000000096000000000000009f00000000",
            INIT_4D => X"0000007a000000000000007f000000000000007a000000000000006900000000",
            INIT_4E => X"0000007a00000000000000800000000000000084000000000000007f00000000",
            INIT_4F => X"00000062000000000000006b0000000000000077000000000000007700000000",
            INIT_50 => X"0000009400000000000000a300000000000000ac00000000000000b800000000",
            INIT_51 => X"000000ca00000000000000ba0000000000000092000000000000008600000000",
            INIT_52 => X"00000058000000000000008200000000000000b200000000000000c000000000",
            INIT_53 => X"00000090000000000000009800000000000000ac000000000000008c00000000",
            INIT_54 => X"00000069000000000000007a0000000000000084000000000000009100000000",
            INIT_55 => X"0000007000000000000000790000000000000077000000000000006400000000",
            INIT_56 => X"0000006c00000000000000640000000000000071000000000000007a00000000",
            INIT_57 => X"000000720000000000000075000000000000007a000000000000007c00000000",
            INIT_58 => X"0000008e000000000000009e00000000000000a900000000000000b700000000",
            INIT_59 => X"000000cc00000000000000b20000000000000084000000000000007e00000000",
            INIT_5A => X"00000090000000000000009d00000000000000af00000000000000c300000000",
            INIT_5B => X"000000830000000000000087000000000000009800000000000000a400000000",
            INIT_5C => X"00000054000000000000006f0000000000000074000000000000007c00000000",
            INIT_5D => X"0000006d00000000000000710000000000000073000000000000006100000000",
            INIT_5E => X"00000064000000000000005f0000000000000066000000000000007200000000",
            INIT_5F => X"0000007b00000000000000820000000000000082000000000000007400000000",
            INIT_60 => X"0000008e000000000000009900000000000000a100000000000000b100000000",
            INIT_61 => X"000000cc00000000000000b2000000000000007a000000000000007700000000",
            INIT_62 => X"000000a800000000000000aa00000000000000b400000000000000c500000000",
            INIT_63 => X"0000007b000000000000007a0000000000000087000000000000009d00000000",
            INIT_64 => X"0000004b000000000000005e000000000000006d000000000000007700000000",
            INIT_65 => X"000000710000000000000070000000000000006f000000000000006800000000",
            INIT_66 => X"00000066000000000000005c0000000000000064000000000000007000000000",
            INIT_67 => X"00000073000000000000007e0000000000000082000000000000007700000000",
            INIT_68 => X"00000091000000000000008d000000000000009000000000000000a300000000",
            INIT_69 => X"000000c800000000000000a9000000000000006b000000000000007400000000",
            INIT_6A => X"000000a300000000000000ac00000000000000b700000000000000c200000000",
            INIT_6B => X"0000007900000000000000730000000000000081000000000000009600000000",
            INIT_6C => X"00000051000000000000004e0000000000000064000000000000007000000000",
            INIT_6D => X"00000072000000000000006a0000000000000065000000000000006800000000",
            INIT_6E => X"0000007000000000000000630000000000000063000000000000007200000000",
            INIT_6F => X"0000006e00000000000000740000000000000075000000000000007600000000",
            INIT_70 => X"0000008f0000000000000083000000000000007e000000000000008e00000000",
            INIT_71 => X"000000c00000000000000091000000000000005f000000000000007c00000000",
            INIT_72 => X"000000a800000000000000b200000000000000b700000000000000be00000000",
            INIT_73 => X"00000065000000000000005c0000000000000062000000000000008200000000",
            INIT_74 => X"0000005f000000000000004b000000000000005c000000000000006800000000",
            INIT_75 => X"00000074000000000000006a0000000000000061000000000000006300000000",
            INIT_76 => X"0000006e0000000000000071000000000000006c000000000000006d00000000",
            INIT_77 => X"000000770000000000000074000000000000006c000000000000006700000000",
            INIT_78 => X"0000007800000000000000700000000000000068000000000000007b00000000",
            INIT_79 => X"000000ae00000000000000760000000000000057000000000000007400000000",
            INIT_7A => X"0000008d00000000000000a400000000000000ae00000000000000b500000000",
            INIT_7B => X"0000004600000000000000390000000000000045000000000000006300000000",
            INIT_7C => X"0000006000000000000000580000000000000051000000000000005700000000",
            INIT_7D => X"00000070000000000000006b000000000000005e000000000000005d00000000",
            INIT_7E => X"0000005d0000000000000061000000000000006c000000000000006b00000000",
            INIT_7F => X"00000076000000000000007b0000000000000076000000000000006500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE53;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE54 : if BRAM_NAME = "sampleifmap_layersamples_instance54" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000c700000000000000cd00000000000000d200000000000000d900000000",
            INIT_01 => X"000000bd00000000000000cf00000000000000d600000000000000da00000000",
            INIT_02 => X"000000a900000000000000a600000000000000ae00000000000000bb00000000",
            INIT_03 => X"0000008f000000000000008c000000000000009a000000000000009600000000",
            INIT_04 => X"000000df00000000000000db00000000000000bf00000000000000a700000000",
            INIT_05 => X"000000e100000000000000e200000000000000d700000000000000db00000000",
            INIT_06 => X"000000bb00000000000000af00000000000000be00000000000000db00000000",
            INIT_07 => X"000000a200000000000000a100000000000000aa00000000000000c800000000",
            INIT_08 => X"000000d700000000000000dc00000000000000dd00000000000000de00000000",
            INIT_09 => X"000000b300000000000000d300000000000000e100000000000000d800000000",
            INIT_0A => X"000000bc00000000000000be00000000000000c000000000000000b400000000",
            INIT_0B => X"000000db00000000000000d100000000000000ce00000000000000c700000000",
            INIT_0C => X"000000ec00000000000000ec00000000000000eb00000000000000e500000000",
            INIT_0D => X"000000e500000000000000e100000000000000e200000000000000e900000000",
            INIT_0E => X"000000cd00000000000000d000000000000000d400000000000000e700000000",
            INIT_0F => X"000000c800000000000000ba00000000000000b700000000000000d800000000",
            INIT_10 => X"000000e800000000000000e700000000000000e900000000000000ea00000000",
            INIT_11 => X"000000ad00000000000000d900000000000000ef00000000000000e900000000",
            INIT_12 => X"000000b700000000000000ad00000000000000b400000000000000a400000000",
            INIT_13 => X"000000e000000000000000d400000000000000bc00000000000000be00000000",
            INIT_14 => X"000000e100000000000000e300000000000000eb00000000000000da00000000",
            INIT_15 => X"000000e100000000000000d600000000000000df00000000000000e500000000",
            INIT_16 => X"000000d800000000000000e600000000000000e800000000000000ea00000000",
            INIT_17 => X"000000d300000000000000d000000000000000ca00000000000000d100000000",
            INIT_18 => X"000000f200000000000000f400000000000000f400000000000000f500000000",
            INIT_19 => X"0000009e00000000000000e400000000000000f300000000000000f400000000",
            INIT_1A => X"0000009f0000000000000083000000000000009d000000000000009200000000",
            INIT_1B => X"0000009f00000000000000a20000000000000088000000000000009100000000",
            INIT_1C => X"000000d300000000000000c300000000000000cb00000000000000a900000000",
            INIT_1D => X"000000e200000000000000d000000000000000cb00000000000000d100000000",
            INIT_1E => X"000000d500000000000000e400000000000000e900000000000000e600000000",
            INIT_1F => X"000000d400000000000000e000000000000000db00000000000000c700000000",
            INIT_20 => X"000000f400000000000000f400000000000000f300000000000000f500000000",
            INIT_21 => X"0000007500000000000000cf00000000000000f100000000000000f500000000",
            INIT_22 => X"0000006b0000000000000059000000000000006c000000000000006300000000",
            INIT_23 => X"0000005c0000000000000064000000000000005b000000000000006400000000",
            INIT_24 => X"00000095000000000000007c000000000000007c000000000000006600000000",
            INIT_25 => X"000000e900000000000000ca00000000000000b900000000000000b600000000",
            INIT_26 => X"000000cd00000000000000e300000000000000e200000000000000e100000000",
            INIT_27 => X"000000de00000000000000e200000000000000d500000000000000c200000000",
            INIT_28 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_29 => X"0000007e00000000000000d800000000000000ed00000000000000f500000000",
            INIT_2A => X"00000066000000000000005b000000000000005a000000000000004800000000",
            INIT_2B => X"00000063000000000000006b0000000000000067000000000000006500000000",
            INIT_2C => X"0000005d000000000000005b0000000000000059000000000000005900000000",
            INIT_2D => X"000000eb00000000000000d800000000000000be000000000000007e00000000",
            INIT_2E => X"000000c400000000000000d800000000000000df00000000000000e700000000",
            INIT_2F => X"000000ec00000000000000d900000000000000bd00000000000000ae00000000",
            INIT_30 => X"000000f400000000000000f300000000000000f300000000000000f500000000",
            INIT_31 => X"0000009e00000000000000d900000000000000db00000000000000f100000000",
            INIT_32 => X"0000009700000000000000840000000000000072000000000000005000000000",
            INIT_33 => X"0000008a000000000000008f0000000000000084000000000000008c00000000",
            INIT_34 => X"000000780000000000000072000000000000007a000000000000008200000000",
            INIT_35 => X"000000e900000000000000dd000000000000009b000000000000006e00000000",
            INIT_36 => X"000000c000000000000000c600000000000000e000000000000000eb00000000",
            INIT_37 => X"000000eb00000000000000cc00000000000000ab00000000000000a700000000",
            INIT_38 => X"000000f600000000000000f300000000000000f300000000000000f400000000",
            INIT_39 => X"0000009900000000000000d700000000000000c700000000000000e300000000",
            INIT_3A => X"000000ca00000000000000bb0000000000000092000000000000005100000000",
            INIT_3B => X"000000830000000000000083000000000000009e00000000000000cf00000000",
            INIT_3C => X"000000840000000000000083000000000000008d000000000000008100000000",
            INIT_3D => X"000000d7000000000000009f0000000000000084000000000000009f00000000",
            INIT_3E => X"000000d100000000000000d400000000000000d700000000000000e500000000",
            INIT_3F => X"000000dd00000000000000b200000000000000ab00000000000000c500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f500000000000000f400000000000000f300000000000000f400000000",
            INIT_41 => X"0000008200000000000000da00000000000000ce00000000000000e300000000",
            INIT_42 => X"0000008100000000000000800000000000000082000000000000005100000000",
            INIT_43 => X"0000007d0000000000000074000000000000009100000000000000b800000000",
            INIT_44 => X"0000007d000000000000008e0000000000000089000000000000007c00000000",
            INIT_45 => X"000000c600000000000000900000000000000093000000000000009900000000",
            INIT_46 => X"000000dc00000000000000e900000000000000db00000000000000d600000000",
            INIT_47 => X"000000c900000000000000a900000000000000a400000000000000b800000000",
            INIT_48 => X"000000f200000000000000f400000000000000f300000000000000f300000000",
            INIT_49 => X"0000006e00000000000000a800000000000000be00000000000000e400000000",
            INIT_4A => X"0000006e00000000000000770000000000000086000000000000005300000000",
            INIT_4B => X"0000007800000000000000730000000000000080000000000000008f00000000",
            INIT_4C => X"0000007d00000000000000920000000000000083000000000000007d00000000",
            INIT_4D => X"000000c4000000000000008c000000000000009b000000000000009500000000",
            INIT_4E => X"000000e900000000000000f000000000000000f000000000000000e900000000",
            INIT_4F => X"000000dc00000000000000d700000000000000c800000000000000c800000000",
            INIT_50 => X"000000f500000000000000f400000000000000f100000000000000ef00000000",
            INIT_51 => X"0000005f0000000000000082000000000000008500000000000000dc00000000",
            INIT_52 => X"0000006c00000000000000740000000000000074000000000000004e00000000",
            INIT_53 => X"0000006c000000000000006d000000000000006b000000000000006d00000000",
            INIT_54 => X"0000007300000000000000780000000000000078000000000000007300000000",
            INIT_55 => X"000000a7000000000000008f0000000000000096000000000000008800000000",
            INIT_56 => X"000000f300000000000000f500000000000000e400000000000000d000000000",
            INIT_57 => X"000000f400000000000000f500000000000000f500000000000000f400000000",
            INIT_58 => X"000000f400000000000000f200000000000000e900000000000000de00000000",
            INIT_59 => X"0000005900000000000000a500000000000000a900000000000000d800000000",
            INIT_5A => X"00000064000000000000005b0000000000000043000000000000003d00000000",
            INIT_5B => X"000000600000000000000062000000000000005f000000000000005f00000000",
            INIT_5C => X"00000061000000000000005a000000000000005f000000000000006000000000",
            INIT_5D => X"0000007e00000000000000810000000000000079000000000000006900000000",
            INIT_5E => X"000000f300000000000000f800000000000000d8000000000000009b00000000",
            INIT_5F => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_60 => X"000000e300000000000000ec00000000000000df00000000000000d000000000",
            INIT_61 => X"0000006400000000000000b500000000000000b700000000000000bf00000000",
            INIT_62 => X"0000006500000000000000580000000000000038000000000000003700000000",
            INIT_63 => X"0000005400000000000000560000000000000063000000000000006f00000000",
            INIT_64 => X"00000071000000000000005d0000000000000054000000000000005200000000",
            INIT_65 => X"0000008100000000000000700000000000000062000000000000006d00000000",
            INIT_66 => X"000000f400000000000000f500000000000000e200000000000000ae00000000",
            INIT_67 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_68 => X"000000c300000000000000db00000000000000cc00000000000000c800000000",
            INIT_69 => X"00000066000000000000009c000000000000009a00000000000000aa00000000",
            INIT_6A => X"00000066000000000000006c0000000000000063000000000000006800000000",
            INIT_6B => X"00000055000000000000005e0000000000000075000000000000007300000000",
            INIT_6C => X"0000008c000000000000007a000000000000006a000000000000005a00000000",
            INIT_6D => X"0000007c000000000000006c0000000000000068000000000000008000000000",
            INIT_6E => X"000000d400000000000000c300000000000000b3000000000000009600000000",
            INIT_6F => X"000000f400000000000000f400000000000000f500000000000000ef00000000",
            INIT_70 => X"000000a900000000000000cf00000000000000d200000000000000c800000000",
            INIT_71 => X"0000008a0000000000000093000000000000009400000000000000a400000000",
            INIT_72 => X"0000005d000000000000006a000000000000005c000000000000008100000000",
            INIT_73 => X"0000004d0000000000000054000000000000005d000000000000005900000000",
            INIT_74 => X"0000005100000000000000510000000000000051000000000000004c00000000",
            INIT_75 => X"00000052000000000000004b000000000000004a000000000000004f00000000",
            INIT_76 => X"0000008f000000000000008c000000000000007b000000000000006500000000",
            INIT_77 => X"000000f400000000000000f400000000000000f400000000000000bf00000000",
            INIT_78 => X"0000007700000000000000c400000000000000e200000000000000d200000000",
            INIT_79 => X"000000c000000000000000ba0000000000000096000000000000007000000000",
            INIT_7A => X"00000037000000000000004d000000000000004d000000000000006c00000000",
            INIT_7B => X"0000003f000000000000003c000000000000002f000000000000002d00000000",
            INIT_7C => X"00000036000000000000003b000000000000003f000000000000003b00000000",
            INIT_7D => X"00000040000000000000003d0000000000000032000000000000003100000000",
            INIT_7E => X"00000067000000000000005b000000000000004b000000000000004700000000",
            INIT_7F => X"000000f400000000000000f600000000000000e1000000000000008700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE54;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE55 : if BRAM_NAME = "sampleifmap_layersamples_instance55" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000006000000000000000b400000000000000c100000000000000c700000000",
            INIT_01 => X"000000a100000000000000c00000000000000091000000000000005d00000000",
            INIT_02 => X"00000062000000000000005c0000000000000049000000000000005600000000",
            INIT_03 => X"00000047000000000000004f000000000000004f000000000000006800000000",
            INIT_04 => X"0000001b000000000000001e000000000000001c000000000000002500000000",
            INIT_05 => X"0000001c00000000000000160000000000000032000000000000003400000000",
            INIT_06 => X"00000068000000000000005b0000000000000035000000000000001800000000",
            INIT_07 => X"000000f300000000000000f700000000000000ce000000000000008000000000",
            INIT_08 => X"0000007100000000000000c200000000000000c700000000000000d300000000",
            INIT_09 => X"00000047000000000000009f000000000000009d000000000000007800000000",
            INIT_0A => X"0000007c0000000000000074000000000000005a000000000000004400000000",
            INIT_0B => X"0000006600000000000000800000000000000079000000000000009500000000",
            INIT_0C => X"0000006400000000000000700000000000000062000000000000004e00000000",
            INIT_0D => X"00000063000000000000005c0000000000000093000000000000009400000000",
            INIT_0E => X"0000008e0000000000000087000000000000006c000000000000005e00000000",
            INIT_0F => X"000000f500000000000000f200000000000000b7000000000000009c00000000",
            INIT_10 => X"0000006600000000000000b700000000000000ca00000000000000dc00000000",
            INIT_11 => X"0000001e000000000000008400000000000000a5000000000000006e00000000",
            INIT_12 => X"00000053000000000000006b0000000000000062000000000000003900000000",
            INIT_13 => X"0000006400000000000000810000000000000065000000000000005200000000",
            INIT_14 => X"0000009f000000000000009e00000000000000ae000000000000009900000000",
            INIT_15 => X"000000a300000000000000a200000000000000a800000000000000ac00000000",
            INIT_16 => X"00000077000000000000009c00000000000000af00000000000000a000000000",
            INIT_17 => X"000000f700000000000000e40000000000000087000000000000007200000000",
            INIT_18 => X"0000006200000000000000bc00000000000000cf00000000000000db00000000",
            INIT_19 => X"0000002a000000000000006f000000000000008d000000000000005300000000",
            INIT_1A => X"0000003e000000000000004c0000000000000048000000000000003a00000000",
            INIT_1B => X"0000005d00000000000000400000000000000038000000000000003500000000",
            INIT_1C => X"00000065000000000000005b000000000000007c00000000000000a000000000",
            INIT_1D => X"000000670000000000000067000000000000006b000000000000007400000000",
            INIT_1E => X"00000043000000000000007e000000000000009b000000000000006300000000",
            INIT_1F => X"000000f800000000000000d90000000000000076000000000000005100000000",
            INIT_20 => X"0000006500000000000000c700000000000000d200000000000000d900000000",
            INIT_21 => X"0000003c000000000000005d0000000000000058000000000000003800000000",
            INIT_22 => X"00000046000000000000003f000000000000002e000000000000003800000000",
            INIT_23 => X"0000004100000000000000400000000000000036000000000000003c00000000",
            INIT_24 => X"0000006700000000000000690000000000000072000000000000006300000000",
            INIT_25 => X"00000061000000000000005d0000000000000060000000000000006400000000",
            INIT_26 => X"000000490000000000000064000000000000006f000000000000006600000000",
            INIT_27 => X"000000f900000000000000d40000000000000072000000000000005200000000",
            INIT_28 => X"0000007500000000000000ca00000000000000cd00000000000000d100000000",
            INIT_29 => X"0000004400000000000000510000000000000046000000000000005300000000",
            INIT_2A => X"00000033000000000000002b0000000000000023000000000000003200000000",
            INIT_2B => X"0000003f0000000000000057000000000000004d000000000000004400000000",
            INIT_2C => X"0000004800000000000000520000000000000047000000000000003400000000",
            INIT_2D => X"0000005d000000000000003e0000000000000043000000000000004000000000",
            INIT_2E => X"0000006c0000000000000053000000000000003c000000000000005800000000",
            INIT_2F => X"000000fa00000000000000cc000000000000006c000000000000007000000000",
            INIT_30 => X"0000006800000000000000c500000000000000ca00000000000000cd00000000",
            INIT_31 => X"000000490000000000000047000000000000006f000000000000005d00000000",
            INIT_32 => X"0000002200000000000000260000000000000029000000000000003f00000000",
            INIT_33 => X"0000004f000000000000008e0000000000000063000000000000004b00000000",
            INIT_34 => X"0000007600000000000000930000000000000056000000000000001e00000000",
            INIT_35 => X"0000009900000000000000660000000000000072000000000000006300000000",
            INIT_36 => X"0000008d000000000000004a000000000000003f00000000000000b200000000",
            INIT_37 => X"000000f600000000000000c3000000000000005a000000000000007700000000",
            INIT_38 => X"0000005700000000000000b900000000000000c200000000000000c600000000",
            INIT_39 => X"000000630000000000000061000000000000006c000000000000003100000000",
            INIT_3A => X"0000002400000000000000270000000000000033000000000000005f00000000",
            INIT_3B => X"0000003700000000000000570000000000000032000000000000002800000000",
            INIT_3C => X"0000007f0000000000000097000000000000004f000000000000002000000000",
            INIT_3D => X"0000009c00000000000000740000000000000088000000000000007a00000000",
            INIT_3E => X"0000004a00000000000000350000000000000037000000000000009f00000000",
            INIT_3F => X"000000f000000000000000c2000000000000004e000000000000003e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004d00000000000000a900000000000000b400000000000000b600000000",
            INIT_41 => X"00000090000000000000006c000000000000003b000000000000002500000000",
            INIT_42 => X"00000020000000000000002b000000000000003c000000000000006a00000000",
            INIT_43 => X"00000021000000000000001e000000000000001c000000000000001d00000000",
            INIT_44 => X"00000058000000000000003a000000000000002a000000000000002700000000",
            INIT_45 => X"00000075000000000000007a0000000000000079000000000000006a00000000",
            INIT_46 => X"000000320000000000000033000000000000002f000000000000004300000000",
            INIT_47 => X"000000e100000000000000ba0000000000000050000000000000003300000000",
            INIT_48 => X"0000007d00000000000000a400000000000000a500000000000000a800000000",
            INIT_49 => X"0000008d000000000000006f0000000000000060000000000000005b00000000",
            INIT_4A => X"000000240000000000000037000000000000004a000000000000006000000000",
            INIT_4B => X"0000001f000000000000001d000000000000001e000000000000001e00000000",
            INIT_4C => X"000000ae00000000000000400000000000000018000000000000002300000000",
            INIT_4D => X"000000b500000000000000b300000000000000cb00000000000000cd00000000",
            INIT_4E => X"00000030000000000000002b0000000000000026000000000000005700000000",
            INIT_4F => X"000000d300000000000000ae000000000000005b000000000000004200000000",
            INIT_50 => X"000000b400000000000000af00000000000000a300000000000000a200000000",
            INIT_51 => X"0000008d000000000000006c0000000000000076000000000000009800000000",
            INIT_52 => X"00000030000000000000004e0000000000000053000000000000005b00000000",
            INIT_53 => X"0000001d00000000000000190000000000000018000000000000001900000000",
            INIT_54 => X"000000a400000000000000470000000000000026000000000000002700000000",
            INIT_55 => X"000000a600000000000000a900000000000000b100000000000000b800000000",
            INIT_56 => X"00000031000000000000001e000000000000001e000000000000005100000000",
            INIT_57 => X"000000ce00000000000000a9000000000000005f000000000000004e00000000",
            INIT_58 => X"000000a600000000000000b300000000000000ac000000000000009a00000000",
            INIT_59 => X"0000009200000000000000670000000000000075000000000000009200000000",
            INIT_5A => X"0000003600000000000000520000000000000055000000000000005700000000",
            INIT_5B => X"000000250000000000000021000000000000001e000000000000002000000000",
            INIT_5C => X"000000650000000000000056000000000000004d000000000000003600000000",
            INIT_5D => X"00000089000000000000008e0000000000000079000000000000006b00000000",
            INIT_5E => X"000000360000000000000021000000000000001e000000000000003c00000000",
            INIT_5F => X"000000c700000000000000a5000000000000005b000000000000004e00000000",
            INIT_60 => X"00000094000000000000009e00000000000000a900000000000000a600000000",
            INIT_61 => X"0000007100000000000000670000000000000085000000000000008f00000000",
            INIT_62 => X"0000003c000000000000004b0000000000000051000000000000004f00000000",
            INIT_63 => X"0000002c000000000000002a0000000000000027000000000000002a00000000",
            INIT_64 => X"0000004d00000000000000410000000000000036000000000000003000000000",
            INIT_65 => X"0000008b0000000000000083000000000000006e000000000000005a00000000",
            INIT_66 => X"000000360000000000000026000000000000001d000000000000003500000000",
            INIT_67 => X"000000c400000000000000a9000000000000005b000000000000004600000000",
            INIT_68 => X"0000008d0000000000000093000000000000009700000000000000a200000000",
            INIT_69 => X"0000004e000000000000006b0000000000000085000000000000008900000000",
            INIT_6A => X"0000003c0000000000000046000000000000004e000000000000004800000000",
            INIT_6B => X"00000030000000000000002e000000000000002a000000000000003200000000",
            INIT_6C => X"00000042000000000000003b0000000000000033000000000000003100000000",
            INIT_6D => X"0000007100000000000000650000000000000059000000000000004c00000000",
            INIT_6E => X"000000340000000000000023000000000000001d000000000000004500000000",
            INIT_6F => X"000000ba00000000000000ae0000000000000062000000000000003f00000000",
            INIT_70 => X"0000008c000000000000008e000000000000008d000000000000009400000000",
            INIT_71 => X"0000003c000000000000006a000000000000008c000000000000008f00000000",
            INIT_72 => X"000000370000000000000042000000000000004a000000000000004200000000",
            INIT_73 => X"0000003a00000000000000360000000000000034000000000000003900000000",
            INIT_74 => X"000000460000000000000041000000000000003a000000000000003a00000000",
            INIT_75 => X"0000005d00000000000000570000000000000050000000000000004900000000",
            INIT_76 => X"0000003700000000000000260000000000000025000000000000004d00000000",
            INIT_77 => X"000000b400000000000000b30000000000000083000000000000004a00000000",
            INIT_78 => X"000000a200000000000000a00000000000000095000000000000009000000000",
            INIT_79 => X"0000003d000000000000007e0000000000000092000000000000009e00000000",
            INIT_7A => X"00000043000000000000003a0000000000000039000000000000003900000000",
            INIT_7B => X"0000004800000000000000490000000000000045000000000000004600000000",
            INIT_7C => X"0000006200000000000000590000000000000049000000000000004400000000",
            INIT_7D => X"0000006100000000000000630000000000000061000000000000005e00000000",
            INIT_7E => X"0000004700000000000000400000000000000045000000000000005200000000",
            INIT_7F => X"000000ba00000000000000b600000000000000a4000000000000007700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE55;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE56 : if BRAM_NAME = "sampleifmap_layersamples_instance56" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ca00000000000000d000000000000000d000000000000000d700000000",
            INIT_01 => X"000000b900000000000000ca00000000000000d100000000000000d700000000",
            INIT_02 => X"000000a0000000000000009800000000000000a800000000000000b800000000",
            INIT_03 => X"0000009d000000000000009a00000000000000a7000000000000009d00000000",
            INIT_04 => X"000000e100000000000000e100000000000000cb00000000000000b500000000",
            INIT_05 => X"000000e400000000000000e500000000000000db00000000000000de00000000",
            INIT_06 => X"000000c400000000000000b800000000000000c500000000000000dd00000000",
            INIT_07 => X"000000a500000000000000b000000000000000b800000000000000d000000000",
            INIT_08 => X"000000d900000000000000e100000000000000e000000000000000e200000000",
            INIT_09 => X"000000ab00000000000000cc00000000000000dd00000000000000d500000000",
            INIT_0A => X"000000b100000000000000b200000000000000bd00000000000000b400000000",
            INIT_0B => X"000000e000000000000000d000000000000000cd00000000000000c400000000",
            INIT_0C => X"000000f300000000000000f200000000000000f000000000000000ec00000000",
            INIT_0D => X"000000e700000000000000e400000000000000e500000000000000ee00000000",
            INIT_0E => X"000000d200000000000000d400000000000000d600000000000000e700000000",
            INIT_0F => X"000000c500000000000000bf00000000000000be00000000000000de00000000",
            INIT_10 => X"000000eb00000000000000ea00000000000000ea00000000000000eb00000000",
            INIT_11 => X"000000a600000000000000d600000000000000ef00000000000000ea00000000",
            INIT_12 => X"000000b100000000000000a800000000000000b100000000000000a600000000",
            INIT_13 => X"000000df00000000000000ce00000000000000b700000000000000b800000000",
            INIT_14 => X"000000e800000000000000e300000000000000ec00000000000000dc00000000",
            INIT_15 => X"000000e000000000000000d900000000000000e400000000000000eb00000000",
            INIT_16 => X"000000dd00000000000000e600000000000000e900000000000000e900000000",
            INIT_17 => X"000000d200000000000000d100000000000000ce00000000000000d900000000",
            INIT_18 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_19 => X"0000009900000000000000e300000000000000f400000000000000f400000000",
            INIT_1A => X"0000009f0000000000000082000000000000009b000000000000009200000000",
            INIT_1B => X"000000a000000000000000a2000000000000008a000000000000009000000000",
            INIT_1C => X"000000dc00000000000000c200000000000000cd00000000000000ac00000000",
            INIT_1D => X"000000e000000000000000d300000000000000d300000000000000de00000000",
            INIT_1E => X"000000db00000000000000e500000000000000e900000000000000e600000000",
            INIT_1F => X"000000d400000000000000e200000000000000df00000000000000cf00000000",
            INIT_20 => X"000000f400000000000000f400000000000000f400000000000000f500000000",
            INIT_21 => X"0000007000000000000000cd00000000000000f000000000000000f500000000",
            INIT_22 => X"0000006d000000000000005b000000000000006d000000000000006200000000",
            INIT_23 => X"0000005c0000000000000064000000000000005c000000000000006500000000",
            INIT_24 => X"0000009a000000000000007c000000000000007d000000000000006800000000",
            INIT_25 => X"000000e300000000000000c900000000000000c200000000000000c200000000",
            INIT_26 => X"000000d300000000000000e300000000000000de00000000000000dc00000000",
            INIT_27 => X"000000e100000000000000e800000000000000dc00000000000000cb00000000",
            INIT_28 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_29 => X"0000007b00000000000000d400000000000000eb00000000000000f600000000",
            INIT_2A => X"00000069000000000000005f000000000000005d000000000000004700000000",
            INIT_2B => X"00000066000000000000006e000000000000006a000000000000006700000000",
            INIT_2C => X"0000005d000000000000005b0000000000000059000000000000005b00000000",
            INIT_2D => X"000000e600000000000000d900000000000000c5000000000000008100000000",
            INIT_2E => X"000000c600000000000000d600000000000000da00000000000000dd00000000",
            INIT_2F => X"000000ed00000000000000e200000000000000c500000000000000b400000000",
            INIT_30 => X"000000f400000000000000f300000000000000f300000000000000f500000000",
            INIT_31 => X"0000009c00000000000000d500000000000000d600000000000000f000000000",
            INIT_32 => X"0000009a00000000000000890000000000000077000000000000004f00000000",
            INIT_33 => X"00000096000000000000009b000000000000008b000000000000009000000000",
            INIT_34 => X"0000007e00000000000000790000000000000080000000000000008e00000000",
            INIT_35 => X"000000e900000000000000e100000000000000a0000000000000007200000000",
            INIT_36 => X"000000ba00000000000000c000000000000000da00000000000000e900000000",
            INIT_37 => X"000000ec00000000000000d400000000000000b000000000000000a500000000",
            INIT_38 => X"000000f700000000000000f300000000000000f300000000000000f400000000",
            INIT_39 => X"0000009600000000000000d300000000000000c100000000000000e200000000",
            INIT_3A => X"000000c800000000000000bc0000000000000098000000000000005100000000",
            INIT_3B => X"00000090000000000000008d00000000000000a500000000000000cd00000000",
            INIT_3C => X"0000008f000000000000008d0000000000000096000000000000008e00000000",
            INIT_3D => X"000000d600000000000000a3000000000000008c00000000000000a700000000",
            INIT_3E => X"000000d200000000000000d300000000000000d100000000000000e000000000",
            INIT_3F => X"000000dc00000000000000af00000000000000ae00000000000000c700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f500000000000000f400000000000000f300000000000000f400000000",
            INIT_41 => X"0000007f00000000000000d800000000000000ca00000000000000e100000000",
            INIT_42 => X"0000008700000000000000840000000000000086000000000000005100000000",
            INIT_43 => X"00000087000000000000007c000000000000009700000000000000b900000000",
            INIT_44 => X"0000008800000000000000960000000000000091000000000000008600000000",
            INIT_45 => X"000000c0000000000000008e000000000000009e00000000000000a400000000",
            INIT_46 => X"000000d700000000000000e700000000000000d800000000000000cf00000000",
            INIT_47 => X"000000c4000000000000009c000000000000009e00000000000000b100000000",
            INIT_48 => X"000000f200000000000000f400000000000000f200000000000000f200000000",
            INIT_49 => X"0000006e00000000000000a800000000000000bd00000000000000e300000000",
            INIT_4A => X"000000760000000000000080000000000000008c000000000000005300000000",
            INIT_4B => X"00000081000000000000007c0000000000000087000000000000009300000000",
            INIT_4C => X"000000860000000000000097000000000000008b000000000000008500000000",
            INIT_4D => X"000000c1000000000000009100000000000000a4000000000000009e00000000",
            INIT_4E => X"000000e600000000000000ef00000000000000ef00000000000000e500000000",
            INIT_4F => X"000000d700000000000000cc00000000000000be00000000000000c100000000",
            INIT_50 => X"000000f400000000000000f300000000000000ef00000000000000e800000000",
            INIT_51 => X"0000005e0000000000000080000000000000008100000000000000da00000000",
            INIT_52 => X"00000070000000000000007a000000000000007a000000000000004f00000000",
            INIT_53 => X"0000007300000000000000730000000000000070000000000000007100000000",
            INIT_54 => X"0000007e000000000000007f0000000000000080000000000000007c00000000",
            INIT_55 => X"000000aa0000000000000099000000000000009e000000000000009000000000",
            INIT_56 => X"000000f400000000000000f600000000000000e300000000000000ce00000000",
            INIT_57 => X"000000f400000000000000f500000000000000f300000000000000f300000000",
            INIT_58 => X"000000f200000000000000f200000000000000e300000000000000cd00000000",
            INIT_59 => X"00000058000000000000009f00000000000000a100000000000000d300000000",
            INIT_5A => X"00000066000000000000005e0000000000000045000000000000003c00000000",
            INIT_5B => X"0000006600000000000000670000000000000061000000000000006200000000",
            INIT_5C => X"00000067000000000000005f0000000000000064000000000000006800000000",
            INIT_5D => X"000000800000000000000089000000000000007f000000000000007100000000",
            INIT_5E => X"000000f300000000000000f800000000000000d7000000000000009900000000",
            INIT_5F => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_60 => X"000000dc00000000000000e400000000000000d500000000000000bc00000000",
            INIT_61 => X"0000006300000000000000ad00000000000000aa00000000000000b400000000",
            INIT_62 => X"00000066000000000000005a0000000000000039000000000000003700000000",
            INIT_63 => X"0000005500000000000000580000000000000067000000000000007200000000",
            INIT_64 => X"00000073000000000000005d0000000000000055000000000000005500000000",
            INIT_65 => X"0000008600000000000000760000000000000065000000000000007000000000",
            INIT_66 => X"000000f400000000000000f500000000000000e100000000000000b000000000",
            INIT_67 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_68 => X"000000b500000000000000ca00000000000000bc00000000000000b800000000",
            INIT_69 => X"00000063000000000000008d0000000000000086000000000000009800000000",
            INIT_6A => X"00000067000000000000006f0000000000000066000000000000006700000000",
            INIT_6B => X"0000005600000000000000600000000000000078000000000000007600000000",
            INIT_6C => X"00000092000000000000007d000000000000006b000000000000005c00000000",
            INIT_6D => X"0000007f000000000000006e000000000000006a000000000000008400000000",
            INIT_6E => X"000000d200000000000000c300000000000000b3000000000000009800000000",
            INIT_6F => X"000000f400000000000000f400000000000000f500000000000000ee00000000",
            INIT_70 => X"0000009800000000000000bd00000000000000c200000000000000b600000000",
            INIT_71 => X"0000007e000000000000007f000000000000007b000000000000009200000000",
            INIT_72 => X"0000005e0000000000000069000000000000005d000000000000007c00000000",
            INIT_73 => X"0000004f0000000000000055000000000000005d000000000000005a00000000",
            INIT_74 => X"0000005500000000000000540000000000000053000000000000004e00000000",
            INIT_75 => X"00000053000000000000004c000000000000004b000000000000005100000000",
            INIT_76 => X"0000008a000000000000008a000000000000007a000000000000006500000000",
            INIT_77 => X"000000f400000000000000f400000000000000f400000000000000bc00000000",
            INIT_78 => X"0000006500000000000000a700000000000000cc00000000000000bd00000000",
            INIT_79 => X"000000ae00000000000000a9000000000000007d000000000000006500000000",
            INIT_7A => X"00000036000000000000004f000000000000004d000000000000006700000000",
            INIT_7B => X"0000003e000000000000003b000000000000002f000000000000002b00000000",
            INIT_7C => X"000000340000000000000039000000000000003e000000000000003b00000000",
            INIT_7D => X"00000040000000000000003d0000000000000030000000000000002f00000000",
            INIT_7E => X"00000061000000000000005a000000000000004a000000000000004600000000",
            INIT_7F => X"000000f400000000000000f600000000000000df000000000000008000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE56;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE57 : if BRAM_NAME = "sampleifmap_layersamples_instance57" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000054000000000000009700000000000000a400000000000000ae00000000",
            INIT_01 => X"0000009200000000000000ac000000000000007c000000000000005200000000",
            INIT_02 => X"0000005a00000000000000570000000000000049000000000000005300000000",
            INIT_03 => X"00000044000000000000004c000000000000004b000000000000006400000000",
            INIT_04 => X"00000017000000000000001a0000000000000017000000000000002100000000",
            INIT_05 => X"000000190000000000000014000000000000002f000000000000003000000000",
            INIT_06 => X"0000006400000000000000560000000000000032000000000000001500000000",
            INIT_07 => X"000000f300000000000000f700000000000000ca000000000000007800000000",
            INIT_08 => X"0000006800000000000000b300000000000000b400000000000000c000000000",
            INIT_09 => X"00000040000000000000008e0000000000000087000000000000006800000000",
            INIT_0A => X"00000078000000000000006c0000000000000057000000000000004100000000",
            INIT_0B => X"00000062000000000000007d0000000000000076000000000000009500000000",
            INIT_0C => X"00000060000000000000006a0000000000000059000000000000004600000000",
            INIT_0D => X"0000006000000000000000590000000000000090000000000000009000000000",
            INIT_0E => X"0000008b00000000000000820000000000000067000000000000005a00000000",
            INIT_0F => X"000000f400000000000000f100000000000000b2000000000000009700000000",
            INIT_10 => X"0000005e00000000000000ab00000000000000bd00000000000000d100000000",
            INIT_11 => X"0000001c00000000000000760000000000000092000000000000006200000000",
            INIT_12 => X"0000004f0000000000000067000000000000005f000000000000003600000000",
            INIT_13 => X"0000005f00000000000000800000000000000064000000000000005300000000",
            INIT_14 => X"0000009e000000000000009b00000000000000aa000000000000009200000000",
            INIT_15 => X"000000a100000000000000a000000000000000a800000000000000ab00000000",
            INIT_16 => X"00000077000000000000009b00000000000000ac000000000000009e00000000",
            INIT_17 => X"000000f700000000000000e20000000000000080000000000000006f00000000",
            INIT_18 => X"0000005b00000000000000b000000000000000c100000000000000d000000000",
            INIT_19 => X"000000280000000000000064000000000000007f000000000000004c00000000",
            INIT_1A => X"0000003900000000000000490000000000000044000000000000003500000000",
            INIT_1B => X"00000059000000000000003d0000000000000035000000000000003200000000",
            INIT_1C => X"0000006200000000000000570000000000000077000000000000009c00000000",
            INIT_1D => X"0000006400000000000000630000000000000068000000000000007100000000",
            INIT_1E => X"0000003f000000000000007a0000000000000098000000000000006000000000",
            INIT_1F => X"000000f800000000000000d60000000000000070000000000000004d00000000",
            INIT_20 => X"0000005f00000000000000be00000000000000c300000000000000ca00000000",
            INIT_21 => X"000000380000000000000053000000000000004e000000000000003300000000",
            INIT_22 => X"00000044000000000000003c0000000000000027000000000000003300000000",
            INIT_23 => X"0000003d000000000000003b0000000000000033000000000000003900000000",
            INIT_24 => X"000000650000000000000066000000000000006e000000000000005f00000000",
            INIT_25 => X"00000060000000000000005c000000000000005f000000000000006300000000",
            INIT_26 => X"000000460000000000000060000000000000006c000000000000006400000000",
            INIT_27 => X"000000f900000000000000d0000000000000006c000000000000004f00000000",
            INIT_28 => X"0000006e00000000000000c000000000000000c000000000000000c200000000",
            INIT_29 => X"0000003f0000000000000049000000000000003e000000000000004c00000000",
            INIT_2A => X"000000300000000000000028000000000000001d000000000000002e00000000",
            INIT_2B => X"0000003b00000000000000530000000000000048000000000000004100000000",
            INIT_2C => X"00000043000000000000004d0000000000000043000000000000003000000000",
            INIT_2D => X"00000058000000000000003b0000000000000040000000000000003c00000000",
            INIT_2E => X"00000069000000000000004e0000000000000036000000000000005200000000",
            INIT_2F => X"000000f900000000000000c90000000000000065000000000000006b00000000",
            INIT_30 => X"0000006100000000000000bb00000000000000be00000000000000c300000000",
            INIT_31 => X"0000004300000000000000410000000000000063000000000000005500000000",
            INIT_32 => X"0000002000000000000000230000000000000026000000000000003a00000000",
            INIT_33 => X"0000004c000000000000008d0000000000000060000000000000004800000000",
            INIT_34 => X"00000071000000000000008c000000000000004f000000000000001900000000",
            INIT_35 => X"000000920000000000000061000000000000006d000000000000005e00000000",
            INIT_36 => X"0000008a0000000000000045000000000000003a00000000000000ab00000000",
            INIT_37 => X"000000f400000000000000c00000000000000053000000000000007400000000",
            INIT_38 => X"0000005200000000000000b000000000000000b700000000000000bd00000000",
            INIT_39 => X"0000005e00000000000000590000000000000063000000000000002c00000000",
            INIT_3A => X"0000002100000000000000240000000000000030000000000000005a00000000",
            INIT_3B => X"000000340000000000000055000000000000002f000000000000002600000000",
            INIT_3C => X"0000007b0000000000000091000000000000004a000000000000001c00000000",
            INIT_3D => X"0000009700000000000000710000000000000086000000000000007700000000",
            INIT_3E => X"0000004700000000000000320000000000000033000000000000009c00000000",
            INIT_3F => X"000000ee00000000000000c00000000000000047000000000000003b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004800000000000000a300000000000000ad00000000000000ae00000000",
            INIT_41 => X"0000008b00000000000000650000000000000036000000000000002200000000",
            INIT_42 => X"0000001e0000000000000028000000000000003a000000000000006600000000",
            INIT_43 => X"0000001e000000000000001a0000000000000019000000000000001a00000000",
            INIT_44 => X"0000005600000000000000350000000000000026000000000000002500000000",
            INIT_45 => X"0000007200000000000000760000000000000075000000000000006800000000",
            INIT_46 => X"0000002e0000000000000030000000000000002b000000000000003e00000000",
            INIT_47 => X"000000df00000000000000b8000000000000004b000000000000002f00000000",
            INIT_48 => X"00000078000000000000009e00000000000000a000000000000000a200000000",
            INIT_49 => X"0000008800000000000000670000000000000059000000000000005700000000",
            INIT_4A => X"0000002200000000000000340000000000000048000000000000005c00000000",
            INIT_4B => X"0000001d000000000000001b000000000000001b000000000000001c00000000",
            INIT_4C => X"000000af000000000000003d0000000000000015000000000000002000000000",
            INIT_4D => X"000000b400000000000000b100000000000000ca00000000000000cf00000000",
            INIT_4E => X"0000002c00000000000000280000000000000022000000000000005400000000",
            INIT_4F => X"000000d100000000000000ab0000000000000057000000000000003e00000000",
            INIT_50 => X"000000b000000000000000a8000000000000009c000000000000009c00000000",
            INIT_51 => X"0000008800000000000000660000000000000070000000000000009300000000",
            INIT_52 => X"0000002d000000000000004b0000000000000051000000000000005600000000",
            INIT_53 => X"0000001a00000000000000170000000000000016000000000000001600000000",
            INIT_54 => X"000000a400000000000000450000000000000022000000000000002300000000",
            INIT_55 => X"000000a500000000000000a900000000000000b100000000000000b900000000",
            INIT_56 => X"0000002d000000000000001a0000000000000019000000000000004e00000000",
            INIT_57 => X"000000cc00000000000000a7000000000000005c000000000000004b00000000",
            INIT_58 => X"000000a100000000000000ad00000000000000a7000000000000009500000000",
            INIT_59 => X"0000008e00000000000000630000000000000071000000000000008d00000000",
            INIT_5A => X"00000033000000000000004f0000000000000053000000000000005300000000",
            INIT_5B => X"00000022000000000000001f000000000000001c000000000000001d00000000",
            INIT_5C => X"0000006100000000000000510000000000000048000000000000003200000000",
            INIT_5D => X"00000085000000000000008a0000000000000074000000000000006600000000",
            INIT_5E => X"00000032000000000000001d000000000000001b000000000000003700000000",
            INIT_5F => X"000000c600000000000000a40000000000000059000000000000004c00000000",
            INIT_60 => X"00000090000000000000009b00000000000000a600000000000000a400000000",
            INIT_61 => X"0000006c00000000000000630000000000000082000000000000008b00000000",
            INIT_62 => X"0000003800000000000000480000000000000050000000000000004c00000000",
            INIT_63 => X"0000002900000000000000270000000000000024000000000000002600000000",
            INIT_64 => X"00000048000000000000003d0000000000000033000000000000002d00000000",
            INIT_65 => X"00000083000000000000007c0000000000000067000000000000005400000000",
            INIT_66 => X"000000320000000000000021000000000000001a000000000000003100000000",
            INIT_67 => X"000000c300000000000000a90000000000000059000000000000004500000000",
            INIT_68 => X"0000008d0000000000000092000000000000009400000000000000a000000000",
            INIT_69 => X"0000004900000000000000660000000000000082000000000000008700000000",
            INIT_6A => X"000000380000000000000042000000000000004d000000000000004500000000",
            INIT_6B => X"0000002d000000000000002b0000000000000028000000000000002f00000000",
            INIT_6C => X"0000003d00000000000000360000000000000030000000000000002e00000000",
            INIT_6D => X"0000006a000000000000005e0000000000000054000000000000004600000000",
            INIT_6E => X"00000030000000000000001f000000000000001a000000000000004000000000",
            INIT_6F => X"000000ba00000000000000af0000000000000062000000000000003d00000000",
            INIT_70 => X"0000008c000000000000008e000000000000008d000000000000009300000000",
            INIT_71 => X"000000390000000000000068000000000000008b000000000000008f00000000",
            INIT_72 => X"00000034000000000000003f000000000000004a000000000000004000000000",
            INIT_73 => X"0000003600000000000000330000000000000031000000000000003700000000",
            INIT_74 => X"00000042000000000000003d0000000000000036000000000000003600000000",
            INIT_75 => X"000000570000000000000051000000000000004a000000000000004400000000",
            INIT_76 => X"0000003400000000000000230000000000000021000000000000004800000000",
            INIT_77 => X"000000b500000000000000b60000000000000084000000000000004800000000",
            INIT_78 => X"000000a300000000000000a10000000000000096000000000000009200000000",
            INIT_79 => X"0000003a000000000000007c0000000000000091000000000000009d00000000",
            INIT_7A => X"0000004100000000000000390000000000000038000000000000003700000000",
            INIT_7B => X"0000004500000000000000460000000000000042000000000000004300000000",
            INIT_7C => X"0000005f00000000000000570000000000000048000000000000004300000000",
            INIT_7D => X"0000005e0000000000000060000000000000005f000000000000005c00000000",
            INIT_7E => X"00000046000000000000003e0000000000000044000000000000005100000000",
            INIT_7F => X"000000b900000000000000b600000000000000a3000000000000007600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE57;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE58 : if BRAM_NAME = "sampleifmap_layersamples_instance58" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b600000000000000bf00000000000000ca00000000000000d100000000",
            INIT_01 => X"000000af00000000000000c600000000000000d100000000000000d100000000",
            INIT_02 => X"000000a0000000000000009d00000000000000a500000000000000ab00000000",
            INIT_03 => X"0000008f000000000000008d000000000000009a000000000000009500000000",
            INIT_04 => X"000000db00000000000000d600000000000000bc00000000000000a400000000",
            INIT_05 => X"000000d600000000000000d900000000000000ca00000000000000d100000000",
            INIT_06 => X"000000ad00000000000000a100000000000000b100000000000000d000000000",
            INIT_07 => X"000000950000000000000095000000000000009d00000000000000b700000000",
            INIT_08 => X"000000cd00000000000000d200000000000000d400000000000000d400000000",
            INIT_09 => X"000000a300000000000000c800000000000000db00000000000000cf00000000",
            INIT_0A => X"000000b600000000000000b800000000000000b600000000000000a500000000",
            INIT_0B => X"000000d700000000000000cd00000000000000c900000000000000c200000000",
            INIT_0C => X"000000e400000000000000e300000000000000e300000000000000df00000000",
            INIT_0D => X"000000d700000000000000d300000000000000d400000000000000dd00000000",
            INIT_0E => X"000000bb00000000000000c300000000000000cd00000000000000df00000000",
            INIT_0F => X"000000ba00000000000000ad00000000000000aa00000000000000c600000000",
            INIT_10 => X"000000e200000000000000e300000000000000e500000000000000e600000000",
            INIT_11 => X"000000a400000000000000d300000000000000ec00000000000000e300000000",
            INIT_12 => X"000000b800000000000000b700000000000000ad000000000000009f00000000",
            INIT_13 => X"000000e000000000000000cf00000000000000bf00000000000000bc00000000",
            INIT_14 => X"000000d600000000000000e000000000000000e500000000000000db00000000",
            INIT_15 => X"000000d300000000000000c800000000000000d000000000000000d600000000",
            INIT_16 => X"000000c500000000000000db00000000000000e000000000000000de00000000",
            INIT_17 => X"000000c600000000000000c500000000000000bc00000000000000b900000000",
            INIT_18 => X"000000f100000000000000f400000000000000f400000000000000f500000000",
            INIT_19 => X"000000af00000000000000e300000000000000f100000000000000f200000000",
            INIT_1A => X"000000bb00000000000000a100000000000000b000000000000000a800000000",
            INIT_1B => X"000000b600000000000000b800000000000000a000000000000000ae00000000",
            INIT_1C => X"000000ca00000000000000d000000000000000d500000000000000b900000000",
            INIT_1D => X"000000d400000000000000c400000000000000ba00000000000000b900000000",
            INIT_1E => X"000000bb00000000000000d500000000000000dc00000000000000d700000000",
            INIT_1F => X"000000c800000000000000d400000000000000c500000000000000a900000000",
            INIT_20 => X"000000f400000000000000f400000000000000f300000000000000f500000000",
            INIT_21 => X"0000008400000000000000cd00000000000000f100000000000000f500000000",
            INIT_22 => X"000000a7000000000000008a00000000000000a1000000000000008b00000000",
            INIT_23 => X"0000008d000000000000009b000000000000008b000000000000009f00000000",
            INIT_24 => X"000000a4000000000000009900000000000000a6000000000000008e00000000",
            INIT_25 => X"000000e000000000000000c400000000000000a900000000000000a900000000",
            INIT_26 => X"000000b100000000000000d400000000000000d100000000000000d100000000",
            INIT_27 => X"000000d200000000000000cc00000000000000b800000000000000a000000000",
            INIT_28 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_29 => X"0000008100000000000000d700000000000000ee00000000000000f600000000",
            INIT_2A => X"000000aa00000000000000a0000000000000009c000000000000007100000000",
            INIT_2B => X"000000a700000000000000b100000000000000aa00000000000000aa00000000",
            INIT_2C => X"0000008f0000000000000098000000000000009d000000000000009d00000000",
            INIT_2D => X"000000e400000000000000cd00000000000000b3000000000000009400000000",
            INIT_2E => X"000000aa00000000000000c100000000000000ce00000000000000da00000000",
            INIT_2F => X"000000df00000000000000c000000000000000a0000000000000009300000000",
            INIT_30 => X"000000f400000000000000f300000000000000f300000000000000f500000000",
            INIT_31 => X"000000b400000000000000dd00000000000000dd00000000000000f100000000",
            INIT_32 => X"000000cf00000000000000c400000000000000b4000000000000008300000000",
            INIT_33 => X"000000d300000000000000d900000000000000cb00000000000000c800000000",
            INIT_34 => X"000000bf00000000000000c000000000000000c300000000000000cc00000000",
            INIT_35 => X"000000e100000000000000cd00000000000000a600000000000000a300000000",
            INIT_36 => X"000000a900000000000000b100000000000000d500000000000000e300000000",
            INIT_37 => X"000000da00000000000000b20000000000000092000000000000009100000000",
            INIT_38 => X"000000f700000000000000f200000000000000f200000000000000f400000000",
            INIT_39 => X"000000c000000000000000d900000000000000ca00000000000000e600000000",
            INIT_3A => X"000000e800000000000000e000000000000000c2000000000000008600000000",
            INIT_3B => X"000000d100000000000000ce00000000000000d700000000000000ea00000000",
            INIT_3C => X"000000cf00000000000000ca00000000000000d000000000000000cf00000000",
            INIT_3D => X"000000cc000000000000009a00000000000000b400000000000000e000000000",
            INIT_3E => X"000000bc00000000000000c400000000000000c900000000000000dc00000000",
            INIT_3F => X"000000c7000000000000009a000000000000009200000000000000ab00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f500000000000000f300000000000000f300000000000000f500000000",
            INIT_41 => X"000000ae00000000000000df00000000000000d100000000000000e300000000",
            INIT_42 => X"000000c100000000000000c100000000000000ba000000000000008700000000",
            INIT_43 => X"000000c900000000000000c100000000000000cc00000000000000dd00000000",
            INIT_44 => X"000000c600000000000000cd00000000000000cd00000000000000ca00000000",
            INIT_45 => X"000000bc00000000000000a300000000000000d000000000000000dc00000000",
            INIT_46 => X"000000cb00000000000000df00000000000000d100000000000000cb00000000",
            INIT_47 => X"000000b20000000000000094000000000000008b00000000000000a100000000",
            INIT_48 => X"000000f200000000000000f300000000000000f100000000000000f200000000",
            INIT_49 => X"000000a400000000000000c200000000000000cd00000000000000e500000000",
            INIT_4A => X"000000b800000000000000bd00000000000000c1000000000000008c00000000",
            INIT_4B => X"000000c400000000000000c000000000000000c400000000000000ca00000000",
            INIT_4C => X"000000c600000000000000d000000000000000ca00000000000000c700000000",
            INIT_4D => X"000000c800000000000000bc00000000000000e000000000000000d700000000",
            INIT_4E => X"000000e300000000000000ed00000000000000ee00000000000000e600000000",
            INIT_4F => X"000000d300000000000000ca00000000000000ba00000000000000bc00000000",
            INIT_50 => X"000000f400000000000000f300000000000000ee00000000000000ea00000000",
            INIT_51 => X"0000009c00000000000000a900000000000000a000000000000000df00000000",
            INIT_52 => X"000000ac00000000000000b300000000000000b1000000000000008600000000",
            INIT_53 => X"000000b700000000000000b400000000000000ae00000000000000ae00000000",
            INIT_54 => X"000000be00000000000000bc00000000000000be00000000000000bb00000000",
            INIT_55 => X"000000c400000000000000d000000000000000dc00000000000000cd00000000",
            INIT_56 => X"000000f400000000000000f600000000000000e600000000000000d900000000",
            INIT_57 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_58 => X"000000f200000000000000f200000000000000e600000000000000d300000000",
            INIT_59 => X"0000009700000000000000be00000000000000b600000000000000d800000000",
            INIT_5A => X"000000a00000000000000093000000000000006e000000000000006a00000000",
            INIT_5B => X"000000aa00000000000000a6000000000000009f000000000000009e00000000",
            INIT_5C => X"000000a6000000000000009e00000000000000a300000000000000a900000000",
            INIT_5D => X"000000af00000000000000c600000000000000bd00000000000000ad00000000",
            INIT_5E => X"000000f300000000000000f800000000000000e000000000000000b700000000",
            INIT_5F => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_60 => X"000000e100000000000000e900000000000000da00000000000000c400000000",
            INIT_61 => X"0000009f00000000000000c300000000000000b400000000000000bd00000000",
            INIT_62 => X"000000a0000000000000008d000000000000005c000000000000005d00000000",
            INIT_63 => X"0000008c000000000000008f00000000000000a800000000000000ba00000000",
            INIT_64 => X"000000a700000000000000920000000000000089000000000000008b00000000",
            INIT_65 => X"00000096000000000000008f0000000000000083000000000000009800000000",
            INIT_66 => X"000000f400000000000000f300000000000000e300000000000000bc00000000",
            INIT_67 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_68 => X"000000c100000000000000d300000000000000c700000000000000c300000000",
            INIT_69 => X"0000008900000000000000a2000000000000009500000000000000a400000000",
            INIT_6A => X"000000a600000000000000b200000000000000aa000000000000009600000000",
            INIT_6B => X"0000009200000000000000a600000000000000cd00000000000000bd00000000",
            INIT_6C => X"000000d300000000000000c000000000000000ac000000000000009900000000",
            INIT_6D => X"0000008a0000000000000080000000000000008000000000000000af00000000",
            INIT_6E => X"000000d300000000000000bf00000000000000b100000000000000a000000000",
            INIT_6F => X"000000f300000000000000f300000000000000f500000000000000ef00000000",
            INIT_70 => X"000000a200000000000000c800000000000000cf00000000000000c200000000",
            INIT_71 => X"00000089000000000000008e0000000000000088000000000000009c00000000",
            INIT_72 => X"0000009f00000000000000b100000000000000b200000000000000a200000000",
            INIT_73 => X"0000008b000000000000009500000000000000a3000000000000009600000000",
            INIT_74 => X"0000009300000000000000920000000000000092000000000000008d00000000",
            INIT_75 => X"00000085000000000000007f000000000000007c000000000000008600000000",
            INIT_76 => X"000000a600000000000000ad00000000000000a3000000000000009500000000",
            INIT_77 => X"000000f400000000000000f300000000000000f500000000000000cc00000000",
            INIT_78 => X"0000006e00000000000000ad00000000000000d000000000000000c300000000",
            INIT_79 => X"000000b900000000000000b4000000000000008b000000000000007100000000",
            INIT_7A => X"00000057000000000000007f000000000000009a000000000000008500000000",
            INIT_7B => X"0000005f0000000000000059000000000000004c000000000000004900000000",
            INIT_7C => X"00000058000000000000005e0000000000000060000000000000005c00000000",
            INIT_7D => X"0000006700000000000000630000000000000056000000000000005600000000",
            INIT_7E => X"0000009b000000000000008f0000000000000074000000000000006d00000000",
            INIT_7F => X"000000f500000000000000f500000000000000e800000000000000af00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE58;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE59 : if BRAM_NAME = "sampleifmap_layersamples_instance59" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000006500000000000000a100000000000000aa00000000000000b700000000",
            INIT_01 => X"000000a100000000000000b50000000000000088000000000000006000000000",
            INIT_02 => X"0000008700000000000000810000000000000084000000000000008000000000",
            INIT_03 => X"0000006a000000000000007d000000000000007d000000000000008c00000000",
            INIT_04 => X"00000027000000000000002c000000000000002b000000000000003500000000",
            INIT_05 => X"0000002800000000000000230000000000000047000000000000004d00000000",
            INIT_06 => X"0000009700000000000000910000000000000050000000000000002000000000",
            INIT_07 => X"000000f300000000000000f600000000000000db00000000000000a700000000",
            INIT_08 => X"0000007c00000000000000c200000000000000c100000000000000ca00000000",
            INIT_09 => X"0000004900000000000000990000000000000092000000000000007800000000",
            INIT_0A => X"0000009400000000000000830000000000000087000000000000006900000000",
            INIT_0B => X"0000008300000000000000a9000000000000009f00000000000000b800000000",
            INIT_0C => X"0000007a00000000000000840000000000000076000000000000006600000000",
            INIT_0D => X"00000073000000000000006f00000000000000aa00000000000000af00000000",
            INIT_0E => X"000000b500000000000000b20000000000000091000000000000006f00000000",
            INIT_0F => X"000000f400000000000000f200000000000000c500000000000000bb00000000",
            INIT_10 => X"0000007200000000000000b800000000000000c800000000000000d800000000",
            INIT_11 => X"000000240000000000000082000000000000009d000000000000007300000000",
            INIT_12 => X"0000006300000000000000810000000000000095000000000000004f00000000",
            INIT_13 => X"00000084000000000000009d0000000000000081000000000000006f00000000",
            INIT_14 => X"000000b900000000000000b700000000000000c100000000000000b100000000",
            INIT_15 => X"000000bd00000000000000ba00000000000000c100000000000000c800000000",
            INIT_16 => X"0000009700000000000000b600000000000000c700000000000000b500000000",
            INIT_17 => X"000000f600000000000000e800000000000000a2000000000000009400000000",
            INIT_18 => X"0000007100000000000000bb00000000000000cc00000000000000d900000000",
            INIT_19 => X"0000003d0000000000000071000000000000008b000000000000006000000000",
            INIT_1A => X"0000005d00000000000000730000000000000070000000000000004e00000000",
            INIT_1B => X"0000007d000000000000005e0000000000000053000000000000005500000000",
            INIT_1C => X"0000008a000000000000007f000000000000009f00000000000000bf00000000",
            INIT_1D => X"0000008f000000000000008c000000000000009500000000000000a000000000",
            INIT_1E => X"00000063000000000000009f00000000000000bd000000000000008a00000000",
            INIT_1F => X"000000f700000000000000e2000000000000009a000000000000007300000000",
            INIT_20 => X"0000007500000000000000c700000000000000d000000000000000d500000000",
            INIT_21 => X"000000540000000000000063000000000000005c000000000000004900000000",
            INIT_22 => X"0000006900000000000000610000000000000041000000000000004b00000000",
            INIT_23 => X"0000005f00000000000000670000000000000057000000000000005f00000000",
            INIT_24 => X"00000097000000000000009900000000000000a2000000000000008600000000",
            INIT_25 => X"0000008f00000000000000890000000000000090000000000000009600000000",
            INIT_26 => X"0000006f000000000000008f0000000000000099000000000000009300000000",
            INIT_27 => X"000000f700000000000000de0000000000000092000000000000007300000000",
            INIT_28 => X"0000008300000000000000cc00000000000000ce00000000000000cc00000000",
            INIT_29 => X"0000005a000000000000005c0000000000000051000000000000006500000000",
            INIT_2A => X"000000450000000000000039000000000000002d000000000000004600000000",
            INIT_2B => X"00000057000000000000007d000000000000006f000000000000006200000000",
            INIT_2C => X"0000006700000000000000700000000000000066000000000000004a00000000",
            INIT_2D => X"0000007d000000000000005e0000000000000065000000000000006200000000",
            INIT_2E => X"0000009500000000000000710000000000000052000000000000007300000000",
            INIT_2F => X"000000f800000000000000d40000000000000089000000000000009a00000000",
            INIT_30 => X"0000007500000000000000ce00000000000000d000000000000000d100000000",
            INIT_31 => X"0000005e0000000000000056000000000000007a000000000000006900000000",
            INIT_32 => X"0000002f00000000000000330000000000000036000000000000005600000000",
            INIT_33 => X"0000006300000000000000ad0000000000000083000000000000006600000000",
            INIT_34 => X"00000082000000000000009e0000000000000064000000000000002d00000000",
            INIT_35 => X"000000ab000000000000007c000000000000008a000000000000007900000000",
            INIT_36 => X"000000ab000000000000005f000000000000004b00000000000000bb00000000",
            INIT_37 => X"000000fa00000000000000cf0000000000000075000000000000009800000000",
            INIT_38 => X"0000006800000000000000cc00000000000000d600000000000000dd00000000",
            INIT_39 => X"0000008000000000000000720000000000000074000000000000003b00000000",
            INIT_3A => X"0000003000000000000000340000000000000041000000000000007c00000000",
            INIT_3B => X"0000004b000000000000006c0000000000000046000000000000003800000000",
            INIT_3C => X"0000008f00000000000000a6000000000000005f000000000000003000000000",
            INIT_3D => X"000000af000000000000008f00000000000000a7000000000000009100000000",
            INIT_3E => X"000000620000000000000048000000000000004a00000000000000af00000000",
            INIT_3F => X"000000fb00000000000000d60000000000000068000000000000005400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006300000000000000c900000000000000d400000000000000d700000000",
            INIT_41 => X"000000b000000000000000800000000000000044000000000000002f00000000",
            INIT_42 => X"0000002d00000000000000380000000000000050000000000000008700000000",
            INIT_43 => X"0000002f000000000000002b0000000000000027000000000000002800000000",
            INIT_44 => X"0000006e0000000000000050000000000000003c000000000000003700000000",
            INIT_45 => X"0000008b00000000000000900000000000000093000000000000007d00000000",
            INIT_46 => X"0000004300000000000000460000000000000043000000000000005c00000000",
            INIT_47 => X"000000fb00000000000000d9000000000000006d000000000000004500000000",
            INIT_48 => X"0000009d00000000000000cb00000000000000cf00000000000000cf00000000",
            INIT_49 => X"000000aa00000000000000850000000000000075000000000000007300000000",
            INIT_4A => X"0000003000000000000000480000000000000065000000000000007e00000000",
            INIT_4B => X"0000002d00000000000000290000000000000029000000000000002800000000",
            INIT_4C => X"000000c000000000000000530000000000000027000000000000003200000000",
            INIT_4D => X"000000c900000000000000c700000000000000dc00000000000000da00000000",
            INIT_4E => X"0000003f00000000000000380000000000000034000000000000006b00000000",
            INIT_4F => X"000000f700000000000000d2000000000000007e000000000000005a00000000",
            INIT_50 => X"000000d800000000000000ce00000000000000c000000000000000bc00000000",
            INIT_51 => X"000000a10000000000000086000000000000009a00000000000000bf00000000",
            INIT_52 => X"0000003e00000000000000680000000000000073000000000000007900000000",
            INIT_53 => X"0000002900000000000000230000000000000022000000000000002100000000",
            INIT_54 => X"000000b300000000000000550000000000000031000000000000003300000000",
            INIT_55 => X"000000bb00000000000000be00000000000000c000000000000000c700000000",
            INIT_56 => X"0000004200000000000000260000000000000027000000000000006000000000",
            INIT_57 => X"000000f500000000000000d10000000000000085000000000000006f00000000",
            INIT_58 => X"000000c600000000000000cd00000000000000c600000000000000bf00000000",
            INIT_59 => X"000000a00000000000000084000000000000009e00000000000000b500000000",
            INIT_5A => X"00000046000000000000006f0000000000000076000000000000007200000000",
            INIT_5B => X"00000031000000000000002c0000000000000026000000000000002700000000",
            INIT_5C => X"0000007e0000000000000069000000000000005d000000000000004400000000",
            INIT_5D => X"000000a600000000000000ad0000000000000096000000000000008700000000",
            INIT_5E => X"00000047000000000000002a0000000000000028000000000000004800000000",
            INIT_5F => X"000000f200000000000000cf0000000000000082000000000000007100000000",
            INIT_60 => X"000000b800000000000000c600000000000000d100000000000000ce00000000",
            INIT_61 => X"00000085000000000000008200000000000000a300000000000000ab00000000",
            INIT_62 => X"0000004d0000000000000068000000000000006f000000000000006b00000000",
            INIT_63 => X"000000390000000000000035000000000000002f000000000000003200000000",
            INIT_64 => X"0000006800000000000000570000000000000048000000000000003f00000000",
            INIT_65 => X"000000b000000000000000a80000000000000091000000000000007800000000",
            INIT_66 => X"0000004700000000000000300000000000000028000000000000004500000000",
            INIT_67 => X"000000ee00000000000000d4000000000000007e000000000000006600000000",
            INIT_68 => X"000000bd00000000000000c200000000000000c200000000000000c700000000",
            INIT_69 => X"00000065000000000000008600000000000000a600000000000000b200000000",
            INIT_6A => X"0000004f00000000000000600000000000000069000000000000006300000000",
            INIT_6B => X"0000003e000000000000003b0000000000000036000000000000003e00000000",
            INIT_6C => X"00000057000000000000004e0000000000000045000000000000004100000000",
            INIT_6D => X"0000008f00000000000000810000000000000074000000000000006400000000",
            INIT_6E => X"00000047000000000000002c0000000000000027000000000000005700000000",
            INIT_6F => X"000000e800000000000000df0000000000000085000000000000005900000000",
            INIT_70 => X"000000bc00000000000000be00000000000000bc00000000000000c100000000",
            INIT_71 => X"00000050000000000000009000000000000000bc00000000000000bd00000000",
            INIT_72 => X"0000004600000000000000580000000000000063000000000000005a00000000",
            INIT_73 => X"0000004e000000000000004a0000000000000045000000000000004900000000",
            INIT_74 => X"0000005d0000000000000056000000000000004e000000000000004e00000000",
            INIT_75 => X"00000072000000000000006d0000000000000066000000000000006100000000",
            INIT_76 => X"0000004a00000000000000300000000000000030000000000000005e00000000",
            INIT_77 => X"000000e700000000000000e800000000000000ad000000000000006400000000",
            INIT_78 => X"000000cd00000000000000d000000000000000c700000000000000c400000000",
            INIT_79 => X"0000005500000000000000a500000000000000bb00000000000000c800000000",
            INIT_7A => X"00000054000000000000004e000000000000004c000000000000004c00000000",
            INIT_7B => X"0000006300000000000000620000000000000059000000000000005400000000",
            INIT_7C => X"0000007c00000000000000720000000000000063000000000000005e00000000",
            INIT_7D => X"0000007f00000000000000800000000000000081000000000000007d00000000",
            INIT_7E => X"000000600000000000000054000000000000005b000000000000007000000000",
            INIT_7F => X"000000df00000000000000e100000000000000cc000000000000009400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE59;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE0 : if BRAM_NAME = "samplegold_layersamples_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000021000000000000001f000000000000002f000000000000001800000000",
            INIT_01 => X"0000002c00000000000000240000000000000028000000000000001900000000",
            INIT_02 => X"0000001900000000000000080000000000000000000000000000001b00000000",
            INIT_03 => X"0000001c0000000000000027000000000000002a000000000000002800000000",
            INIT_04 => X"000000190000000000000021000000000000001d000000000000003b00000000",
            INIT_05 => X"0000001300000000000000100000000000000013000000000000001b00000000",
            INIT_06 => X"0000000b00000000000000080000000000000000000000000000000f00000000",
            INIT_07 => X"000000000000000000000000000000000000001b000000000000001000000000",
            INIT_08 => X"000000220000000000000014000000000000002b000000000000002100000000",
            INIT_09 => X"000000000000000000000009000000000000002c000000000000003400000000",
            INIT_0A => X"0000000000000000000000030000000000000012000000000000000700000000",
            INIT_0B => X"0000001b00000000000000000000000000000030000000000000002000000000",
            INIT_0C => X"0000000c000000000000000f0000000000000012000000000000001d00000000",
            INIT_0D => X"0000003200000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000100000000000000030000000000000000e00000000",
            INIT_0F => X"0000000000000000000000120000000000000000000000000000002000000000",
            INIT_10 => X"0000002a00000000000000370000000000000000000000000000000000000000",
            INIT_11 => X"0000001c000000000000001b0000000000000000000000000000001d00000000",
            INIT_12 => X"0000000000000000000000000000000000000021000000000000000e00000000",
            INIT_13 => X"0000002f000000000000000f0000000000000032000000000000000000000000",
            INIT_14 => X"00000034000000000000002b0000000000000041000000000000003000000000",
            INIT_15 => X"0000000000000000000000350000000000000005000000000000000000000000",
            INIT_16 => X"00000002000000000000000b0000000000000015000000000000001200000000",
            INIT_17 => X"000000000000000000000000000000000000005c000000000000001900000000",
            INIT_18 => X"0000000000000000000000380000000000000019000000000000000000000000",
            INIT_19 => X"0000000400000000000000080000000000000025000000000000002f00000000",
            INIT_1A => X"0000000000000000000000320000000000000000000000000000000f00000000",
            INIT_1B => X"0000001900000000000000000000000000000000000000000000002000000000",
            INIT_1C => X"000000260000000000000000000000000000003b000000000000001400000000",
            INIT_1D => X"0000003d00000000000000040000000000000000000000000000003700000000",
            INIT_1E => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_1F => X"0000000f00000000000000420000000000000028000000000000000000000000",
            INIT_20 => X"0000004200000000000000110000000000000019000000000000000000000000",
            INIT_21 => X"0000000c00000000000000020000000000000027000000000000001900000000",
            INIT_22 => X"0000000c0000000000000000000000000000003b000000000000000000000000",
            INIT_23 => X"0000000000000000000000190000000000000006000000000000000000000000",
            INIT_24 => X"00000000000000000000001e0000000000000023000000000000000300000000",
            INIT_25 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_26 => X"0000000000000000000000020000000000000000000000000000004000000000",
            INIT_27 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"00000008000000000000002b0000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_3F => X"0000001e00000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000100000000000000000000000000000000000000000000001300000000",
            INIT_41 => X"00000000000000000000000a000000000000000e00000000000000b700000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000022000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000023000000000000000000000000",
            INIT_4A => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000008700000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"000000000000000000000000000000000000001500000000000000a700000000",
            INIT_4D => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000004e00000000000000000000000000000000000000000000000b00000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"000000480000000000000000000000000000005a000000000000005f00000000",
            INIT_55 => X"0000002300000000000000000000000000000002000000000000000300000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_57 => X"0000000000000000000000990000000000000000000000000000000000000000",
            INIT_58 => X"0000003e00000000000000240000000000000000000000000000000000000000",
            INIT_59 => X"000000000000000000000000000000000000003a000000000000006d00000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"000000000000000000000047000000000000003f000000000000000c00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000860000000000000000000000000000000000000000",
            INIT_62 => X"0000007500000000000000bf0000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000050000000000000006300000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000740000000000000000000000000000000000000000",
            INIT_66 => X"000000000000000000000000000000000000005c000000000000002e00000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000005f00000000000000590000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000590000000000000000000000000000000000000000",
            INIT_6D => X"0000001a000000000000006e000000000000000d000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000013000000000000002100000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"00000020000000000000002e0000000000000000000000000000000000000000",
            INIT_71 => X"0000002700000000000000250000000000000023000000000000003600000000",
            INIT_72 => X"0000000d0000000000000025000000000000002d000000000000002800000000",
            INIT_73 => X"0000001700000000000000240000000000000028000000000000001100000000",
            INIT_74 => X"0000003a00000000000000240000000000000028000000000000001300000000",
            INIT_75 => X"0000000000000000000000000000000000000042000000000000001c00000000",
            INIT_76 => X"0000000000000000000000150000000000000001000000000000000000000000",
            INIT_77 => X"0000000c0000000000000025000000000000000d000000000000000000000000",
            INIT_78 => X"00000022000000000000002b0000000000000063000000000000000000000000",
            INIT_79 => X"000000000000000000000000000000000000000b000000000000003b00000000",
            INIT_7A => X"000000000000000000000000000000000000003d000000000000002100000000",
            INIT_7B => X"00000000000000000000001b0000000000000021000000000000000000000000",
            INIT_7C => X"0000000000000000000000360000000000000004000000000000006200000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000004800000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000009700000000",
            INIT_7F => X"000000000000000000000000000000000000006f000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE0;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE1 : if BRAM_NAME = "samplegold_layersamples_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001e000000000000000000000000000000f0000000000000000000000000",
            INIT_01 => X"000000e800000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000005100000000",
            INIT_04 => X"0000000000000000000000540000000000000044000000000000007000000000",
            INIT_05 => X"00000000000000000000012e0000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_07 => X"0000000000000000000000060000000000000000000000000000002b00000000",
            INIT_08 => X"0000000000000000000000000000000000000063000000000000005b00000000",
            INIT_09 => X"00000000000000000000000000000000000000bd000000000000000000000000",
            INIT_0A => X"0000001100000000000000000000000000000002000000000000000000000000",
            INIT_0B => X"0000008000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_0D => X"0000002800000000000000000000000000000000000000000000008700000000",
            INIT_0E => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_0F => X"0000003800000000000000070000000000000000000000000000000000000000",
            INIT_10 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_11 => X"0000001e000000000000002f0000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_13 => X"0000006d000000000000006a0000000000000000000000000000003d00000000",
            INIT_14 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_15 => X"00000004000000000000002d000000000000001a000000000000000000000000",
            INIT_16 => X"000000fb00000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"00000000000000000000003f0000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000002000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"00000000000000000000005d0000000000000000000000000000002a00000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000003f00000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"000000000000000000000000000000000000000000000000000000d800000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"000000fa00000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000100000000000000000000000000000000000000000000000700000000",
            INIT_29 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000700000000000000040000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000060000000000000001000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000003700000000000000000000000000000000000000000000000500000000",
            INIT_2F => X"0000000000000000000000560000000000000053000000000000001c00000000",
            INIT_30 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000003500000000000000500000000000000005000000000000000500000000",
            INIT_32 => X"000000000000000000000000000000000000002500000000000000a700000000",
            INIT_33 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_34 => X"00000008000000000000000c0000000000000052000000000000000f00000000",
            INIT_35 => X"000000000000000000000000000000000000003e000000000000000300000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000120000000000000000000000000000000800000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000023000000000000004100000000",
            INIT_3B => X"000000000000000000000000000000000000002a000000000000000000000000",
            INIT_3C => X"00000000000000000000004b0000000000000001000000000000000000000000",
            INIT_3D => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_3F => X"0000003900000000000000000000000000000015000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_41 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000020000000000000032000000000000002300000000",
            INIT_43 => X"0000001000000000000000190000000000000006000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000004a00000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"00000000000000000000001d0000000000000071000000000000006300000000",
            INIT_49 => X"000000310000000000000003000000000000003b000000000000008200000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_4B => X"0000000000000000000000000000000000000055000000000000000000000000",
            INIT_4C => X"0000000000000000000000170000000000000000000000000000003400000000",
            INIT_4D => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_4E => X"0000001f00000000000000050000000000000009000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_50 => X"00000034000000000000001d0000000000000000000000000000000000000000",
            INIT_51 => X"0000003300000000000000320000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_53 => X"000000aa00000000000000b1000000000000009c000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000003600000000",
            INIT_55 => X"0000000000000000000000000000000000000009000000000000000700000000",
            INIT_56 => X"0000006200000000000000000000000000000017000000000000002e00000000",
            INIT_57 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_5A => X"0000000200000000000000000000000000000000000000000000000b00000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_5D => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"000000000000000000000007000000000000001e000000000000009c00000000",
            INIT_5F => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000330000000000000023000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"000000a000000000000000060000000000000011000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"00000000000000000000004a0000000000000000000000000000000000000000",
            INIT_69 => X"0000007800000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"000000000000000000000000000000000000000a000000000000000900000000",
            INIT_6B => X"0000000000000000000000500000000000000000000000000000000c00000000",
            INIT_6C => X"0000000000000000000000000000000000000080000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000001900000000000000000000000000000002000000000000001400000000",
            INIT_6F => X"000000000000000000000000000000000000000d000000000000002600000000",
            INIT_70 => X"00000000000000000000001d0000000000000000000000000000004f00000000",
            INIT_71 => X"0000000000000000000000320000000000000015000000000000000000000000",
            INIT_72 => X"0000003400000000000000000000000000000000000000000000002a00000000",
            INIT_73 => X"0000004300000000000000000000000000000019000000000000000000000000",
            INIT_74 => X"0000000000000000000000190000000000000000000000000000000000000000",
            INIT_75 => X"0000002c000000000000000a0000000000000000000000000000000000000000",
            INIT_76 => X"00000000000000000000003d0000000000000062000000000000000000000000",
            INIT_77 => X"0000004b00000000000000000000000000000000000000000000000f00000000",
            INIT_78 => X"0000000000000000000000000000000000000039000000000000000000000000",
            INIT_79 => X"0000000000000000000000680000000000000000000000000000005e00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000005200000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"000000bd00000000000000000000000000000009000000000000000000000000",
            INIT_7D => X"0000000b00000000000000000000000000000000000000000000002e00000000",
            INIT_7E => X"0000000000000000000000120000000000000000000000000000000d00000000",
            INIT_7F => X"0000000000000000000000230000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE1;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE2 : if BRAM_NAME = "samplegold_layersamples_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000056000000000000000000000000",
            INIT_01 => X"0000008100000000000000000000000000000064000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000002900000000000000000000000000000044000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"00000000000000000000001400000000000000bd000000000000004500000000",
            INIT_06 => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000007000000000",
            INIT_08 => X"00000038000000000000008b0000000000000088000000000000000e00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000100000000000000000000000000000035000000000000000f00000000",
            INIT_0B => X"0000000000000000000000200000000000000178000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000005900000000000000000000000000000000000000000000001700000000",
            INIT_0F => X"0000000000000000000000120000000000000000000000000000009c00000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000f00000000000000000000000000000012000000000000001900000000",
            INIT_12 => X"0000000f00000000000000c70000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000020000000000000003000000000000000000000000",
            INIT_15 => X"00000000000000000000002a0000000000000098000000000000000000000000",
            INIT_16 => X"00000000000000000000002b0000000000000055000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_18 => X"0000000a00000000000000000000000000000000000000000000000900000000",
            INIT_19 => X"0000004f00000000000000560000000000000042000000000000005200000000",
            INIT_1A => X"0000005400000000000000450000000000000058000000000000005800000000",
            INIT_1B => X"0000003e0000000000000047000000000000005f000000000000005c00000000",
            INIT_1C => X"0000005a00000000000000510000000000000049000000000000003700000000",
            INIT_1D => X"0000005e00000000000000450000000000000050000000000000005700000000",
            INIT_1E => X"0000006800000000000000640000000000000097000000000000003c00000000",
            INIT_1F => X"000000320000000000000045000000000000001e000000000000004000000000",
            INIT_20 => X"0000007e00000000000000570000000000000023000000000000001400000000",
            INIT_21 => X"0000004800000000000000610000000000000056000000000000000000000000",
            INIT_22 => X"000000000000000000000017000000000000008d000000000000000000000000",
            INIT_23 => X"00000053000000000000001c000000000000001d000000000000000000000000",
            INIT_24 => X"0000000000000000000000b50000000000000031000000000000000000000000",
            INIT_25 => X"0000000500000000000000960000000000000047000000000000004b00000000",
            INIT_26 => X"0000000000000000000000280000000000000027000000000000004e00000000",
            INIT_27 => X"00000045000000000000004d0000000000000000000000000000008500000000",
            INIT_28 => X"0000007000000000000000000000000000000066000000000000000000000000",
            INIT_29 => X"0000005f000000000000000a0000000000000069000000000000000000000000",
            INIT_2A => X"0000001600000000000000000000000000000047000000000000006b00000000",
            INIT_2B => X"000000000000000000000063000000000000001e000000000000006400000000",
            INIT_2C => X"00000043000000000000008c000000000000000c000000000000000000000000",
            INIT_2D => X"0000003200000000000000a50000000000000000000000000000000000000000",
            INIT_2E => X"00000065000000000000006a000000000000000000000000000000a600000000",
            INIT_2F => X"00000000000000000000003d000000000000002e000000000000000000000000",
            INIT_30 => X"0000000000000000000000b80000000000000016000000000000007900000000",
            INIT_31 => X"000000720000000000000064000000000000001f000000000000000000000000",
            INIT_32 => X"000000010000000000000056000000000000006d000000000000000000000000",
            INIT_33 => X"000000400000000000000017000000000000003b000000000000000000000000",
            INIT_34 => X"000000000000000000000000000000000000006e000000000000000000000000",
            INIT_35 => X"0000000000000000000000530000000000000010000000000000008300000000",
            INIT_36 => X"0000000000000000000000000000000000000058000000000000006300000000",
            INIT_37 => X"000000a10000000000000000000000000000003b000000000000003200000000",
            INIT_38 => X"0000002700000000000000000000000000000049000000000000000000000000",
            INIT_39 => X"0000000000000000000000430000000000000000000000000000004d00000000",
            INIT_3A => X"0000003000000000000000030000000000000000000000000000006700000000",
            INIT_3B => X"0000000000000000000000c40000000000000000000000000000001a00000000",
            INIT_3C => X"0000005200000000000000000000000000000000000000000000002400000000",
            INIT_3D => X"000000000000000000000065000000000000001a000000000000000300000000",
            INIT_3E => X"00000000000000000000004f000000000000000d000000000000000000000000",
            INIT_3F => X"000000f800000000000000000000000000000098000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006e00000000000000090000000000000000000000000000001000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_42 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_43 => X"0000002500000000000000850000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"000000000000000000000000000000000000006d000000000000003e00000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"000000b800000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000040000000000000033000000000000003d00000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"000000000000000000000000000000000000005f000000000000000000000000",
            INIT_58 => X"0000000000000000000000340000000000000000000000000000000000000000",
            INIT_59 => X"00000000000000000000000000000000000000a8000000000000001000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"00000000000000000000001d0000000000000017000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000005b00000000",
            INIT_60 => X"000000000000000000000000000000000000004c000000000000000000000000",
            INIT_61 => X"000000000000000000000000000000000000004d000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"000000000000000000000054000000000000005a000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_68 => X"00000000000000000000004a0000000000000000000000000000000000000000",
            INIT_69 => X"00000000000000000000002d0000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"000000070000000000000016000000000000002b000000000000008000000000",
            INIT_6E => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_70 => X"0000002600000000000000000000000000000022000000000000000000000000",
            INIT_71 => X"0000000000000000000000280000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000029000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"000000000000000000000010000000000000001b000000000000000000000000",
            INIT_75 => X"0000005500000000000000a10000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000030000000000000002600000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_78 => X"000000b5000000000000006b0000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000008b00000000",
            INIT_7A => X"0000008500000000000000130000000000000017000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000043000000000000008700000000",
            INIT_7C => X"0000000300000000000000000000000000000000000000000000001e00000000",
            INIT_7D => X"0000000000000000000000000000000000000001000000000000000300000000",
            INIT_7E => X"0000003500000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000330000000000000000000000000000006500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE2;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE3 : if BRAM_NAME = "samplegold_layersamples_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000001a00000000000000040000000000000000000000000000000000000000",
            INIT_02 => X"0000007200000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"000000000000000000000000000000000000001d000000000000004f00000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"000000170000000000000048000000000000000b000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000002300000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000024000000000000001400000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000003100000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"00000000000000000000001e0000000000000000000000000000001600000000",
            INIT_18 => X"0000003c0000000000000000000000000000000f000000000000001a00000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_1A => X"000000230000000000000017000000000000000d000000000000000000000000",
            INIT_1B => X"0000001000000000000000130000000000000005000000000000000000000000",
            INIT_1C => X"0000002c00000000000000180000000000000000000000000000002700000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"00000000000000000000004d0000000000000000000000000000002f00000000",
            INIT_1F => X"000000190000000000000000000000000000000e000000000000001900000000",
            INIT_20 => X"00000000000000000000007a0000000000000007000000000000001400000000",
            INIT_21 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"000000260000000000000000000000000000002e000000000000000d00000000",
            INIT_23 => X"0000000600000000000000100000000000000011000000000000002300000000",
            INIT_24 => X"0000000000000000000000000000000000000058000000000000002200000000",
            INIT_25 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_26 => X"0000002500000000000000200000000000000000000000000000000000000000",
            INIT_27 => X"0000005400000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"00000000000000000000000d0000000000000053000000000000004400000000",
            INIT_29 => X"0000000000000000000000270000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_2B => X"0000003800000000000000380000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000100000000000000029000000000000007900000000",
            INIT_2D => X"0000000000000000000000010000000000000049000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000004000000000000001300000000",
            INIT_2F => X"0000006700000000000000240000000000000044000000000000000000000000",
            INIT_30 => X"00000031000000000000004000000000000000a6000000000000000000000000",
            INIT_31 => X"000000560000000000000041000000000000004b000000000000003d00000000",
            INIT_32 => X"0000005000000000000000500000000000000079000000000000007300000000",
            INIT_33 => X"0000002600000000000000200000000000000043000000000000006a00000000",
            INIT_34 => X"0000007f00000000000000840000000000000081000000000000008d00000000",
            INIT_35 => X"000000ba00000000000000b10000000000000098000000000000009b00000000",
            INIT_36 => X"000000f900000000000000cc00000000000000cc00000000000000cc00000000",
            INIT_37 => X"0000007e00000000000000780000000000000000000000000000006900000000",
            INIT_38 => X"000000af00000000000000a800000000000000af00000000000000ae00000000",
            INIT_39 => X"000000cf00000000000000d300000000000000cd00000000000000ba00000000",
            INIT_3A => X"000000db000000000000010400000000000000e100000000000000ca00000000",
            INIT_3B => X"000000ac000000000000009600000000000000bf000000000000002200000000",
            INIT_3C => X"000000c200000000000000b000000000000000ae00000000000000bf00000000",
            INIT_3D => X"000000f200000000000000e700000000000000db00000000000000da00000000",
            INIT_3E => X"000000cd00000000000000f1000000000000010200000000000000fc00000000",
            INIT_3F => X"000000a600000000000000a600000000000000a6000000000000009100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d600000000000000d200000000000000b600000000000000ab00000000",
            INIT_41 => X"00000103000000000000011300000000000000cd00000000000000c800000000",
            INIT_42 => X"000000e200000000000000e100000000000000e300000000000000d500000000",
            INIT_43 => X"000000fd00000000000000eb00000000000000d500000000000000e100000000",
            INIT_44 => X"00000095000000000000008800000000000000a900000000000000e100000000",
            INIT_45 => X"000000dd00000000000000c400000000000000c700000000000000ae00000000",
            INIT_46 => X"000000df00000000000000ea00000000000000ee00000000000000f200000000",
            INIT_47 => X"0000008100000000000000b500000000000000c000000000000000e800000000",
            INIT_48 => X"0000004c00000000000000300000000000000027000000000000003d00000000",
            INIT_49 => X"00000090000000000000008400000000000000b4000000000000008400000000",
            INIT_4A => X"000000d600000000000000f300000000000000f200000000000000ea00000000",
            INIT_4B => X"0000003b00000000000000170000000000000033000000000000006f00000000",
            INIT_4C => X"0000002f000000000000002c0000000000000010000000000000001c00000000",
            INIT_4D => X"000000ce0000000000000066000000000000002f000000000000009600000000",
            INIT_4E => X"0000005a000000000000006e00000000000000c100000000000000e600000000",
            INIT_4F => X"0000003a000000000000002a000000000000001c000000000000001c00000000",
            INIT_50 => X"0000006800000000000000190000000000000012000000000000002f00000000",
            INIT_51 => X"0000007f00000000000000a7000000000000005d000000000000000000000000",
            INIT_52 => X"0000002200000000000000400000000000000067000000000000006e00000000",
            INIT_53 => X"0000002700000000000000370000000000000025000000000000002200000000",
            INIT_54 => X"00000000000000000000003a0000000000000018000000000000002200000000",
            INIT_55 => X"0000005100000000000000d40000000000000093000000000000002b00000000",
            INIT_56 => X"00000032000000000000002f000000000000005d000000000000003500000000",
            INIT_57 => X"000000160000000000000004000000000000002c000000000000003d00000000",
            INIT_58 => X"0000004c00000000000000000000000000000016000000000000000f00000000",
            INIT_59 => X"00000054000000000000008e00000000000000b7000000000000004800000000",
            INIT_5A => X"000000550000000000000019000000000000002d000000000000003d00000000",
            INIT_5B => X"00000015000000000000001b0000000000000010000000000000000f00000000",
            INIT_5C => X"00000008000000000000000e0000000000000000000000000000002800000000",
            INIT_5D => X"000000220000000000000042000000000000006b000000000000005900000000",
            INIT_5E => X"000000320000000000000082000000000000001d000000000000002a00000000",
            INIT_5F => X"000000680000000000000034000000000000000d000000000000001500000000",
            INIT_60 => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"00000037000000000000002d0000000000000033000000000000003f00000000",
            INIT_62 => X"0000000e00000000000000260000000000000083000000000000001200000000",
            INIT_63 => X"0000001600000000000000b90000000000000068000000000000002500000000",
            INIT_64 => X"0000000000000000000000200000000000000000000000000000000d00000000",
            INIT_65 => X"00000021000000000000003d000000000000001b000000000000001b00000000",
            INIT_66 => X"000000250000000000000000000000000000000d000000000000001400000000",
            INIT_67 => X"0000000b000000000000000500000000000000a200000000000000a300000000",
            INIT_68 => X"00000000000000000000001e0000000000000012000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000006a00000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000003b00000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000006700000000000000760000000000000066000000000000000000000000",
            INIT_7B => X"0000007300000000000000610000000000000064000000000000006300000000",
            INIT_7C => X"000000680000000000000070000000000000007e000000000000008f00000000",
            INIT_7D => X"0000005b000000000000004e000000000000004d000000000000006500000000",
            INIT_7E => X"0000006e00000000000000740000000000000075000000000000006200000000",
            INIT_7F => X"0000007500000000000000220000000000000000000000000000006600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE3;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE4 : if BRAM_NAME = "samplegold_layersamples_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000009300000000",
            INIT_01 => X"0000006f00000000000000470000000000000050000000000000001400000000",
            INIT_02 => X"0000008000000000000000790000000000000070000000000000009a00000000",
            INIT_03 => X"00000000000000000000000c000000000000003400000000000000c200000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"000000000000000000000000000000000000003b000000000000000000000000",
            INIT_06 => X"00000004000000000000004b0000000000000077000000000000004b00000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000003d00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000002900000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000006d00000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000005200000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000002e000000000000004a0000000000000007000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_1A => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_1F => X"00000000000000000000003e0000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000002400000000000000230000000000000000000000000000000000000000",
            INIT_33 => X"0000001c00000000000000230000000000000024000000000000001900000000",
            INIT_34 => X"0000002c00000000000000250000000000000024000000000000002100000000",
            INIT_35 => X"0000001a00000000000000120000000000000011000000000000001800000000",
            INIT_36 => X"0000001c00000000000000260000000000000026000000000000002a00000000",
            INIT_37 => X"000000020000000000000050000000000000001e000000000000002800000000",
            INIT_38 => X"00000028000000000000001c0000000000000015000000000000001d00000000",
            INIT_39 => X"0000002e00000000000000270000000000000013000000000000001c00000000",
            INIT_3A => X"0000002800000000000000270000000000000026000000000000002f00000000",
            INIT_3B => X"00000011000000000000000f0000000000000060000000000000002d00000000",
            INIT_3C => X"000000000000000000000014000000000000002c000000000000000200000000",
            INIT_3D => X"0000004900000000000000380000000000000016000000000000002800000000",
            INIT_3E => X"0000002b00000000000000230000000000000035000000000000002e00000000",
            INIT_3F => X"0000001d00000000000000000000000000000042000000000000000600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000019000000000000000f000000000000000a000000000000000d00000000",
            INIT_41 => X"000000560000000000000000000000000000002d000000000000001c00000000",
            INIT_42 => X"0000000000000000000000350000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000290000000000000000000000000000000000000000",
            INIT_44 => X"0000002a00000000000000260000000000000000000000000000001800000000",
            INIT_45 => X"0000000000000000000000340000000000000000000000000000000000000000",
            INIT_46 => X"0000002800000000000000000000000000000049000000000000000000000000",
            INIT_47 => X"00000000000000000000000d000000000000004b000000000000000700000000",
            INIT_48 => X"000000000000000000000011000000000000001f000000000000000000000000",
            INIT_49 => X"000000420000000000000000000000000000006d000000000000000000000000",
            INIT_4A => X"0000000000000000000000440000000000000000000000000000004e00000000",
            INIT_4B => X"0000000300000000000000000000000000000044000000000000003600000000",
            INIT_4C => X"0000000000000000000000110000000000000025000000000000001100000000",
            INIT_4D => X"0000000d000000000000004b0000000000000000000000000000002b00000000",
            INIT_4E => X"0000001b00000000000000040000000000000000000000000000004000000000",
            INIT_4F => X"0000001100000000000000150000000000000009000000000000003800000000",
            INIT_50 => X"0000000100000000000000000000000000000000000000000000001a00000000",
            INIT_51 => X"0000000000000000000000000000000000000034000000000000000000000000",
            INIT_52 => X"0000003300000000000000070000000000000048000000000000001800000000",
            INIT_53 => X"0000002f00000000000000150000000000000000000000000000005300000000",
            INIT_54 => X"0000001200000000000000000000000000000000000000000000002900000000",
            INIT_55 => X"0000000000000000000000000000000000000009000000000000001900000000",
            INIT_56 => X"0000000a00000000000000030000000000000000000000000000006300000000",
            INIT_57 => X"0000001900000000000000340000000000000031000000000000001300000000",
            INIT_58 => X"0000000000000000000000170000000000000000000000000000006600000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000001700000000000000220000000000000000000000000000000000000000",
            INIT_5B => X"000000430000000000000034000000000000003d000000000000000b00000000",
            INIT_5C => X"0000002e00000000000000400000000000000000000000000000000000000000",
            INIT_5D => X"0000001a0000000000000016000000000000001d000000000000000000000000",
            INIT_5E => X"000000270000000000000023000000000000002b000000000000002300000000",
            INIT_5F => X"0000001a0000000000000027000000000000001d000000000000002300000000",
            INIT_60 => X"0000001200000000000000000000000000000068000000000000000000000000",
            INIT_61 => X"000000280000000000000025000000000000001a000000000000001900000000",
            INIT_62 => X"0000001400000000000000210000000000000023000000000000002800000000",
            INIT_63 => X"00000000000000000000001f0000000000000025000000000000001800000000",
            INIT_64 => X"0000001a0000000000000014000000000000000c000000000000008b00000000",
            INIT_65 => X"0000002000000000000000170000000000000014000000000000001d00000000",
            INIT_66 => X"0000003d00000000000000280000000000000021000000000000003100000000",
            INIT_67 => X"0000007300000000000000190000000000000023000000000000001800000000",
            INIT_68 => X"000000100000000000000023000000000000002c000000000000002f00000000",
            INIT_69 => X"0000001800000000000000260000000000000022000000000000001800000000",
            INIT_6A => X"0000004e0000000000000028000000000000003b000000000000001d00000000",
            INIT_6B => X"0000004d0000000000000052000000000000004f000000000000005900000000",
            INIT_6C => X"0000004b0000000000000056000000000000005a000000000000005400000000",
            INIT_6D => X"0000003d00000000000000410000000000000045000000000000004e00000000",
            INIT_6E => X"0000005600000000000000490000000000000033000000000000003f00000000",
            INIT_6F => X"00000082000000000000004b0000000000000059000000000000005300000000",
            INIT_70 => X"0000001d000000000000003c0000000000000060000000000000005900000000",
            INIT_71 => X"00000037000000000000002e000000000000002a000000000000002900000000",
            INIT_72 => X"00000057000000000000003c0000000000000063000000000000003d00000000",
            INIT_73 => X"0000003e00000000000000910000000000000056000000000000005400000000",
            INIT_74 => X"00000054000000000000003f0000000000000000000000000000000d00000000",
            INIT_75 => X"0000003f00000000000000180000000000000029000000000000002100000000",
            INIT_76 => X"00000054000000000000005d0000000000000029000000000000003900000000",
            INIT_77 => X"00000019000000000000005a0000000000000021000000000000006200000000",
            INIT_78 => X"0000003b00000000000000570000000000000046000000000000001d00000000",
            INIT_79 => X"0000003300000000000000250000000000000003000000000000001300000000",
            INIT_7A => X"000000ac00000000000000210000000000000059000000000000008c00000000",
            INIT_7B => X"00000024000000000000002d0000000000000071000000000000006200000000",
            INIT_7C => X"0000002100000000000000330000000000000062000000000000000000000000",
            INIT_7D => X"000000a900000000000000400000000000000004000000000000000800000000",
            INIT_7E => X"0000006400000000000000bb0000000000000055000000000000006000000000",
            INIT_7F => X"00000046000000000000002e000000000000003b000000000000009300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE4;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE5 : if BRAM_NAME = "samplegold_layersamples_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001200000000000000290000000000000026000000000000008a00000000",
            INIT_01 => X"0000005300000000000000ca0000000000000023000000000000000000000000",
            INIT_02 => X"000000c60000000000000074000000000000006d000000000000004c00000000",
            INIT_03 => X"0000006c000000000000007e0000000000000041000000000000005500000000",
            INIT_04 => X"0000002a0000000000000027000000000000001a000000000000002c00000000",
            INIT_05 => X"00000054000000000000002e0000000000000090000000000000005f00000000",
            INIT_06 => X"00000060000000000000007b00000000000000cb000000000000002f00000000",
            INIT_07 => X"000000350000000000000066000000000000007a000000000000003100000000",
            INIT_08 => X"0000008d000000000000001e000000000000004b000000000000002100000000",
            INIT_09 => X"000000470000000000000067000000000000004b00000000000000a800000000",
            INIT_0A => X"0000002a000000000000004e0000000000000042000000000000004600000000",
            INIT_0B => X"0000000900000000000000170000000000000069000000000000005700000000",
            INIT_0C => X"0000009f00000000000000a00000000000000050000000000000002800000000",
            INIT_0D => X"00000012000000000000006a0000000000000053000000000000007000000000",
            INIT_0E => X"0000004d00000000000000480000000000000087000000000000002300000000",
            INIT_0F => X"0000005d00000000000000200000000000000000000000000000001a00000000",
            INIT_10 => X"00000073000000000000009b00000000000000b3000000000000005200000000",
            INIT_11 => X"00000094000000000000005e0000000000000096000000000000006f00000000",
            INIT_12 => X"000000000000000000000000000000000000004800000000000000a100000000",
            INIT_13 => X"00000030000000000000003e000000000000001e000000000000000000000000",
            INIT_14 => X"000000fb00000000000000640000000000000089000000000000008400000000",
            INIT_15 => X"000000280000000000000033000000000000002d00000000000000fb00000000",
            INIT_16 => X"000000150000000000000016000000000000000a000000000000001500000000",
            INIT_17 => X"00000020000000000000001d0000000000000025000000000000001a00000000",
            INIT_18 => X"00000026000000000000012e000000000000004e000000000000006000000000",
            INIT_19 => X"0000000900000000000000100000000000000018000000000000001500000000",
            INIT_1A => X"00000030000000000000001e000000000000000c000000000000000800000000",
            INIT_1B => X"0000001900000000000000170000000000000021000000000000001e00000000",
            INIT_1C => X"00000017000000000000001600000000000000dd000000000000006500000000",
            INIT_1D => X"00000015000000000000000d0000000000000014000000000000001400000000",
            INIT_1E => X"0000002600000000000000110000000000000026000000000000001b00000000",
            INIT_1F => X"0000002a00000000000000160000000000000021000000000000005700000000",
            INIT_20 => X"0000001b0000000000000015000000000000000d000000000000004800000000",
            INIT_21 => X"0000001e00000000000000210000000000000018000000000000000f00000000",
            INIT_22 => X"000000100000000000000051000000000000001b000000000000000700000000",
            INIT_23 => X"0000000300000000000000080000000000000007000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_26 => X"0000000a00000000000000010000000000000000000000000000000000000000",
            INIT_27 => X"000000080000000000000000000000000000000b000000000000001a00000000",
            INIT_28 => X"000000000000000000000021000000000000000000000000000000ac00000000",
            INIT_29 => X"00000000000000000000000e0000000000000020000000000000001e00000000",
            INIT_2A => X"000000000000000000000015000000000000000c000000000000000000000000",
            INIT_2B => X"00000000000000000000000e0000000000000000000000000000000b00000000",
            INIT_2C => X"0000005a000000000000001f0000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000a30000000000000000000000000000001e00000000",
            INIT_2F => X"0000004200000000000000000000000000000035000000000000001400000000",
            INIT_30 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_31 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"000000040000000000000000000000000000008e000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000008500000000",
            INIT_34 => X"0000000000000000000000000000000000000035000000000000000000000000",
            INIT_35 => X"0000000000000000000000110000000000000000000000000000001600000000",
            INIT_36 => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000012c00000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"00000069000000000000003c0000000000000000000000000000000000000000",
            INIT_3B => X"000000cc00000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000830000000000000011000000000000000000000000",
            INIT_3F => X"0000000000000000000000700000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_41 => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000003e00000000000000000000000000000000000000000000000d00000000",
            INIT_43 => X"0000000000000000000000270000000000000000000000000000000000000000",
            INIT_44 => X"00000000000000000000003f0000000000000008000000000000000000000000",
            INIT_45 => X"0000000000000000000000200000000000000000000000000000000000000000",
            INIT_46 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_47 => X"0000004a00000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000470000000000000000000000000000005500000000",
            INIT_49 => X"0000003d000000000000000000000000000000eb000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000006100000000",
            INIT_4B => X"000000000000000000000025000000000000005f000000000000002e00000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"000000000000000000000000000000000000000000000000000000ba00000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000025000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_62 => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000005400000000",
            INIT_64 => X"000000000000000000000000000000000000000000000000000000c500000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000002f00000000",
            INIT_66 => X"000000000000000000000000000000000000002d000000000000001300000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"000000af00000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"00000000000000000000000f0000000000000000000000000000009200000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000003b00000000",
            INIT_6C => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"000000000000000000000000000000000000002d000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000015a00000000",
            INIT_70 => X"0000000000000000000000000000000000000092000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000003600000000",
            INIT_72 => X"000000d700000000000000000000000000000004000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000059000000000000000000000000",
            INIT_74 => X"000000000000000000000000000000000000000000000000000000be00000000",
            INIT_75 => X"0000001900000000000000000000000000000000000000000000000400000000",
            INIT_76 => X"000000d4000000000000003e0000000000000000000000000000000000000000",
            INIT_77 => X"0000008700000000000000000000000000000007000000000000000000000000",
            INIT_78 => X"0000000700000000000000360000000000000000000000000000000000000000",
            INIT_79 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_7A => X"00000011000000000000005f0000000000000000000000000000006100000000",
            INIT_7B => X"000000b60000000000000000000000000000002d000000000000000000000000",
            INIT_7C => X"000000000000000000000043000000000000001d000000000000000000000000",
            INIT_7D => X"0000004d00000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"000000220000000000000000000000000000002a000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE5;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE6 : if BRAM_NAME = "samplegold_layersamples_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b400000000000000000000000000000002000000000000004400000000",
            INIT_01 => X"0000000000000000000000850000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000003a00000000000001000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000051000000000000000000000000",
            INIT_06 => X"000000000000000000000007000000000000003d000000000000003c00000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"00000000000000000000008b0000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000004300000000000000820000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000001000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000030000000000000003200000000",
            INIT_12 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000009000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000009200000000000000970000000000000093000000000000008b00000000",
            INIT_4D => X"0000009b00000000000000ab000000000000009c000000000000008300000000",
            INIT_4E => X"000000710000000000000066000000000000005a000000000000007400000000",
            INIT_4F => X"00000099000000000000009a000000000000007f000000000000007900000000",
            INIT_50 => X"00000066000000000000009e0000000000000098000000000000009a00000000",
            INIT_51 => X"0000002a0000000000000039000000000000006e000000000000007600000000",
            INIT_52 => X"0000006e00000000000000200000000000000000000000000000000000000000",
            INIT_53 => X"000000a1000000000000007c0000000000000037000000000000007d00000000",
            INIT_54 => X"00000039000000000000004d000000000000009f00000000000000a000000000",
            INIT_55 => X"0000000000000000000000000000000000000022000000000000001500000000",
            INIT_56 => X"0000006200000000000000260000000000000000000000000000000000000000",
            INIT_57 => X"0000009f00000000000000910000000000000032000000000000000000000000",
            INIT_58 => X"000000000000000000000014000000000000005a000000000000006600000000",
            INIT_59 => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_5A => X"0000000000000000000000460000000000000000000000000000000000000000",
            INIT_5B => X"00000017000000000000009f0000000000000069000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_5E => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_5F => X"000000120000000000000006000000000000002f000000000000006e00000000",
            INIT_60 => X"0000002c00000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000005e00000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000250000000000000000000000000000006200000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_66 => X"0000003700000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000011000000000000003600000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_69 => X"0000000000000000000000470000000000000000000000000000000000000000",
            INIT_6A => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000002000000000000000000000000000000012000000000000000000000000",
            INIT_6C => X"000000000000000000000000000000000000002f000000000000000000000000",
            INIT_6D => X"000000000000000000000000000000000000005e000000000000003700000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000001a00000000000000000000000000000000000000000000000e00000000",
            INIT_70 => X"0000004b00000000000000020000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000006a00000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE6;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE7 : if BRAM_NAME = "samplegold_layersamples_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"00000009000000000000000d0000000000000000000000000000000000000000",
            INIT_1B => X"0000002d00000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"000000000000000000000000000000000000000e000000000000000b00000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"000000080000000000000000000000000000000e000000000000000000000000",
            INIT_1F => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_20 => X"0000002b000000000000002e0000000000000003000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_26 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000600000000000000130000000000000012000000000000000300000000",
            INIT_28 => X"0000000000000000000000200000000000000000000000000000001800000000",
            INIT_29 => X"0000005200000000000000500000000000000000000000000000000000000000",
            INIT_2A => X"0000003f000000000000004d000000000000005b000000000000006500000000",
            INIT_2B => X"0000003d000000000000002f000000000000002e000000000000003b00000000",
            INIT_2C => X"0000001100000000000000210000000000000026000000000000002d00000000",
            INIT_2D => X"000000300000000000000000000000000000002f000000000000000000000000",
            INIT_2E => X"0000003500000000000000310000000000000036000000000000003100000000",
            INIT_2F => X"0000004100000000000000450000000000000041000000000000003600000000",
            INIT_30 => X"0000000000000000000000290000000000000009000000000000001600000000",
            INIT_31 => X"0000005b000000000000005d0000000000000018000000000000002a00000000",
            INIT_32 => X"00000119000000000000001c000000000000002f000000000000003a00000000",
            INIT_33 => X"00000088000000000000009000000000000000c700000000000000f700000000",
            INIT_34 => X"0000003a00000000000000000000000000000000000000000000002400000000",
            INIT_35 => X"0000002e0000000000000039000000000000002f000000000000002b00000000",
            INIT_36 => X"00000136000000000000018e0000000000000065000000000000002b00000000",
            INIT_37 => X"000000000000000000000000000000000000002f00000000000000ae00000000",
            INIT_38 => X"0000001a00000000000000360000000000000000000000000000000000000000",
            INIT_39 => X"0000001d0000000000000025000000000000001c000000000000001200000000",
            INIT_3A => X"0000000000000000000000370000000000000086000000000000001300000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"00000000000000000000001d000000000000002e000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000004c00000000000000050000000000000000000000000000000000000000",
            INIT_46 => X"000000000000000000000000000000000000002e000000000000000c00000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000d1000000000000010a000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000004c00000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"00000000000000000000005300000000000000d400000000000000ae00000000",
            INIT_4F => X"0000004600000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"000000ae00000000000000e000000000000000d4000000000000003300000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000004d00000000",
            INIT_52 => X"0000011f00000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000062000000000000010e00000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000008800000000000000ba0000000000000076000000000000000e00000000",
            INIT_56 => X"000000000000000000000005000000000000007400000000000000ba00000000",
            INIT_57 => X"000000000000000000000000000000000000004f000000000000003d00000000",
            INIT_58 => X"0000003e0000000000000098000000000000000f000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000002d00000000000000050000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000006d00000000000000bb0000000000000077000000000000002b00000000",
            INIT_5E => X"000000bf00000000000000d600000000000000d3000000000000008c00000000",
            INIT_5F => X"00000018000000000000003b000000000000006800000000000000a300000000",
            INIT_60 => X"00000028000000000000004f0000000000000003000000000000002600000000",
            INIT_61 => X"000000d500000000000000010000000000000000000000000000000000000000",
            INIT_62 => X"00000154000000000000012b00000000000000ef00000000000000bc00000000",
            INIT_63 => X"000000d700000000000001040000000000000132000000000000015a00000000",
            INIT_64 => X"000000000000000000000043000000000000007b00000000000000ba00000000",
            INIT_65 => X"0000001200000000000000110000000000000000000000000000000000000000",
            INIT_66 => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000c000000000000000c0000000000000000000000000000000000000000",
            INIT_69 => X"00000071000000000000003b0000000000000000000000000000000000000000",
            INIT_6A => X"000000d500000000000000060000000000000006000000000000003900000000",
            INIT_6B => X"000000e400000000000000900000000000000069000000000000008e00000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000007800000000",
            INIT_6D => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_6E => X"00000060000000000000003b0000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000008b00000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000003b00000000000000260000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE7;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE8 : if BRAM_NAME = "samplegold_layersamples_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000020000000000000000000000000",
            INIT_02 => X"0000000000000000000000220000000000000000000000000000000000000000",
            INIT_03 => X"0000004600000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000008300000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000003100000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000041000000000000003100000000",
            INIT_0A => X"0000000000000000000000480000000000000000000000000000000000000000",
            INIT_0B => X"0000002d000000000000000a0000000000000069000000000000000000000000",
            INIT_0C => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000004600000000",
            INIT_0E => X"000000a300000000000000610000000000000000000000000000000f00000000",
            INIT_0F => X"0000000000000000000000630000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000001710000000000000003000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000200000000000000060000000000000050000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000001a00000000000000000000000000000022000000000000000000000000",
            INIT_1B => X"0000002200000000000000270000000000000053000000000000003600000000",
            INIT_1C => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"00000000000000000000001b0000000000000000000000000000001500000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000007900000000",
            INIT_1F => X"000000000000000000000000000000000000004a000000000000003700000000",
            INIT_20 => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000002b0000000000000000000000000000002c000000000000000f00000000",
            INIT_22 => X"0000000800000000000000000000000000000000000000000000001800000000",
            INIT_23 => X"00000050000000000000006d000000000000005e000000000000014400000000",
            INIT_24 => X"0000001e000000000000001a000000000000003a000000000000004100000000",
            INIT_25 => X"0000000900000000000000000000000000000000000000000000002b00000000",
            INIT_26 => X"000000c000000000000000010000000000000000000000000000000000000000",
            INIT_27 => X"00000027000000000000004c0000000000000066000000000000007300000000",
            INIT_28 => X"0000002200000000000000250000000000000000000000000000001f00000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000001700000000000000320000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000040000000000000047000000000000002600000000",
            INIT_2C => X"0000000000000000000000190000000000000017000000000000000a00000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000000000001a000000000000003200000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"00000000000000000000000f000000000000001d000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_39 => X"0000000d00000000000000120000000000000000000000000000000000000000",
            INIT_3A => X"0000003f00000000000000320000000000000004000000000000000000000000",
            INIT_3B => X"000000e800000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"000000000000000000000000000000000000001000000000000000b600000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_3E => X"0000004000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000003a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_43 => X"0000004200000000000000a50000000000000076000000000000000000000000",
            INIT_44 => X"000000f4000000000000009b0000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000069000000000000015400000000",
            INIT_46 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000007700000000000000680000000000000000000000000000001100000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000006300000000",
            INIT_49 => X"000000cc000000000000010600000000000000ec000000000000007800000000",
            INIT_4A => X"0000002200000000000000000000000000000052000000000000009e00000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000061000000000000000000000000",
            INIT_4F => X"0000006300000000000000520000000000000037000000000000002400000000",
            INIT_50 => X"0000003b000000000000005b000000000000008d000000000000007100000000",
            INIT_51 => X"0000000000000000000000000000000000000033000000000000003600000000",
            INIT_52 => X"000000b600000000000000c700000000000000c8000000000000000000000000",
            INIT_53 => X"000000200000000000000048000000000000006a000000000000008f00000000",
            INIT_54 => X"00000023000000000000001d0000000000000004000000000000000700000000",
            INIT_55 => X"00000000000000000000001b0000000000000053000000000000002400000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000009900000000000000120000000000000000000000000000000000000000",
            INIT_58 => X"00000000000000000000005b000000000000009300000000000000b400000000",
            INIT_59 => X"00000000000000000000000b000000000000000a000000000000000000000000",
            INIT_5A => X"0000000000000000000000200000000000000043000000000000000b00000000",
            INIT_5B => X"0000000000000000000000000000000000000018000000000000000000000000",
            INIT_5C => X"0000003b00000000000000920000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_5F => X"0000008e00000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000003f00000000",
            INIT_61 => X"000000040000000000000000000000000000000c000000000000000000000000",
            INIT_62 => X"000000260000000000000012000000000000000d000000000000000900000000",
            INIT_63 => X"000000000000000000000000000000000000003b000000000000009200000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"000000100000000000000036000000000000000d000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000007c00000000000000770000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000004e00000000",
            INIT_78 => X"00000000000000000000002b0000000000000018000000000000000000000000",
            INIT_79 => X"00000036000000000000008800000000000000b2000000000000010200000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000002400000000000000580000000000000000000000000000000000000000",
            INIT_7C => X"0000001c00000000000000440000000000000000000000000000000000000000",
            INIT_7D => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"000000b2000000000000006500000000000000a5000000000000008500000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE8;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE9 : if BRAM_NAME = "samplegold_layersamples_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000035000000000000009400000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"000000000000000000000000000000000000003d000000000000000000000000",
            INIT_04 => X"0000004100000000000000190000000000000037000000000000001600000000",
            INIT_05 => X"000000a900000000000000410000000000000093000000000000000b00000000",
            INIT_06 => X"000000d200000000000000000000000000000082000000000000009f00000000",
            INIT_07 => X"000000250000000000000042000000000000005f000000000000007700000000",
            INIT_08 => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_09 => X"0000000000000000000000010000000000000027000000000000000000000000",
            INIT_0A => X"0000000000000000000000300000000000000000000000000000000000000000",
            INIT_0B => X"0000007200000000000000640000000000000049000000000000002d00000000",
            INIT_0C => X"00000063000000000000006b0000000000000080000000000000007800000000",
            INIT_0D => X"0000000000000000000000000000000000000002000000000000003000000000",
            INIT_0E => X"0000001c00000000000000000000000000000031000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000028000000000000003500000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000050000000000000000000000000",
            INIT_12 => X"0000002b00000000000000180000000000000008000000000000004300000000",
            INIT_13 => X"000000010000000000000000000000000000000b000000000000000a00000000",
            INIT_14 => X"0000000000000000000000bb0000000000000074000000000000002b00000000",
            INIT_15 => X"0000007500000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"000000090000000000000010000000000000000c000000000000000a00000000",
            INIT_17 => X"000000a900000000000000000000000000000000000000000000000900000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"00000000000000000000005c0000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000029000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000003700000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000024000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000020000000000000010000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000004c00000000",
            INIT_34 => X"0000003c00000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000007a00000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000003500000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000390000000000000000000000000000000000000000",
            INIT_47 => X"00000000000000000000001c000000000000004c000000000000004700000000",
            INIT_48 => X"0000000000000000000000000000000000000029000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000059000000000000000000000000",
            INIT_4B => X"00000000000000000000000f000000000000001e000000000000002600000000",
            INIT_4C => X"00000010000000000000002b000000000000001f000000000000001b00000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"000000190000000000000009000000000000001600000000000000d000000000",
            INIT_4F => X"0000003100000000000000000000000000000012000000000000001500000000",
            INIT_50 => X"000000000000000000000000000000000000000c000000000000004000000000",
            INIT_51 => X"0000009400000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000001a000000000000001c0000000000000020000000000000003200000000",
            INIT_53 => X"0000000200000000000000000000000000000000000000000000001400000000",
            INIT_54 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"000000420000000000000048000000000000001d000000000000001400000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000003e00000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000008000000000000000450000000000000057000000000000005200000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000014800000000000000ef000000000000001e000000000000001f00000000",
            INIT_6A => X"00000000000000000000000000000000000000c9000000000000012800000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000002e000000000000005c0000000000000072000000000000005c00000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"000000c100000000000000960000000000000018000000000000000000000000",
            INIT_6F => X"0000007a0000000000000089000000000000008900000000000000f700000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"00000020000000000000002e000000000000000f000000000000000300000000",
            INIT_75 => X"000000c4000000000000006c00000000000000c9000000000000004e00000000",
            INIT_76 => X"0000006e00000000000000d800000000000000bd00000000000000ce00000000",
            INIT_77 => X"0000007300000000000000af0000000000000094000000000000000e00000000",
            INIT_78 => X"0000000000000000000000240000000000000041000000000000007100000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000220000000000000000000000000000000500000000",
            INIT_7B => X"0000002000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"000000c200000000000000a8000000000000008d000000000000005a00000000",
            INIT_7D => X"0000001b000000000000004d000000000000006a000000000000008f00000000",
            INIT_7E => X"0000002d00000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"000000000000000000000000000000000000002a000000000000005f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE9;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE10 : if BRAM_NAME = "samplegold_layersamples_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000003200000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"000000000000000000000000000000000000000e000000000000001100000000",
            INIT_04 => X"00000072000000000000006d00000000000000a3000000000000006b00000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000006b00000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"00000000000000000000000e000000000000007e000000000000004700000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000003900000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000003700000000000000380000000000000038000000000000003800000000",
            INIT_0F => X"0000003300000000000000370000000000000037000000000000003800000000",
            INIT_10 => X"000000380000000000000037000000000000003f000000000000003d00000000",
            INIT_11 => X"0000003800000000000000380000000000000038000000000000003800000000",
            INIT_12 => X"0000003900000000000000380000000000000039000000000000003800000000",
            INIT_13 => X"00000062000000000000003e0000000000000038000000000000003700000000",
            INIT_14 => X"0000003900000000000000380000000000000033000000000000003800000000",
            INIT_15 => X"0000003700000000000000340000000000000033000000000000003900000000",
            INIT_16 => X"00000035000000000000003e0000000000000037000000000000003900000000",
            INIT_17 => X"0000002f00000000000000620000000000000048000000000000005300000000",
            INIT_18 => X"0000003900000000000000370000000000000037000000000000002800000000",
            INIT_19 => X"00000035000000000000003a0000000000000047000000000000004900000000",
            INIT_1A => X"000000580000000000000027000000000000005c000000000000003700000000",
            INIT_1B => X"00000044000000000000007b000000000000007f000000000000006400000000",
            INIT_1C => X"00000045000000000000003d0000000000000041000000000000004600000000",
            INIT_1D => X"00000036000000000000002c0000000000000038000000000000001c00000000",
            INIT_1E => X"0000004b00000000000000410000000000000037000000000000004b00000000",
            INIT_1F => X"0000003d00000000000000520000000000000060000000000000005f00000000",
            INIT_20 => X"00000068000000000000006a0000000000000043000000000000000700000000",
            INIT_21 => X"0000001800000000000000380000000000000018000000000000005300000000",
            INIT_22 => X"000000710000000000000022000000000000001a000000000000001800000000",
            INIT_23 => X"00000049000000000000008e000000000000006e000000000000007200000000",
            INIT_24 => X"0000002e000000000000001d000000000000004f000000000000004100000000",
            INIT_25 => X"00000068000000000000007d0000000000000088000000000000003500000000",
            INIT_26 => X"000000370000000000000045000000000000003c000000000000006500000000",
            INIT_27 => X"00000018000000000000003e0000000000000021000000000000002d00000000",
            INIT_28 => X"0000001500000000000000340000000000000084000000000000001200000000",
            INIT_29 => X"0000006c00000000000000640000000000000070000000000000004a00000000",
            INIT_2A => X"00000066000000000000006b0000000000000058000000000000004700000000",
            INIT_2B => X"0000000000000000000000570000000000000066000000000000005c00000000",
            INIT_2C => X"0000004c00000000000000430000000000000058000000000000006500000000",
            INIT_2D => X"00000062000000000000005c0000000000000051000000000000005900000000",
            INIT_2E => X"0000005a000000000000006f000000000000006d000000000000005e00000000",
            INIT_2F => X"000000620000000000000055000000000000005a000000000000005400000000",
            INIT_30 => X"00000083000000000000007e0000000000000078000000000000007400000000",
            INIT_31 => X"0000008a0000000000000089000000000000008f00000000000000a000000000",
            INIT_32 => X"0000005f00000000000000760000000000000082000000000000008800000000",
            INIT_33 => X"0000005100000000000000460000000000000031000000000000005100000000",
            INIT_34 => X"0000006700000000000000370000000000000034000000000000004300000000",
            INIT_35 => X"0000006d00000000000000720000000000000074000000000000006300000000",
            INIT_36 => X"00000035000000000000005d0000000000000069000000000000006900000000",
            INIT_37 => X"0000003200000000000000330000000000000000000000000000001700000000",
            INIT_38 => X"000000a6000000000000006d0000000000000009000000000000001900000000",
            INIT_39 => X"00000055000000000000006a0000000000000084000000000000009200000000",
            INIT_3A => X"0000001b00000000000000180000000000000022000000000000002c00000000",
            INIT_3B => X"0000000500000000000000000000000000000000000000000000000200000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000400000000000000430000000000000023000000000000001000000000",
            INIT_3F => X"0000000100000000000000020000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"00000011000000000000000d0000000000000000000000000000000000000000",
            INIT_42 => X"000000090000000000000005000000000000001f000000000000002800000000",
            INIT_43 => X"00000000000000000000000a0000000000000006000000000000000a00000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000002f000000000000001c000000000000000d000000000000000900000000",
            INIT_46 => X"0000001400000000000000140000000000000014000000000000001200000000",
            INIT_47 => X"0000001800000000000000140000000000000014000000000000001400000000",
            INIT_48 => X"00000012000000000000000d0000000000000011000000000000001900000000",
            INIT_49 => X"0000001200000000000000150000000000000014000000000000001500000000",
            INIT_4A => X"0000001400000000000000150000000000000014000000000000001400000000",
            INIT_4B => X"0000001100000000000000160000000000000014000000000000001400000000",
            INIT_4C => X"00000015000000000000000b0000000000000000000000000000000900000000",
            INIT_4D => X"0000001400000000000000120000000000000015000000000000001400000000",
            INIT_4E => X"0000001400000000000000160000000000000016000000000000001600000000",
            INIT_4F => X"000000000000000000000000000000000000000b000000000000000b00000000",
            INIT_50 => X"0000001500000000000000130000000000000002000000000000000000000000",
            INIT_51 => X"0000000d00000000000000000000000000000000000000000000001400000000",
            INIT_52 => X"0000000c00000000000000220000000000000018000000000000001700000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_54 => X"0000000e00000000000000060000000000000000000000000000000300000000",
            INIT_55 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"00000006000000000000001f0000000000000008000000000000001300000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_58 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_59 => X"000000040000000000000003000000000000002d000000000000000700000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000001000000000000001800000000",
            INIT_5D => X"00000000000000000000000c0000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000400000000000000190000000000000000000000000000000000000000",
            INIT_61 => X"0000001200000000000000000000000000000000000000000000002700000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000900000000000000000000000000000000000000000000000400000000",
            INIT_70 => X"0000000f00000000000000000000000000000007000000000000001100000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000001300000000000000170000000000000029000000000000000900000000",
            INIT_73 => X"0000000d000000000000001b0000000000000018000000000000001400000000",
            INIT_74 => X"0000009900000000000000570000000000000011000000000000000600000000",
            INIT_75 => X"0000003d000000000000007a00000000000000a100000000000000b500000000",
            INIT_76 => X"0000000700000000000000100000000000000022000000000000001b00000000",
            INIT_77 => X"0000000e000000000000000d0000000000000015000000000000001100000000",
            INIT_78 => X"000000df0000000000000114000000000000006f000000000000000e00000000",
            INIT_79 => X"000000230000000000000045000000000000003c000000000000006a00000000",
            INIT_7A => X"0000002300000000000000000000000000000009000000000000000f00000000",
            INIT_7B => X"0000001200000000000000180000000000000013000000000000001900000000",
            INIT_7C => X"00000063000000000000003c000000000000005f000000000000003800000000",
            INIT_7D => X"0000000e00000000000000120000000000000015000000000000004600000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE10;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE11 : if BRAM_NAME = "samplegold_layersamples_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"00000046000000000000001e0000000000000000000000000000000000000000",
            INIT_25 => X"000000000000000000000000000000000000000e000000000000004700000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000003900000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000005400000000000000000000000000000000000000000000001200000000",
            INIT_2D => X"00000062000000000000002b000000000000000b000000000000003000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000013400000000000000350000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000071000000000000015300000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"00000000000000000000003f0000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"00000008000000000000000b0000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_44 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_46 => X"0000000700000000000000000000000000000000000000000000002400000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000500000000000000150000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_4E => X"00000018000000000000001e0000000000000000000000000000004400000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000001000000000000000110000000000000000000000000000003f00000000",
            INIT_52 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_53 => X"0000000b00000000000000110000000000000005000000000000000000000000",
            INIT_54 => X"0000002a00000000000000000000000000000000000000000000001300000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000019000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000300000000000000000000000000000006000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000030000000000000018000000000000000f00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000e00000000000000050000000000000006000000000000001300000000",
            INIT_61 => X"0000000e00000000000000040000000000000023000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000001c000000000000001e0000000000000002000000000000000000000000",
            INIT_64 => X"0000001e00000000000000160000000000000005000000000000001100000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000001d00000000000000240000000000000038000000000000001900000000",
            INIT_68 => X"0000000000000000000000220000000000000020000000000000001800000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"000000250000000000000018000000000000001a000000000000001300000000",
            INIT_6B => X"00000039000000000000003d0000000000000038000000000000003100000000",
            INIT_6C => X"000000000000000000000009000000000000002f000000000000002f00000000",
            INIT_6D => X"000000260000000000000018000000000000000b000000000000000000000000",
            INIT_6E => X"000000eb0000000000000021000000000000001c000000000000002600000000",
            INIT_6F => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_70 => X"000000ea00000000000000ee00000000000000ec00000000000000ed00000000",
            INIT_71 => X"000000ec00000000000000ec00000000000000ec00000000000000ed00000000",
            INIT_72 => X"000000ed00000000000000ec00000000000000ed00000000000000ec00000000",
            INIT_73 => X"000000ed00000000000000ec00000000000000ed00000000000000ed00000000",
            INIT_74 => X"000000f400000000000000ef00000000000000ec00000000000000ec00000000",
            INIT_75 => X"000000ec00000000000000ec00000000000000e500000000000000d000000000",
            INIT_76 => X"000000ed00000000000000ec00000000000000eb00000000000000ee00000000",
            INIT_77 => X"000000e700000000000000f200000000000000ed00000000000000ed00000000",
            INIT_78 => X"000000bb00000000000000ac00000000000000cc00000000000000f600000000",
            INIT_79 => X"000000ef00000000000000ee00000000000000ef00000000000000d400000000",
            INIT_7A => X"000000ef00000000000000f100000000000000ea00000000000000e500000000",
            INIT_7B => X"000000d200000000000000d7000000000000010000000000000000f100000000",
            INIT_7C => X"000000d10000000000000092000000000000009e00000000000000a300000000",
            INIT_7D => X"0000009800000000000000f100000000000000ef00000000000000f000000000",
            INIT_7E => X"000000ee00000000000000ea00000000000000e3000000000000009900000000",
            INIT_7F => X"000000e100000000000000e400000000000000e600000000000000e300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE11;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE12 : if BRAM_NAME = "samplegold_layersamples_instance12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bd00000000000000c900000000000000e600000000000000e900000000",
            INIT_01 => X"0000009f000000000000008900000000000000f100000000000000a900000000",
            INIT_02 => X"000000d900000000000000e700000000000000d400000000000000f200000000",
            INIT_03 => X"000000d500000000000000c900000000000000d200000000000000cd00000000",
            INIT_04 => X"000000bc0000000000000091000000000000009900000000000000a300000000",
            INIT_05 => X"000000b00000000000000078000000000000008300000000000000ec00000000",
            INIT_06 => X"0000001d000000000000002300000000000000e1000000000000009600000000",
            INIT_07 => X"000000e500000000000000f400000000000000ac000000000000003e00000000",
            INIT_08 => X"000000b100000000000000ca00000000000000c000000000000000cd00000000",
            INIT_09 => X"0000009e000000000000005a0000000000000078000000000000000000000000",
            INIT_0A => X"000000da00000000000000a1000000000000008000000000000000a700000000",
            INIT_0B => X"000000540000000000000062000000000000008300000000000000aa00000000",
            INIT_0C => X"0000000300000000000000a30000000000000075000000000000005c00000000",
            INIT_0D => X"000000e200000000000000c6000000000000009600000000000000cc00000000",
            INIT_0E => X"0000009900000000000000b000000000000000ef00000000000000ed00000000",
            INIT_0F => X"0000009c00000000000000ac00000000000000a600000000000000a500000000",
            INIT_10 => X"00000088000000000000009d000000000000007e000000000000009200000000",
            INIT_11 => X"0000008a000000000000008e0000000000000090000000000000009000000000",
            INIT_12 => X"0000004e00000000000000790000000000000068000000000000008600000000",
            INIT_13 => X"000000450000000000000039000000000000003d000000000000005d00000000",
            INIT_14 => X"0000000700000000000000000000000000000000000000000000005600000000",
            INIT_15 => X"0000002f00000000000000180000000000000011000000000000000500000000",
            INIT_16 => X"0000001300000000000000200000000000000034000000000000003000000000",
            INIT_17 => X"00000055000000000000003d0000000000000014000000000000001100000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000003100000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000570000000000000041000000000000005800000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000005a0000000000000066000000000000002a000000000000000000000000",
            INIT_1E => X"0000002f0000000000000022000000000000004d000000000000005b00000000",
            INIT_1F => X"000000000000000000000000000000000000007f000000000000005300000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"000000000000000000000028000000000000005c000000000000000000000000",
            INIT_22 => X"0000006100000000000000510000000000000047000000000000000b00000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000009100000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"00000053000000000000002f0000000000000000000000000000000000000000",
            INIT_26 => X"00000098000000000000006f000000000000005b000000000000004b00000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000009000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000910000000000000030000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000e70000000000000000000000000000000000000000",
            INIT_42 => X"00000084000000000000000d0000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000003100000000000000230000000000000000000000000000000000000000",
            INIT_45 => X"00000029000000000000002c0000000000000000000000000000017700000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000600000000000000300000000000000000000000000000000000000000",
            INIT_51 => X"000000af00000000000000260000000000000009000000000000000500000000",
            INIT_52 => X"0000006800000000000000500000000000000042000000000000005a00000000",
            INIT_53 => X"0000001200000000000000000000000000000000000000000000008f00000000",
            INIT_54 => X"0000000000000000000000000000000000000027000000000000000000000000",
            INIT_55 => X"0000000000000000000000620000000000000027000000000000000800000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000270000000000000012000000000000002500000000",
            INIT_58 => X"0000002400000000000000150000000000000029000000000000002500000000",
            INIT_59 => X"0000000000000000000000380000000000000054000000000000002600000000",
            INIT_5A => X"00000000000000000000006a0000000000000069000000000000000000000000",
            INIT_5B => X"0000002c00000000000000000000000000000000000000000000000400000000",
            INIT_5C => X"000000370000000000000035000000000000002d000000000000003900000000",
            INIT_5D => X"0000008700000000000000790000000000000024000000000000005400000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000001100000000000000500000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"000000000000000000000037000000000000003c000000000000000b00000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000007e00000000000000bd0000000000000085000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000b0000000000000004c000000000000001400000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000007200000000000000850000000000000041000000000000001600000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000005200000000",
            INIT_75 => X"0000007b00000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"00000000000000000000000000000000000000ac00000000000000d000000000",
            INIT_77 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"00000075000000000000001c000000000000000e000000000000000300000000",
            INIT_79 => X"0000000000000000000000ad000000000000007c000000000000002b00000000",
            INIT_7A => X"000000000000000000000045000000000000008c000000000000000000000000",
            INIT_7B => X"0000001000000000000000180000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000320000000000000021000000000000000000000000",
            INIT_7E => X"0000002c00000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE12;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE13 : if BRAM_NAME = "samplegold_layersamples_instance13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003c0000000000000034000000000000001e000000000000000000000000",
            INIT_01 => X"0000007200000000000000770000000000000068000000000000006d00000000",
            INIT_02 => X"0000000200000000000000280000000000000057000000000000005700000000",
            INIT_03 => X"0000001b00000000000000310000000000000000000000000000003a00000000",
            INIT_04 => X"0000003f000000000000000f0000000000000006000000000000000b00000000",
            INIT_05 => X"000000c2000000000000009c0000000000000068000000000000007d00000000",
            INIT_06 => X"0000007a00000000000000a400000000000000c100000000000000d500000000",
            INIT_07 => X"0000002700000000000000340000000000000051000000000000005800000000",
            INIT_08 => X"0000007d00000000000000000000000000000008000000000000000000000000",
            INIT_09 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000006700000000000000000000000000000000000000000000000500000000",
            INIT_0D => X"0000015900000000000000000000000000000000000000000000001f00000000",
            INIT_0E => X"0000000c00000000000000010000000000000010000000000000006300000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000004d00000000",
            INIT_10 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_11 => X"0000003d000000000000000e0000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000018000000000000000d00000000",
            INIT_13 => X"00000000000000000000001c0000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000410000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"000000000000000000000008000000000000000f000000000000000000000000",
            INIT_7F => X"0000000b00000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE13;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE14 : if BRAM_NAME = "samplegold_layersamples_instance14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_04 => X"0000000000000000000000020000000000000001000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"000000000000000000000010000000000000001f000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000002800000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000003000000000000000900000000",
            INIT_15 => X"0000000000000000000000520000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_17 => X"00000000000000000000001a0000000000000002000000000000001f00000000",
            INIT_18 => X"0000000600000000000000000000000000000005000000000000001800000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"000000000000000000000000000000000000002a000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000003000000000000001900000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000380000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000003900000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000002d00000000000000400000000000000001000000000000000200000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_29 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"000000000000000000000000000000000000000f000000000000001700000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000027000000000000000000000000",
            INIT_30 => X"0000000100000000000000000000000000000010000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000002800000000000000070000000000000011000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000120000000000000014000000000000000000000000",
            INIT_37 => X"0000000000000000000000060000000000000002000000000000000000000000",
            INIT_38 => X"00000021000000000000000e0000000000000011000000000000001b00000000",
            INIT_39 => X"000000000000000000000000000000000000000c000000000000002200000000",
            INIT_3A => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_3B => X"0000001300000000000000100000000000000013000000000000000000000000",
            INIT_3C => X"0000000800000000000000150000000000000010000000000000000a00000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"000000220000000000000000000000000000000d000000000000000000000000",
            INIT_3F => X"000000090000000000000009000000000000001d000000000000001500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000002c00000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"000000000000000000000019000000000000003a000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000002200000000000000520000000000000000000000000000000000000000",
            INIT_4A => X"000000030000000000000030000000000000001e000000000000004700000000",
            INIT_4B => X"0000000300000000000000200000000000000000000000000000000800000000",
            INIT_4C => X"000000060000000000000023000000000000002a000000000000003a00000000",
            INIT_4D => X"0000007a00000000000000ab0000000000000000000000000000000100000000",
            INIT_4E => X"00000059000000000000009d0000000000000111000000000000007300000000",
            INIT_4F => X"00000094000000000000008900000000000000a9000000000000007400000000",
            INIT_50 => X"0000007600000000000000ad00000000000000ae00000000000000b300000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000005300000000",
            INIT_52 => X"0000007400000000000000290000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000043000000000000005e00000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000005500000000000000080000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000002000000000000005e00000000",
            INIT_5E => X"0000001c00000000000000610000000000000007000000000000000000000000",
            INIT_5F => X"0000003100000000000000350000000000000008000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000004c00000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000800000000000000000000000000000000000000000000003a00000000",
            INIT_65 => X"00000000000000000000005d000000000000007d000000000000006600000000",
            INIT_66 => X"0000007000000000000000220000000000000000000000000000000000000000",
            INIT_67 => X"00000001000000000000003f0000000000000021000000000000002d00000000",
            INIT_68 => X"000000310000000000000069000000000000007f000000000000004000000000",
            INIT_69 => X"0000000800000000000000150000000000000035000000000000001b00000000",
            INIT_6A => X"000000000000000000000000000000000000000a000000000000001500000000",
            INIT_6B => X"0000002200000000000000190000000000000004000000000000004300000000",
            INIT_6C => X"0000001a00000000000000050000000000000032000000000000003200000000",
            INIT_6D => X"00000077000000000000006f0000000000000037000000000000000a00000000",
            INIT_6E => X"0000000e0000000000000076000000000000007a000000000000004e00000000",
            INIT_6F => X"0000000000000000000000400000000000000043000000000000000000000000",
            INIT_70 => X"000000000000000000000000000000000000001c000000000000001800000000",
            INIT_71 => X"0000001b00000000000000350000000000000066000000000000007800000000",
            INIT_72 => X"0000001a000000000000002e0000000000000031000000000000001f00000000",
            INIT_73 => X"0000000700000000000000110000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000001d000000000000001d0000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000004000000000000000800000000",
            INIT_78 => X"0000003c0000000000000000000000000000002e000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000200000000000000440000000000000000000000000000000300000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000007700000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000001800000000000000000000000000000000000000000000000500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE14;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE15 : if BRAM_NAME = "samplegold_layersamples_instance15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000001e000000000000005c000000000000000000000000",
            INIT_01 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000004100000000000000aa0000000000000000000000000000003900000000",
            INIT_03 => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_04 => X"00000000000000000000002c0000000000000015000000000000007300000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_06 => X"0000007b00000000000000300000000000000000000000000000000000000000",
            INIT_07 => X"0000002700000000000000000000000000000063000000000000000000000000",
            INIT_08 => X"00000022000000000000000c0000000000000024000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_0A => X"0000000000000000000000500000000000000022000000000000000000000000",
            INIT_0B => X"00000000000000000000001d0000000000000000000000000000002800000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_0D => X"0000006100000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000002f00000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000600000000000000350000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000170000000000000033000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000003400000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000026000000000000000000000000",
            INIT_1D => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_1F => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000005f00000000",
            INIT_21 => X"0000002800000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000280000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_2B => X"0000000000000000000000000000000000000024000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000006300000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000006500000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000400000000000000070000000000000000000000000000000e00000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000014500000000000000ef000000000000010a000000000000004400000000",
            INIT_3F => X"0000004500000000000000000000000000000000000000000000003900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005900000000000000610000000000000093000000000000003600000000",
            INIT_41 => X"00000000000000000000001a0000000000000045000000000000003900000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000260000000000000076000000000000005a00000000",
            INIT_44 => X"0000001300000000000000130000000000000039000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000003b00000000000000040000000000000000000000000000000000000000",
            INIT_48 => X"0000003f000000000000002c0000000000000065000000000000002300000000",
            INIT_49 => X"0000000000000000000000160000000000000028000000000000002c00000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000002400000000000000430000000000000000000000000000000000000000",
            INIT_4E => X"00000000000000000000006e000000000000003d000000000000000400000000",
            INIT_4F => X"0000000000000000000000000000000000000065000000000000000000000000",
            INIT_50 => X"0000001400000000000000560000000000000031000000000000000000000000",
            INIT_51 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"00000000000000000000007e0000000000000000000000000000000000000000",
            INIT_53 => X"00000000000000000000004c000000000000000a000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000004600000000",
            INIT_57 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"000000000000000000000000000000000000007900000000000000a200000000",
            INIT_59 => X"0000000000000000000000030000000000000000000000000000004400000000",
            INIT_5A => X"0000008400000000000000250000000000000010000000000000000900000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000005c00000000",
            INIT_5C => X"0000002100000000000000000000000000000039000000000000000000000000",
            INIT_5D => X"00000000000000000000001a0000000000000000000000000000002500000000",
            INIT_5E => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000032000000000000007700000000",
            INIT_60 => X"000000000000000000000000000000000000000c000000000000002700000000",
            INIT_61 => X"00000050000000000000004b0000000000000000000000000000000500000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_63 => X"0000000000000000000000000000000000000031000000000000002a00000000",
            INIT_64 => X"0000000000000000000000020000000000000000000000000000000700000000",
            INIT_65 => X"0000001300000000000000030000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000005000000000000001a00000000",
            INIT_67 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000005900000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"000000b000000000000000000000000000000015000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"000000010000000000000000000000000000003a000000000000000000000000",
            INIT_75 => X"0000001700000000000000000000000000000011000000000000000000000000",
            INIT_76 => X"00000000000000000000000000000000000000a3000000000000000d00000000",
            INIT_77 => X"0000001a000000000000002f0000000000000000000000000000000000000000",
            INIT_78 => X"00000021000000000000000d0000000000000028000000000000003300000000",
            INIT_79 => X"000000650000000000000016000000000000003c000000000000002300000000",
            INIT_7A => X"0000000000000000000000100000000000000026000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_7C => X"000000000000000000000000000000000000002c000000000000000000000000",
            INIT_7D => X"00000000000000000000001b0000000000000000000000000000000000000000",
            INIT_7E => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000090000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE15;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE16 : if BRAM_NAME = "samplegold_layersamples_instance16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000007c00000000000000080000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000006d00000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"00000000000000000000006b0000000000000006000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000063000000000000000500000000",
            INIT_08 => X"0000000000000000000000000000000000000030000000000000001300000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"00000000000000000000005e0000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000150000000000000012000000000000000000000000",
            INIT_0C => X"0000003500000000000000550000000000000000000000000000000000000000",
            INIT_0D => X"0000007c00000000000000190000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000003000000000000005d00000000",
            INIT_0F => X"0000000000000000000000540000000000000045000000000000000000000000",
            INIT_10 => X"0000002600000000000000000000000000000005000000000000003200000000",
            INIT_11 => X"00000023000000000000002e0000000000000037000000000000006f00000000",
            INIT_12 => X"0000002600000000000000000000000000000000000000000000005800000000",
            INIT_13 => X"0000008300000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000004700000000000000000000000000000007000000000000004600000000",
            INIT_15 => X"0000000a000000000000001e0000000000000000000000000000003000000000",
            INIT_16 => X"00000056000000000000007e000000000000006b000000000000001000000000",
            INIT_17 => X"0000000900000000000000000000000000000000000000000000004100000000",
            INIT_18 => X"0000000e0000000000000000000000000000001b000000000000005600000000",
            INIT_19 => X"0000001800000000000000020000000000000000000000000000004100000000",
            INIT_1A => X"0000002400000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000009000000000000003400000000",
            INIT_1C => X"000000010000000000000011000000000000000b000000000000005200000000",
            INIT_1D => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000003d00000000000000000000000000000029000000000000001500000000",
            INIT_20 => X"0000000000000000000000010000000000000000000000000000001000000000",
            INIT_21 => X"0000000000000000000000000000000000000006000000000000006c00000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000048000000000000000000000000",
            INIT_28 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_2B => X"000000070000000000000000000000000000000000000000000000b300000000",
            INIT_2C => X"0000000000000000000000180000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"000000000000000000000011000000000000003d000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_33 => X"0000000000000000000000680000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000270000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"00000000000000000000001b000000000000000000000000000000ac00000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000004400000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000088000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000003200000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000008f00000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000004400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000390000000000000000000000000000000000000000",
            INIT_42 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000019000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000034000000000000000000000000",
            INIT_49 => X"0000000e00000000000000080000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_4C => X"0000000000000000000000000000000000000009000000000000000600000000",
            INIT_4D => X"00000007000000000000000b0000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000050000000000000000000000000000001c000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000023000000000000000000000000",
            INIT_55 => X"0000000a000000000000000c0000000000000000000000000000000400000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000030000000000000000000000000000003e00000000",
            INIT_59 => X"0000000000000000000000000000000000000033000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_62 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000006f000000000000003c0000000000000000000000000000002900000000",
            INIT_64 => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"00000010000000000000004a0000000000000038000000000000002000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"000000c300000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"00000032000000000000005a0000000000000070000000000000006700000000",
            INIT_69 => X"0000005e00000000000000500000000000000034000000000000000200000000",
            INIT_6A => X"00000008000000000000002a0000000000000037000000000000005200000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000007000000000000001000000000",
            INIT_6F => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"000000000000000000000039000000000000000c000000000000000700000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000002f00000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_77 => X"00000042000000000000001c0000000000000000000000000000000000000000",
            INIT_78 => X"00000028000000000000000c0000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000700000000000000000000000000000000000000000000003d00000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"000000000000000000000000000000000000007e000000000000003f00000000",
            INIT_7E => X"0000000d00000000000000270000000000000047000000000000000600000000",
            INIT_7F => X"0000004500000000000000000000000000000000000000000000002100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE16;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE17 : if BRAM_NAME = "samplegold_layersamples_instance17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000000000003e000000000000005e00000000",
            INIT_01 => X"0000001300000000000000470000000000000039000000000000000000000000",
            INIT_02 => X"0000000000000000000000150000000000000020000000000000002400000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"00000000000000000000005d0000000000000086000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000028000000000000000000000000",
            INIT_06 => X"0000007a000000000000004d0000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000110000000000000068000000000000009500000000",
            INIT_08 => X"000000010000000000000031000000000000000e000000000000000000000000",
            INIT_09 => X"00000000000000000000000a0000000000000006000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000250000000000000028000000000000000e00000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_11 => X"000000b400000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"00000079000000000000007b000000000000008e000000000000006600000000",
            INIT_13 => X"0000004800000000000000620000000000000053000000000000005700000000",
            INIT_14 => X"00000042000000000000003d0000000000000033000000000000004c00000000",
            INIT_15 => X"0000004500000000000000950000000000000032000000000000005500000000",
            INIT_16 => X"0000004000000000000000570000000000000056000000000000005c00000000",
            INIT_17 => X"00000077000000000000003a000000000000004d000000000000004900000000",
            INIT_18 => X"000000460000000000000037000000000000002d000000000000000000000000",
            INIT_19 => X"00000030000000000000001c0000000000000072000000000000002800000000",
            INIT_1A => X"0000004f00000000000000310000000000000037000000000000003400000000",
            INIT_1B => X"0000000100000000000000910000000000000010000000000000001c00000000",
            INIT_1C => X"0000001e000000000000002a0000000000000034000000000000001200000000",
            INIT_1D => X"0000000000000000000000100000000000000000000000000000004400000000",
            INIT_1E => X"0000004f000000000000001f000000000000000d000000000000000500000000",
            INIT_1F => X"0000000e00000000000000560000000000000055000000000000005600000000",
            INIT_20 => X"000000250000000000000000000000000000000c000000000000000000000000",
            INIT_21 => X"0000000000000000000000020000000000000020000000000000001900000000",
            INIT_22 => X"0000006000000000000000520000000000000012000000000000000000000000",
            INIT_23 => X"00000004000000000000002a000000000000005f000000000000007300000000",
            INIT_24 => X"00000034000000000000005f0000000000000000000000000000004c00000000",
            INIT_25 => X"0000005a0000000000000071000000000000003b000000000000006e00000000",
            INIT_26 => X"0000006e00000000000000660000000000000081000000000000008100000000",
            INIT_27 => X"0000001400000000000000650000000000000044000000000000002d00000000",
            INIT_28 => X"0000005f000000000000005d0000000000000075000000000000002700000000",
            INIT_29 => X"000000a10000000000000094000000000000006f000000000000006200000000",
            INIT_2A => X"0000003a0000000000000087000000000000009c000000000000009c00000000",
            INIT_2B => X"000000260000000000000000000000000000002c000000000000001800000000",
            INIT_2C => X"0000009700000000000000870000000000000086000000000000008900000000",
            INIT_2D => X"00000094000000000000009b0000000000000099000000000000009700000000",
            INIT_2E => X"0000000700000000000000160000000000000074000000000000007500000000",
            INIT_2F => X"0000008f00000000000000510000000000000053000000000000001c00000000",
            INIT_30 => X"0000009b0000000000000092000000000000006d000000000000007800000000",
            INIT_31 => X"00000055000000000000007d000000000000008d000000000000009200000000",
            INIT_32 => X"0000003900000000000000340000000000000039000000000000006d00000000",
            INIT_33 => X"0000008b00000000000000a00000000000000009000000000000003000000000",
            INIT_34 => X"0000008a000000000000008f0000000000000093000000000000009700000000",
            INIT_35 => X"0000005600000000000000370000000000000065000000000000007b00000000",
            INIT_36 => X"000000330000000000000039000000000000004c000000000000004b00000000",
            INIT_37 => X"0000009800000000000000a20000000000000099000000000000001b00000000",
            INIT_38 => X"0000009d000000000000006a000000000000006a000000000000008400000000",
            INIT_39 => X"00000048000000000000004b000000000000002b000000000000006100000000",
            INIT_3A => X"0000003a00000000000000350000000000000042000000000000004900000000",
            INIT_3B => X"0000007900000000000000b5000000000000008b000000000000007800000000",
            INIT_3C => X"0000005800000000000000640000000000000060000000000000007c00000000",
            INIT_3D => X"0000004e0000000000000049000000000000004e000000000000004f00000000",
            INIT_3E => X"0000005800000000000000300000000000000042000000000000004b00000000",
            INIT_3F => X"0000005a00000000000000600000000000000066000000000000006600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000049000000000000004f000000000000004d000000000000004f00000000",
            INIT_41 => X"0000004400000000000000370000000000000046000000000000004c00000000",
            INIT_42 => X"0000003d00000000000000460000000000000038000000000000003800000000",
            INIT_43 => X"0000003e0000000000000040000000000000003d000000000000004300000000",
            INIT_44 => X"0000005b00000000000000330000000000000049000000000000004600000000",
            INIT_45 => X"000000390000000000000039000000000000003a000000000000003c00000000",
            INIT_46 => X"00000039000000000000002d000000000000002e000000000000003900000000",
            INIT_47 => X"000000450000000000000042000000000000003f000000000000003b00000000",
            INIT_48 => X"0000003800000000000000500000000000000018000000000000003a00000000",
            INIT_49 => X"0000003200000000000000340000000000000037000000000000003400000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000001100000000000000060000000000000006000000000000000900000000",
            INIT_4D => X"0000000000000000000000060000000000000012000000000000000200000000",
            INIT_4E => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000b000000000000000f0000000000000012000000000000000800000000",
            INIT_50 => X"0000000b00000000000000140000000000000000000000000000001400000000",
            INIT_51 => X"0000000000000000000000000000000000000011000000000000001b00000000",
            INIT_52 => X"00000014000000000000002b0000000000000010000000000000000a00000000",
            INIT_53 => X"000000050000000000000000000000000000000f000000000000002400000000",
            INIT_54 => X"0000002a00000000000000130000000000000002000000000000000000000000",
            INIT_55 => X"0000002a00000000000000000000000000000002000000000000001f00000000",
            INIT_56 => X"0000001f0000000000000032000000000000003e000000000000002c00000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_58 => X"0000002c00000000000000260000000000000000000000000000000000000000",
            INIT_59 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"00000000000000000000000b0000000000000048000000000000002700000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000004400000000000000230000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000003900000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000001c000000000000000d000000000000002a000000000000000700000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"000000220000000000000000000000000000000f000000000000001600000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000c00000000000000100000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE17;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE18 : if BRAM_NAME = "samplegold_layersamples_instance18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"000000000000000000000006000000000000000a000000000000000300000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_3C => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000005000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000230000000000000000000000000000000900000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_43 => X"0000000000000000000000230000000000000000000000000000001a00000000",
            INIT_44 => X"000000000000000000000000000000000000002e000000000000000000000000",
            INIT_45 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000200000000000000150000000000000002000000000000000000000000",
            INIT_48 => X"0000001c00000000000000000000000000000018000000000000001900000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_4A => X"0000000000000000000000000000000000000007000000000000000f00000000",
            INIT_4B => X"0000001600000000000000000000000000000029000000000000000000000000",
            INIT_4C => X"0000003700000000000000000000000000000000000000000000000700000000",
            INIT_4D => X"0000002200000000000000000000000000000022000000000000000000000000",
            INIT_4E => X"0000001400000000000000070000000000000031000000000000000000000000",
            INIT_4F => X"000000000000000000000024000000000000000b000000000000000600000000",
            INIT_50 => X"000000000000000000000079000000000000000b000000000000000f00000000",
            INIT_51 => X"0000000000000000000000040000000000000000000000000000001f00000000",
            INIT_52 => X"0000000000000000000000150000000000000003000000000000000e00000000",
            INIT_53 => X"0000000000000000000000000000000000000029000000000000001d00000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_58 => X"000000000000000000000000000000000000003c000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000001000000000000000040000000000000020000000000000001400000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"00000004000000000000000a0000000000000000000000000000000a00000000",
            INIT_5D => X"0000000d00000000000000120000000000000001000000000000000000000000",
            INIT_5E => X"0000000000000000000000120000000000000000000000000000000500000000",
            INIT_5F => X"0000000000000000000000080000000000000004000000000000000300000000",
            INIT_60 => X"0000000100000000000000060000000000000006000000000000000700000000",
            INIT_61 => X"00000001000000000000003b0000000000000006000000000000000500000000",
            INIT_62 => X"00000016000000000000000d0000000000000030000000000000000000000000",
            INIT_63 => X"000000320000000000000034000000000000001a000000000000002300000000",
            INIT_64 => X"0000001c00000000000000080000000000000037000000000000000700000000",
            INIT_65 => X"0000000e0000000000000000000000000000000c000000000000002600000000",
            INIT_66 => X"0000002f000000000000002f000000000000002d000000000000002800000000",
            INIT_67 => X"000000040000000000000013000000000000001f000000000000002400000000",
            INIT_68 => X"00000026000000000000001b0000000000000001000000000000001100000000",
            INIT_69 => X"0000002a00000000000000220000000000000023000000000000001a00000000",
            INIT_6A => X"0000001e00000000000000200000000000000018000000000000002a00000000",
            INIT_6B => X"0000002c000000000000001c0000000000000020000000000000002100000000",
            INIT_6C => X"0000002c000000000000002b0000000000000028000000000000002500000000",
            INIT_6D => X"00000021000000000000002d0000000000000018000000000000003600000000",
            INIT_6E => X"000000270000000000000025000000000000001f000000000000001c00000000",
            INIT_6F => X"0000003000000000000000320000000000000026000000000000002600000000",
            INIT_70 => X"0000002e0000000000000033000000000000002e000000000000003200000000",
            INIT_71 => X"0000001500000000000000250000000000000017000000000000001300000000",
            INIT_72 => X"000000af00000000000000350000000000000022000000000000002200000000",
            INIT_73 => X"000000e100000000000000ce00000000000000c7000000000000007a00000000",
            INIT_74 => X"000000e900000000000000f300000000000000ec00000000000000d600000000",
            INIT_75 => X"000000e600000000000000f100000000000000e700000000000000fc00000000",
            INIT_76 => X"0000008100000000000000b900000000000000e400000000000000fd00000000",
            INIT_77 => X"000000d700000000000000ea00000000000000d100000000000000cd00000000",
            INIT_78 => X"0000010400000000000000e500000000000000f200000000000000f000000000",
            INIT_79 => X"0000010300000000000000eb00000000000000f200000000000000a100000000",
            INIT_7A => X"000000c7000000000000007700000000000000bc00000000000000e500000000",
            INIT_7B => X"000000ef00000000000000d000000000000000ef00000000000000cd00000000",
            INIT_7C => X"0000009500000000000000cd00000000000000ca00000000000000cf00000000",
            INIT_7D => X"000000e500000000000000f300000000000000e900000000000000dc00000000",
            INIT_7E => X"000000c500000000000000cf000000000000006f00000000000000b400000000",
            INIT_7F => X"000000c400000000000000cb00000000000000c900000000000000dc00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE18;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE19 : if BRAM_NAME = "samplegold_layersamples_instance19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000060000000000000004a000000000000004d000000000000009400000000",
            INIT_01 => X"0000006200000000000000bd00000000000000de00000000000000a100000000",
            INIT_02 => X"0000008c0000000000000082000000000000006c000000000000004d00000000",
            INIT_03 => X"0000003e000000000000008c0000000000000081000000000000009000000000",
            INIT_04 => X"0000005d0000000000000020000000000000002f000000000000004400000000",
            INIT_05 => X"0000001f000000000000001b000000000000006b00000000000000a200000000",
            INIT_06 => X"0000004700000000000000500000000000000015000000000000004a00000000",
            INIT_07 => X"00000039000000000000003e000000000000004f000000000000005f00000000",
            INIT_08 => X"00000099000000000000008f0000000000000085000000000000002000000000",
            INIT_09 => X"00000025000000000000002a0000000000000040000000000000003400000000",
            INIT_0A => X"0000005d0000000000000055000000000000005d000000000000002f00000000",
            INIT_0B => X"0000007f000000000000005d000000000000004c000000000000004200000000",
            INIT_0C => X"000000100000000000000083000000000000009500000000000000b100000000",
            INIT_0D => X"0000006c000000000000004b0000000000000041000000000000003d00000000",
            INIT_0E => X"000000950000000000000094000000000000008f000000000000008500000000",
            INIT_0F => X"0000008d000000000000006d0000000000000095000000000000009100000000",
            INIT_10 => X"0000006500000000000000300000000000000031000000000000008d00000000",
            INIT_11 => X"0000009b00000000000000880000000000000058000000000000005900000000",
            INIT_12 => X"0000007600000000000000730000000000000083000000000000009000000000",
            INIT_13 => X"00000086000000000000008a0000000000000074000000000000006e00000000",
            INIT_14 => X"0000004c0000000000000028000000000000008a000000000000007c00000000",
            INIT_15 => X"000000780000000000000062000000000000007e000000000000007700000000",
            INIT_16 => X"0000008a00000000000000650000000000000092000000000000008c00000000",
            INIT_17 => X"00000055000000000000007b0000000000000098000000000000008d00000000",
            INIT_18 => X"0000007500000000000000680000000000000051000000000000002e00000000",
            INIT_19 => X"00000088000000000000006a0000000000000075000000000000006d00000000",
            INIT_1A => X"0000007300000000000000880000000000000025000000000000002a00000000",
            INIT_1B => X"0000001e000000000000000c0000000000000031000000000000005000000000",
            INIT_1C => X"0000001e0000000000000067000000000000005b000000000000005100000000",
            INIT_1D => X"0000002f0000000000000068000000000000006d000000000000002300000000",
            INIT_1E => X"0000000f000000000000002f0000000000000039000000000000002f00000000",
            INIT_1F => X"0000003f00000000000000000000000000000000000000000000000900000000",
            INIT_20 => X"0000002a00000000000000290000000000000043000000000000005200000000",
            INIT_21 => X"0000001f00000000000000200000000000000017000000000000002400000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000200000000000000040000000000000000000000000000000000000000",
            INIT_25 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000002000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000002e00000000000000000000000000000000000000000000000200000000",
            INIT_3F => X"0000000000000000000000000000000000000004000000000000000200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000570000000000000015000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_42 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_43 => X"00000014000000000000001d0000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000003f00000000",
            INIT_45 => X"00000046000000000000000f0000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000003d00000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000008e00000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"00000000000000000000003b0000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000005c00000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_55 => X"0000000000000000000000330000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000d00000000000000000000000000000016000000000000000a00000000",
            INIT_60 => X"00000010000000000000000e000000000000000b000000000000000800000000",
            INIT_61 => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_62 => X"0000000700000000000000060000000000000000000000000000000300000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_68 => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"000000090000000000000000000000000000000c000000000000000000000000",
            INIT_6C => X"0000001b000000000000003f0000000000000000000000000000000000000000",
            INIT_6D => X"000000000000000000000035000000000000007d000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_6F => X"000000000000000000000015000000000000000f000000000000000c00000000",
            INIT_70 => X"0000006300000000000000000000000000000000000000000000001400000000",
            INIT_71 => X"000000470000000000000156000000000000005f000000000000000500000000",
            INIT_72 => X"0000005b0000000000000009000000000000006d000000000000003100000000",
            INIT_73 => X"0000004200000000000000690000000000000069000000000000007b00000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000004c00000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"00000008000000000000000000000000000000ff000000000000000000000000",
            INIT_7A => X"0000002900000000000000000000000000000002000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"00000000000000000000000d0000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE19;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE20 : if BRAM_NAME = "samplegold_layersamples_instance20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000032000000000000004c00000000",
            INIT_01 => X"0000002d00000000000000170000000000000000000000000000000000000000",
            INIT_02 => X"0000000300000000000000030000000000000000000000000000001e00000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000004800000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"000000000000000000000000000000000000000b000000000000001200000000",
            INIT_08 => X"00000017000000000000000c0000000000000006000000000000000000000000",
            INIT_09 => X"0000004000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000400000000000000000000000000000000000000000000004300000000",
            INIT_0B => X"00000005000000000000001d0000000000000013000000000000005700000000",
            INIT_0C => X"000000030000000000000075000000000000000a000000000000000300000000",
            INIT_0D => X"0000004a00000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000001c00000000000000000000000000000000000000000000002d00000000",
            INIT_0F => X"0000000000000000000000090000000000000002000000000000000f00000000",
            INIT_10 => X"0000005400000000000000240000000000000054000000000000000100000000",
            INIT_11 => X"0000002700000000000000430000000000000016000000000000000300000000",
            INIT_12 => X"0000000800000000000000160000000000000004000000000000000000000000",
            INIT_13 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_14 => X"0000002400000000000000280000000000000045000000000000002800000000",
            INIT_15 => X"0000001400000000000000100000000000000011000000000000001100000000",
            INIT_16 => X"0000000000000000000000070000000000000000000000000000001900000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000003c00000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE20;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE21 : if BRAM_NAME = "samplegold_layersamples_instance21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000200000000000000070000000000000001000000000000000000000000",
            INIT_0E => X"0000000100000000000000030000000000000005000000000000000100000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"000000a500000000000000bd0000000000000000000000000000000000000000",
            INIT_11 => X"0000009e000000000000009a000000000000009b000000000000009d00000000",
            INIT_12 => X"0000000000000000000000670000000000000082000000000000008400000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000003f0000000000000063000000000000008b000000000000000b00000000",
            INIT_15 => X"0000003400000000000000320000000000000050000000000000007600000000",
            INIT_16 => X"0000000000000000000000000000000000000018000000000000002400000000",
            INIT_17 => X"0000004e00000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000006a0000000000000078000000000000007f00000000000000b300000000",
            INIT_19 => X"0000009c00000000000000b8000000000000008b000000000000008c00000000",
            INIT_1A => X"0000000000000000000000000000000000000039000000000000007f00000000",
            INIT_1B => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000a00000000000000010000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000010000000000000019000000000000002e00000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"00000011000000000000000a0000000000000018000000000000004e00000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000008400000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000001400000000000000250000000000000023000000000000002400000000",
            INIT_30 => X"00000000000000000000000a0000000000000022000000000000003c00000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"00000027000000000000003d0000000000000038000000000000000000000000",
            INIT_33 => X"0000001e00000000000000000000000000000000000000000000003600000000",
            INIT_34 => X"000000000000000000000000000000000000001c000000000000000400000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_37 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_38 => X"0000000900000000000000190000000000000000000000000000000000000000",
            INIT_39 => X"0000000400000000000000110000000000000021000000000000000100000000",
            INIT_3A => X"0000000400000000000000030000000000000003000000000000000000000000",
            INIT_3B => X"000000230000000000000021000000000000001d000000000000002200000000",
            INIT_3C => X"0000003200000000000000340000000000000037000000000000002700000000",
            INIT_3D => X"0000002900000000000000300000000000000044000000000000004600000000",
            INIT_3E => X"0000001b0000000000000025000000000000002c000000000000002f00000000",
            INIT_3F => X"0000001100000000000000100000000000000013000000000000001600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000019000000000000001f0000000000000000000000000000000200000000",
            INIT_41 => X"0000001e0000000000000015000000000000000e000000000000001800000000",
            INIT_42 => X"000000120000000000000014000000000000000d000000000000001900000000",
            INIT_43 => X"0000000000000000000000000000000000000003000000000000000800000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000002d00000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000009400000000000000b000000000000000b5000000000000005800000000",
            INIT_4A => X"000000630000000000000092000000000000009900000000000000a100000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000040000000000000001000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000480000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"000000b700000000000000fb0000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"000000dd00000000000000230000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000007100000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"000000c600000000000000170000000000000000000000000000000000000000",
            INIT_64 => X"00000000000000000000006200000000000000df000000000000012d00000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"00000000000000000000000c000000000000003f000000000000004d00000000",
            INIT_68 => X"00000149000000000000015e00000000000000f1000000000000004300000000",
            INIT_69 => X"000000000000000000000000000000000000003800000000000000cc00000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"000000de00000000000000c90000000000000000000000000000000000000000",
            INIT_6E => X"000000b20000000000000119000000000000010700000000000000f700000000",
            INIT_6F => X"0000003100000000000000a30000000000000088000000000000006700000000",
            INIT_70 => X"00000071000000000000004f000000000000000f000000000000005700000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000005d00000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"000000a300000000000000900000000000000074000000000000004800000000",
            INIT_74 => X"000000e100000000000000d800000000000000cc00000000000000bb00000000",
            INIT_75 => X"0000005400000000000000720000000000000080000000000000007200000000",
            INIT_76 => X"000000300000000000000033000000000000003e000000000000004500000000",
            INIT_77 => X"0000000000000000000000070000000000000010000000000000001800000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000190000000000000070000000000000000000000000",
            INIT_7D => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE21;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE22 : if BRAM_NAME = "samplegold_layersamples_instance22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_01 => X"0000003100000000000000560000000000000030000000000000000000000000",
            INIT_02 => X"00000041000000000000003c000000000000003c000000000000005b00000000",
            INIT_03 => X"0000000000000000000000000000000000000009000000000000007800000000",
            INIT_04 => X"0000003900000000000000000000000000000000000000000000001400000000",
            INIT_05 => X"0000003e0000000000000005000000000000000d000000000000000000000000",
            INIT_06 => X"0000003400000000000000020000000000000000000000000000000100000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000003a00000000",
            INIT_08 => X"0000000700000000000000120000000000000000000000000000000000000000",
            INIT_09 => X"0000001100000000000000100000000000000000000000000000000b00000000",
            INIT_0A => X"0000006a00000000000000000000000000000002000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000002400000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000019000000000000008400000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000075000000000000009600000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"00000026000000000000006d000000000000006f000000000000005800000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000001d00000000000000080000000000000000000000000000000000000000",
            INIT_20 => X"000000890000000000000000000000000000000b000000000000001000000000",
            INIT_21 => X"000000000000000000000032000000000000006f000000000000006600000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_23 => X"0000004a00000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000003f00000000000000000000000000000000000000000000003c00000000",
            INIT_26 => X"00000032000000000000001f0000000000000019000000000000001800000000",
            INIT_27 => X"0000000000000000000000510000000000000022000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_29 => X"0000000000000000000000060000000000000007000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000001700000000000000000000000000000026000000000000000a00000000",
            INIT_2C => X"0000000f00000000000000260000000000000025000000000000001300000000",
            INIT_2D => X"0000000000000000000000040000000000000005000000000000003200000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_30 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_35 => X"0000002500000000000000230000000000000024000000000000000000000000",
            INIT_36 => X"0000004a000000000000004d0000000000000048000000000000003900000000",
            INIT_37 => X"00000033000000000000004c0000000000000048000000000000005b00000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000110000000000000034000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000058000000000000000f0000000000000000000000000000000000000000",
            INIT_41 => X"00000054000000000000002b0000000000000058000000000000004b00000000",
            INIT_42 => X"0000005e00000000000000810000000000000084000000000000007900000000",
            INIT_43 => X"0000000000000000000000040000000000000006000000000000007700000000",
            INIT_44 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000210000000000000034000000000000001800000000",
            INIT_46 => X"0000000000000000000000120000000000000027000000000000001e00000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"000000b500000000000000640000000000000000000000000000000800000000",
            INIT_4C => X"000000030000000000000000000000000000000000000000000000a900000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000018000000000000002b00000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"000000000000000000000051000000000000007c000000000000000e00000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000002d00000000000000060000000000000000000000000000000000000000",
            INIT_58 => X"000000ed000000000000004c0000000000000000000000000000000300000000",
            INIT_59 => X"000000000000000000000000000000000000000000000000000000c800000000",
            INIT_5A => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_5B => X"000000e700000000000000050000000000000033000000000000003e00000000",
            INIT_5C => X"00000008000000000000006a0000000000000000000000000000007e00000000",
            INIT_5D => X"000000370000000000000021000000000000004400000000000000b600000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"000000000000000000000000000000000000001b000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000007b00000000000000730000000000000000000000000000000000000000",
            INIT_66 => X"0000005600000000000000530000000000000060000000000000006e00000000",
            INIT_67 => X"0000001b00000000000000230000000000000036000000000000004000000000",
            INIT_68 => X"00000026000000000000000d0000000000000004000000000000001a00000000",
            INIT_69 => X"000000120000000000000010000000000000000b000000000000003800000000",
            INIT_6A => X"0000001500000000000000290000000000000011000000000000000b00000000",
            INIT_6B => X"0000000000000000000000210000000000000026000000000000001900000000",
            INIT_6C => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000250000000000000000000000000000000000000000",
            INIT_72 => X"000000100000000000000000000000000000001f000000000000001000000000",
            INIT_73 => X"0000000000000000000000000000000000000016000000000000001200000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE22;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE23 : if BRAM_NAME = "samplegold_layersamples_instance23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000000000004f000000000000000500000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"00000000000000000000000c000000000000002b000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000059000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000001f000000000000000b0000000000000000000000000000009800000000",
            INIT_0D => X"0000000000000000000000000000000000000030000000000000004f00000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"000000f100000000000000010000000000000000000000000000000000000000",
            INIT_10 => X"0000000b00000000000000000000000000000000000000000000001f00000000",
            INIT_11 => X"0000005a0000000000000060000000000000000f000000000000002c00000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"000000bf00000000000000b1000000000000009a000000000000000000000000",
            INIT_17 => X"000000ac00000000000000b200000000000000c000000000000000ba00000000",
            INIT_18 => X"0000005c00000000000000340000000000000068000000000000007c00000000",
            INIT_19 => X"0000001f00000000000000250000000000000060000000000000003300000000",
            INIT_1A => X"0000001e00000000000000000000000000000000000000000000000a00000000",
            INIT_1B => X"0000004200000000000000340000000000000022000000000000001f00000000",
            INIT_1C => X"0000005b00000000000000680000000000000056000000000000005900000000",
            INIT_1D => X"0000002000000000000000640000000000000077000000000000006100000000",
            INIT_1E => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_21 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"000000140000000000000000000000000000000000000000000000c200000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000002400000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000002000000000000000e00000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"000000000000000000000000000000000000002c000000000000002400000000",
            INIT_32 => X"0000001e00000000000000000000000000000000000000000000001100000000",
            INIT_33 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"000000000000000000000000000000000000005c000000000000002e00000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000000000000000000000000000000000000db000000000000000c00000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000118000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"000000000000000000000000000000000000000000000000000000ff00000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000005200000000000000410000000000000000000000000000000000000000",
            INIT_4C => X"000000580000000000000000000000000000000c00000000000000db00000000",
            INIT_4D => X"00000000000000000000002d000000000000003e000000000000003900000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_58 => X"0000000900000000000000010000000000000010000000000000000900000000",
            INIT_59 => X"0000001f00000000000000000000000000000000000000000000000700000000",
            INIT_5A => X"0000000f0000000000000006000000000000000b000000000000000a00000000",
            INIT_5B => X"0000001700000000000000030000000000000015000000000000000700000000",
            INIT_5C => X"0000000000000000000000160000000000000011000000000000001500000000",
            INIT_5D => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000001a00000000000000340000000000000000000000000000000000000000",
            INIT_63 => X"000000360000000000000031000000000000002c000000000000002000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000003900000000",
            INIT_65 => X"0000005400000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000001700000000000000150000000000000005000000000000001200000000",
            INIT_67 => X"0000000d000000000000000e000000000000000b000000000000001f00000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000002900000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000005a00000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"000000000000000000000000000000000000003400000000000000f900000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"00000000000000000000000000000000000000d1000000000000007c00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000009f000000000000011d0000000000000084000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE23;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE24 : if BRAM_NAME = "samplegold_layersamples_instance24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001300000000000000020000000000000000000000000000000000000000",
            INIT_01 => X"0000004000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000910000000000000131000000000000011400000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"000000e400000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000011a0000000000000113000000000000010e000000000000010300000000",
            INIT_08 => X"0000009400000000000000c8000000000000012f000000000000014900000000",
            INIT_09 => X"0000005000000000000000b6000000000000009500000000000000c300000000",
            INIT_0A => X"0000000a0000000000000000000000000000006e000000000000004500000000",
            INIT_0B => X"000000540000000000000044000000000000003e000000000000001900000000",
            INIT_0C => X"0000007500000000000000610000000000000050000000000000005c00000000",
            INIT_0D => X"0000007c00000000000000840000000000000076000000000000007500000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000006700000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000005700000000000000040000000000000000000000000000000000000000",
            INIT_16 => X"0000004c000000000000004d000000000000007b000000000000007500000000",
            INIT_17 => X"00000054000000000000004a000000000000005b000000000000005a00000000",
            INIT_18 => X"0000004400000000000000510000000000000056000000000000005200000000",
            INIT_19 => X"000000800000000000000067000000000000004b000000000000004d00000000",
            INIT_1A => X"000000000000000000000000000000000000000b000000000000007b00000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000004f00000000000000520000000000000000000000000000000000000000",
            INIT_1D => X"0000007500000000000000850000000000000065000000000000004e00000000",
            INIT_1E => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_1F => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_20 => X"00000055000000000000005a000000000000002d000000000000000000000000",
            INIT_21 => X"0000000000000000000000740000000000000083000000000000007000000000",
            INIT_22 => X"0000000000000000000000020000000000000003000000000000000000000000",
            INIT_23 => X"0000001d00000000000000000000000000000008000000000000000200000000",
            INIT_24 => X"00000081000000000000005e000000000000005c000000000000000000000000",
            INIT_25 => X"0000005900000000000000780000000000000077000000000000008300000000",
            INIT_26 => X"0000005700000000000000540000000000000057000000000000005500000000",
            INIT_27 => X"0000005c0000000000000040000000000000004a000000000000005500000000",
            INIT_28 => X"0000007700000000000000720000000000000067000000000000006900000000",
            INIT_29 => X"0000007200000000000000790000000000000074000000000000005400000000",
            INIT_2A => X"0000006f000000000000006f000000000000006d000000000000006c00000000",
            INIT_2B => X"00000065000000000000006a0000000000000069000000000000006700000000",
            INIT_2C => X"0000008200000000000000970000000000000063000000000000006600000000",
            INIT_2D => X"00000068000000000000005c000000000000000f000000000000000700000000",
            INIT_2E => X"00000061000000000000006a0000000000000068000000000000006c00000000",
            INIT_2F => X"0000005f00000000000000630000000000000065000000000000006600000000",
            INIT_30 => X"0000008e00000000000000630000000000000075000000000000005f00000000",
            INIT_31 => X"00000059000000000000001c0000000000000000000000000000002800000000",
            INIT_32 => X"00000063000000000000005c000000000000005e000000000000006100000000",
            INIT_33 => X"00000059000000000000006c000000000000006a000000000000006900000000",
            INIT_34 => X"0000007b00000000000000520000000000000058000000000000005b00000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_36 => X"000000670000000000000068000000000000004e000000000000003800000000",
            INIT_37 => X"0000004c00000000000000510000000000000069000000000000006500000000",
            INIT_38 => X"0000000000000000000000620000000000000063000000000000005400000000",
            INIT_39 => X"00000018000000000000000f0000000000000002000000000000000000000000",
            INIT_3A => X"0000003900000000000000050000000000000000000000000000000000000000",
            INIT_3B => X"000000530000000000000052000000000000004e000000000000005f00000000",
            INIT_3C => X"0000005100000000000000960000000000000054000000000000007a00000000",
            INIT_3D => X"0000006400000000000000420000000000000069000000000000000d00000000",
            INIT_3E => X"0000004c000000000000004d000000000000002a000000000000005300000000",
            INIT_3F => X"0000001a000000000000001e0000000000000023000000000000001700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003100000000000000260000000000000023000000000000001400000000",
            INIT_41 => X"00000053000000000000004d000000000000004f000000000000004700000000",
            INIT_42 => X"0000002c00000000000000540000000000000060000000000000006300000000",
            INIT_43 => X"0000002c0000000000000033000000000000003f000000000000003c00000000",
            INIT_44 => X"00000036000000000000002c000000000000002d000000000000002d00000000",
            INIT_45 => X"000000280000000000000028000000000000002e000000000000002b00000000",
            INIT_46 => X"0000000a00000000000000050000000000000024000000000000002f00000000",
            INIT_47 => X"0000000800000000000000030000000000000004000000000000001100000000",
            INIT_48 => X"0000000500000000000000070000000000000003000000000000000800000000",
            INIT_49 => X"0000000900000000000000070000000000000006000000000000000100000000",
            INIT_4A => X"0000000d00000000000000090000000000000000000000000000001800000000",
            INIT_4B => X"00000012000000000000000e0000000000000003000000000000000600000000",
            INIT_4C => X"00000007000000000000000e000000000000000f000000000000000400000000",
            INIT_4D => X"0000003800000000000000360000000000000006000000000000000000000000",
            INIT_4E => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000010000000000000000000000000000000100000000",
            INIT_51 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_52 => X"0000007300000000000000520000000000000000000000000000000000000000",
            INIT_53 => X"0000006600000000000000660000000000000065000000000000006700000000",
            INIT_54 => X"0000000c00000000000000390000000000000056000000000000006100000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000005600000000000000560000000000000029000000000000000000000000",
            INIT_57 => X"0000004c0000000000000042000000000000005a000000000000006200000000",
            INIT_58 => X"0000000000000000000000230000000000000038000000000000004200000000",
            INIT_59 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000003c000000000000003b0000000000000049000000000000005100000000",
            INIT_5B => X"000000600000000000000057000000000000004b000000000000005700000000",
            INIT_5C => X"0000000000000000000000000000000000000025000000000000005d00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_69 => X"000000000000000000000000000000000000001e000000000000001900000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_6D => X"0000000000000000000000320000000000000026000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000020000000000000000000000000000000200000000",
            INIT_71 => X"0000003300000000000000250000000000000012000000000000000900000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_73 => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_74 => X"0000003b00000000000000000000000000000008000000000000000000000000",
            INIT_75 => X"00000002000000000000002f0000000000000009000000000000002900000000",
            INIT_76 => X"0000001e00000000000000180000000000000023000000000000002c00000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000001700000000000000110000000000000010000000000000001300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE24;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE25 : if BRAM_NAME = "samplegold_layersamples_instance25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001300000000000000170000000000000011000000000000001300000000",
            INIT_01 => X"0000001500000000000000150000000000000014000000000000001600000000",
            INIT_02 => X"00000015000000000000001a0000000000000000000000000000000c00000000",
            INIT_03 => X"0000001e00000000000000160000000000000017000000000000001300000000",
            INIT_04 => X"0000001c00000000000000220000000000000021000000000000001f00000000",
            INIT_05 => X"0000000000000000000000080000000000000019000000000000001a00000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"000000000000000000000000000000000000000a000000000000004d00000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000006a000000000000006c0000000000000007000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000140000000000000006000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000150000000000000000000000000000000e00000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_5D => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_61 => X"0000000700000000000000090000000000000000000000000000000000000000",
            INIT_62 => X"00000000000000000000001a0000000000000009000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000300000000000000000000000000000000000000000000000b00000000",
            INIT_65 => X"00000000000000000000001d0000000000000000000000000000000000000000",
            INIT_66 => X"00000006000000000000001c0000000000000000000000000000000e00000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000001100000000000000080000000000000000000000000000000000000000",
            INIT_70 => X"0000001700000000000000180000000000000020000000000000000d00000000",
            INIT_71 => X"0000002700000000000000250000000000000029000000000000001a00000000",
            INIT_72 => X"0000004c00000000000000280000000000000020000000000000002800000000",
            INIT_73 => X"0000001f000000000000001c0000000000000017000000000000000000000000",
            INIT_74 => X"0000001f000000000000001b000000000000001b000000000000002100000000",
            INIT_75 => X"0000002b00000000000000240000000000000024000000000000002500000000",
            INIT_76 => X"00000096000000000000006b0000000000000072000000000000003000000000",
            INIT_77 => X"000000960000000000000097000000000000009c00000000000000b200000000",
            INIT_78 => X"0000009f000000000000009c00000000000000a800000000000000a900000000",
            INIT_79 => X"000000a300000000000000a300000000000000aa00000000000000a100000000",
            INIT_7A => X"000000b4000000000000009900000000000000c300000000000000c400000000",
            INIT_7B => X"0000009c00000000000000a7000000000000009c00000000000000bb00000000",
            INIT_7C => X"000000a900000000000000a8000000000000009c000000000000009d00000000",
            INIT_7D => X"000000c700000000000000c0000000000000008e00000000000000a400000000",
            INIT_7E => X"000000c900000000000000ad000000000000009600000000000000c600000000",
            INIT_7F => X"0000008d0000000000000092000000000000009d000000000000007500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE25;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE26 : if BRAM_NAME = "samplegold_layersamples_instance26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a300000000000000ae0000000000000099000000000000008800000000",
            INIT_01 => X"000000c800000000000000cd00000000000000b900000000000000a500000000",
            INIT_02 => X"0000008400000000000000c100000000000000a8000000000000009800000000",
            INIT_03 => X"0000009a000000000000008c000000000000008e000000000000008900000000",
            INIT_04 => X"000000a8000000000000009800000000000000a1000000000000009400000000",
            INIT_05 => X"000000a700000000000000c100000000000000c3000000000000009200000000",
            INIT_06 => X"0000009600000000000000b400000000000000a800000000000000ab00000000",
            INIT_07 => X"000000a1000000000000009b000000000000008c000000000000009400000000",
            INIT_08 => X"000000bd00000000000000a1000000000000009a000000000000009700000000",
            INIT_09 => X"000000c000000000000000b800000000000000be00000000000000c100000000",
            INIT_0A => X"000000a200000000000000a8000000000000009f00000000000000a000000000",
            INIT_0B => X"000000a900000000000000ab00000000000000b100000000000000aa00000000",
            INIT_0C => X"000000be00000000000000bf00000000000000b800000000000000ab00000000",
            INIT_0D => X"00000081000000000000009800000000000000bf00000000000000be00000000",
            INIT_0E => X"000000be00000000000000ac000000000000008d000000000000008700000000",
            INIT_0F => X"000000be00000000000000c200000000000000c300000000000000c600000000",
            INIT_10 => X"000000c200000000000000c500000000000000c100000000000000c100000000",
            INIT_11 => X"0000007c00000000000000b000000000000000ca00000000000000c900000000",
            INIT_12 => X"000000c300000000000000a6000000000000007c000000000000005000000000",
            INIT_13 => X"000000bd00000000000000be00000000000000c100000000000000ca00000000",
            INIT_14 => X"000000d300000000000000ba00000000000000bc00000000000000be00000000",
            INIT_15 => X"0000005f00000000000000c400000000000000d200000000000000d400000000",
            INIT_16 => X"0000009f0000000000000088000000000000004e000000000000002a00000000",
            INIT_17 => X"000000c100000000000000c000000000000000ab00000000000000af00000000",
            INIT_18 => X"000000d400000000000000d600000000000000ba00000000000000be00000000",
            INIT_19 => X"00000006000000000000004b00000000000000ec00000000000000d300000000",
            INIT_1A => X"00000046000000000000002e000000000000001b000000000000001200000000",
            INIT_1B => X"000000aa000000000000009d0000000000000096000000000000005900000000",
            INIT_1C => X"000000d000000000000000ce00000000000000cb00000000000000b800000000",
            INIT_1D => X"0000000d0000000000000031000000000000004900000000000000b600000000",
            INIT_1E => X"0000002b00000000000000150000000000000066000000000000002600000000",
            INIT_1F => X"000000b50000000000000099000000000000005f000000000000001c00000000",
            INIT_20 => X"000000af00000000000000b400000000000000ba00000000000000b200000000",
            INIT_21 => X"00000094000000000000007f000000000000008f00000000000000aa00000000",
            INIT_22 => X"0000008b00000000000000940000000000000088000000000000009f00000000",
            INIT_23 => X"00000042000000000000009c000000000000009a000000000000009a00000000",
            INIT_24 => X"0000003b000000000000003c0000000000000043000000000000004400000000",
            INIT_25 => X"0000004b00000000000000430000000000000032000000000000003300000000",
            INIT_26 => X"0000004a00000000000000460000000000000044000000000000004400000000",
            INIT_27 => X"000000200000000000000015000000000000003e000000000000004e00000000",
            INIT_28 => X"0000000900000000000000120000000000000011000000000000001c00000000",
            INIT_29 => X"00000000000000000000000c0000000000000009000000000000000900000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000200000000000000000000000000000000000000000000000100000000",
            INIT_2D => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_2E => X"00000044000000000000002b0000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000002e00000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000001600000000000000000000000000000018000000000000000000000000",
            INIT_39 => X"000000000000000000000000000000000000001f000000000000001700000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000003e000000000000000f0000000000000000000000000000000000000000",
            INIT_56 => X"00000000000000000000006f00000000000000c5000000000000006600000000",
            INIT_57 => X"0000000e00000000000000d4000000000000003f000000000000009800000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"000000000000000000000000000000000000006b000000000000000000000000",
            INIT_64 => X"0000001c00000000000000000000000000000008000000000000000000000000",
            INIT_65 => X"0000001700000000000000070000000000000018000000000000001400000000",
            INIT_66 => X"0000009c00000000000000070000000000000005000000000000000b00000000",
            INIT_67 => X"0000000000000000000000000000000000000025000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_6C => X"0000004500000000000000320000000000000057000000000000005f00000000",
            INIT_6D => X"0000003b00000000000000410000000000000044000000000000003900000000",
            INIT_6E => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_7A => X"0000000700000000000000010000000000000000000000000000001100000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"000000f300000000000000990000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE26;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE27 : if BRAM_NAME = "samplegold_layersamples_instance27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000250000000000000000000000000000000000000000",
            INIT_02 => X"000000ea00000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"000000000000000000000000000000000000000000000000000000a800000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"000000000000000000000000000000000000002b000000000000000000000000",
            INIT_06 => X"00000038000000000000000c0000000000000000000000000000000000000000",
            INIT_07 => X"00000009000000000000003800000000000000d3000000000000010600000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000003100000000",
            INIT_0A => X"00000000000000000000002e0000000000000042000000000000000000000000",
            INIT_0B => X"0000011700000000000000f60000000000000044000000000000000000000000",
            INIT_0C => X"0000003a0000000000000000000000000000003000000000000000b800000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_0F => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000006500000000000000ac0000000000000000000000000000000000000000",
            INIT_11 => X"0000008c0000000000000084000000000000007c000000000000006e00000000",
            INIT_12 => X"0000001c000000000000005b0000000000000026000000000000003600000000",
            INIT_13 => X"000000390000000000000000000000000000001f000000000000002d00000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000004700000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000003d00000000000000410000000000000021000000000000000d00000000",
            INIT_17 => X"000000590000000000000054000000000000005e000000000000005500000000",
            INIT_18 => X"00000026000000000000003a0000000000000038000000000000000000000000",
            INIT_19 => X"0000001700000000000000190000000000000017000000000000001800000000",
            INIT_1A => X"0000000000000000000000050000000000000000000000000000001400000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000001100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE27;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE28 : if BRAM_NAME = "samplegold_layersamples_instance28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000140000000000000000000000000000000100000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000270000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"000000000000000000000000000000000000002d000000000000000000000000",
            INIT_27 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"000000100000000000000021000000000000000a000000000000002000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_2B => X"0000001300000000000000080000000000000011000000000000000000000000",
            INIT_2C => X"000000170000000000000020000000000000001c000000000000001600000000",
            INIT_2D => X"0000000d0000000000000000000000000000000c000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"000000200000000000000003000000000000002d000000000000000000000000",
            INIT_30 => X"00000000000000000000001f000000000000002a000000000000001300000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000002e00000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000001c000000000000000b0000000000000013000000000000000000000000",
            INIT_34 => X"0000003500000000000000190000000000000019000000000000001800000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000002e000000000000001a000000000000000c000000000000000000000000",
            INIT_38 => X"0000000000000000000000130000000000000033000000000000002900000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"00000023000000000000002d000000000000001a000000000000002700000000",
            INIT_3C => X"0000000000000000000000000000000000000002000000000000002300000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000003f0000000000000018000000000000002e000000000000000a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000002e00000000000000270000000000000018000000000000001700000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_4A => X"0000000000000000000000160000000000000012000000000000000000000000",
            INIT_4B => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"000000000000000000000017000000000000001b000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000005100000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000100000000000000000000000000000002000000000",
            INIT_51 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"000000000000000000000000000000000000004c000000000000000e00000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000002e00000000000000000000000000000000000000000000001b00000000",
            INIT_5B => X"0000000000000000000000000000000000000010000000000000001300000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_60 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000003000000000000000000000000000000000000000000000004500000000",
            INIT_67 => X"0000000000000000000000000000000000000048000000000000001700000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"00000000000000000000004a000000000000004a000000000000000000000000",
            INIT_6A => X"0000000400000000000000110000000000000041000000000000000000000000",
            INIT_6B => X"000000000000000000000000000000000000006a000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000003b00000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"00000000000000000000007600000000000000a0000000000000000000000000",
            INIT_76 => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000063000000000000009300000000",
            INIT_78 => X"0000000400000000000000220000000000000000000000000000000000000000",
            INIT_79 => X"00000000000000000000008200000000000000e0000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000001900000000000000000000000000000010000000000000000000000000",
            INIT_7C => X"0000000200000000000000000000000000000000000000000000006200000000",
            INIT_7D => X"000000000000000000000063000000000000007e000000000000000000000000",
            INIT_7E => X"0000003900000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000085000000000000004600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE28;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE29 : if BRAM_NAME = "samplegold_layersamples_instance29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000007100000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000001a0000000000000000000000000000003f000000000000000000000000",
            INIT_03 => X"0000003a000000000000000000000000000000be000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000380000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000060000000000000000000000000000005300000000",
            INIT_07 => X"000000000000000000000026000000000000000000000000000000d300000000",
            INIT_08 => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000042000000000000000000000000",
            INIT_0A => X"000000cd00000000000000000000000000000000000000000000002400000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000004100000000000000000000000000000000000000000000002100000000",
            INIT_0D => X"0000005000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000630000000000000000000000000000000000000000",
            INIT_0F => X"0000005900000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000830000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000067000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000073000000000000000000000000",
            INIT_13 => X"00000000000000000000006d0000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000009400000000",
            INIT_17 => X"0000000000000000000000440000000000000026000000000000000000000000",
            INIT_18 => X"000000000000000000000007000000000000001a000000000000000000000000",
            INIT_19 => X"000000240000000000000028000000000000001f000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000016000000000000001f00000000",
            INIT_1C => X"0000000000000000000000040000000000000029000000000000000c00000000",
            INIT_1D => X"0000000000000000000000400000000000000004000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000400000000000000000000000000000000000000000",
            INIT_20 => X"000000000000000000000000000000000000000a000000000000003600000000",
            INIT_21 => X"0000000b0000000000000000000000000000002d000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000002700000000000000490000000000000000000000000000000300000000",
            INIT_24 => X"0000000f00000000000000000000000000000007000000000000000100000000",
            INIT_25 => X"0000003900000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000025000000000000000000000000",
            INIT_27 => X"00000000000000000000005f0000000000000000000000000000000500000000",
            INIT_28 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_29 => X"0000000700000000000000000000000000000019000000000000000000000000",
            INIT_2A => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_2B => X"000000030000000000000000000000000000001c000000000000001d00000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000007a00000000000000190000000000000000000000000000004a00000000",
            INIT_2E => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"00000000000000000000008f0000000000000000000000000000000000000000",
            INIT_30 => X"0000008f00000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000008e00000000000000770000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000600000000000000080000000000000047000000000000000000000000",
            INIT_34 => X"00000012000000000000004a0000000000000000000000000000000000000000",
            INIT_35 => X"0000008d00000000000000a50000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000150000000000000015000000000000000000000000",
            INIT_38 => X"0000000000000000000000550000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_3C => X"00000000000000000000000f0000000000000025000000000000003000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000022000000000000001900000000",
            INIT_3F => X"000000000000000000000000000000000000000b000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000260000000000000000000000000000000000000000",
            INIT_42 => X"0000001200000000000000160000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_44 => X"000000000000000000000002000000000000001f000000000000001f00000000",
            INIT_45 => X"0000005100000000000000000000000000000000000000000000003b00000000",
            INIT_46 => X"00000000000000000000000d0000000000000000000000000000004200000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_49 => X"000000000000000000000018000000000000003a000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000001d000000000000000e0000000000000006000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_4F => X"0000001000000000000000030000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000000000000000000000000000000000003b000000000000003c00000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_53 => X"0000000000000000000000100000000000000010000000000000001200000000",
            INIT_54 => X"000000000000000000000023000000000000005f000000000000000000000000",
            INIT_55 => X"00000000000000000000004e000000000000002c000000000000000000000000",
            INIT_56 => X"00000000000000000000003a0000000000000000000000000000000000000000",
            INIT_57 => X"00000018000000000000000a0000000000000000000000000000000000000000",
            INIT_58 => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000001200000000000000000000000000000012000000000000005900000000",
            INIT_5A => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000003100000000000000000000000000000000000000000000000600000000",
            INIT_5C => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_5D => X"0000003300000000000000000000000000000000000000000000001c00000000",
            INIT_5E => X"0000000000000000000000000000000000000008000000000000004b00000000",
            INIT_5F => X"0000002b0000000000000000000000000000002d000000000000000000000000",
            INIT_60 => X"0000000400000000000000230000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000150000000000000005000000000000001e00000000",
            INIT_62 => X"0000002000000000000000000000000000000000000000000000003800000000",
            INIT_63 => X"0000000000000000000000000000000000000044000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_65 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_66 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_69 => X"0000004d00000000000000000000000000000000000000000000004600000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_6B => X"000000000000000000000028000000000000001f000000000000002200000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000004400000000000000000000000000000000000000000000005700000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000001000000000000003e00000000",
            INIT_70 => X"000000000000000000000080000000000000004b000000000000002800000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"00000000000000000000000f0000000000000000000000000000007500000000",
            INIT_73 => X"0000000000000000000000280000000000000000000000000000002400000000",
            INIT_74 => X"000000000000000000000000000000000000000000000000000000a800000000",
            INIT_75 => X"0000006600000000000000000000000000000034000000000000000000000000",
            INIT_76 => X"0000000a00000000000000000000000000000015000000000000000500000000",
            INIT_77 => X"0000003700000000000000000000000000000040000000000000000000000000",
            INIT_78 => X"00000000000000000000002e0000000000000023000000000000000000000000",
            INIT_79 => X"000000000000000000000040000000000000002b000000000000000000000000",
            INIT_7A => X"000000780000000000000000000000000000003a000000000000000000000000",
            INIT_7B => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_7C => X"000000080000000000000000000000000000003b000000000000000000000000",
            INIT_7D => X"0000003300000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000007000000000",
            INIT_7F => X"000000b100000000000000000000000000000022000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE29;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE30 : if BRAM_NAME = "samplegold_layersamples_instance30" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003900000000000000130000000000000000000000000000002500000000",
            INIT_01 => X"0000000000000000000000740000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_03 => X"0000006f00000000000000de0000000000000000000000000000000800000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000003300000000000000000000000000000013000000000000000000000000",
            INIT_07 => X"00000000000000000000000000000000000000bc000000000000000000000000",
            INIT_08 => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000280000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000007000000000",
            INIT_0C => X"0000000000000000000000390000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"000000c200000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"00000010000000000000003f0000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"000000000000000000000000000000000000008b000000000000001f00000000",
            INIT_13 => X"000000230000000000000000000000000000000b000000000000004600000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000003000000000",
            INIT_15 => X"0000004600000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"00000000000000000000008d0000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_18 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"000000000000000000000000000000000000002f000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000021000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000003800000000",
            INIT_1F => X"000000b300000000000000160000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_21 => X"0000003700000000000000000000000000000002000000000000003600000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000003600000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"000000d9000000000000001f0000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000760000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"00000006000000000000000f0000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000003000000000000008c00000000",
            INIT_29 => X"0000000b000000000000001f0000000000000031000000000000000000000000",
            INIT_2A => X"000000320000000000000000000000000000007a000000000000000100000000",
            INIT_2B => X"0000006f00000000000000000000000000000009000000000000000000000000",
            INIT_2C => X"000000110000000000000000000000000000010c000000000000000000000000",
            INIT_2D => X"0000000300000000000000180000000000000010000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000007000000000",
            INIT_2F => X"00000000000000000000006a0000000000000000000000000000002f00000000",
            INIT_30 => X"0000002f0000000000000046000000000000000000000000000000f100000000",
            INIT_31 => X"0000005b00000000000000000000000000000014000000000000001b00000000",
            INIT_32 => X"0000000000000000000000260000000000000000000000000000000000000000",
            INIT_33 => X"0000009c0000000000000000000000000000000c000000000000003c00000000",
            INIT_34 => X"0000000000000000000000490000000000000049000000000000000c00000000",
            INIT_35 => X"000000000000000000000000000000000000005b000000000000002b00000000",
            INIT_36 => X"0000005900000000000000000000000000000037000000000000005d00000000",
            INIT_37 => X"0000000d00000000000000490000000000000000000000000000000000000000",
            INIT_38 => X"000000ac0000000000000000000000000000003f00000000000000bc00000000",
            INIT_39 => X"000000a200000000000000090000000000000000000000000000001000000000",
            INIT_3A => X"0000003a00000000000000000000000000000008000000000000000000000000",
            INIT_3B => X"000000fc000000000000000e0000000000000025000000000000000000000000",
            INIT_3C => X"000000ad00000000000000000000000000000000000000000000005400000000",
            INIT_3D => X"0000000000000000000000220000000000000000000000000000000000000000",
            INIT_3E => X"000000000000000000000023000000000000000f000000000000003300000000",
            INIT_3F => X"0000005e00000000000001160000000000000000000000000000005400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002e000000000000002e0000000000000000000000000000000000000000",
            INIT_41 => X"00000014000000000000000e0000000000000030000000000000001800000000",
            INIT_42 => X"00000016000000000000000d000000000000000e000000000000000500000000",
            INIT_43 => X"00000000000000000000003f00000000000000c9000000000000000000000000",
            INIT_44 => X"0000000000000000000000520000000000000010000000000000000000000000",
            INIT_45 => X"0000002600000000000000310000000000000010000000000000000000000000",
            INIT_46 => X"0000000000000000000000970000000000000000000000000000001700000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000008e00000000",
            INIT_48 => X"0000000000000000000000c90000000000000000000000000000000000000000",
            INIT_49 => X"0000000a000000000000000e0000000000000029000000000000000300000000",
            INIT_4A => X"000000ac00000000000000080000000000000024000000000000000800000000",
            INIT_4B => X"0000000000000000000000370000000000000001000000000000000600000000",
            INIT_4C => X"0000001700000000000000400000000000000000000000000000001900000000",
            INIT_4D => X"0000003200000000000000100000000000000045000000000000000000000000",
            INIT_4E => X"0000006e0000000000000000000000000000002f000000000000008200000000",
            INIT_4F => X"0000000000000000000000000000000000000052000000000000000000000000",
            INIT_50 => X"00000035000000000000001c0000000000000000000000000000006800000000",
            INIT_51 => X"0000004400000000000000260000000000000022000000000000001200000000",
            INIT_52 => X"0000002c00000000000000000000000000000002000000000000000000000000",
            INIT_53 => X"0000000000000000000000260000000000000000000000000000009100000000",
            INIT_54 => X"0000003e0000000000000000000000000000000b000000000000000000000000",
            INIT_55 => X"00000000000000000000004b0000000000000028000000000000002c00000000",
            INIT_56 => X"0000006400000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000059000000000000006000000000",
            INIT_58 => X"0000000000000000000000250000000000000000000000000000003a00000000",
            INIT_59 => X"0000001a00000000000000000000000000000070000000000000004e00000000",
            INIT_5A => X"0000001d00000000000000000000000000000000000000000000007e00000000",
            INIT_5B => X"00000058000000000000000c0000000000000036000000000000007b00000000",
            INIT_5C => X"00000040000000000000001d0000000000000000000000000000000000000000",
            INIT_5D => X"0000008500000000000000000000000000000000000000000000008900000000",
            INIT_5E => X"0000001900000000000000000000000000000000000000000000008100000000",
            INIT_5F => X"0000000b000000000000002a0000000000000059000000000000006d00000000",
            INIT_60 => X"00000067000000000000002c0000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000002700000000000000000000000000000022000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000019000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"00000005000000000000000a0000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"000000000000000000000000000000000000004b000000000000000400000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000002f00000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000230000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"000000000000000000000000000000000000004e000000000000000000000000",
            INIT_74 => X"0000000b00000000000000190000000000000000000000000000000000000000",
            INIT_75 => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_77 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_78 => X"00000000000000000000000c0000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000060000000000000011000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000410000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE30;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE31 : if BRAM_NAME = "samplegold_layersamples_instance31" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000090000000000000014000000000000000f00000000",
            INIT_01 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_02 => X"0000006000000000000000270000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_04 => X"00000000000000000000006e000000000000000f000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"000000c800000000000000220000000000000000000000000000001500000000",
            INIT_0F => X"0000004100000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"000000000000000000000093000000000000003e000000000000002000000000",
            INIT_11 => X"0000002400000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"000000a500000000000000170000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_16 => X"0000008c000000000000000a0000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000003f00000000",
            INIT_18 => X"0000002b000000000000009a0000000000000050000000000000000000000000",
            INIT_19 => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"000000430000000000000028000000000000001d000000000000000000000000",
            INIT_1B => X"0000000100000000000000000000000000000019000000000000000000000000",
            INIT_1C => X"0000005400000000000000000000000000000030000000000000000000000000",
            INIT_1D => X"0000000000000000000000110000000000000004000000000000000000000000",
            INIT_1E => X"000000000000000000000027000000000000002d000000000000001f00000000",
            INIT_1F => X"0000000000000000000000150000000000000000000000000000000800000000",
            INIT_20 => X"00000000000000000000004b0000000000000000000000000000002b00000000",
            INIT_21 => X"0000001e00000000000000000000000000000013000000000000003300000000",
            INIT_22 => X"0000000b00000000000000000000000000000013000000000000001600000000",
            INIT_23 => X"0000000a000000000000001d0000000000000002000000000000001b00000000",
            INIT_24 => X"00000033000000000000001d0000000000000043000000000000000000000000",
            INIT_25 => X"000000270000000000000020000000000000000e000000000000002d00000000",
            INIT_26 => X"00000000000000000000001b0000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000050000000000000016000000000000000000000000",
            INIT_28 => X"00000023000000000000006f000000000000001d000000000000002f00000000",
            INIT_29 => X"0000000000000000000000000000000000000063000000000000000600000000",
            INIT_2A => X"0000000900000000000000000000000000000033000000000000000300000000",
            INIT_2B => X"0000001100000000000000000000000000000009000000000000000000000000",
            INIT_2C => X"0000000000000000000000100000000000000077000000000000002c00000000",
            INIT_2D => X"00000000000000000000000a0000000000000048000000000000002500000000",
            INIT_2E => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_2F => X"0000002400000000000000110000000000000000000000000000000000000000",
            INIT_30 => X"00000000000000000000000b000000000000001b000000000000006d00000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000004500000000000000140000000000000000000000000000000000000000",
            INIT_34 => X"0000001a00000000000000120000000000000007000000000000001700000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"00000007000000000000002e0000000000000011000000000000001300000000",
            INIT_38 => X"0000000000000000000000030000000000000000000000000000001300000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"00000002000000000000001d0000000000000039000000000000000000000000",
            INIT_3C => X"0000000000000000000000170000000000000010000000000000001800000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000001e00000000000000110000000000000000000000000000000000000000",
            INIT_3F => X"0000001a00000000000000000000000000000038000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000290000000000000000000000000000000c00000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000003200000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"000000050000000000000018000000000000001e000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000002a00000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_47 => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"00000000000000000000003a0000000000000021000000000000000000000000",
            INIT_4B => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"00000000000000000000001a000000000000002c000000000000000b00000000",
            INIT_4F => X"0000000a000000000000000a0000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_51 => X"00000000000000000000001c000000000000000d000000000000000000000000",
            INIT_52 => X"0000000000000000000000180000000000000000000000000000001700000000",
            INIT_53 => X"00000000000000000000000f0000000000000006000000000000000000000000",
            INIT_54 => X"0000000200000000000000060000000000000000000000000000001900000000",
            INIT_55 => X"0000000600000000000000000000000000000019000000000000003200000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000400000000000000000000000000000000000000000000001a00000000",
            INIT_58 => X"00000020000000000000001b000000000000000b000000000000000800000000",
            INIT_59 => X"000000000000000000000001000000000000001a000000000000001b00000000",
            INIT_5A => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000009000000000000001600000000",
            INIT_5C => X"000000080000000000000025000000000000001d000000000000000800000000",
            INIT_5D => X"0000000e000000000000001e0000000000000000000000000000000200000000",
            INIT_5E => X"0000000f000000000000002d0000000000000000000000000000001100000000",
            INIT_5F => X"000000450000000000000000000000000000001a000000000000000000000000",
            INIT_60 => X"0000002100000000000000090000000000000015000000000000002a00000000",
            INIT_61 => X"0000000000000000000000050000000000000018000000000000000000000000",
            INIT_62 => X"000000000000000000000019000000000000001b000000000000001200000000",
            INIT_63 => X"0000000000000000000000260000000000000020000000000000002500000000",
            INIT_64 => X"0000000000000000000000030000000000000000000000000000002400000000",
            INIT_65 => X"0000003b00000000000000000000000000000000000000000000001700000000",
            INIT_66 => X"000000260000000000000045000000000000001a000000000000003d00000000",
            INIT_67 => X"0000001b00000000000000220000000000000028000000000000003400000000",
            INIT_68 => X"0000002100000000000000000000000000000008000000000000000000000000",
            INIT_69 => X"0000006c000000000000003f0000000000000003000000000000000000000000",
            INIT_6A => X"00000052000000000000004c0000000000000079000000000000006200000000",
            INIT_6B => X"0000000300000000000000170000000000000062000000000000004d00000000",
            INIT_6C => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_6D => X"00000065000000000000003f000000000000005c000000000000000800000000",
            INIT_6E => X"0000006c000000000000007b0000000000000071000000000000005800000000",
            INIT_6F => X"0000000000000000000000140000000000000055000000000000004800000000",
            INIT_70 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_71 => X"0000005a00000000000000620000000000000046000000000000002200000000",
            INIT_72 => X"0000006d000000000000004b000000000000006b000000000000007c00000000",
            INIT_73 => X"0000000000000000000000000000000000000016000000000000002900000000",
            INIT_74 => X"0000002000000000000000050000000000000000000000000000000000000000",
            INIT_75 => X"0000005000000000000000660000000000000052000000000000001800000000",
            INIT_76 => X"0000004f000000000000005c000000000000004d000000000000007000000000",
            INIT_77 => X"0000001000000000000000090000000000000000000000000000001300000000",
            INIT_78 => X"0000002400000000000000000000000000000007000000000000000300000000",
            INIT_79 => X"0000004c000000000000005d0000000000000065000000000000004400000000",
            INIT_7A => X"00000004000000000000004b0000000000000062000000000000006500000000",
            INIT_7B => X"0000003500000000000000670000000000000000000000000000001200000000",
            INIT_7C => X"00000065000000000000000b0000000000000000000000000000001900000000",
            INIT_7D => X"0000007700000000000000420000000000000051000000000000006b00000000",
            INIT_7E => X"0000000000000000000000220000000000000053000000000000006600000000",
            INIT_7F => X"0000002d000000000000002a000000000000000d000000000000001700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE31;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE32 : if BRAM_NAME = "samplegold_layersamples_instance32" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000057000000000000003d000000000000000b000000000000002600000000",
            INIT_01 => X"0000006000000000000000670000000000000055000000000000003400000000",
            INIT_02 => X"0000001d00000000000000000000000000000000000000000000005a00000000",
            INIT_03 => X"0000003100000000000000210000000000000017000000000000001600000000",
            INIT_04 => X"000000390000000000000019000000000000002d000000000000002e00000000",
            INIT_05 => X"000000340000000000000053000000000000005b000000000000006800000000",
            INIT_06 => X"0000002600000000000000070000000000000000000000000000000000000000",
            INIT_07 => X"0000002d000000000000001f000000000000002a000000000000002100000000",
            INIT_08 => X"00000042000000000000002e0000000000000039000000000000002100000000",
            INIT_09 => X"0000002d000000000000000e0000000000000026000000000000004a00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000004700000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000020000000000000002500000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"000000000000000000000036000000000000004d000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_3F => X"000000000000000000000006000000000000001e000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000031000000000000000400000000",
            INIT_42 => X"0000003700000000000000860000000000000000000000000000000000000000",
            INIT_43 => X"0000005a000000000000008a000000000000008a000000000000009a00000000",
            INIT_44 => X"0000007400000000000000a00000000000000045000000000000008800000000",
            INIT_45 => X"0000007000000000000000ce000000000000002f00000000000000a400000000",
            INIT_46 => X"0000009300000000000000310000000000000058000000000000005300000000",
            INIT_47 => X"0000007a000000000000006d000000000000004f000000000000008800000000",
            INIT_48 => X"000000af0000000000000073000000000000009e000000000000004700000000",
            INIT_49 => X"00000098000000000000006f00000000000000c3000000000000003900000000",
            INIT_4A => X"0000005100000000000000700000000000000058000000000000006d00000000",
            INIT_4B => X"0000009d00000000000000a2000000000000006a000000000000002c00000000",
            INIT_4C => X"0000003400000000000000be000000000000006d000000000000007000000000",
            INIT_4D => X"0000009900000000000000aa000000000000008500000000000000bb00000000",
            INIT_4E => X"00000008000000000000004e000000000000007600000000000000af00000000",
            INIT_4F => X"00000085000000000000005600000000000000ec00000000000000dc00000000",
            INIT_50 => X"000000c2000000000000008f00000000000000ca000000000000003e00000000",
            INIT_51 => X"000000b0000000000000005e00000000000000cc000000000000007900000000",
            INIT_52 => X"0000009b000000000000003c000000000000005200000000000000a500000000",
            INIT_53 => X"0000009f00000000000000cd000000000000004d000000000000009300000000",
            INIT_54 => X"0000007900000000000000aa000000000000006600000000000000c300000000",
            INIT_55 => X"0000009100000000000000a2000000000000002500000000000000b500000000",
            INIT_56 => X"00000000000000000000004c00000000000000d1000000000000005300000000",
            INIT_57 => X"0000007b00000000000000760000000000000072000000000000005e00000000",
            INIT_58 => X"000000a9000000000000008f00000000000000a0000000000000004800000000",
            INIT_59 => X"0000007e00000000000000640000000000000091000000000000003e00000000",
            INIT_5A => X"0000002700000000000000000000000000000005000000000000001c00000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_5C => X"000000510000000000000078000000000000008b000000000000006c00000000",
            INIT_5D => X"0000003b00000000000000850000000000000058000000000000008900000000",
            INIT_5E => X"0000000000000000000000010000000000000014000000000000000000000000",
            INIT_5F => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000007200000000000000550000000000000052000000000000007800000000",
            INIT_61 => X"000000000000000000000020000000000000006f000000000000004e00000000",
            INIT_62 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000006800000000000000460000000000000065000000000000006400000000",
            INIT_65 => X"00000000000000000000002d0000000000000087000000000000008a00000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"00000059000000000000005e0000000000000031000000000000000e00000000",
            INIT_68 => X"0000009500000000000000700000000000000086000000000000007500000000",
            INIT_69 => X"00000000000000000000003b000000000000004b000000000000005800000000",
            INIT_6A => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000003800000000000000b70000000000000026000000000000002200000000",
            INIT_6C => X"0000009e000000000000009100000000000000b3000000000000009c00000000",
            INIT_6D => X"00000000000000000000000b000000000000002e000000000000005200000000",
            INIT_6E => X"0000002200000000000000000000000000000008000000000000000000000000",
            INIT_6F => X"00000071000000000000006800000000000000ab000000000000004400000000",
            INIT_70 => X"0000008a00000000000000a900000000000000bb000000000000009d00000000",
            INIT_71 => X"000000000000000000000000000000000000000a000000000000003100000000",
            INIT_72 => X"0000000b00000000000000320000000000000000000000000000000400000000",
            INIT_73 => X"000000af000000000000005600000000000000a800000000000000d400000000",
            INIT_74 => X"000000c100000000000000cc00000000000000c300000000000000ae00000000",
            INIT_75 => X"00000000000000000000000a0000000000000020000000000000008000000000",
            INIT_76 => X"0000008f000000000000007d000000000000001f000000000000000000000000",
            INIT_77 => X"000000b40000000000000074000000000000009900000000000000ac00000000",
            INIT_78 => X"000000e100000000000000e700000000000000ae00000000000000a100000000",
            INIT_79 => X"000000080000000000000009000000000000001d000000000000006200000000",
            INIT_7A => X"0000001d00000000000000d800000000000000a6000000000000004400000000",
            INIT_7B => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_7C => X"0000003a0000000000000000000000000000000f000000000000000000000000",
            INIT_7D => X"000000600000000000000000000000000000002f000000000000001a00000000",
            INIT_7E => X"0000000000000000000000190000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000010000000000000001700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE32;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE33 : if BRAM_NAME = "samplegold_layersamples_instance33" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001b00000000000000240000000000000000000000000000000000000000",
            INIT_01 => X"0000001100000000000000510000000000000012000000000000002a00000000",
            INIT_02 => X"0000000a000000000000000b000000000000003f000000000000003a00000000",
            INIT_03 => X"0000000700000000000000000000000000000000000000000000000c00000000",
            INIT_04 => X"00000017000000000000001d0000000000000002000000000000003000000000",
            INIT_05 => X"0000005c000000000000003c000000000000008e000000000000001d00000000",
            INIT_06 => X"0000000100000000000000350000000000000010000000000000000200000000",
            INIT_07 => X"0000000000000000000000500000000000000038000000000000000000000000",
            INIT_08 => X"0000004b00000000000000410000000000000000000000000000001100000000",
            INIT_09 => X"0000000700000000000000820000000000000058000000000000009700000000",
            INIT_0A => X"0000000000000000000000190000000000000051000000000000004b00000000",
            INIT_0B => X"0000003a0000000000000000000000000000001b000000000000004500000000",
            INIT_0C => X"0000007b0000000000000028000000000000006f000000000000003900000000",
            INIT_0D => X"0000004e00000000000000000000000000000053000000000000006700000000",
            INIT_0E => X"00000049000000000000004d000000000000000e000000000000005d00000000",
            INIT_0F => X"0000004e00000000000000520000000000000051000000000000001e00000000",
            INIT_10 => X"0000005e000000000000007a0000000000000034000000000000004000000000",
            INIT_11 => X"0000004b000000000000003a0000000000000001000000000000004100000000",
            INIT_12 => X"0000003c000000000000004c0000000000000059000000000000007400000000",
            INIT_13 => X"0000004800000000000000540000000000000051000000000000005c00000000",
            INIT_14 => X"0000002b000000000000005d0000000000000056000000000000005d00000000",
            INIT_15 => X"00000078000000000000004a0000000000000030000000000000001600000000",
            INIT_16 => X"00000070000000000000005e0000000000000031000000000000006e00000000",
            INIT_17 => X"0000007100000000000000630000000000000058000000000000005b00000000",
            INIT_18 => X"0000001d0000000000000017000000000000005b000000000000007e00000000",
            INIT_19 => X"00000079000000000000004a0000000000000044000000000000004800000000",
            INIT_1A => X"00000082000000000000006d0000000000000067000000000000005e00000000",
            INIT_1B => X"0000007e0000000000000076000000000000006f000000000000008200000000",
            INIT_1C => X"00000036000000000000005b0000000000000004000000000000004000000000",
            INIT_1D => X"0000007300000000000000470000000000000048000000000000002a00000000",
            INIT_1E => X"0000009800000000000000850000000000000089000000000000006200000000",
            INIT_1F => X"000000250000000000000056000000000000007b000000000000006900000000",
            INIT_20 => X"0000001f000000000000002c0000000000000046000000000000000b00000000",
            INIT_21 => X"0000007f0000000000000036000000000000003b000000000000002a00000000",
            INIT_22 => X"0000006f000000000000008e000000000000009900000000000000a000000000",
            INIT_23 => X"0000006e00000000000000170000000000000054000000000000007000000000",
            INIT_24 => X"0000003900000000000000510000000000000088000000000000001b00000000",
            INIT_25 => X"000000a3000000000000008d0000000000000045000000000000004f00000000",
            INIT_26 => X"0000008000000000000000850000000000000076000000000000008700000000",
            INIT_27 => X"0000007c0000000000000048000000000000003c000000000000005e00000000",
            INIT_28 => X"00000048000000000000006c000000000000008f000000000000008600000000",
            INIT_29 => X"0000005600000000000000910000000000000087000000000000005f00000000",
            INIT_2A => X"0000006600000000000000690000000000000096000000000000007600000000",
            INIT_2B => X"000000290000000000000044000000000000005a000000000000000000000000",
            INIT_2C => X"000000540000000000000079000000000000008b000000000000006f00000000",
            INIT_2D => X"0000009000000000000000480000000000000032000000000000006100000000",
            INIT_2E => X"0000002100000000000000310000000000000078000000000000007e00000000",
            INIT_2F => X"000000270000000000000000000000000000003d000000000000000300000000",
            INIT_30 => X"00000070000000000000007e0000000000000099000000000000007e00000000",
            INIT_31 => X"0000007e0000000000000071000000000000005c000000000000006b00000000",
            INIT_32 => X"0000007e0000000000000014000000000000000a000000000000003000000000",
            INIT_33 => X"0000000600000000000000750000000000000000000000000000002400000000",
            INIT_34 => X"00000000000000000000001d0000000000000072000000000000000000000000",
            INIT_35 => X"0000002a00000000000000000000000000000000000000000000000500000000",
            INIT_36 => X"00000000000000000000001c0000000000000010000000000000000000000000",
            INIT_37 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_38 => X"00000000000000000000003e0000000000000000000000000000003f00000000",
            INIT_39 => X"0000000000000000000000650000000000000000000000000000001c00000000",
            INIT_3A => X"0000000000000000000000000000000000000004000000000000009200000000",
            INIT_3B => X"0000006600000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000016000000000000006500000000",
            INIT_3D => X"0000000000000000000000000000000000000039000000000000003a00000000",
            INIT_3E => X"0000000100000000000000a00000000000000000000000000000002300000000",
            INIT_3F => X"00000000000000000000008f0000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007b000000000000000000000000000000ac000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000005700000000",
            INIT_42 => X"0000000000000000000000000000000000000089000000000000000000000000",
            INIT_43 => X"0000009900000000000000000000000000000000000000000000006000000000",
            INIT_44 => X"0000000000000000000000110000000000000052000000000000000600000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000008e00000000000000000000000000000000000000000000007100000000",
            INIT_47 => X"00000000000000000000004a0000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000630000000000000000000000000000000000000000",
            INIT_49 => X"0000005500000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000300000000000000000000000000000007000000000000000000000000",
            INIT_4D => X"00000016000000000000001e0000000000000000000000000000000000000000",
            INIT_4E => X"0000001100000000000000000000000000000014000000000000000000000000",
            INIT_4F => X"0000001000000000000000130000000000000000000000000000001000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000320000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000180000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000004b00000000000000000000000000000011000000000000001500000000",
            INIT_59 => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000004b00000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"00000000000000000000009a0000000000000000000000000000004100000000",
            INIT_5D => X"0000001b00000000000000000000000000000000000000000000002500000000",
            INIT_5E => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"000000000000000000000000000000000000001e000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000004c00000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000002700000000000000000000000000000000000000000000009f00000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000003c00000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"000000000000000000000000000000000000000000000000000000cf00000000",
            INIT_6C => X"0000000000000000000000310000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000190000000000000009000000000000000000000000",
            INIT_6E => X"0000000000000000000000580000000000000000000000000000001d00000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"00000000000000000000003c0000000000000046000000000000000000000000",
            INIT_71 => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_74 => X"0000003500000000000000000000000000000000000000000000000100000000",
            INIT_75 => X"00000000000000000000000d0000000000000086000000000000000000000000",
            INIT_76 => X"0000003a00000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000250000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000450000000000000000000000000000006100000000",
            INIT_7A => X"00000000000000000000009b0000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000003000000000000001c00000000",
            INIT_7E => X"00000000000000000000001f00000000000000c6000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000001800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE33;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE34 : if BRAM_NAME = "samplegold_layersamples_instance34" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_01 => X"000000000000000000000000000000000000002b000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000051000000000000004700000000",
            INIT_03 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000003800000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000003000000000000000d00000000",
            INIT_08 => X"0000001b00000000000000000000000000000052000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"000000050000000000000000000000000000002b000000000000002400000000",
            INIT_0B => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000037000000000000000000000000",
            INIT_0D => X"0000002400000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000107000000000000000200000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000560000000000000000000000000000004600000000",
            INIT_12 => X"00000000000000000000000000000000000000b5000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"00000012000000000000000b0000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000024000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000f00000000000000017000000000000000000000000",
            INIT_19 => X"0000000000000000000000640000000000000000000000000000000000000000",
            INIT_1A => X"0000003100000000000000000000000000000079000000000000000000000000",
            INIT_1B => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_1C => X"00000019000000000000010e0000000000000050000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_20 => X"0000002100000000000000ba000000000000009f000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"000000000000000000000000000000000000003f000000000000003d00000000",
            INIT_23 => X"0000000000000000000000000000000000000062000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000150000000000000013000000000000001a00000000",
            INIT_5D => X"00000029000000000000002c0000000000000018000000000000003300000000",
            INIT_5E => X"00000000000000000000004c0000000000000019000000000000003900000000",
            INIT_5F => X"0000002e000000000000000e000000000000002f000000000000001d00000000",
            INIT_60 => X"0000001300000000000000060000000000000010000000000000001500000000",
            INIT_61 => X"0000002700000000000000240000000000000038000000000000001000000000",
            INIT_62 => X"0000002600000000000000160000000000000041000000000000001800000000",
            INIT_63 => X"0000001f0000000000000033000000000000000a000000000000000000000000",
            INIT_64 => X"00000037000000000000002e0000000000000011000000000000000300000000",
            INIT_65 => X"0000004100000000000000000000000000000024000000000000001b00000000",
            INIT_66 => X"0000002e000000000000001f000000000000000d000000000000003e00000000",
            INIT_67 => X"00000002000000000000000e000000000000002e000000000000000e00000000",
            INIT_68 => X"0000002200000000000000490000000000000040000000000000003600000000",
            INIT_69 => X"0000005a00000000000000190000000000000026000000000000003600000000",
            INIT_6A => X"0000001600000000000000000000000000000020000000000000001d00000000",
            INIT_6B => X"0000004400000000000000120000000000000000000000000000002300000000",
            INIT_6C => X"0000002b000000000000005c0000000000000006000000000000003f00000000",
            INIT_6D => X"0000002800000000000000700000000000000042000000000000004900000000",
            INIT_6E => X"0000001f00000000000000050000000000000000000000000000000b00000000",
            INIT_6F => X"000000400000000000000034000000000000000b000000000000002600000000",
            INIT_70 => X"0000004400000000000000370000000000000016000000000000003b00000000",
            INIT_71 => X"00000012000000000000002b0000000000000066000000000000003b00000000",
            INIT_72 => X"0000002b000000000000000d000000000000001c000000000000000000000000",
            INIT_73 => X"00000036000000000000001b0000000000000031000000000000002d00000000",
            INIT_74 => X"0000001b000000000000001c000000000000002d000000000000000a00000000",
            INIT_75 => X"0000001000000000000000280000000000000038000000000000001a00000000",
            INIT_76 => X"00000023000000000000001d0000000000000020000000000000001c00000000",
            INIT_77 => X"00000039000000000000001e0000000000000008000000000000001100000000",
            INIT_78 => X"00000018000000000000000f0000000000000016000000000000001400000000",
            INIT_79 => X"0000002c0000000000000000000000000000001f000000000000000000000000",
            INIT_7A => X"0000001500000000000000200000000000000016000000000000001d00000000",
            INIT_7B => X"00000000000000000000000f0000000000000008000000000000001100000000",
            INIT_7C => X"0000000f00000000000000020000000000000032000000000000001100000000",
            INIT_7D => X"0000000a00000000000000110000000000000019000000000000000400000000",
            INIT_7E => X"000000280000000000000007000000000000002a000000000000001c00000000",
            INIT_7F => X"0000000000000000000000170000000000000000000000000000000500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE34;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE35 : if BRAM_NAME = "samplegold_layersamples_instance35" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000c0000000000000000000000000000000c000000000000001800000000",
            INIT_01 => X"0000002400000000000000450000000000000000000000000000004700000000",
            INIT_02 => X"0000002e000000000000000a0000000000000026000000000000001700000000",
            INIT_03 => X"0000000200000000000000020000000000000000000000000000000000000000",
            INIT_04 => X"0000000500000000000000210000000000000010000000000000001700000000",
            INIT_05 => X"00000034000000000000003f000000000000001d000000000000005400000000",
            INIT_06 => X"0000001300000000000000070000000000000026000000000000001c00000000",
            INIT_07 => X"0000000f00000000000000000000000000000007000000000000000000000000",
            INIT_08 => X"0000000b000000000000003d0000000000000024000000000000003100000000",
            INIT_09 => X"0000003900000000000000620000000000000064000000000000005e00000000",
            INIT_0A => X"0000002500000000000000000000000000000007000000000000003e00000000",
            INIT_0B => X"0000000c00000000000000010000000000000000000000000000000b00000000",
            INIT_0C => X"0000002a00000000000000030000000000000042000000000000003700000000",
            INIT_0D => X"00000052000000000000005e000000000000007d000000000000007200000000",
            INIT_0E => X"00000000000000000000001e0000000000000034000000000000004f00000000",
            INIT_0F => X"0000005100000000000000000000000000000009000000000000001300000000",
            INIT_10 => X"0000004100000000000000250000000000000016000000000000004300000000",
            INIT_11 => X"00000060000000000000005b0000000000000070000000000000007300000000",
            INIT_12 => X"00000000000000000000000d000000000000004b000000000000004a00000000",
            INIT_13 => X"0000005f0000000000000014000000000000002e000000000000001400000000",
            INIT_14 => X"00000074000000000000007a0000000000000027000000000000008000000000",
            INIT_15 => X"0000007200000000000000940000000000000084000000000000008800000000",
            INIT_16 => X"0000007100000000000000710000000000000054000000000000007700000000",
            INIT_17 => X"0000003d0000000000000079000000000000005d000000000000007900000000",
            INIT_18 => X"0000007f00000000000000790000000000000075000000000000005600000000",
            INIT_19 => X"0000009f00000000000000980000000000000091000000000000008400000000",
            INIT_1A => X"0000007c00000000000000790000000000000067000000000000005600000000",
            INIT_1B => X"0000004f0000000000000045000000000000007a000000000000007f00000000",
            INIT_1C => X"00000081000000000000006b000000000000006f000000000000006000000000",
            INIT_1D => X"000000820000000000000089000000000000007b000000000000009400000000",
            INIT_1E => X"0000008600000000000000870000000000000081000000000000006600000000",
            INIT_1F => X"00000066000000000000003d0000000000000058000000000000007600000000",
            INIT_20 => X"00000098000000000000008c000000000000006d000000000000005f00000000",
            INIT_21 => X"00000083000000000000009a0000000000000074000000000000007a00000000",
            INIT_22 => X"00000080000000000000007f000000000000008d000000000000008600000000",
            INIT_23 => X"00000062000000000000005d0000000000000052000000000000004100000000",
            INIT_24 => X"0000006a000000000000006f000000000000005e000000000000007400000000",
            INIT_25 => X"0000006b00000000000000650000000000000085000000000000007500000000",
            INIT_26 => X"0000003c000000000000007b000000000000006b000000000000006200000000",
            INIT_27 => X"000000530000000000000053000000000000005a000000000000006b00000000",
            INIT_28 => X"0000006900000000000000280000000000000020000000000000001700000000",
            INIT_29 => X"0000004c0000000000000082000000000000006a000000000000005700000000",
            INIT_2A => X"0000004200000000000000000000000000000075000000000000006700000000",
            INIT_2B => X"0000001000000000000000370000000000000050000000000000004200000000",
            INIT_2C => X"00000025000000000000002a000000000000006c000000000000006a00000000",
            INIT_2D => X"000000640000000000000045000000000000006c000000000000006c00000000",
            INIT_2E => X"0000005500000000000000220000000000000087000000000000007000000000",
            INIT_2F => X"0000004e0000000000000049000000000000000f000000000000003c00000000",
            INIT_30 => X"00000061000000000000003b000000000000002a000000000000003800000000",
            INIT_31 => X"000000610000000000000053000000000000003b000000000000005000000000",
            INIT_32 => X"0000002f000000000000004c000000000000002c00000000000000ac00000000",
            INIT_33 => X"0000005c00000000000000700000000000000058000000000000002300000000",
            INIT_34 => X"000000730000000000000093000000000000004c000000000000005f00000000",
            INIT_35 => X"000000be00000000000000770000000000000039000000000000002800000000",
            INIT_36 => X"000000150000000000000078000000000000002e000000000000003100000000",
            INIT_37 => X"00000089000000000000006b00000000000000b1000000000000001900000000",
            INIT_38 => X"0000003800000000000000630000000000000070000000000000006e00000000",
            INIT_39 => X"0000005100000000000000aa000000000000007a000000000000001900000000",
            INIT_3A => X"00000052000000000000003400000000000000c5000000000000004200000000",
            INIT_3B => X"0000005100000000000000a30000000000000086000000000000009a00000000",
            INIT_3C => X"0000000e00000000000000490000000000000072000000000000004a00000000",
            INIT_3D => X"00000052000000000000008100000000000000ba000000000000007b00000000",
            INIT_3E => X"00000075000000000000008b0000000000000085000000000000008000000000",
            INIT_3F => X"0000003600000000000000420000000000000053000000000000007b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000750000000000000039000000000000005c000000000000002100000000",
            INIT_41 => X"0000004a000000000000006600000000000000b0000000000000009f00000000",
            INIT_42 => X"000000a100000000000000af000000000000007a000000000000004500000000",
            INIT_43 => X"0000004300000000000000530000000000000055000000000000007500000000",
            INIT_44 => X"0000009b0000000000000042000000000000006d000000000000002800000000",
            INIT_45 => X"0000008c0000000000000064000000000000009f000000000000009000000000",
            INIT_46 => X"0000009000000000000000c30000000000000092000000000000009600000000",
            INIT_47 => X"00000075000000000000006e000000000000008b000000000000008300000000",
            INIT_48 => X"0000008f00000000000000c7000000000000007e000000000000005e00000000",
            INIT_49 => X"000000a7000000000000008d000000000000009300000000000000be00000000",
            INIT_4A => X"000000b3000000000000009c00000000000000a7000000000000009600000000",
            INIT_4B => X"0000009600000000000000980000000000000096000000000000009900000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000007900000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"00000000000000000000000c000000000000000c000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000800000000000000080000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_5E => X"00000000000000000000000c0000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000006000000000000000000000000000000000000000000000000500000000",
            INIT_61 => X"0000002300000000000000010000000000000000000000000000000e00000000",
            INIT_62 => X"0000000400000000000000010000000000000000000000000000000500000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000021000000000000000800000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"000000000000000000000006000000000000000e000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000001900000000000000260000000000000035000000000000001800000000",
            INIT_6C => X"000000c700000000000000cb000000000000008300000000000000a400000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000002d00000000",
            INIT_6E => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000210000000000000022000000000000008900000000",
            INIT_70 => X"000000000000000000000000000000000000002a000000000000000d00000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000001c000000000000001a0000000000000042000000000000001c00000000",
            INIT_73 => X"0000005f00000000000000ac000000000000007300000000000000cf00000000",
            INIT_74 => X"000000000000000000000000000000000000004d000000000000001f00000000",
            INIT_75 => X"00000000000000000000000f0000000000000000000000000000002a00000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_77 => X"00000007000000000000000d000000000000001c000000000000000000000000",
            INIT_78 => X"0000006d000000000000000c0000000000000037000000000000000200000000",
            INIT_79 => X"0000000f00000000000000000000000000000000000000000000000e00000000",
            INIT_7A => X"0000000000000000000000010000000000000000000000000000002800000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000004800000000000000000000000000000006000000000000000000000000",
            INIT_7D => X"0000001e000000000000000c0000000000000011000000000000000a00000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE35;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE36 : if BRAM_NAME = "samplegold_layersamples_instance36" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000e000000000000000b0000000000000012000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000002a00000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"000000230000000000000012000000000000002d000000000000002400000000",
            INIT_06 => X"0000003200000000000000000000000000000051000000000000001d00000000",
            INIT_07 => X"0000004300000000000000210000000000000008000000000000002100000000",
            INIT_08 => X"000000460000000000000000000000000000002b000000000000000000000000",
            INIT_09 => X"0000001e0000000000000022000000000000001f000000000000001e00000000",
            INIT_0A => X"0000003d00000000000000120000000000000000000000000000003600000000",
            INIT_0B => X"0000002e00000000000000070000000000000038000000000000003500000000",
            INIT_0C => X"000000340000000000000033000000000000000d000000000000000000000000",
            INIT_0D => X"0000005600000000000000030000000000000023000000000000002c00000000",
            INIT_0E => X"0000001b00000000000000300000000000000000000000000000002f00000000",
            INIT_0F => X"00000019000000000000002c0000000000000036000000000000002e00000000",
            INIT_10 => X"0000002700000000000000450000000000000024000000000000001600000000",
            INIT_11 => X"0000004c00000000000000380000000000000021000000000000004300000000",
            INIT_12 => X"0000001300000000000000000000000000000037000000000000002f00000000",
            INIT_13 => X"00000027000000000000003b000000000000002f000000000000003f00000000",
            INIT_14 => X"0000002c0000000000000025000000000000003a000000000000002300000000",
            INIT_15 => X"0000006200000000000000000000000000000001000000000000000a00000000",
            INIT_16 => X"0000002c00000000000000400000000000000000000000000000005600000000",
            INIT_17 => X"000000140000000000000002000000000000011d000000000000002800000000",
            INIT_18 => X"0000000000000000000000680000000000000020000000000000001c00000000",
            INIT_19 => X"0000000000000000000000450000000000000000000000000000000200000000",
            INIT_1A => X"00000038000000000000002c0000000000000031000000000000000000000000",
            INIT_1B => X"000000000000000000000000000000000000009d00000000000000b300000000",
            INIT_1C => X"000000000000000000000008000000000000000b000000000000005a00000000",
            INIT_1D => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_1E => X"00000000000000000000001f0000000000000021000000000000002800000000",
            INIT_1F => X"00000053000000000000003a000000000000000000000000000000cf00000000",
            INIT_20 => X"0000000000000000000000290000000000000026000000000000000000000000",
            INIT_21 => X"0000006400000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"000000b400000000000000110000000000000000000000000000001c00000000",
            INIT_23 => X"0000007c00000000000000000000000000000013000000000000000000000000",
            INIT_24 => X"0000001f00000000000000300000000000000039000000000000000000000000",
            INIT_25 => X"0000006a00000000000000980000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000c10000000000000000000000000000000000000000",
            INIT_27 => X"00000000000000000000006800000000000000ae000000000000000000000000",
            INIT_28 => X"0000000200000000000000110000000000000000000000000000002800000000",
            INIT_29 => X"0000000000000000000000af0000000000000088000000000000000000000000",
            INIT_2A => X"00000000000000000000000000000000000000b0000000000000000000000000",
            INIT_2B => X"0000006600000000000000210000000000000037000000000000003c00000000",
            INIT_2C => X"0000001f0000000000000015000000000000001b000000000000000000000000",
            INIT_2D => X"00000035000000000000000000000000000000ed000000000000005900000000",
            INIT_2E => X"000000000000000000000000000000000000002a000000000000003f00000000",
            INIT_2F => X"0000000000000000000000000000000000000034000000000000002900000000",
            INIT_30 => X"00000075000000000000002b0000000000000000000000000000000100000000",
            INIT_31 => X"0000003300000000000000550000000000000004000000000000009700000000",
            INIT_32 => X"0000000a00000000000000000000000000000056000000000000003400000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000003800000000",
            INIT_34 => X"0000004700000000000000340000000000000005000000000000000000000000",
            INIT_35 => X"0000000000000000000000920000000000000000000000000000003b00000000",
            INIT_36 => X"0000004e000000000000001d0000000000000000000000000000007300000000",
            INIT_37 => X"0000001500000000000000060000000000000023000000000000000000000000",
            INIT_38 => X"0000000000000000000000350000000000000008000000000000002000000000",
            INIT_39 => X"00000047000000000000001c000000000000003a000000000000002500000000",
            INIT_3A => X"0000002c0000000000000031000000000000000a000000000000002a00000000",
            INIT_3B => X"0000003f000000000000003f0000000000000038000000000000002900000000",
            INIT_3C => X"0000001e00000000000000580000000000000000000000000000002100000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_3F => X"00000044000000000000001a0000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000008000000000000000300000000",
            INIT_42 => X"0000002600000000000000140000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_44 => X"00000000000000000000000d0000000000000000000000000000000d00000000",
            INIT_45 => X"0000000300000000000000030000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000003000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000001000000000000000300000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000070000000000000028000000000000001400000000",
            INIT_4C => X"00000004000000000000001d0000000000000000000000000000000000000000",
            INIT_4D => X"000000170000000000000012000000000000000e000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000005200000000000000600000000000000000000000000000000000000000",
            INIT_50 => X"0000000200000000000000170000000000000000000000000000004d00000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000049000000000000000900000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000c0000000000000000000000000000002e000000000000000000000000",
            INIT_55 => X"0000000200000000000000090000000000000013000000000000000000000000",
            INIT_56 => X"00000000000000000000000a0000000000000017000000000000001500000000",
            INIT_57 => X"0000000300000000000000000000000000000001000000000000000d00000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000008500000000",
            INIT_5D => X"00000022000000000000003a000000000000000d000000000000000000000000",
            INIT_5E => X"0000003000000000000000290000000000000000000000000000000300000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000003b00000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_62 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_63 => X"0000004c00000000000000be000000000000007b000000000000002b00000000",
            INIT_64 => X"0000000b00000000000000000000000000000003000000000000007100000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"00000000000000000000000f0000000000000000000000000000000100000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000002d00000000000000000000000000000035000000000000006a00000000",
            INIT_69 => X"0000000000000000000000000000000000000002000000000000003700000000",
            INIT_6A => X"000000000000000000000000000000000000002b000000000000001a00000000",
            INIT_6B => X"000000000000000000000000000000000000001d000000000000000000000000",
            INIT_6C => X"00000000000000000000001e0000000000000024000000000000000000000000",
            INIT_6D => X"0000001a0000000000000000000000000000006d000000000000005100000000",
            INIT_6E => X"0000002b00000000000000000000000000000003000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"000000000000000000000000000000000000003a000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000180000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000006000000000000001600000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_7C => X"0000000000000000000000470000000000000000000000000000000200000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE36;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE37 : if BRAM_NAME = "samplegold_layersamples_instance37" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000003100000000",
            INIT_05 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_06 => X"0000007500000000000000000000000000000000000000000000000700000000",
            INIT_07 => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_08 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"000000340000000000000063000000000000003a000000000000000000000000",
            INIT_0A => X"000000000000000000000051000000000000001a000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000022000000000000004300000000",
            INIT_0F => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_11 => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000004100000000000000000000000000000000000000000000004900000000",
            INIT_13 => X"0000003a00000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000003e000000000000002d0000000000000000000000000000000000000000",
            INIT_15 => X"0000000a00000000000000ed00000000000000a0000000000000002300000000",
            INIT_16 => X"00000006000000000000004c0000000000000000000000000000000000000000",
            INIT_17 => X"0000001500000000000000bc0000000000000000000000000000000000000000",
            INIT_18 => X"000000780000000000000000000000000000005b000000000000001200000000",
            INIT_19 => X"0000000000000000000000060000000000000000000000000000002b00000000",
            INIT_1A => X"0000000000000000000000070000000000000075000000000000000000000000",
            INIT_1B => X"0000000b000000000000000000000000000000bf000000000000001e00000000",
            INIT_1C => X"0000003a00000000000000820000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_1E => X"0000000000000000000000000000000000000015000000000000006e00000000",
            INIT_1F => X"0000000000000000000000000000000000000053000000000000000000000000",
            INIT_20 => X"0000002200000000000000000000000000000000000000000000007b00000000",
            INIT_21 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_22 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000052000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"000000330000000000000000000000000000002b000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"000000000000000000000000000000000000005d000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000070000000000000011000000000000000000000000",
            INIT_2C => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"00000037000000000000002f000000000000006e000000000000000000000000",
            INIT_2E => X"0000005100000000000000440000000000000059000000000000004400000000",
            INIT_2F => X"0000001f0000000000000012000000000000006c000000000000001f00000000",
            INIT_30 => X"000000510000000000000000000000000000001a000000000000003f00000000",
            INIT_31 => X"0000003d00000000000000340000000000000069000000000000004400000000",
            INIT_32 => X"0000004b0000000000000063000000000000004f000000000000004000000000",
            INIT_33 => X"000000070000000000000000000000000000002d000000000000008800000000",
            INIT_34 => X"0000006400000000000000170000000000000046000000000000001d00000000",
            INIT_35 => X"0000003d0000000000000033000000000000003d000000000000003300000000",
            INIT_36 => X"00000050000000000000001f0000000000000072000000000000004400000000",
            INIT_37 => X"0000002100000000000000440000000000000013000000000000009d00000000",
            INIT_38 => X"000000130000000000000049000000000000002d000000000000001b00000000",
            INIT_39 => X"0000004b00000000000000410000000000000028000000000000003900000000",
            INIT_3A => X"0000003e000000000000001e0000000000000054000000000000004c00000000",
            INIT_3B => X"00000010000000000000002e0000000000000076000000000000003a00000000",
            INIT_3C => X"0000004100000000000000260000000000000000000000000000001c00000000",
            INIT_3D => X"000000470000000000000048000000000000003e000000000000003700000000",
            INIT_3E => X"0000002e00000000000000080000000000000057000000000000005500000000",
            INIT_3F => X"000000200000000000000019000000000000001400000000000000b600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003a00000000000000240000000000000037000000000000000000000000",
            INIT_41 => X"00000000000000000000006a0000000000000000000000000000003600000000",
            INIT_42 => X"0000006900000000000000450000000000000005000000000000007c00000000",
            INIT_43 => X"0000000000000000000000100000000000000022000000000000000000000000",
            INIT_44 => X"00000006000000000000005c000000000000003b000000000000000000000000",
            INIT_45 => X"0000001500000000000000940000000000000036000000000000001400000000",
            INIT_46 => X"0000000000000000000000530000000000000077000000000000002500000000",
            INIT_47 => X"00000000000000000000004f000000000000001b000000000000002100000000",
            INIT_48 => X"0000003a00000000000000000000000000000000000000000000004c00000000",
            INIT_49 => X"000000330000000000000014000000000000000b000000000000004100000000",
            INIT_4A => X"000000120000000000000000000000000000006200000000000000be00000000",
            INIT_4B => X"000000320000000000000000000000000000004d000000000000004f00000000",
            INIT_4C => X"0000008200000000000000000000000000000039000000000000004100000000",
            INIT_4D => X"0000007200000000000000100000000000000020000000000000001400000000",
            INIT_4E => X"000000e800000000000000000000000000000000000000000000004300000000",
            INIT_4F => X"0000013000000000000000270000000000000000000000000000006100000000",
            INIT_50 => X"0000001900000000000000830000000000000000000000000000000000000000",
            INIT_51 => X"00000050000000000000002f000000000000002b000000000000009000000000",
            INIT_52 => X"0000006300000000000001320000000000000000000000000000000000000000",
            INIT_53 => X"0000001000000000000000d8000000000000002e000000000000000000000000",
            INIT_54 => X"0000005a00000000000000000000000000000012000000000000000000000000",
            INIT_55 => X"000000000000000000000004000000000000000c000000000000003e00000000",
            INIT_56 => X"0000002c000000000000002100000000000000e5000000000000000000000000",
            INIT_57 => X"00000039000000000000003f0000000000000094000000000000000000000000",
            INIT_58 => X"00000010000000000000003c000000000000006c000000000000002900000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_5A => X"0000002e0000000000000018000000000000002b000000000000001500000000",
            INIT_5B => X"00000024000000000000005f0000000000000081000000000000000000000000",
            INIT_5C => X"0000003d00000000000000410000000000000065000000000000006c00000000",
            INIT_5D => X"00000000000000000000000f0000000000000000000000000000001600000000",
            INIT_5E => X"0000001c00000000000000530000000000000000000000000000005100000000",
            INIT_5F => X"0000007800000000000000000000000000000031000000000000004f00000000",
            INIT_60 => X"0000002f00000000000000430000000000000046000000000000003100000000",
            INIT_61 => X"0000002100000000000000280000000000000026000000000000004f00000000",
            INIT_62 => X"00000044000000000000001e0000000000000045000000000000002600000000",
            INIT_63 => X"0000003800000000000000280000000000000033000000000000003300000000",
            INIT_64 => X"0000003d000000000000001b0000000000000028000000000000002d00000000",
            INIT_65 => X"0000000000000000000000000000000000000010000000000000005a00000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000008000000000000001900000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000370000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000001300000000000000120000000000000000000000000000000c00000000",
            INIT_78 => X"000000000000000000000000000000000000005b000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000065000000000000006900000000",
            INIT_7B => X"0000000000000000000000000000000000000018000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000058000000000000000000000000",
            INIT_7D => X"0000000000000000000000130000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE37;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE38 : if BRAM_NAME = "samplegold_layersamples_instance38" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000100000000000000000000000000000001200000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000002900000000000000090000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000007f00000000000000610000000000000044000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000008900000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000003a000000000000004b000000000000011b000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000002500000000",
            INIT_0A => X"000000000000000000000000000000000000001b000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_0C => X"00000000000000000000004a0000000000000000000000000000000000000000",
            INIT_0D => X"0000004d000000000000001f000000000000000e000000000000009d00000000",
            INIT_0E => X"0000002200000000000000000000000000000040000000000000000000000000",
            INIT_0F => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000055000000000000001000000000",
            INIT_13 => X"0000001a000000000000001c0000000000000081000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000e00000000000000260000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000024000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000002e00000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000007000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000004a00000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"000000cb00000000000000c300000000000000cc000000000000008900000000",
            INIT_57 => X"000000b700000000000000c500000000000000d900000000000000d100000000",
            INIT_58 => X"0000007b00000000000000730000000000000067000000000000008400000000",
            INIT_59 => X"000000a300000000000000620000000000000081000000000000006e00000000",
            INIT_5A => X"000000df00000000000000d700000000000000be00000000000000b800000000",
            INIT_5B => X"000000bf00000000000000ea00000000000000e300000000000000db00000000",
            INIT_5C => X"000000920000000000000076000000000000006f000000000000006700000000",
            INIT_5D => X"000000aa00000000000000a20000000000000074000000000000009300000000",
            INIT_5E => X"000000e300000000000000d700000000000000d200000000000000c800000000",
            INIT_5F => X"000000ac00000000000000ce00000000000000d800000000000000e600000000",
            INIT_60 => X"00000089000000000000009c000000000000009c00000000000000ab00000000",
            INIT_61 => X"000000c400000000000000b30000000000000069000000000000008e00000000",
            INIT_62 => X"000000de00000000000000e700000000000000da00000000000000cf00000000",
            INIT_63 => X"000000c400000000000000d100000000000000c700000000000000d100000000",
            INIT_64 => X"0000008e000000000000008f0000000000000090000000000000009e00000000",
            INIT_65 => X"000000d400000000000000c600000000000000a8000000000000008300000000",
            INIT_66 => X"000000ae00000000000000a500000000000000d200000000000000d600000000",
            INIT_67 => X"0000008300000000000000ab00000000000000c000000000000000b100000000",
            INIT_68 => X"00000054000000000000008d0000000000000087000000000000007900000000",
            INIT_69 => X"000000b900000000000000c200000000000000ba00000000000000bc00000000",
            INIT_6A => X"0000007600000000000000640000000000000083000000000000008800000000",
            INIT_6B => X"0000006600000000000000480000000000000093000000000000009b00000000",
            INIT_6C => X"00000085000000000000009b0000000000000089000000000000007c00000000",
            INIT_6D => X"000000ab000000000000008800000000000000a800000000000000a500000000",
            INIT_6E => X"0000008500000000000000820000000000000088000000000000007900000000",
            INIT_6F => X"0000007900000000000000540000000000000043000000000000006a00000000",
            INIT_70 => X"0000009b0000000000000099000000000000009f000000000000008300000000",
            INIT_71 => X"000000b500000000000000900000000000000097000000000000008400000000",
            INIT_72 => X"00000069000000000000007f0000000000000078000000000000009e00000000",
            INIT_73 => X"0000006d00000000000000870000000000000047000000000000003e00000000",
            INIT_74 => X"00000075000000000000008c00000000000000b000000000000000a700000000",
            INIT_75 => X"0000009b0000000000000098000000000000007a00000000000000a800000000",
            INIT_76 => X"0000003300000000000000400000000000000070000000000000008800000000",
            INIT_77 => X"000000bb00000000000000560000000000000087000000000000005000000000",
            INIT_78 => X"0000004000000000000000710000000000000075000000000000009e00000000",
            INIT_79 => X"000000b100000000000000bb0000000000000076000000000000008e00000000",
            INIT_7A => X"0000006800000000000000680000000000000039000000000000004700000000",
            INIT_7B => X"0000009c00000000000000bb000000000000005d000000000000008700000000",
            INIT_7C => X"0000003b000000000000007c0000000000000047000000000000008300000000",
            INIT_7D => X"00000047000000000000004500000000000000a6000000000000005a00000000",
            INIT_7E => X"000000830000000000000079000000000000004a000000000000003900000000",
            INIT_7F => X"0000007f00000000000000bb00000000000000a3000000000000005b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE38;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE39 : if BRAM_NAME = "samplegold_layersamples_instance39" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a4000000000000008e00000000000000a1000000000000007a00000000",
            INIT_01 => X"0000001a0000000000000019000000000000002d000000000000008d00000000",
            INIT_02 => X"0000006f000000000000007c000000000000004d000000000000002d00000000",
            INIT_03 => X"0000007700000000000000a400000000000000bb00000000000000bf00000000",
            INIT_04 => X"0000009300000000000000a300000000000000ae000000000000007400000000",
            INIT_05 => X"0000004100000000000000410000000000000053000000000000006d00000000",
            INIT_06 => X"000000b2000000000000007b0000000000000056000000000000006200000000",
            INIT_07 => X"0000007c00000000000000a000000000000000a1000000000000009900000000",
            INIT_08 => X"0000008e00000000000000b300000000000000bf000000000000009f00000000",
            INIT_09 => X"0000009200000000000000a2000000000000008b000000000000008d00000000",
            INIT_0A => X"000000d100000000000000ae0000000000000088000000000000009b00000000",
            INIT_0B => X"000000cc00000000000000a900000000000000b300000000000000ae00000000",
            INIT_0C => X"000000a000000000000000b700000000000000a700000000000000c100000000",
            INIT_0D => X"000000aa00000000000000b000000000000000ba00000000000000b800000000",
            INIT_0E => X"0000003b00000000000000000000000000000000000000000000009200000000",
            INIT_0F => X"00000052000000000000004b000000000000003b000000000000003a00000000",
            INIT_10 => X"00000010000000000000001c0000000000000010000000000000002e00000000",
            INIT_11 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_12 => X"000000270000000000000029000000000000001e000000000000000600000000",
            INIT_13 => X"0000005000000000000000470000000000000034000000000000004100000000",
            INIT_14 => X"0000002e00000000000000250000000000000008000000000000002d00000000",
            INIT_15 => X"00000000000000000000000b000000000000000e000000000000001900000000",
            INIT_16 => X"000000360000000000000042000000000000001f000000000000001700000000",
            INIT_17 => X"0000004000000000000000630000000000000044000000000000004600000000",
            INIT_18 => X"0000003600000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000c00000000000000000000000000000009000000000000003b00000000",
            INIT_1A => X"00000064000000000000003a000000000000003b000000000000003100000000",
            INIT_1B => X"000000450000000000000067000000000000005d000000000000006500000000",
            INIT_1C => X"0000002000000000000000330000000000000018000000000000001a00000000",
            INIT_1D => X"0000001a0000000000000008000000000000001f000000000000002000000000",
            INIT_1E => X"0000001300000000000000540000000000000039000000000000002d00000000",
            INIT_1F => X"00000043000000000000007d0000000000000011000000000000000000000000",
            INIT_20 => X"000000240000000000000034000000000000002e000000000000001e00000000",
            INIT_21 => X"0000001c00000000000000000000000000000000000000000000004600000000",
            INIT_22 => X"0000004700000000000000000000000000000000000000000000004600000000",
            INIT_23 => X"000000210000000000000025000000000000001b000000000000002b00000000",
            INIT_24 => X"000000000000000000000029000000000000002a000000000000002a00000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000003500000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000002b0000000000000000000000000000002b000000000000000f00000000",
            INIT_29 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_2D => X"000000110000000000000008000000000000001e000000000000000000000000",
            INIT_2E => X"0000009000000000000000990000000000000076000000000000008900000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000002500000000",
            INIT_30 => X"000000000000000000000000000000000000001b000000000000002400000000",
            INIT_31 => X"00000000000000000000001f000000000000001700000000000000bb00000000",
            INIT_32 => X"000000000000000000000000000000000000002a000000000000000000000000",
            INIT_33 => X"0000001d00000000000000000000000000000000000000000000001300000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000003a00000000",
            INIT_35 => X"000000a100000000000000bc0000000000000089000000000000009100000000",
            INIT_36 => X"00000000000000000000002f000000000000003a000000000000002900000000",
            INIT_37 => X"0000001300000000000000430000000000000000000000000000004500000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_39 => X"000000060000000000000004000000000000001c000000000000000000000000",
            INIT_3A => X"0000005a0000000000000034000000000000001c000000000000000000000000",
            INIT_3B => X"00000000000000000000002d000000000000002f000000000000002d00000000",
            INIT_3C => X"0000001100000000000000270000000000000000000000000000004e00000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000003300000000000000080000000000000000000000000000000000000000",
            INIT_3F => X"00000021000000000000002c0000000000000052000000000000003e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000020000000000000002a0000000000000000000000000000003200000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000001d000000000000001a0000000000000000000000000000000000000000",
            INIT_43 => X"000000000000000000000006000000000000001a000000000000000000000000",
            INIT_44 => X"0000003a0000000000000059000000000000004d000000000000000900000000",
            INIT_45 => X"0000000d00000000000000230000000000000028000000000000002f00000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_65 => X"00000000000000000000004b0000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000020000000000000000100000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000003500000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"00000000000000000000003f0000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000140000000000000019000000000000001200000000",
            INIT_73 => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"00000000000000000000000a000000000000001a000000000000000c00000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000004e0000000000000056000000000000004a000000000000004b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE39;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE40 : if BRAM_NAME = "samplegold_layersamples_instance40" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002200000000000000260000000000000036000000000000004b00000000",
            INIT_01 => X"000000000000000000000009000000000000000d000000000000000000000000",
            INIT_02 => X"0000006f000000000000006c000000000000000b000000000000002000000000",
            INIT_03 => X"00000055000000000000005f000000000000005b000000000000004000000000",
            INIT_04 => X"0000000000000000000000240000000000000044000000000000004900000000",
            INIT_05 => X"0000002900000000000000270000000000000018000000000000000c00000000",
            INIT_06 => X"0000005d000000000000006b0000000000000078000000000000000c00000000",
            INIT_07 => X"0000005b00000000000000640000000000000068000000000000006300000000",
            INIT_08 => X"0000002500000000000000130000000000000041000000000000004900000000",
            INIT_09 => X"000000220000000000000020000000000000002d000000000000001900000000",
            INIT_0A => X"0000006900000000000000660000000000000071000000000000003b00000000",
            INIT_0B => X"0000004c00000000000000690000000000000066000000000000007600000000",
            INIT_0C => X"0000002f00000000000000340000000000000053000000000000005900000000",
            INIT_0D => X"000000470000000000000029000000000000001b000000000000001800000000",
            INIT_0E => X"000000740000000000000065000000000000006d000000000000006800000000",
            INIT_0F => X"00000055000000000000005e000000000000005d000000000000006c00000000",
            INIT_10 => X"000000180000000000000046000000000000004d000000000000005800000000",
            INIT_11 => X"0000005e0000000000000000000000000000002a000000000000002500000000",
            INIT_12 => X"0000005700000000000000680000000000000079000000000000007c00000000",
            INIT_13 => X"0000004700000000000000440000000000000087000000000000008a00000000",
            INIT_14 => X"0000001400000000000000140000000000000008000000000000005700000000",
            INIT_15 => X"0000009200000000000000580000000000000048000000000000002500000000",
            INIT_16 => X"0000006000000000000000a6000000000000004a000000000000007f00000000",
            INIT_17 => X"0000004100000000000000620000000000000058000000000000004100000000",
            INIT_18 => X"0000002200000000000000110000000000000000000000000000000000000000",
            INIT_19 => X"00000066000000000000008b0000000000000059000000000000002b00000000",
            INIT_1A => X"0000008f00000000000000760000000000000094000000000000008500000000",
            INIT_1B => X"0000000600000000000000650000000000000085000000000000008e00000000",
            INIT_1C => X"00000040000000000000001d000000000000002a000000000000000000000000",
            INIT_1D => X"000000b6000000000000005e000000000000008a000000000000005800000000",
            INIT_1E => X"0000007c000000000000007e00000000000000a1000000000000005d00000000",
            INIT_1F => X"0000000000000000000000000000000000000031000000000000007800000000",
            INIT_20 => X"0000005d00000000000000440000000000000031000000000000004900000000",
            INIT_21 => X"0000007e00000000000000530000000000000072000000000000009700000000",
            INIT_22 => X"0000000000000000000000540000000000000065000000000000005a00000000",
            INIT_23 => X"0000004d00000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000009200000000000000540000000000000062000000000000006400000000",
            INIT_25 => X"0000001f000000000000001e0000000000000000000000000000002200000000",
            INIT_26 => X"000000000000000000000000000000000000001d000000000000005f00000000",
            INIT_27 => X"0000007900000000000000520000000000000000000000000000000000000000",
            INIT_28 => X"0000003b00000000000000550000000000000062000000000000004000000000",
            INIT_29 => X"0000001a00000000000000150000000000000000000000000000001400000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000004e00000000000000510000000000000030000000000000000000000000",
            INIT_2C => X"0000004a000000000000005f0000000000000058000000000000005400000000",
            INIT_2D => X"00000000000000000000001e0000000000000032000000000000004400000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000004600000000000000610000000000000048000000000000000000000000",
            INIT_30 => X"0000003400000000000000470000000000000035000000000000005f00000000",
            INIT_31 => X"0000001b000000000000001c0000000000000045000000000000005700000000",
            INIT_32 => X"0000001c00000000000000080000000000000016000000000000000000000000",
            INIT_33 => X"000000490000000000000063000000000000003c000000000000002600000000",
            INIT_34 => X"0000005500000000000000630000000000000038000000000000004700000000",
            INIT_35 => X"0000003b00000000000000290000000000000040000000000000004900000000",
            INIT_36 => X"0000001c000000000000003a0000000000000041000000000000004600000000",
            INIT_37 => X"0000002c00000000000000000000000000000085000000000000000000000000",
            INIT_38 => X"0000000e00000000000000000000000000000010000000000000000100000000",
            INIT_39 => X"00000016000000000000000e0000000000000000000000000000000000000000",
            INIT_3A => X"0000000700000000000000000000000000000041000000000000001e00000000",
            INIT_3B => X"0000001200000000000000010000000000000000000000000000000000000000",
            INIT_3C => X"00000000000000000000001e0000000000000006000000000000001700000000",
            INIT_3D => X"0000002100000000000000040000000000000022000000000000000000000000",
            INIT_3E => X"0000001b00000000000000000000000000000000000000000000000600000000",
            INIT_3F => X"0000000000000000000000080000000000000000000000000000000700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001300000000000000040000000000000007000000000000000500000000",
            INIT_41 => X"0000000000000000000000180000000000000009000000000000006d00000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_44 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_45 => X"0000001000000000000000340000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000021000000000000000000000000",
            INIT_47 => X"0000003e00000000000000000000000000000001000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000019000000000000000000000000",
            INIT_49 => X"0000002900000000000000080000000000000000000000000000002500000000",
            INIT_4A => X"0000000000000000000000000000000000000042000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000003e00000000",
            INIT_4C => X"0000002600000000000000000000000000000000000000000000002b00000000",
            INIT_4D => X"0000000000000000000000e0000000000000001b000000000000000900000000",
            INIT_4E => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000004300000000000000900000000000000004000000000000000000000000",
            INIT_50 => X"0000002e00000000000000200000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000720000000000000000000000000000001400000000",
            INIT_52 => X"000000000000000000000000000000000000002a000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_54 => X"00000000000000000000005f0000000000000000000000000000000000000000",
            INIT_55 => X"000000000000000000000000000000000000005b000000000000001400000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000004100000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"000000000000000000000000000000000000005d000000000000005400000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000006c00000000",
            INIT_5A => X"0000000000000000000000830000000000000000000000000000000000000000",
            INIT_5B => X"00000040000000000000004a0000000000000010000000000000000000000000",
            INIT_5C => X"0000001800000000000000000000000000000000000000000000007f00000000",
            INIT_5D => X"0000000000000000000000740000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_5F => X"00000051000000000000004e0000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000410000000000000000000000000000000000000000",
            INIT_61 => X"0000006200000000000000580000000000000000000000000000001d00000000",
            INIT_62 => X"0000000d000000000000000e0000000000000000000000000000000000000000",
            INIT_63 => X"000000000000000000000012000000000000001e000000000000002600000000",
            INIT_64 => X"00000000000000000000000d0000000000000000000000000000002100000000",
            INIT_65 => X"00000007000000000000002a0000000000000000000000000000000000000000",
            INIT_66 => X"0000004f0000000000000033000000000000002a000000000000001700000000",
            INIT_67 => X"00000012000000000000005c0000000000000000000000000000006600000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000001a00000000000000000000000000000033000000000000003300000000",
            INIT_6A => X"00000034000000000000006e0000000000000021000000000000002300000000",
            INIT_6B => X"0000006400000000000000000000000000000000000000000000006300000000",
            INIT_6C => X"0000001e00000000000000010000000000000027000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_6E => X"0000000000000000000000020000000000000019000000000000002700000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000003500000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000001c000000000000001f0000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000b00000000000000000000000000000000000000000000000f00000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE40;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE41 : if BRAM_NAME = "samplegold_layersamples_instance41" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000010000000000000002000000000000000000000000",
            INIT_02 => X"0000000000000000000000050000000000000000000000000000007900000000",
            INIT_03 => X"0000004f0000000000000000000000000000000a000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000002400000000000000050000000000000000000000000000003b00000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000008000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_0B => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_0C => X"0000000f00000000000000080000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000130000000000000000000000000000000000000000",
            INIT_0E => X"000000000000000000000008000000000000004b000000000000000000000000",
            INIT_0F => X"0000003f000000000000003b0000000000000047000000000000003f00000000",
            INIT_10 => X"00000000000000000000003f0000000000000017000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000063000000000000000000000000",
            INIT_12 => X"0000005d0000000000000000000000000000000000000000000001b900000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000082000000000000002700000000",
            INIT_15 => X"000000000000000000000000000000000000000d000000000000002300000000",
            INIT_16 => X"00000031000000000000007d0000000000000056000000000000009200000000",
            INIT_17 => X"00000000000000000000005b0000000000000020000000000000000000000000",
            INIT_18 => X"000000000000000000000000000000000000000000000000000000b000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000004500000000",
            INIT_1A => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"00000008000000000000004d000000000000000e000000000000000700000000",
            INIT_1C => X"000000000000000000000010000000000000000000000000000000b200000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000009e00000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"000000380000000000000000000000000000000f000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000025000000000000000000000000",
            INIT_21 => X"0000000000000000000000210000000000000000000000000000003000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000002600000000000000410000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000004f00000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000003f00000000000000380000000000000037000000000000003e00000000",
            INIT_61 => X"0000001d00000000000000350000000000000047000000000000003e00000000",
            INIT_62 => X"000000190000000000000006000000000000000a000000000000001000000000",
            INIT_63 => X"000000440000000000000046000000000000000b000000000000000c00000000",
            INIT_64 => X"000000510000000000000045000000000000003e000000000000004f00000000",
            INIT_65 => X"0000001300000000000000300000000000000040000000000000004600000000",
            INIT_66 => X"00000001000000000000000d0000000000000018000000000000001000000000",
            INIT_67 => X"00000046000000000000004d000000000000001b000000000000001b00000000",
            INIT_68 => X"0000004800000000000000530000000000000048000000000000004f00000000",
            INIT_69 => X"00000025000000000000002d0000000000000057000000000000005500000000",
            INIT_6A => X"0000000f00000000000000180000000000000000000000000000000d00000000",
            INIT_6B => X"0000004f0000000000000048000000000000002f000000000000003f00000000",
            INIT_6C => X"0000004500000000000000470000000000000053000000000000004e00000000",
            INIT_6D => X"00000023000000000000002f0000000000000047000000000000004200000000",
            INIT_6E => X"0000002700000000000000100000000000000016000000000000000b00000000",
            INIT_6F => X"0000005d00000000000000460000000000000045000000000000004200000000",
            INIT_70 => X"0000001a00000000000000260000000000000027000000000000003600000000",
            INIT_71 => X"0000001e0000000000000011000000000000003d000000000000003a00000000",
            INIT_72 => X"00000016000000000000006d000000000000000c000000000000000d00000000",
            INIT_73 => X"0000006400000000000000410000000000000044000000000000004c00000000",
            INIT_74 => X"000000160000000000000019000000000000000c000000000000000000000000",
            INIT_75 => X"00000015000000000000000e000000000000000e000000000000000400000000",
            INIT_76 => X"00000021000000000000004c000000000000000c000000000000001100000000",
            INIT_77 => X"0000003c0000000000000018000000000000004f000000000000002100000000",
            INIT_78 => X"0000000000000000000000050000000000000012000000000000000600000000",
            INIT_79 => X"0000000400000000000000190000000000000009000000000000000000000000",
            INIT_7A => X"0000002e000000000000001e0000000000000030000000000000000000000000",
            INIT_7B => X"0000001900000000000000320000000000000038000000000000002f00000000",
            INIT_7C => X"0000000000000000000000000000000000000009000000000000001000000000",
            INIT_7D => X"0000001e0000000000000000000000000000001a000000000000001400000000",
            INIT_7E => X"000000050000000000000017000000000000001f000000000000000f00000000",
            INIT_7F => X"0000001b00000000000000180000000000000012000000000000003b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE41;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE42 : if BRAM_NAME = "samplegold_layersamples_instance42" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002000000000000000050000000000000000000000000000000300000000",
            INIT_01 => X"0000002c00000000000000000000000000000000000000000000001800000000",
            INIT_02 => X"0000000800000000000000380000000000000000000000000000000800000000",
            INIT_03 => X"000000020000000000000000000000000000002a000000000000001f00000000",
            INIT_04 => X"0000002a000000000000000f0000000000000000000000000000000f00000000",
            INIT_05 => X"00000000000000000000001b0000000000000004000000000000000000000000",
            INIT_06 => X"0000000c00000000000000010000000000000000000000000000000000000000",
            INIT_07 => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_08 => X"0000000000000000000000230000000000000007000000000000001200000000",
            INIT_09 => X"0000003c000000000000001b0000000000000000000000000000001800000000",
            INIT_0A => X"0000000000000000000000090000000000000024000000000000001000000000",
            INIT_0B => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_0C => X"0000001e00000000000000270000000000000009000000000000001f00000000",
            INIT_0D => X"000000390000000000000038000000000000000a000000000000000e00000000",
            INIT_0E => X"0000000500000000000000140000000000000016000000000000000000000000",
            INIT_0F => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_10 => X"0000001e00000000000000000000000000000000000000000000000a00000000",
            INIT_11 => X"00000017000000000000001d000000000000000b000000000000001000000000",
            INIT_12 => X"0000000e0000000000000020000000000000000a000000000000000d00000000",
            INIT_13 => X"00000016000000000000001a0000000000000019000000000000001f00000000",
            INIT_14 => X"0000001900000000000000020000000000000022000000000000000000000000",
            INIT_15 => X"0000001100000000000000070000000000000017000000000000001900000000",
            INIT_16 => X"0000001b0000000000000019000000000000000e000000000000001700000000",
            INIT_17 => X"00000029000000000000000f0000000000000018000000000000001e00000000",
            INIT_18 => X"0000015600000000000001580000000000000155000000000000015e00000000",
            INIT_19 => X"00000137000000000000013a0000000000000149000000000000015a00000000",
            INIT_1A => X"000000dd0000000000000107000000000000010a000000000000011f00000000",
            INIT_1B => X"0000015600000000000000e60000000000000084000000000000004b00000000",
            INIT_1C => X"0000015300000000000001610000000000000155000000000000014600000000",
            INIT_1D => X"0000011800000000000001230000000000000132000000000000013c00000000",
            INIT_1E => X"00000085000000000000008e00000000000000e0000000000000010900000000",
            INIT_1F => X"0000013e00000000000001090000000000000103000000000000009700000000",
            INIT_20 => X"0000012f000000000000012f0000000000000140000000000000014500000000",
            INIT_21 => X"000001090000000000000110000000000000011a000000000000012d00000000",
            INIT_22 => X"000000b60000000000000082000000000000004d000000000000003800000000",
            INIT_23 => X"0000012d0000000000000130000000000000012900000000000000f000000000",
            INIT_24 => X"0000013200000000000001380000000000000130000000000000012b00000000",
            INIT_25 => X"0000005800000000000000c100000000000000fc000000000000011400000000",
            INIT_26 => X"0000011000000000000000fc00000000000000ee000000000000006200000000",
            INIT_27 => X"00000137000000000000013c000000000000013c000000000000012c00000000",
            INIT_28 => X"000000ef00000000000000c900000000000000fa000000000000013300000000",
            INIT_29 => X"00000029000000000000004600000000000000a000000000000000d700000000",
            INIT_2A => X"0000013e00000000000000f900000000000000f800000000000000c000000000",
            INIT_2B => X"0000010f000000000000012e0000000000000135000000000000013d00000000",
            INIT_2C => X"000000000000000000000000000000000000000000000000000000ab00000000",
            INIT_2D => X"0000002600000000000000390000000000000000000000000000000000000000",
            INIT_2E => X"00000141000000000000013a00000000000000ef00000000000000ba00000000",
            INIT_2F => X"0000003000000000000000700000000000000112000000000000013300000000",
            INIT_30 => X"0000000000000000000000780000000000000075000000000000005800000000",
            INIT_31 => X"00000048000000000000000c0000000000000089000000000000000000000000",
            INIT_32 => X"000000d00000000000000139000000000000013c00000000000000a900000000",
            INIT_33 => X"00000032000000000000002e000000000000004f000000000000006e00000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000003e00000000",
            INIT_35 => X"0000003200000000000000280000000000000079000000000000003b00000000",
            INIT_36 => X"00000029000000000000003e00000000000000fb000000000000013f00000000",
            INIT_37 => X"0000000000000000000000000000000000000003000000000000002200000000",
            INIT_38 => X"000000fb00000000000000210000000000000000000000000000000000000000",
            INIT_39 => X"0000011c00000000000000000000000000000000000000000000009d00000000",
            INIT_3A => X"0000004b0000000000000012000000000000002f000000000000001a00000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_3D => X"00000000000000000000008f0000000000000000000000000000000000000000",
            INIT_3E => X"0000000100000000000000450000000000000020000000000000005600000000",
            INIT_3F => X"0000008d00000000000000010000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000300000000000000000000000000000000000000000000000300000000",
            INIT_41 => X"00000011000000000000002200000000000000ad000000000000007700000000",
            INIT_42 => X"0000000000000000000000000000000000000012000000000000003e00000000",
            INIT_43 => X"0000003700000000000000270000000000000076000000000000000000000000",
            INIT_44 => X"0000005f0000000000000055000000000000000b000000000000000000000000",
            INIT_45 => X"000000360000000000000000000000000000001b000000000000009300000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000700000000000000350000000000000001000000000000006e00000000",
            INIT_48 => X"0000009b00000000000000420000000000000074000000000000000000000000",
            INIT_49 => X"00000000000000000000000a0000000000000000000000000000002e00000000",
            INIT_4A => X"00000084000000000000001a0000000000000004000000000000000700000000",
            INIT_4B => X"0000002300000000000000410000000000000055000000000000000000000000",
            INIT_4C => X"0000004a00000000000000880000000000000029000000000000005400000000",
            INIT_4D => X"0000000a00000000000000050000000000000013000000000000002b00000000",
            INIT_4E => X"000000020000000000000031000000000000002c000000000000001800000000",
            INIT_4F => X"0000002000000000000000270000000000000049000000000000002500000000",
            INIT_50 => X"0000002800000000000000230000000000000008000000000000001300000000",
            INIT_51 => X"000000230000000000000027000000000000002b000000000000003000000000",
            INIT_52 => X"0000002d0000000000000088000000000000002e000000000000001900000000",
            INIT_53 => X"0000000200000000000000130000000000000016000000000000000000000000",
            INIT_54 => X"00000020000000000000001e0000000000000000000000000000000000000000",
            INIT_55 => X"0000000c00000000000000140000000000000013000000000000001800000000",
            INIT_56 => X"0000000000000000000000000000000000000001000000000000000c00000000",
            INIT_57 => X"0000003e00000000000000000000000000000000000000000000000600000000",
            INIT_58 => X"000000100000000000000014000000000000001e000000000000005100000000",
            INIT_59 => X"0000000000000000000000000000000000000006000000000000000300000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000600000000000000120000000000000004000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"000000390000000000000029000000000000003b000000000000005200000000",
            INIT_5F => X"0000000c00000000000000080000000000000005000000000000000f00000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000700000000000000050000000000000001000000000000000b00000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000067000000000000004a00000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_67 => X"000000000000000000000000000000000000000b000000000000000600000000",
            INIT_68 => X"0000009600000000000000fc00000000000000d8000000000000009900000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000200000000000000080000000000000000000000000000004200000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000077000000000000000000000000",
            INIT_6E => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_6F => X"00000000000000000000003f000000000000004c000000000000000b00000000",
            INIT_70 => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_72 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000019000000000000002b00000000",
            INIT_74 => X"00000000000000000000008900000000000000cb000000000000000000000000",
            INIT_75 => X"00000000000000000000004b0000000000000000000000000000000000000000",
            INIT_76 => X"0000000300000000000000120000000000000000000000000000011e00000000",
            INIT_77 => X"000000a300000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000003f00000000000000c200000000000000fc00000000000000d900000000",
            INIT_79 => X"0000000000000000000000290000000000000106000000000000008000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"00000000000000000000003c0000000000000000000000000000000000000000",
            INIT_7C => X"0000006e00000000000000050000000000000093000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE42;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE43 : if BRAM_NAME = "samplegold_layersamples_instance43" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000019000000000000005f000000000000009e000000000000001700000000",
            INIT_01 => X"0000009b00000000000000ab0000000000000024000000000000000000000000",
            INIT_02 => X"000001d100000000000001c500000000000001b4000000000000013700000000",
            INIT_03 => X"0000000f0000000000000034000000000000002a00000000000000e800000000",
            INIT_04 => X"000000000000000000000000000000000000001f00000000000000ac00000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"00000000000000000000000f0000000000000048000000000000005700000000",
            INIT_08 => X"0000009d00000000000000ae0000000000000000000000000000000000000000",
            INIT_09 => X"00000087000000000000008500000000000000a4000000000000009b00000000",
            INIT_0A => X"00000040000000000000008c000000000000006b000000000000008a00000000",
            INIT_0B => X"000000340000000000000000000000000000005b000000000000005100000000",
            INIT_0C => X"000000720000000000000077000000000000009d000000000000003900000000",
            INIT_0D => X"000000720000000000000071000000000000007b000000000000008500000000",
            INIT_0E => X"0000006b000000000000005a0000000000000065000000000000006300000000",
            INIT_0F => X"0000003e00000000000000560000000000000000000000000000000100000000",
            INIT_10 => X"0000006a000000000000006e0000000000000064000000000000007000000000",
            INIT_11 => X"0000005f00000000000000670000000000000067000000000000007100000000",
            INIT_12 => X"0000000000000000000000340000000000000079000000000000006200000000",
            INIT_13 => X"0000005f000000000000002c000000000000003d000000000000000600000000",
            INIT_14 => X"000000730000000000000068000000000000006e000000000000007100000000",
            INIT_15 => X"0000005600000000000000540000000000000068000000000000007200000000",
            INIT_16 => X"0000004a000000000000005c0000000000000000000000000000006e00000000",
            INIT_17 => X"0000007600000000000000670000000000000045000000000000005000000000",
            INIT_18 => X"0000006b0000000000000083000000000000006f000000000000007600000000",
            INIT_19 => X"000000000000000000000049000000000000005e000000000000004f00000000",
            INIT_1A => X"0000003a00000000000000070000000000000019000000000000000000000000",
            INIT_1B => X"0000006a00000000000000740000000000000076000000000000004e00000000",
            INIT_1C => X"00000017000000000000007a0000000000000093000000000000006700000000",
            INIT_1D => X"000000000000000000000008000000000000003a000000000000001300000000",
            INIT_1E => X"0000003e0000000000000000000000000000006a000000000000000000000000",
            INIT_1F => X"0000008100000000000000590000000000000071000000000000007700000000",
            INIT_20 => X"000000000000000000000000000000000000004d000000000000006700000000",
            INIT_21 => X"000000000000000000000001000000000000014b000000000000000000000000",
            INIT_22 => X"0000007a000000000000001a0000000000000000000000000000000000000000",
            INIT_23 => X"000000000000000000000025000000000000008f000000000000006e00000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000004200000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000003e00000000",
            INIT_26 => X"0000009d00000000000000720000000000000000000000000000005400000000",
            INIT_27 => X"000000360000000000000000000000000000001f000000000000000b00000000",
            INIT_28 => X"0000000000000000000000000000000000000035000000000000010e00000000",
            INIT_29 => X"0000005b00000000000000230000000000000000000000000000000000000000",
            INIT_2A => X"00000000000000000000008500000000000000cb000000000000000000000000",
            INIT_2B => X"0000017400000000000000740000000000000000000000000000002800000000",
            INIT_2C => X"0000006000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000042000000000000015700000000",
            INIT_2F => X"0000000000000000000001220000000000000058000000000000000000000000",
            INIT_30 => X"000000f900000000000000510000000000000000000000000000000000000000",
            INIT_31 => X"000000a900000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000002e00000000000000000000000000000000000000000000004700000000",
            INIT_33 => X"00000000000000000000000000000000000000ee000000000000003d00000000",
            INIT_34 => X"00000000000000000000011e0000000000000000000000000000000000000000",
            INIT_35 => X"000000260000000000000083000000000000000d000000000000000000000000",
            INIT_36 => X"0000000000000000000000530000000000000000000000000000000000000000",
            INIT_37 => X"0000004400000000000000000000000000000000000000000000003300000000",
            INIT_38 => X"00000000000000000000003d0000000000000030000000000000000000000000",
            INIT_39 => X"00000000000000000000003f000000000000004e000000000000002500000000",
            INIT_3A => X"000000470000000000000049000000000000006b000000000000001a00000000",
            INIT_3B => X"0000000000000000000000590000000000000000000000000000003900000000",
            INIT_3C => X"000000160000000000000000000000000000000f000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"000000000000000000000000000000000000005b000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000000000000000000001a0000000000000001000000000000000000000000",
            INIT_41 => X"0000000700000000000000020000000000000000000000000000000000000000",
            INIT_42 => X"0000000d000000000000000a0000000000000010000000000000000f00000000",
            INIT_43 => X"0000000000000000000000000000000000000022000000000000006f00000000",
            INIT_44 => X"0000000c00000000000000300000000000000000000000000000002300000000",
            INIT_45 => X"0000001000000000000000150000000000000015000000000000000800000000",
            INIT_46 => X"000000000000000000000009000000000000000d000000000000000f00000000",
            INIT_47 => X"000000000000000000000011000000000000000d000000000000002b00000000",
            INIT_48 => X"00000021000000000000002e0000000000000000000000000000000000000000",
            INIT_49 => X"0000000e000000000000000c0000000000000015000000000000001400000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_4B => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_4C => X"000000020000000000000000000000000000000a000000000000002100000000",
            INIT_4D => X"00000012000000000000000c0000000000000000000000000000000000000000",
            INIT_4E => X"0000004a00000000000000210000000000000000000000000000000100000000",
            INIT_4F => X"00000000000000000000000d0000000000000005000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000bd00000000000000330000000000000000000000000000000000000000",
            INIT_52 => X"000000040000000000000000000000000000003f00000000000000b900000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_54 => X"0000007200000000000000150000000000000001000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"00000000000000000000001d0000000000000012000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_58 => X"000000a200000000000000000000000000000000000000000000000e00000000",
            INIT_59 => X"0000000f00000000000000db00000000000000a000000000000000f300000000",
            INIT_5A => X"0000000300000000000000040000000000000023000000000000000000000000",
            INIT_5B => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_5C => X"000000cf00000000000000070000000000000000000000000000005600000000",
            INIT_5D => X"000000000000000000000000000000000000000000000000000000c500000000",
            INIT_5E => X"00000000000000000000001c000000000000001e000000000000000000000000",
            INIT_5F => X"0000000000000000000000440000000000000060000000000000002a00000000",
            INIT_60 => X"0000000000000000000000000000000000000076000000000000004c00000000",
            INIT_61 => X"0000009500000000000000fe000000000000001a000000000000000500000000",
            INIT_62 => X"00000000000000000000002a0000000000000000000000000000000000000000",
            INIT_63 => X"00000000000000000000000a0000000000000018000000000000000000000000",
            INIT_64 => X"000000000000000000000005000000000000000d000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000003d0000000000000042000000000000001a000000000000000000000000",
            INIT_68 => X"000000bc00000000000000d00000000000000000000000000000000000000000",
            INIT_69 => X"0000003400000000000000000000000000000000000000000000002f00000000",
            INIT_6A => X"0000000a00000000000000000000000000000030000000000000000600000000",
            INIT_6B => X"0000000000000000000000050000000000000000000000000000000e00000000",
            INIT_6C => X"0000002a00000000000000250000000000000010000000000000000000000000",
            INIT_6D => X"0000001900000000000000120000000000000006000000000000000200000000",
            INIT_6E => X"00000047000000000000004b0000000000000001000000000000000000000000",
            INIT_6F => X"00000000000000000000004b000000000000002f000000000000003e00000000",
            INIT_70 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_71 => X"0000000000000000000000010000000000000001000000000000000b00000000",
            INIT_72 => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000025000000000000001200000000",
            INIT_74 => X"0000002800000000000000560000000000000019000000000000005100000000",
            INIT_75 => X"00000096000000000000002c0000000000000000000000000000000000000000",
            INIT_76 => X"00000015000000000000000d0000000000000001000000000000001600000000",
            INIT_77 => X"0000000000000000000000250000000000000022000000000000001d00000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_79 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"000000130000000000000000000000000000000b000000000000001300000000",
            INIT_7B => X"0000000000000000000000000000000000000039000000000000000800000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000009900000000",
            INIT_7D => X"00000009000000000000000a0000000000000021000000000000000000000000",
            INIT_7E => X"0000000000000000000000010000000000000000000000000000000900000000",
            INIT_7F => X"0000000c000000000000003c0000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE43;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE44 : if BRAM_NAME = "samplegold_layersamples_instance44" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002b00000000000000410000000000000000000000000000000000000000",
            INIT_01 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000053000000000000001000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"000000d600000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000010d00000000000000870000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000a50000000000000000000000000000012100000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"000000af00000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000041000000000000005600000000",
            INIT_12 => X"0000003300000000000000400000000000000027000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"000000410000000000000000000000000000000b000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"000000000000000000000000000000000000000a000000000000018400000000",
            INIT_17 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_18 => X"000000000000000000000000000000000000000000000000000000c700000000",
            INIT_19 => X"0000002000000000000000470000000000000000000000000000004200000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"00000065000000000000000000000000000000dc000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000073000000000000010100000000",
            INIT_1E => X"000001720000000000000000000000000000004a000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000032000000000000002f00000000",
            INIT_20 => X"0000005d00000000000000c50000000000000000000000000000000000000000",
            INIT_21 => X"0000005800000000000000690000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000016000000000000013b00000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000008100000000",
            INIT_24 => X"0000000000000000000000000000000000000158000000000000000000000000",
            INIT_25 => X"0000000000000000000001150000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"000000000000000000000000000000000000000000000000000000bb00000000",
            INIT_29 => X"00000000000000000000000000000000000000b0000000000000000900000000",
            INIT_2A => X"000000a70000000000000077000000000000009d000000000000001d00000000",
            INIT_2B => X"000000cf00000000000000df00000000000000d900000000000000ce00000000",
            INIT_2C => X"0000005b00000000000000400000000000000042000000000000000000000000",
            INIT_2D => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000024000000000000007200000000",
            INIT_31 => X"0000008700000000000000900000000000000080000000000000000000000000",
            INIT_32 => X"000000740000000000000088000000000000009b000000000000008e00000000",
            INIT_33 => X"0000005e00000000000000420000000000000056000000000000008b00000000",
            INIT_34 => X"0000005000000000000000000000000000000056000000000000003c00000000",
            INIT_35 => X"0000007d0000000000000084000000000000008d000000000000007a00000000",
            INIT_36 => X"0000006b0000000000000060000000000000006a000000000000007100000000",
            INIT_37 => X"0000005700000000000000370000000000000061000000000000005900000000",
            INIT_38 => X"0000005d00000000000000570000000000000000000000000000004d00000000",
            INIT_39 => X"000000500000000000000060000000000000005d000000000000006200000000",
            INIT_3A => X"0000005600000000000000590000000000000056000000000000005700000000",
            INIT_3B => X"0000002b0000000000000043000000000000002e000000000000003b00000000",
            INIT_3C => X"0000004600000000000000490000000000000067000000000000002200000000",
            INIT_3D => X"00000051000000000000004c0000000000000054000000000000004b00000000",
            INIT_3E => X"0000004000000000000000520000000000000063000000000000005800000000",
            INIT_3F => X"0000004d000000000000003c0000000000000000000000000000006400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004a00000000000000490000000000000042000000000000005700000000",
            INIT_41 => X"00000041000000000000004e000000000000003e000000000000005400000000",
            INIT_42 => X"0000007400000000000000a00000000000000034000000000000003800000000",
            INIT_43 => X"0000004800000000000000530000000000000055000000000000000000000000",
            INIT_44 => X"000000530000000000000054000000000000004d000000000000004800000000",
            INIT_45 => X"0000000800000000000000000000000000000000000000000000002200000000",
            INIT_46 => X"000000f5000000000000006c0000000000000000000000000000000000000000",
            INIT_47 => X"000000480000000000000043000000000000008b000000000000000000000000",
            INIT_48 => X"00000011000000000000002c0000000000000064000000000000004d00000000",
            INIT_49 => X"00000011000000000000000d000000000000001a000000000000000000000000",
            INIT_4A => X"0000000e00000000000001c40000000000000000000000000000000000000000",
            INIT_4B => X"0000005500000000000000450000000000000030000000000000000000000000",
            INIT_4C => X"000000000000000000000046000000000000003b000000000000000700000000",
            INIT_4D => X"000000000000000000000000000000000000002e000000000000002400000000",
            INIT_4E => X"0000000000000000000000de00000000000000ba000000000000000000000000",
            INIT_4F => X"0000001b0000000000000017000000000000004f000000000000001b00000000",
            INIT_50 => X"000000000000000000000000000000000000003c000000000000000000000000",
            INIT_51 => X"0000007300000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"000000000000000000000000000000000000000000000000000000d400000000",
            INIT_53 => X"0000000000000000000000f60000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000004f00000000",
            INIT_55 => X"000000b500000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"00000000000000000000003b0000000000000000000000000000000000000000",
            INIT_57 => X"00000031000000000000003c00000000000000e7000000000000000000000000",
            INIT_58 => X"000000a100000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000001c00000000000000000000000000000000000000000000005500000000",
            INIT_5A => X"000000000000000000000000000000000000006e000000000000003500000000",
            INIT_5B => X"0000000000000000000000000000000000000063000000000000001e00000000",
            INIT_5C => X"0000001000000000000001350000000000000000000000000000000000000000",
            INIT_5D => X"000000ac00000000000000000000000000000000000000000000002500000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000002500000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000005600000000",
            INIT_60 => X"0000007600000000000000000000000000000140000000000000000000000000",
            INIT_61 => X"0000000000000000000000a10000000000000000000000000000000000000000",
            INIT_62 => X"0000000100000000000000000000000000000000000000000000000d00000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000004200000000000000190000000000000000000000000000006a00000000",
            INIT_65 => X"000000150000000000000000000000000000002f000000000000000000000000",
            INIT_66 => X"0000000400000000000000490000000000000003000000000000002600000000",
            INIT_67 => X"0000001d00000000000000190000000000000012000000000000000f00000000",
            INIT_68 => X"0000001100000000000000510000000000000030000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_6A => X"00000016000000000000001b000000000000001b000000000000001200000000",
            INIT_6B => X"0000000500000000000000000000000000000011000000000000001d00000000",
            INIT_6C => X"00000052000000000000000b0000000000000003000000000000000000000000",
            INIT_6D => X"000000140000000000000000000000000000000e000000000000000000000000",
            INIT_6E => X"00000014000000000000001b0000000000000022000000000000001a00000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000001400000000000000260000000000000031000000000000005000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_73 => X"0000006f00000000000000070000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000001ad0000000000000164000000000000010400000000",
            INIT_7F => X"000000000000000000000000000000000000008b000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE44;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE45 : if BRAM_NAME = "samplegold_layersamples_instance45" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000049000000000000000800000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"000000000000000000000036000000000000005d000000000000000000000000",
            INIT_04 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_06 => X"0000001f00000000000000660000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000220000000000000041000000000000000000000000",
            INIT_09 => X"0000000700000000000000290000000000000004000000000000002900000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000006500000000000000340000000000000004000000000000000000000000",
            INIT_0D => X"000001aa000000000000009b0000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_0F => X"00000000000000000000002a0000000000000103000000000000003500000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_11 => X"0000010800000000000000000000000000000025000000000000000000000000",
            INIT_12 => X"0000000000000000000000670000000000000026000000000000003700000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000002400000000000000120000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000020000000000000012000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000004500000000000000530000000000000000000000000000000000000000",
            INIT_1A => X"0000006d00000000000000290000000000000000000000000000000900000000",
            INIT_1B => X"0000010e00000000000000eb00000000000000a100000000000000b200000000",
            INIT_1C => X"0000000000000000000000000000000000000102000000000000010a00000000",
            INIT_1D => X"00000000000000000000001e0000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000001f00000000000000730000000000000005000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000000000002c000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"000000000000000000000000000000000000004d000000000000008a00000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"000000550000000000000000000000000000000e000000000000001100000000",
            INIT_3B => X"000000000000000000000000000000000000000c00000000000000da00000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000005300000000000000210000000000000000000000000000000000000000",
            INIT_3E => X"000000840000000000000071000000000000005c000000000000003d00000000",
            INIT_3F => X"00000000000000000000001f0000000000000000000000000000004600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003900000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000004e00000000000000500000000000000000000000000000000100000000",
            INIT_42 => X"00000000000000000000003000000000000000a1000000000000005400000000",
            INIT_43 => X"0000000000000000000000000000000000000032000000000000001100000000",
            INIT_44 => X"000000000000000000000020000000000000001e000000000000007400000000",
            INIT_45 => X"0000004b0000000000000066000000000000006b000000000000000000000000",
            INIT_46 => X"0000005f000000000000005a0000000000000078000000000000000000000000",
            INIT_47 => X"0000009d00000000000000000000000000000000000000000000005000000000",
            INIT_48 => X"000000040000000000000022000000000000000b000000000000004800000000",
            INIT_49 => X"00000017000000000000003000000000000000b6000000000000007100000000",
            INIT_4A => X"0000002b00000000000000630000000000000079000000000000000000000000",
            INIT_4B => X"000000420000000000000084000000000000001d000000000000000000000000",
            INIT_4C => X"0000006d0000000000000022000000000000003d000000000000001300000000",
            INIT_4D => X"000000000000000000000028000000000000003100000000000000ba00000000",
            INIT_4E => X"000000000000000000000000000000000000007a000000000000006100000000",
            INIT_4F => X"0000003a000000000000004c000000000000006d000000000000002100000000",
            INIT_50 => X"000000b5000000000000006f0000000000000060000000000000008100000000",
            INIT_51 => X"0000002b000000000000000e000000000000005e000000000000001800000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000003f00000000",
            INIT_53 => X"0000001300000000000000160000000000000020000000000000003800000000",
            INIT_54 => X"0000002b000000000000003c0000000000000014000000000000001200000000",
            INIT_55 => X"0000000c000000000000000d0000000000000025000000000000003e00000000",
            INIT_56 => X"00000039000000000000000d0000000000000000000000000000000000000000",
            INIT_57 => X"00000032000000000000003a0000000000000033000000000000005600000000",
            INIT_58 => X"0000002d0000000000000000000000000000001b000000000000002c00000000",
            INIT_59 => X"0000000000000000000000060000000000000009000000000000001000000000",
            INIT_5A => X"000001ce00000000000001d800000000000001d600000000000001e900000000",
            INIT_5B => X"0000016a0000000000000186000000000000019300000000000001b500000000",
            INIT_5C => X"000000c9000000000000010a0000000000000115000000000000014c00000000",
            INIT_5D => X"000001a800000000000000cc0000000000000051000000000000006900000000",
            INIT_5E => X"0000015f000000000000017b0000000000000189000000000000018900000000",
            INIT_5F => X"0000011d000000000000012e0000000000000142000000000000014400000000",
            INIT_60 => X"00000038000000000000009800000000000000e9000000000000011100000000",
            INIT_61 => X"00000129000000000000013400000000000000eb000000000000009500000000",
            INIT_62 => X"000001200000000000000125000000000000012e000000000000012800000000",
            INIT_63 => X"0000010b00000000000001180000000000000120000000000000012400000000",
            INIT_64 => X"000000d5000000000000006d0000000000000012000000000000009600000000",
            INIT_65 => X"0000011b0000000000000114000000000000010400000000000000f300000000",
            INIT_66 => X"0000012b000000000000012b0000000000000123000000000000011900000000",
            INIT_67 => X"0000004d00000000000000ea0000000000000117000000000000012900000000",
            INIT_68 => X"000000f300000000000000fd00000000000000d2000000000000003000000000",
            INIT_69 => X"0000011f00000000000001210000000000000120000000000000010e00000000",
            INIT_6A => X"000000f600000000000000fa000000000000010d000000000000011f00000000",
            INIT_6B => X"00000045000000000000001000000000000000a700000000000000e300000000",
            INIT_6C => X"0000012000000000000000e900000000000000e400000000000000b800000000",
            INIT_6D => X"00000106000000000000011a000000000000011e000000000000011f00000000",
            INIT_6E => X"00000024000000000000002f000000000000005700000000000000b400000000",
            INIT_6F => X"00000008000000000000001e0000000000000010000000000000000000000000",
            INIT_70 => X"00000120000000000000012200000000000000d2000000000000009a00000000",
            INIT_71 => X"0000005d00000000000000a400000000000000f6000000000000011800000000",
            INIT_72 => X"0000000000000000000000140000000000000000000000000000001900000000",
            INIT_73 => X"0000002200000000000000100000000000000000000000000000001a00000000",
            INIT_74 => X"000000c30000000000000119000000000000011c000000000000007600000000",
            INIT_75 => X"0000001f00000000000000240000000000000032000000000000008b00000000",
            INIT_76 => X"0000000000000000000000430000000000000025000000000000001a00000000",
            INIT_77 => X"000000410000000000000018000000000000000a000000000000000000000000",
            INIT_78 => X"00000000000000000000006100000000000000e6000000000000011a00000000",
            INIT_79 => X"0000002e00000000000000000000000000000000000000000000000200000000",
            INIT_7A => X"0000000000000000000000270000000000000000000000000000000200000000",
            INIT_7B => X"000000f600000000000000320000000000000018000000000000004a00000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000008600000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000001600000000000000a50000000000000007000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE45;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE46 : if BRAM_NAME = "samplegold_layersamples_instance46" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_01 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_03 => X"00000000000000000000000000000000000000ae000000000000000000000000",
            INIT_04 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_07 => X"0000000000000000000000000000000000000003000000000000007100000000",
            INIT_08 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_09 => X"0000000500000000000000010000000000000000000000000000000000000000",
            INIT_0A => X"0000007b000000000000002a0000000000000000000000000000000b00000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000001800000000000000000000000000000000000000000000001900000000",
            INIT_0E => X"0000002c00000000000000690000000000000016000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000800000000000000050000000000000001000000000000000000000000",
            INIT_11 => X"0000000c000000000000000c0000000000000000000000000000000000000000",
            INIT_12 => X"000001c800000000000001960000000000000154000000000000000b00000000",
            INIT_13 => X"0000019f00000000000001af00000000000001d500000000000001e000000000",
            INIT_14 => X"000000fb0000000000000127000000000000015e000000000000017c00000000",
            INIT_15 => X"0000008e0000000000000047000000000000006700000000000000cc00000000",
            INIT_16 => X"000001a1000000000000018d000000000000017b00000000000001b900000000",
            INIT_17 => X"0000013100000000000001490000000000000156000000000000018500000000",
            INIT_18 => X"0000006600000000000000b100000000000000ec000000000000010e00000000",
            INIT_19 => X"0000016100000000000000a30000000000000004000000000000000000000000",
            INIT_1A => X"0000011d0000000000000138000000000000014b000000000000016100000000",
            INIT_1B => X"000000df00000000000000e900000000000000fb00000000000000fa00000000",
            INIT_1C => X"000000000000000000000000000000000000006d00000000000000ce00000000",
            INIT_1D => X"000000ee00000000000000f000000000000000aa000000000000004200000000",
            INIT_1E => X"000000ec00000000000000e800000000000000e500000000000000e800000000",
            INIT_1F => X"000000a900000000000000ae00000000000000b800000000000000cd00000000",
            INIT_20 => X"000000c900000000000000650000000000000000000000000000003100000000",
            INIT_21 => X"000000f100000000000000ee00000000000000d000000000000000d800000000",
            INIT_22 => X"000000a900000000000000da00000000000000f000000000000000f100000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000009100000000",
            INIT_24 => X"000000c300000000000000be0000000000000068000000000000000000000000",
            INIT_25 => X"000000ee00000000000000ea00000000000000ec00000000000000e800000000",
            INIT_26 => X"000000000000000000000000000000000000001500000000000000d800000000",
            INIT_27 => X"0000000000000000000000000000000000000005000000000000000d00000000",
            INIT_28 => X"000000ee00000000000000a50000000000000019000000000000003e00000000",
            INIT_29 => X"0000006d00000000000000d500000000000000f400000000000000ea00000000",
            INIT_2A => X"0000003700000000000000270000000000000025000000000000005100000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"000000ee00000000000000ed000000000000005b000000000000004200000000",
            INIT_2D => X"0000000000000000000000000000000000000003000000000000009000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000001100000000000000b300000000000000f0000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"000000000000000000000000000000000000000000000000000000d300000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"000000c400000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000006400000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"00000000000000000000003c0000000000000013000000000000000000000000",
            INIT_3B => X"0000000000000000000000c4000000000000000b000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000077000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"000000090000000000000000000000000000000c000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000003400000000",
            INIT_44 => X"000000a600000000000000a60000000000000094000000000000004300000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000003500000000",
            INIT_46 => X"0000001b00000000000000000000000000000000000000000000002700000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000004600000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000200000000000000000000000000000000000000000",
            INIT_63 => X"0000001800000000000000650000000000000000000000000000002800000000",
            INIT_64 => X"000000000000000000000000000000000000002b000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000002b000000000000001a000000000000000d000000000000000000000000",
            INIT_67 => X"00000000000000000000003d0000000000000000000000000000002500000000",
            INIT_68 => X"0000000000000000000000000000000000000029000000000000000000000000",
            INIT_69 => X"0000001500000000000000330000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000052000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000003000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000003800000000",
            INIT_6F => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000002700000000000000300000000000000000000000000000000000000000",
            INIT_71 => X"0000001c00000000000000000000000000000019000000000000000000000000",
            INIT_72 => X"0000002600000000000000130000000000000000000000000000006a00000000",
            INIT_73 => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_74 => X"0000000e00000000000000090000000000000094000000000000000000000000",
            INIT_75 => X"0000005a00000000000000000000000000000000000000000000004a00000000",
            INIT_76 => X"0000001e0000000000000000000000000000001f000000000000001d00000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_78 => X"0000003100000000000000230000000000000000000000000000007700000000",
            INIT_79 => X"0000000f000000000000002d0000000000000000000000000000002e00000000",
            INIT_7A => X"00000000000000000000006b0000000000000000000000000000001600000000",
            INIT_7B => X"0000003f00000000000000000000000000000000000000000000000400000000",
            INIT_7C => X"0000000a00000000000000120000000000000019000000000000000000000000",
            INIT_7D => X"0000002300000000000000200000000000000016000000000000000000000000",
            INIT_7E => X"00000013000000000000000c0000000000000047000000000000001600000000",
            INIT_7F => X"0000004000000000000000220000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE46;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE47 : if BRAM_NAME = "samplegold_layersamples_instance47" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000024000000000000002d000000000000002e000000000000002500000000",
            INIT_01 => X"000000000000000000000015000000000000001c000000000000002700000000",
            INIT_02 => X"0000005a00000000000000230000000000000024000000000000002800000000",
            INIT_03 => X"0000005a0000000000000063000000000000006f000000000000005b00000000",
            INIT_04 => X"0000002e0000000000000036000000000000004b000000000000004900000000",
            INIT_05 => X"0000000600000000000000000000000000000018000000000000003000000000",
            INIT_06 => X"0000005200000000000000550000000000000000000000000000000000000000",
            INIT_07 => X"000000280000000000000035000000000000003d000000000000004d00000000",
            INIT_08 => X"0000000f0000000000000017000000000000001e000000000000002c00000000",
            INIT_09 => X"0000000000000000000000000000000000000006000000000000000300000000",
            INIT_0A => X"0000002300000000000000310000000000000043000000000000000200000000",
            INIT_0B => X"0000001600000000000000140000000000000015000000000000001c00000000",
            INIT_0C => X"0000003600000000000000080000000000000012000000000000001400000000",
            INIT_0D => X"0000001300000000000000170000000000000000000000000000000000000000",
            INIT_0E => X"0000000c000000000000000d0000000000000009000000000000000a00000000",
            INIT_0F => X"00000021000000000000001d0000000000000017000000000000001000000000",
            INIT_10 => X"000000000000000000000010000000000000001b000000000000002200000000",
            INIT_11 => X"0000000b0000000000000007000000000000000f000000000000000c00000000",
            INIT_12 => X"000000150000000000000011000000000000000f000000000000000c00000000",
            INIT_13 => X"0000001f000000000000002f000000000000003c000000000000002b00000000",
            INIT_14 => X"0000002000000000000000000000000000000000000000000000004900000000",
            INIT_15 => X"0000000e000000000000000c0000000000000003000000000000000d00000000",
            INIT_16 => X"00000014000000000000000b0000000000000013000000000000001200000000",
            INIT_17 => X"0000007b00000000000000b00000000000000092000000000000007000000000",
            INIT_18 => X"0000002600000000000000000000000000000019000000000000007700000000",
            INIT_19 => X"000000170000000000000014000000000000000f000000000000000000000000",
            INIT_1A => X"0000005100000000000000450000000000000036000000000000000300000000",
            INIT_1B => X"000000e200000000000000000000000000000000000000000000000500000000",
            INIT_1C => X"00000000000000000000000d0000000000000000000000000000006800000000",
            INIT_1D => X"0000002b00000000000000000000000000000012000000000000001300000000",
            INIT_1E => X"0000000000000000000000010000000000000005000000000000002000000000",
            INIT_1F => X"000000ce00000000000000d400000000000000a6000000000000000600000000",
            INIT_20 => X"0000001400000000000000110000000000000000000000000000000000000000",
            INIT_21 => X"00000020000000000000000c000000000000001b000000000000000000000000",
            INIT_22 => X"000000f000000000000000dd0000000000000000000000000000000000000000",
            INIT_23 => X"00000000000000000000000b00000000000000fa00000000000000db00000000",
            INIT_24 => X"0000006100000000000000000000000000000081000000000000000500000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000003400000000",
            INIT_26 => X"000000ec00000000000000b800000000000000d2000000000000000000000000",
            INIT_27 => X"0000009100000000000000830000000000000063000000000000009400000000",
            INIT_28 => X"0000003f00000000000000920000000000000000000000000000009f00000000",
            INIT_29 => X"0000001700000000000000000000000000000000000000000000000600000000",
            INIT_2A => X"00000020000000000000000000000000000000f800000000000000b400000000",
            INIT_2B => X"0000001d000000000000009400000000000000a4000000000000006b00000000",
            INIT_2C => X"0000000000000000000000550000000000000000000000000000000000000000",
            INIT_2D => X"000000b900000000000000460000000000000024000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000008a00000000",
            INIT_2F => X"000000000000000000000000000000000000004c000000000000006200000000",
            INIT_30 => X"000000000000000000000000000000000000004c000000000000000000000000",
            INIT_31 => X"0000006300000000000000a70000000000000099000000000000003900000000",
            INIT_32 => X"0000005600000000000000000000000000000005000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"00000056000000000000002e0000000000000000000000000000003d00000000",
            INIT_35 => X"0000000700000000000000110000000000000063000000000000006200000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"000000190000000000000034000000000000002a000000000000006300000000",
            INIT_3C => X"0000000f00000000000000240000000000000017000000000000001000000000",
            INIT_3D => X"0000002500000000000000080000000000000000000000000000002d00000000",
            INIT_3E => X"0000001f00000000000000260000000000000000000000000000000f00000000",
            INIT_3F => X"00000020000000000000001f000000000000000c000000000000003400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002a0000000000000021000000000000002c000000000000001c00000000",
            INIT_41 => X"000000000000000000000033000000000000003b000000000000002900000000",
            INIT_42 => X"00000000000000000000000b0000000000000033000000000000005c00000000",
            INIT_43 => X"000000320000000000000029000000000000001b000000000000001300000000",
            INIT_44 => X"00000032000000000000003c0000000000000038000000000000003300000000",
            INIT_45 => X"00000073000000000000000f000000000000000000000000000000a800000000",
            INIT_46 => X"000000320000000000000035000000000000002a000000000000002d00000000",
            INIT_47 => X"0000004b000000000000003a000000000000003e000000000000003000000000",
            INIT_48 => X"0000000000000000000000550000000000000050000000000000005300000000",
            INIT_49 => X"0000001900000000000000120000000000000029000000000000000000000000",
            INIT_4A => X"0000003000000000000000300000000000000036000000000000003c00000000",
            INIT_4B => X"0000001700000000000000350000000000000064000000000000003a00000000",
            INIT_4C => X"0000002d000000000000001800000000000000ab000000000000004e00000000",
            INIT_4D => X"0000003a000000000000002f0000000000000029000000000000003000000000",
            INIT_4E => X"0000003800000000000000300000000000000033000000000000003500000000",
            INIT_4F => X"00000000000000000000005300000000000000e9000000000000007500000000",
            INIT_50 => X"0000000000000000000000000000000000000069000000000000000000000000",
            INIT_51 => X"0000003000000000000000370000000000000026000000000000002500000000",
            INIT_52 => X"0000000000000000000000bc000000000000002a000000000000003400000000",
            INIT_53 => X"0000002f00000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000030000000000000000000000000000007a00000000",
            INIT_55 => X"00000046000000000000002b000000000000002c000000000000000000000000",
            INIT_56 => X"0000000000000000000000260000000000000000000000000000007600000000",
            INIT_57 => X"0000000000000000000001860000000000000132000000000000006e00000000",
            INIT_58 => X"000000de00000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000260000000000000031000000000000003000000000",
            INIT_5A => X"000000fd00000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"00000018000000000000003700000000000000fc000000000000004c00000000",
            INIT_5D => X"0000000000000000000000110000000000000000000000000000019900000000",
            INIT_5E => X"0000000000000000000000000000000000000069000000000000003a00000000",
            INIT_5F => X"0000007c00000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000ae0000000000000000000000000000000000000000",
            INIT_61 => X"0000007d00000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"000000000000000000000000000000000000000000000000000000d300000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"000000340000000000000001000000000000004f000000000000000000000000",
            INIT_65 => X"0000007300000000000000a10000000000000044000000000000000000000000",
            INIT_66 => X"00000000000000000000002e0000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_68 => X"0000000000000000000000220000000000000017000000000000003e00000000",
            INIT_69 => X"00000000000000000000008e000000000000007d00000000000000b500000000",
            INIT_6A => X"00000021000000000000000f0000000000000035000000000000000000000000",
            INIT_6B => X"0000004600000000000000210000000000000000000000000000003300000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000002e00000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000005200000000",
            INIT_6F => X"000000000000000000000034000000000000002c000000000000000000000000",
            INIT_70 => X"0000003c000000000000002f0000000000000068000000000000000500000000",
            INIT_71 => X"0000003200000000000000190000000000000020000000000000003000000000",
            INIT_72 => X"0000002b000000000000002a0000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000003800000000",
            INIT_74 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"00000002000000000000005e0000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000340000000000000000000000000000000900000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_7E => X"0000000000000000000000030000000000000000000000000000000400000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE47;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE48 : if BRAM_NAME = "samplegold_layersamples_instance48" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000030000000000000027000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"000000000000000000000000000000000000009f000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000008a00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"000000740000000000000030000000000000005e000000000000000a00000000",
            INIT_0C => X"00000000000000000000000000000000000000e0000000000000004e00000000",
            INIT_0D => X"000000000000000000000000000000000000000000000000000000ad00000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000005100000000000000300000000000000009000000000000007300000000",
            INIT_13 => X"0000000000000000000000020000000000000000000000000000005b00000000",
            INIT_14 => X"0000000f00000000000000000000000000000035000000000000000000000000",
            INIT_15 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000006200000000000000100000000000000034000000000000000000000000",
            INIT_17 => X"0000000000000000000000ff0000000000000014000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000011700000000",
            INIT_1A => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000001fa0000000000000025000000000000000000000000",
            INIT_1C => X"00000000000000000000002e0000000000000000000000000000000000000000",
            INIT_1D => X"0000004900000000000000000000000000000000000000000000009800000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000003600000000",
            INIT_1F => X"0000000000000000000000660000000000000053000000000000000000000000",
            INIT_20 => X"0000009e00000000000000210000000000000019000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"00000000000000000000003e0000000000000000000000000000000000000000",
            INIT_23 => X"0000001a0000000000000000000000000000011f000000000000000000000000",
            INIT_24 => X"00000004000000000000008a0000000000000056000000000000000000000000",
            INIT_25 => X"000000f000000000000000ff0000000000000102000000000000009500000000",
            INIT_26 => X"00000000000000000000003d0000000000000034000000000000009c00000000",
            INIT_27 => X"000000000000000000000001000000000000000d000000000000008600000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"000000000000000000000000000000000000000c000000000000008400000000",
            INIT_2B => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000009b00000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000009a00000000000000ac00000000000000a5000000000000009a00000000",
            INIT_65 => X"000000570000000000000074000000000000007f000000000000008400000000",
            INIT_66 => X"000000000000000000000031000000000000004d000000000000003a00000000",
            INIT_67 => X"0000008400000000000000890000000000000022000000000000002600000000",
            INIT_68 => X"00000045000000000000004f000000000000005b000000000000006600000000",
            INIT_69 => X"0000003d000000000000003e0000000000000045000000000000004300000000",
            INIT_6A => X"0000001300000000000000070000000000000004000000000000002700000000",
            INIT_6B => X"0000003e0000000000000032000000000000003d000000000000001e00000000",
            INIT_6C => X"0000002c00000000000000310000000000000037000000000000002d00000000",
            INIT_6D => X"00000000000000000000003c0000000000000038000000000000003e00000000",
            INIT_6E => X"0000001d00000000000000220000000000000015000000000000000000000000",
            INIT_6F => X"0000002b000000000000002a000000000000002d000000000000002d00000000",
            INIT_70 => X"00000033000000000000002c000000000000002c000000000000003300000000",
            INIT_71 => X"0000002400000000000000000000000000000025000000000000004000000000",
            INIT_72 => X"0000001f000000000000002d0000000000000024000000000000003200000000",
            INIT_73 => X"0000002a00000000000000260000000000000027000000000000002500000000",
            INIT_74 => X"0000001a00000000000000170000000000000023000000000000002a00000000",
            INIT_75 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000002100000000000000240000000000000028000000000000002800000000",
            INIT_77 => X"0000001600000000000000150000000000000025000000000000002400000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_79 => X"00000000000000000000001e0000000000000000000000000000000000000000",
            INIT_7A => X"0000001700000000000000220000000000000025000000000000001d00000000",
            INIT_7B => X"0000000000000000000000000000000000000005000000000000001b00000000",
            INIT_7C => X"00000000000000000000001e0000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"00000000000000000000001a0000000000000019000000000000002500000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE48;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE49 : if BRAM_NAME = "samplegold_layersamples_instance49" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_01 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_03 => X"0000000000000000000000000000000000000038000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000400000000000000130000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000018000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000b00000000000000040000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000220000000000000018000000000000001200000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000c00000000000000120000000000000011000000000000000500000000",
            INIT_23 => X"0000000000000000000000000000000000000018000000000000000f00000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000001b000000000000000b0000000000000000000000000000000000000000",
            INIT_27 => X"0000003300000000000000000000000000000000000000000000002d00000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000002e00000000000000260000000000000028000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"000000000000000000000030000000000000003d000000000000001c00000000",
            INIT_2F => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000036000000000000003b00000000",
            INIT_33 => X"000000000000000000000000000000000000002a000000000000000500000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000002c00000000",
            INIT_37 => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000003600000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000510000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000075000000000000002900000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000003400000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000c00000000000000150000000000000000000000000000005f00000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000006000000000000000260000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000900000000000000430000000000000030000000000000000000000000",
            INIT_4D => X"0000004e000000000000002d0000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000003400000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"000000410000000000000014000000000000003d000000000000004a00000000",
            INIT_51 => X"0000002e000000000000004a0000000000000058000000000000005900000000",
            INIT_52 => X"0000002c00000000000000470000000000000052000000000000001b00000000",
            INIT_53 => X"0000005b000000000000003d0000000000000011000000000000000300000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000006300000000",
            INIT_55 => X"0000000100000000000000000000000000000010000000000000000a00000000",
            INIT_56 => X"0000000500000000000000000000000000000000000000000000000100000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_58 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000800000000000000030000000000000030000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000f0000000000000014000000000000002a000000000000000000000000",
            INIT_5D => X"000000000000000000000000000000000000001b000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"00000038000000000000001d0000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000015000000000000000700000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000002300000000000000050000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000a00000000000000000000000000000000000000000000000200000000",
            INIT_6B => X"0000000900000000000000000000000000000000000000000000000300000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000002c00000000",
            INIT_6D => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"000000000000000000000000000000000000001e000000000000001400000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000005700000000000000060000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000330000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000110000000000000000000000000000004800000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000017000000000000000000000000",
            INIT_7A => X"0000006c000000000000009b000000000000009e000000000000000800000000",
            INIT_7B => X"00000000000000000000000f0000000000000034000000000000008800000000",
            INIT_7C => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_7D => X"000000ec00000000000001070000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"00000000000000000000000f0000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE49;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE50 : if BRAM_NAME = "samplegold_layersamples_instance50" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000001e00000000000000480000000000000048000000000000000000000000",
            INIT_02 => X"0000002300000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_05 => X"00000078000000000000003a0000000000000000000000000000000000000000",
            INIT_06 => X"0000000600000000000000000000000000000000000000000000005100000000",
            INIT_07 => X"000000000000000000000054000000000000004d000000000000000e00000000",
            INIT_08 => X"000000480000000000000022000000000000000c000000000000000900000000",
            INIT_09 => X"0000000000000000000000030000000000000036000000000000006f00000000",
            INIT_0A => X"0000000500000000000000110000000000000000000000000000000200000000",
            INIT_0B => X"0000002300000000000000410000000000000028000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000010000000000000000f00000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000190000000000000000000000000000002200000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_19 => X"0000001800000000000000030000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000003000000000000001e00000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000080000000000000000000000000000001900000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_20 => X"0000000000000000000000260000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"00000000000000000000000e0000000000000028000000000000001100000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000045000000000000000000000000",
            INIT_25 => X"0000003000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"00000000000000000000000e0000000000000000000000000000002800000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000b00000000000000010000000000000000000000000000000800000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_2D => X"0000000200000000000000040000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000200000000000000000000000000000009000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000003700000000000000070000000000000000000000000000001e00000000",
            INIT_3C => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000020000000000000000000000000000001200000000",
            INIT_3E => X"0000001600000000000000000000000000000029000000000000000000000000",
            INIT_3F => X"0000000200000000000000300000000000000015000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000041000000000000001a0000000000000000000000000000000000000000",
            INIT_41 => X"0000000d00000000000000100000000000000007000000000000000000000000",
            INIT_42 => X"000000040000000000000000000000000000001e000000000000005300000000",
            INIT_43 => X"00000016000000000000002d000000000000000e000000000000002000000000",
            INIT_44 => X"000000000000000000000024000000000000002a000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000015000000000000000600000000",
            INIT_49 => X"000000000000000000000000000000000000002c000000000000000000000000",
            INIT_4A => X"0000000f00000000000000040000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000011000000000000002300000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000e00000000000000000000000000000018000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"00000033000000000000004b000000000000000d000000000000000000000000",
            INIT_51 => X"0000000000000000000000250000000000000032000000000000001600000000",
            INIT_52 => X"0000000200000000000000000000000000000001000000000000000700000000",
            INIT_53 => X"0000001400000000000000000000000000000000000000000000000500000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000001d00000000000000000000000000000015000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_5A => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_5B => X"0000000a00000000000000080000000000000000000000000000000000000000",
            INIT_5C => X"000000000000000000000000000000000000001e000000000000000f00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"000000000000000000000000000000000000000a000000000000000d00000000",
            INIT_60 => X"000000000000000000000004000000000000005e000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000130000000000000028000000000000000000000000",
            INIT_63 => X"000000000000000000000012000000000000004c000000000000003b00000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_69 => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000007b00000000000000000000000000000000000000000000000e00000000",
            INIT_6B => X"000000000000000000000021000000000000000000000000000000ce00000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_6E => X"0000000000000000000000000000000000000080000000000000000000000000",
            INIT_6F => X"000000220000000000000000000000000000002b000000000000004100000000",
            INIT_70 => X"0000000000000000000000000000000000000034000000000000006400000000",
            INIT_71 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"000000000000000000000000000000000000003e000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000270000000000000000000000000000000200000000",
            INIT_76 => X"0000000100000000000000370000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_78 => X"0000000000000000000000000000000000000002000000000000000500000000",
            INIT_79 => X"0000003000000000000000080000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_7B => X"0000000900000000000000030000000000000004000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_7D => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_7F => X"00000014000000000000000c0000000000000004000000000000000100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE50;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE51 : if BRAM_NAME = "samplegold_layersamples_instance51" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_01 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000400000000000000090000000000000012000000000000001000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000001000000000000003a00000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_07 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_0C => X"0000002600000000000000220000000000000000000000000000000000000000",
            INIT_0D => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"000000000000000000000010000000000000005d000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_16 => X"0000000700000000000000000000000000000000000000000000000800000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000003900000000",
            INIT_18 => X"0000000000000000000000000000000000000025000000000000000600000000",
            INIT_19 => X"0000000400000000000000070000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"000000000000000000000060000000000000000d000000000000000000000000",
            INIT_1F => X"0000003d000000000000007c000000000000007e000000000000000000000000",
            INIT_20 => X"0000000000000000000000090000000000000000000000000000008000000000",
            INIT_21 => X"0000000300000000000000140000000000000000000000000000000000000000",
            INIT_22 => X"0000001c00000000000000000000000000000000000000000000000d00000000",
            INIT_23 => X"0000005a000000000000001a000000000000000200000000000000b900000000",
            INIT_24 => X"0000000400000000000000000000000000000018000000000000000700000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_26 => X"00000000000000000000006a00000000000000f6000000000000001200000000",
            INIT_27 => X"0000000000000000000000000000000000000017000000000000004b00000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_29 => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000028000000000000000000000000",
            INIT_2B => X"0000000000000000000000340000000000000008000000000000001200000000",
            INIT_2C => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_2E => X"0000000000000000000000540000000000000032000000000000000000000000",
            INIT_2F => X"0000000500000000000000030000000000000000000000000000000000000000",
            INIT_30 => X"0000001b00000000000000000000000000000022000000000000000e00000000",
            INIT_31 => X"0000004100000000000000490000000000000000000000000000000400000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_34 => X"000000000000000000000007000000000000000e000000000000000000000000",
            INIT_35 => X"00000000000000000000000d0000000000000005000000000000000600000000",
            INIT_36 => X"0000001e0000000000000020000000000000000b000000000000000000000000",
            INIT_37 => X"000000150000000000000018000000000000001b000000000000001200000000",
            INIT_38 => X"0000001f000000000000000c0000000000000019000000000000001a00000000",
            INIT_39 => X"000000000000000000000002000000000000001b000000000000000600000000",
            INIT_3A => X"0000002b000000000000003e0000000000000000000000000000002c00000000",
            INIT_3B => X"00000020000000000000001b0000000000000015000000000000001100000000",
            INIT_3C => X"000000030000000000000026000000000000001a000000000000001900000000",
            INIT_3D => X"0000002a000000000000000c000000000000001c000000000000000c00000000",
            INIT_3E => X"00000009000000000000002a0000000000000024000000000000002d00000000",
            INIT_3F => X"000000170000000000000026000000000000001d000000000000002400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000800000000000000070000000000000026000000000000001f00000000",
            INIT_41 => X"0000003b00000000000000260000000000000000000000000000006700000000",
            INIT_42 => X"00000000000000000000002c0000000000000025000000000000003400000000",
            INIT_43 => X"00000024000000000000001c0000000000000031000000000000001300000000",
            INIT_44 => X"000000a300000000000000000000000000000000000000000000002800000000",
            INIT_45 => X"000000420000000000000006000000000000001d000000000000005600000000",
            INIT_46 => X"0000001500000000000000380000000000000044000000000000005700000000",
            INIT_47 => X"0000002f000000000000002e0000000000000014000000000000002f00000000",
            INIT_48 => X"0000002f000000000000009a0000000000000000000000000000000000000000",
            INIT_49 => X"0000006100000000000000280000000000000000000000000000004500000000",
            INIT_4A => X"0000000e00000000000000550000000000000047000000000000004600000000",
            INIT_4B => X"000000000000000000000032000000000000002b000000000000000000000000",
            INIT_4C => X"0000000000000000000000e50000000000000016000000000000000000000000",
            INIT_4D => X"000000280000000000000037000000000000005a000000000000000000000000",
            INIT_4E => X"0000003700000000000000090000000000000057000000000000005200000000",
            INIT_4F => X"000000000000000000000000000000000000002f000000000000000e00000000",
            INIT_50 => X"0000000000000000000000c90000000000000000000000000000001d00000000",
            INIT_51 => X"0000005d000000000000001e000000000000001d000000000000005c00000000",
            INIT_52 => X"0000000500000000000000310000000000000042000000000000005700000000",
            INIT_53 => X"0000001800000000000000000000000000000000000000000000002400000000",
            INIT_54 => X"0000003b00000000000000b60000000000000074000000000000004700000000",
            INIT_55 => X"0000005600000000000000460000000000000012000000000000004600000000",
            INIT_56 => X"00000043000000000000001d000000000000000c000000000000005800000000",
            INIT_57 => X"000000d500000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000007200000000000000000000000000000096000000000000000000000000",
            INIT_59 => X"000000630000000000000046000000000000002b000000000000001d00000000",
            INIT_5A => X"000000000000000000000036000000000000005a000000000000002500000000",
            INIT_5B => X"00000010000000000000000e000000000000008a000000000000002000000000",
            INIT_5C => X"000000290000000000000011000000000000002e000000000000002600000000",
            INIT_5D => X"00000033000000000000005e0000000000000043000000000000002a00000000",
            INIT_5E => X"000000000000000000000000000000000000003a000000000000004800000000",
            INIT_5F => X"000000130000000000000079000000000000003d000000000000004c00000000",
            INIT_60 => X"0000000700000000000000000000000000000068000000000000000800000000",
            INIT_61 => X"00000000000000000000003e000000000000005c000000000000002b00000000",
            INIT_62 => X"0000000000000000000000000000000000000001000000000000008600000000",
            INIT_63 => X"0000000000000000000000570000000000000047000000000000000a00000000",
            INIT_64 => X"000000440000000000000000000000000000000e000000000000005900000000",
            INIT_65 => X"0000001d00000000000000200000000000000079000000000000003b00000000",
            INIT_66 => X"00000025000000000000001a0000000000000008000000000000000300000000",
            INIT_67 => X"00000027000000000000001e000000000000002d000000000000000e00000000",
            INIT_68 => X"0000004400000000000000000000000000000000000000000000002a00000000",
            INIT_69 => X"0000001f000000000000000c0000000000000033000000000000004a00000000",
            INIT_6A => X"0000000000000000000000340000000000000027000000000000002100000000",
            INIT_6B => X"0000003400000000000000440000000000000045000000000000001600000000",
            INIT_6C => X"0000004c000000000000001d000000000000000d000000000000003400000000",
            INIT_6D => X"0000000000000000000000000000000000000031000000000000002900000000",
            INIT_6E => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"00000015000000000000001b0000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000003700000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE51;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE52 : if BRAM_NAME = "samplegold_layersamples_instance52" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000200000000000000078000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"00000000000000000000000a000000000000000b000000000000000000000000",
            INIT_08 => X"0000000000000000000000660000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000005600000000000000000000000000000000000000000000001700000000",
            INIT_10 => X"00000000000000000000000c000000000000001e000000000000005b00000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000005000000000000000000000000000000040000000000000002300000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"000000ad00000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000220000000000000041000000000000004000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000001000000000000000190000000000000000000000000000000400000000",
            INIT_1B => X"0000000000000000000000310000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000001100000000000000000000000000000000000000000000001000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_20 => X"0000003c00000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"000000000000000000000000000000000000001c000000000000002300000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"00000000000000000000000c000000000000000b000000000000001800000000",
            INIT_27 => X"00000013000000000000000b0000000000000000000000000000000000000000",
            INIT_28 => X"0000000c000000000000000e000000000000000c000000000000000d00000000",
            INIT_29 => X"0000001f000000000000001a000000000000000d000000000000000700000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_2B => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000300000000000000000000000000000001000000000000000000000000",
            INIT_2D => X"0000000900000000000000170000000000000014000000000000000400000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"00000000000000000000002a0000000000000013000000000000000e00000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"000000000000000000000000000000000000004e000000000000001b00000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000001400000000000000130000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000005100000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000001b00000000000000120000000000000012000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000003f00000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000000000000000000015000000000000000e000000000000001200000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000002d00000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"000000170000000000000006000000000000002f000000000000000f00000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000002d000000000000002a0000000000000000000000000000000000000000",
            INIT_48 => X"000000100000000000000000000000000000004a000000000000000800000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000001800000000000000450000000000000036000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"000000080000000000000014000000000000001b000000000000002100000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000002000000000000000900000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000f000000000000000f0000000000000005000000000000000300000000",
            INIT_5F => X"00000018000000000000002a0000000000000032000000000000002300000000",
            INIT_60 => X"0000000b00000000000000100000000000000012000000000000000d00000000",
            INIT_61 => X"0000000300000000000000140000000000000015000000000000000f00000000",
            INIT_62 => X"0000003800000000000000040000000000000019000000000000000800000000",
            INIT_63 => X"00000028000000000000004e0000000000000045000000000000004100000000",
            INIT_64 => X"0000002d000000000000002b000000000000002a000000000000001e00000000",
            INIT_65 => X"0000000900000000000000050000000000000030000000000000003300000000",
            INIT_66 => X"000000510000000000000036000000000000001e000000000000001000000000",
            INIT_67 => X"0000003e00000000000000510000000000000066000000000000006300000000",
            INIT_68 => X"0000002f00000000000000310000000000000040000000000000003500000000",
            INIT_69 => X"000000230000000000000015000000000000000c000000000000003100000000",
            INIT_6A => X"0000005b0000000000000052000000000000003b000000000000002d00000000",
            INIT_6B => X"0000004600000000000000550000000000000084000000000000007200000000",
            INIT_6C => X"000000460000000000000035000000000000003a000000000000004c00000000",
            INIT_6D => X"0000001a00000000000000430000000000000025000000000000001f00000000",
            INIT_6E => X"0000006000000000000000530000000000000042000000000000003700000000",
            INIT_6F => X"000000600000000000000072000000000000007e000000000000007600000000",
            INIT_70 => X"0000002a00000000000000690000000000000063000000000000006300000000",
            INIT_71 => X"0000003c0000000000000007000000000000001b000000000000001f00000000",
            INIT_72 => X"0000006200000000000000470000000000000041000000000000005300000000",
            INIT_73 => X"000000700000000000000068000000000000007b000000000000006b00000000",
            INIT_74 => X"0000001400000000000000130000000000000062000000000000007400000000",
            INIT_75 => X"00000032000000000000002a0000000000000030000000000000001200000000",
            INIT_76 => X"00000053000000000000005c000000000000005a000000000000004500000000",
            INIT_77 => X"0000005c000000000000006a0000000000000065000000000000006800000000",
            INIT_78 => X"000000310000000000000025000000000000001e000000000000003b00000000",
            INIT_79 => X"000000580000000000000042000000000000005a000000000000001000000000",
            INIT_7A => X"0000005900000000000000480000000000000056000000000000005f00000000",
            INIT_7B => X"000000460000000000000053000000000000005d000000000000006800000000",
            INIT_7C => X"0000002d00000000000000300000000000000035000000000000002c00000000",
            INIT_7D => X"0000005e00000000000000520000000000000067000000000000005100000000",
            INIT_7E => X"0000005b000000000000004f000000000000003d000000000000004b00000000",
            INIT_7F => X"0000002e000000000000006c0000000000000052000000000000005500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE52;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE53 : if BRAM_NAME = "samplegold_layersamples_instance53" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000370000000000000020000000000000001d000000000000003a00000000",
            INIT_01 => X"0000004d00000000000000530000000000000053000000000000004f00000000",
            INIT_02 => X"000000560000000000000053000000000000004d000000000000003f00000000",
            INIT_03 => X"0000001c000000000000001b0000000000000068000000000000005c00000000",
            INIT_04 => X"0000003a000000000000002d0000000000000018000000000000000700000000",
            INIT_05 => X"0000004d00000000000000510000000000000032000000000000004b00000000",
            INIT_06 => X"00000070000000000000005a0000000000000053000000000000005700000000",
            INIT_07 => X"0000000000000000000000000000000000000002000000000000007600000000",
            INIT_08 => X"0000003f000000000000002f0000000000000028000000000000001f00000000",
            INIT_09 => X"00000042000000000000003e0000000000000039000000000000004a00000000",
            INIT_0A => X"00000078000000000000007b000000000000006a000000000000005900000000",
            INIT_0B => X"0000002900000000000000190000000000000015000000000000000000000000",
            INIT_0C => X"0000003c0000000000000055000000000000003e000000000000002400000000",
            INIT_0D => X"000000420000000000000042000000000000003a000000000000004000000000",
            INIT_0E => X"0000001f0000000000000073000000000000008b000000000000007400000000",
            INIT_0F => X"0000005400000000000000520000000000000044000000000000003200000000",
            INIT_10 => X"0000005000000000000000560000000000000056000000000000005a00000000",
            INIT_11 => X"0000005d0000000000000036000000000000002e000000000000004900000000",
            INIT_12 => X"0000005200000000000000420000000000000083000000000000007e00000000",
            INIT_13 => X"000000750000000000000075000000000000006b000000000000005f00000000",
            INIT_14 => X"0000007100000000000000800000000000000075000000000000006800000000",
            INIT_15 => X"00000086000000000000006e0000000000000065000000000000006900000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000008500000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"000000000000000000000001000000000000000b000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000800000000000000160000000000000008000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"00000014000000000000000c000000000000000b000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000800000000000000110000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_2F => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000003500000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000260000000000000000000000000000000000000000",
            INIT_3C => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"000000000000000000000018000000000000000c000000000000002900000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_42 => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000001e00000000000000290000000000000000000000000000000000000000",
            INIT_47 => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000002600000000",
            INIT_49 => X"0000000000000000000000140000000000000017000000000000000200000000",
            INIT_4A => X"000000000000000000000044000000000000003c000000000000000000000000",
            INIT_4B => X"0000002c000000000000001e000000000000002a000000000000002d00000000",
            INIT_4C => X"0000003000000000000000200000000000000000000000000000001500000000",
            INIT_4D => X"0000003100000000000000360000000000000021000000000000001b00000000",
            INIT_4E => X"0000003200000000000000370000000000000051000000000000004a00000000",
            INIT_4F => X"0000006900000000000000440000000000000026000000000000002700000000",
            INIT_50 => X"0000003e00000000000000330000000000000038000000000000004f00000000",
            INIT_51 => X"00000024000000000000002f000000000000002e000000000000003100000000",
            INIT_52 => X"00000042000000000000003e0000000000000038000000000000002300000000",
            INIT_53 => X"0000008c00000000000000840000000000000078000000000000000400000000",
            INIT_54 => X"0000003100000000000000360000000000000038000000000000007a00000000",
            INIT_55 => X"0000001300000000000000170000000000000024000000000000002b00000000",
            INIT_56 => X"0000003400000000000000380000000000000042000000000000003b00000000",
            INIT_57 => X"000000b100000000000000bc00000000000000ac000000000000009000000000",
            INIT_58 => X"0000002b000000000000002f0000000000000037000000000000006100000000",
            INIT_59 => X"0000003f000000000000000d000000000000000d000000000000000d00000000",
            INIT_5A => X"000000b600000000000000420000000000000037000000000000004100000000",
            INIT_5B => X"0000009600000000000000b200000000000000b500000000000000c400000000",
            INIT_5C => X"000000110000000000000044000000000000005f000000000000008100000000",
            INIT_5D => X"0000002b000000000000002c000000000000000f000000000000001000000000",
            INIT_5E => X"000000b200000000000000a3000000000000000c000000000000007500000000",
            INIT_5F => X"000000b900000000000000c100000000000000a200000000000000b000000000",
            INIT_60 => X"000000000000000000000027000000000000009100000000000000ae00000000",
            INIT_61 => X"0000007400000000000000180000000000000016000000000000000000000000",
            INIT_62 => X"000000ad00000000000000ae0000000000000092000000000000000000000000",
            INIT_63 => X"000000c700000000000000b400000000000000c200000000000000bd00000000",
            INIT_64 => X"000000000000000000000000000000000000004000000000000000be00000000",
            INIT_65 => X"0000000300000000000000280000000000000011000000000000001700000000",
            INIT_66 => X"000000c000000000000000b20000000000000073000000000000005900000000",
            INIT_67 => X"000000af00000000000000c900000000000000aa00000000000000c000000000",
            INIT_68 => X"0000002700000000000000050000000000000020000000000000007400000000",
            INIT_69 => X"0000003200000000000000020000000000000029000000000000001700000000",
            INIT_6A => X"000000c1000000000000009b000000000000007f000000000000003300000000",
            INIT_6B => X"000000bf00000000000000ca00000000000000c300000000000000bd00000000",
            INIT_6C => X"0000000a000000000000001d0000000000000013000000000000004e00000000",
            INIT_6D => X"0000004d000000000000006b0000000000000000000000000000001e00000000",
            INIT_6E => X"000000c800000000000000c30000000000000073000000000000006800000000",
            INIT_6F => X"0000005500000000000000c200000000000000df00000000000000c900000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000005300000000000000a3000000000000005d000000000000005200000000",
            INIT_72 => X"000000c600000000000000c700000000000000cd000000000000007c00000000",
            INIT_73 => X"00000000000000000000004200000000000000bc00000000000000d800000000",
            INIT_74 => X"000000900000000000000000000000000000000a000000000000000000000000",
            INIT_75 => X"0000006c000000000000009500000000000000a1000000000000009000000000",
            INIT_76 => X"000000ca00000000000000a800000000000000b600000000000000b600000000",
            INIT_77 => X"0000000900000000000000000000000000000036000000000000009900000000",
            INIT_78 => X"00000069000000000000004c0000000000000004000000000000001100000000",
            INIT_79 => X"000000b2000000000000004300000000000000a800000000000000b200000000",
            INIT_7A => X"0000005a00000000000000b300000000000000a400000000000000b800000000",
            INIT_7B => X"0000002900000000000000280000000000000000000000000000001200000000",
            INIT_7C => X"00000035000000000000002e000000000000001e000000000000002000000000",
            INIT_7D => X"000000a3000000000000009b0000000000000082000000000000006b00000000",
            INIT_7E => X"0000000d000000000000007100000000000000ad00000000000000ba00000000",
            INIT_7F => X"0000002d00000000000000240000000000000027000000000000001300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE53;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE54 : if BRAM_NAME = "samplegold_layersamples_instance54" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002200000000000000280000000000000000000000000000001500000000",
            INIT_01 => X"000000a10000000000000076000000000000005d000000000000006d00000000",
            INIT_02 => X"000000000000000000000004000000000000009400000000000000a800000000",
            INIT_03 => X"0000000000000000000000050000000000000005000000000000001700000000",
            INIT_04 => X"00000000000000000000001c0000000000000011000000000000000000000000",
            INIT_05 => X"0000003c00000000000000320000000000000027000000000000000000000000",
            INIT_06 => X"0000002300000000000000000000000000000000000000000000002700000000",
            INIT_07 => X"0000002c000000000000002c0000000000000020000000000000001e00000000",
            INIT_08 => X"0000000c00000000000000130000000000000022000000000000002500000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_0A => X"0000001e00000000000000200000000000000000000000000000000000000000",
            INIT_0B => X"00000028000000000000002e0000000000000000000000000000002600000000",
            INIT_0C => X"0000000000000000000000020000000000000013000000000000002200000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"00000020000000000000001a000000000000001a000000000000000000000000",
            INIT_0F => X"00000015000000000000000b000000000000000e000000000000000000000000",
            INIT_10 => X"0000002700000000000000260000000000000004000000000000001100000000",
            INIT_11 => X"0000001200000000000000210000000000000022000000000000002d00000000",
            INIT_12 => X"0000000000000000000000000000000000000012000000000000001100000000",
            INIT_13 => X"0000001d00000000000000080000000000000005000000000000000000000000",
            INIT_14 => X"0000002f0000000000000033000000000000002b000000000000002100000000",
            INIT_15 => X"0000002300000000000000090000000000000015000000000000001a00000000",
            INIT_16 => X"0000000000000000000000000000000000000080000000000000004300000000",
            INIT_17 => X"000000220000000000000022000000000000002e000000000000001800000000",
            INIT_18 => X"00000029000000000000002a0000000000000028000000000000001e00000000",
            INIT_19 => X"00000088000000000000007b0000000000000023000000000000002400000000",
            INIT_1A => X"0000002400000000000000000000000000000000000000000000007f00000000",
            INIT_1B => X"0000001f00000000000000250000000000000026000000000000003700000000",
            INIT_1C => X"0000003d0000000000000033000000000000001d000000000000002200000000",
            INIT_1D => X"000000670000000000000076000000000000007b000000000000003900000000",
            INIT_1E => X"0000003300000000000000290000000000000023000000000000001c00000000",
            INIT_1F => X"000000230000000000000029000000000000002d000000000000002000000000",
            INIT_20 => X"0000002d000000000000003b0000000000000034000000000000001400000000",
            INIT_21 => X"00000049000000000000008a000000000000006d000000000000006400000000",
            INIT_22 => X"0000002500000000000000320000000000000009000000000000002900000000",
            INIT_23 => X"0000001900000000000000200000000000000039000000000000003c00000000",
            INIT_24 => X"0000007500000000000000130000000000000015000000000000002600000000",
            INIT_25 => X"00000094000000000000007d000000000000008b000000000000007c00000000",
            INIT_26 => X"00000035000000000000002f0000000000000051000000000000007c00000000",
            INIT_27 => X"00000018000000000000001d0000000000000027000000000000003800000000",
            INIT_28 => X"000000ed00000000000000bc0000000000000023000000000000002400000000",
            INIT_29 => X"00000096000000000000009000000000000000d600000000000000fc00000000",
            INIT_2A => X"0000003600000000000000310000000000000033000000000000004c00000000",
            INIT_2B => X"0000000b00000000000000150000000000000024000000000000003500000000",
            INIT_2C => X"0000008000000000000001140000000000000105000000000000000000000000",
            INIT_2D => X"0000003a00000000000000470000000000000058000000000000007600000000",
            INIT_2E => X"0000003500000000000000380000000000000035000000000000002100000000",
            INIT_2F => X"000000040000000000000011000000000000000f000000000000001d00000000",
            INIT_30 => X"0000004b0000000000000057000000000000009c00000000000000e100000000",
            INIT_31 => X"0000000e00000000000000130000000000000001000000000000001e00000000",
            INIT_32 => X"00000031000000000000002f0000000000000019000000000000001600000000",
            INIT_33 => X"0000004f0000000000000012000000000000001e000000000000001100000000",
            INIT_34 => X"0000002c000000000000003d0000000000000038000000000000004500000000",
            INIT_35 => X"0000000f00000000000000150000000000000027000000000000001500000000",
            INIT_36 => X"00000021000000000000003c000000000000004f000000000000001a00000000",
            INIT_37 => X"000000320000000000000024000000000000001e000000000000001a00000000",
            INIT_38 => X"0000001b000000000000000a000000000000002d000000000000004000000000",
            INIT_39 => X"0000002000000000000000090000000000000024000000000000000200000000",
            INIT_3A => X"0000000b000000000000002b0000000000000025000000000000003400000000",
            INIT_3B => X"000000040000000000000018000000000000002e000000000000001600000000",
            INIT_3C => X"0000001f00000000000000220000000000000000000000000000000000000000",
            INIT_3D => X"0000000500000000000000010000000000000000000000000000000800000000",
            INIT_3E => X"0000000500000000000000000000000000000005000000000000001300000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"00000000000000000000000d000000000000000f000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000003a000000000000002c000000000000000e000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000027000000000000003f00000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000003300000000000000230000000000000004000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000013000000000000000f00000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"00000025000000000000001b0000000000000000000000000000000900000000",
            INIT_4C => X"0000000000000000000000000000000000000002000000000000001700000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"00000000000000000000003a0000000000000060000000000000004d00000000",
            INIT_4F => X"0000000000000000000000290000000000000034000000000000001a00000000",
            INIT_50 => X"0000000000000000000000000000000000000002000000000000000c00000000",
            INIT_51 => X"00000000000000000000001b0000000000000008000000000000000500000000",
            INIT_52 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000001900000000000000000000000000000000000000000000005700000000",
            INIT_54 => X"0000000c00000000000000000000000000000011000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000330000000000000000000000000000000000000000",
            INIT_57 => X"00000000000000000000001b0000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000080000000000000013000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000c00000000000000620000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000019000000000000001400000000",
            INIT_5C => X"000000050000000000000000000000000000000b000000000000001200000000",
            INIT_5D => X"0000001300000000000000170000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000190000000000000026000000000000000e00000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000005f00000000000000000000000000000004000000000000000f00000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000002a00000000",
            INIT_62 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000002100000000000000090000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_69 => X"0000003b00000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"00000000000000000000001b0000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_6E => X"000000000000000000000015000000000000001e000000000000000d00000000",
            INIT_6F => X"000000000000000000000006000000000000001e000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_71 => X"0000000000000000000000010000000000000000000000000000000f00000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_74 => X"00000019000000000000001c0000000000000000000000000000000000000000",
            INIT_75 => X"0000001500000000000000000000000000000000000000000000000a00000000",
            INIT_76 => X"0000001200000000000000000000000000000000000000000000000400000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000023000000000000000200000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000c00000000000000000000000000000000000000000000000100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE54;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE55 : if BRAM_NAME = "samplegold_layersamples_instance55" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000004000000000000000e000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_04 => X"0000004b00000000000000000000000000000005000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"00000000000000000000002f0000000000000000000000000000000000000000",
            INIT_08 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000020000000000000000000000000",
            INIT_0C => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_0E => X"0000004300000000000000000000000000000007000000000000000000000000",
            INIT_0F => X"0000000100000000000000000000000000000000000000000000004600000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_12 => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000002300000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000260000000000000028000000000000004800000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000002400000000000000960000000000000000000000000000000000000000",
            INIT_1E => X"0000000300000000000000230000000000000000000000000000005400000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000004f00000000000000220000000000000000000000000000000000000000",
            INIT_21 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"00000018000000000000004c0000000000000000000000000000002a00000000",
            INIT_23 => X"0000002f00000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000d000000000000000b000000000000002b000000000000000000000000",
            INIT_25 => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_27 => X"0000003700000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000d00000000000000000000000000000000000000000000000400000000",
            INIT_29 => X"0000002500000000000000000000000000000021000000000000001c00000000",
            INIT_2A => X"000000000000000000000075000000000000000c000000000000000000000000",
            INIT_2B => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_2C => X"000000000000000000000000000000000000001f000000000000001700000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000002500000000",
            INIT_2E => X"00000005000000000000002f0000000000000016000000000000000300000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000030000000000000013000000000000003400000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000005e00000000000000360000000000000016000000000000000000000000",
            INIT_6D => X"0000000400000000000000130000000000000042000000000000005b00000000",
            INIT_6E => X"00000000000000000000000f0000000000000011000000000000000c00000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"00000088000000000000007d000000000000005a000000000000001e00000000",
            INIT_71 => X"0000000f000000000000000e000000000000006400000000000000a000000000",
            INIT_72 => X"0000000000000000000000000000000000000005000000000000000c00000000",
            INIT_73 => X"0000002e00000000000000000000000000000000000000000000000300000000",
            INIT_74 => X"0000009e00000000000000960000000000000084000000000000007e00000000",
            INIT_75 => X"00000021000000000000003c0000000000000060000000000000007e00000000",
            INIT_76 => X"0000000e00000000000000100000000000000001000000000000000300000000",
            INIT_77 => X"0000007b00000000000000340000000000000000000000000000000800000000",
            INIT_78 => X"000000a600000000000000860000000000000070000000000000007800000000",
            INIT_79 => X"00000021000000000000006f0000000000000095000000000000009e00000000",
            INIT_7A => X"000000000000000000000000000000000000001f000000000000001e00000000",
            INIT_7B => X"0000006a0000000000000057000000000000002c000000000000000000000000",
            INIT_7C => X"000000a20000000000000091000000000000008e000000000000006c00000000",
            INIT_7D => X"0000001d0000000000000054000000000000009500000000000000a100000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_7F => X"0000007c000000000000005e000000000000003a000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE55;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE56 : if BRAM_NAME = "samplegold_layersamples_instance56" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000096000000000000007e0000000000000079000000000000009300000000",
            INIT_01 => X"000000000000000000000019000000000000005800000000000000a600000000",
            INIT_02 => X"0000002d00000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000008c00000000000000560000000000000043000000000000000000000000",
            INIT_04 => X"0000009a00000000000000950000000000000077000000000000007f00000000",
            INIT_05 => X"0000000000000000000000210000000000000033000000000000007200000000",
            INIT_06 => X"0000001a000000000000000e0000000000000002000000000000000000000000",
            INIT_07 => X"00000080000000000000006d0000000000000044000000000000000000000000",
            INIT_08 => X"00000089000000000000009a0000000000000090000000000000007c00000000",
            INIT_09 => X"0000000000000000000000000000000000000008000000000000005400000000",
            INIT_0A => X"0000001300000000000000240000000000000000000000000000000000000000",
            INIT_0B => X"000000830000000000000086000000000000007a000000000000004100000000",
            INIT_0C => X"0000003d000000000000008b000000000000009a000000000000008b00000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_0E => X"0000007400000000000000630000000000000061000000000000003200000000",
            INIT_0F => X"0000007600000000000000850000000000000085000000000000007d00000000",
            INIT_10 => X"0000001300000000000000370000000000000088000000000000009900000000",
            INIT_11 => X"0000000600000000000000200000000000000000000000000000000000000000",
            INIT_12 => X"000000100000000000000073000000000000008c000000000000002800000000",
            INIT_13 => X"000000720000000000000071000000000000008c000000000000006d00000000",
            INIT_14 => X"0000000c000000000000001a000000000000003c000000000000006900000000",
            INIT_15 => X"0000002800000000000000120000000000000000000000000000000000000000",
            INIT_16 => X"00000069000000000000005a0000000000000039000000000000002900000000",
            INIT_17 => X"0000006500000000000000730000000000000051000000000000008600000000",
            INIT_18 => X"0000001300000000000000110000000000000037000000000000003700000000",
            INIT_19 => X"0000002d00000000000000260000000000000014000000000000001400000000",
            INIT_1A => X"0000005a00000000000000680000000000000055000000000000003300000000",
            INIT_1B => X"00000043000000000000006d000000000000007a000000000000006100000000",
            INIT_1C => X"0000002d00000000000000100000000000000007000000000000002d00000000",
            INIT_1D => X"000000360000000000000022000000000000002b000000000000002b00000000",
            INIT_1E => X"0000004b000000000000003f0000000000000038000000000000003b00000000",
            INIT_1F => X"0000002100000000000000340000000000000049000000000000004f00000000",
            INIT_20 => X"0000002400000000000000240000000000000000000000000000003000000000",
            INIT_21 => X"0000000200000000000000190000000000000013000000000000000a00000000",
            INIT_22 => X"0000000b0000000000000000000000000000002f000000000000003100000000",
            INIT_23 => X"0000002f00000000000000290000000000000017000000000000002600000000",
            INIT_24 => X"000000010000000000000029000000000000001c000000000000000000000000",
            INIT_25 => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000800000000000000000000000000000000000000000000006e00000000",
            INIT_27 => X"0000001400000000000000330000000000000022000000000000001300000000",
            INIT_28 => X"0000002f0000000000000000000000000000001a000000000000000000000000",
            INIT_29 => X"0000001c000000000000002e0000000000000010000000000000002500000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"00000000000000000000000c0000000000000035000000000000000000000000",
            INIT_2C => X"0000001a000000000000002d0000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000027000000000000002b00000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"00000036000000000000001c000000000000000a000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_34 => X"00000010000000000000003c0000000000000033000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000001800000000000000110000000000000012000000000000001000000000",
            INIT_38 => X"0000000000000000000000000000000000000003000000000000002300000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000006c00000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000011000000000000000500000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000580000000000000000000000000000000000000000",
            INIT_3F => X"0000004800000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002400000000000000140000000000000019000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000b00000000000000120000000000000005000000000000000000000000",
            INIT_44 => X"0000001200000000000000320000000000000025000000000000000800000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_46 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000001a000000000000001e0000000000000000000000000000000000000000",
            INIT_48 => X"00000031000000000000000c0000000000000004000000000000002b00000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_4A => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_4B => X"000000000000000000000048000000000000000d000000000000000400000000",
            INIT_4C => X"00000030000000000000001d0000000000000013000000000000001100000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000f00000000000000080000000000000065000000000000003f00000000",
            INIT_4F => X"0000001b0000000000000006000000000000002f000000000000002c00000000",
            INIT_50 => X"000000000000000000000023000000000000002d000000000000001800000000",
            INIT_51 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000003300000000000000270000000000000012000000000000001a00000000",
            INIT_53 => X"00000034000000000000001f000000000000000f000000000000002c00000000",
            INIT_54 => X"0000000000000000000000000000000000000018000000000000001000000000",
            INIT_55 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"00000012000000000000003e0000000000000029000000000000002800000000",
            INIT_57 => X"00000006000000000000002b000000000000001c000000000000001a00000000",
            INIT_58 => X"00000000000000000000001f0000000000000000000000000000001900000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"000000000000000000000024000000000000001c000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_61 => X"0000006100000000000000680000000000000040000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000047000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"00000012000000000000002a00000000000000c5000000000000002200000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"000000000000000000000000000000000000001b000000000000000000000000",
            INIT_79 => X"00000020000000000000008d00000000000000ad000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000042000000000000001200000000",
            INIT_7C => X"0000000000000000000000300000000000000000000000000000000000000000",
            INIT_7D => X"00000000000000000000005b0000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"00000000000000000000000f0000000000000018000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE56;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE57 : if BRAM_NAME = "samplegold_layersamples_instance57" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"000000000000000000000048000000000000002e000000000000000000000000",
            INIT_07 => X"000000000000000000000001000000000000002c000000000000001c00000000",
            INIT_08 => X"0000000000000000000000110000000000000045000000000000000000000000",
            INIT_09 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_0A => X"0000002700000000000000230000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000011000000000000002700000000",
            INIT_0C => X"0000002700000000000000000000000000000000000000000000000200000000",
            INIT_0D => X"0000000000000000000000000000000000000019000000000000000000000000",
            INIT_0E => X"0000001d000000000000001f0000000000000036000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_10 => X"0000013b00000000000000000000000000000014000000000000000000000000",
            INIT_11 => X"0000001e00000000000000000000000000000000000000000000002100000000",
            INIT_12 => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_13 => X"000000060000000000000000000000000000000000000000000000ee00000000",
            INIT_14 => X"0000003f00000000000000c70000000000000000000000000000000000000000",
            INIT_15 => X"0000001800000000000000000000000000000000000000000000006500000000",
            INIT_16 => X"000000e600000000000000000000000000000000000000000000001b00000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"00000054000000000000009a0000000000000040000000000000000100000000",
            INIT_19 => X"0000002b00000000000000000000000000000000000000000000002a00000000",
            INIT_1A => X"0000000600000000000000150000000000000032000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000006300000000000000000000000000000031000000000000006f00000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"000000000000000000000051000000000000000000000000000000ad00000000",
            INIT_1F => X"0000003700000000000000000000000000000025000000000000000000000000",
            INIT_20 => X"0000000000000000000000660000000000000000000000000000000000000000",
            INIT_21 => X"0000007e00000000000000090000000000000000000000000000000000000000",
            INIT_22 => X"000000000000000000000000000000000000002b000000000000001f00000000",
            INIT_23 => X"0000000000000000000000080000000000000000000000000000003300000000",
            INIT_24 => X"000000000000000000000000000000000000002a000000000000000000000000",
            INIT_25 => X"0000002800000000000000520000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000003d00000000",
            INIT_27 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_28 => X"0000005100000000000000000000000000000014000000000000000000000000",
            INIT_29 => X"0000003d000000000000002e000000000000000e000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"00000000000000000000006d0000000000000000000000000000001200000000",
            INIT_2C => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000005900000000000000800000000000000000000000000000003900000000",
            INIT_2E => X"0000001300000000000000000000000000000010000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000057000000000000000000000000",
            INIT_30 => X"0000001500000000000000890000000000000000000000000000000000000000",
            INIT_31 => X"00000000000000000000008b0000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000050000000000000000000000000000008000000000",
            INIT_33 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_34 => X"0000000000000000000000130000000000000000000000000000000000000000",
            INIT_35 => X"0000004600000000000000000000000000000031000000000000000000000000",
            INIT_36 => X"00000000000000000000001c0000000000000000000000000000000000000000",
            INIT_37 => X"0000001b00000000000000290000000000000000000000000000000000000000",
            INIT_38 => X"0000000d00000000000000270000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000050000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_3C => X"000000000000000000000000000000000000004a000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000008c00000000000000000000000000000000000000000000005100000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000c00000000000000000000000000000008000000000000002a00000000",
            INIT_41 => X"0000006500000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000270000000000000000000000000000000000000000",
            INIT_43 => X"0000000e000000000000001e0000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000460000000000000000000000000000000700000000",
            INIT_45 => X"00000018000000000000005a0000000000000000000000000000000000000000",
            INIT_46 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000140000000000000047000000000000000000000000",
            INIT_48 => X"0000000000000000000000120000000000000014000000000000000000000000",
            INIT_49 => X"0000000e00000000000000000000000000000000000000000000001300000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"000000000000000000000000000000000000002e000000000000002200000000",
            INIT_4C => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000600000000000000100000000000000000000000000000000000000000",
            INIT_50 => X"0000003d00000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000004000000000000000000000000000000000000000000000001f00000000",
            INIT_52 => X"0000000000000000000000070000000000000004000000000000002d00000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_54 => X"000000000000000000000000000000000000007e000000000000005a00000000",
            INIT_55 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000002a00000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000100000000000000000000000000000000000000000000000f00000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_5B => X"000000000000000000000000000000000000000d000000000000001200000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"000000060000000000000000000000000000003e000000000000001000000000",
            INIT_5E => X"0000000000000000000000000000000000000007000000000000000d00000000",
            INIT_5F => X"0000000800000000000000050000000000000000000000000000000700000000",
            INIT_60 => X"0000000c00000000000000880000000000000068000000000000000000000000",
            INIT_61 => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000030000000000000000000000000000003100000000",
            INIT_68 => X"0000002300000000000000150000000000000005000000000000000000000000",
            INIT_69 => X"00000099000000000000001c0000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000003600000000",
            INIT_6B => X"0000000a000000000000002f0000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_6E => X"0000000400000000000000000000000000000000000000000000002900000000",
            INIT_6F => X"0000002700000000000000030000000000000000000000000000000f00000000",
            INIT_70 => X"0000001b00000000000000000000000000000000000000000000000600000000",
            INIT_71 => X"00000000000000000000001b0000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_75 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_76 => X"0000001300000000000000030000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000008900000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000003000000000000000500000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_7B => X"0000001c000000000000000c000000000000000b000000000000000000000000",
            INIT_7C => X"00000010000000000000000a0000000000000009000000000000000300000000",
            INIT_7D => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000600000000000000050000000000000004000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE57;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE58 : if BRAM_NAME = "samplegold_layersamples_instance58" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000300000000000000000000000000000004000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000024000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000003f00000000",
            INIT_08 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_09 => X"0000002e00000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000330000000000000000000000000000001d00000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000003b00000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_0F => X"00000000000000000000003a0000000000000000000000000000000000000000",
            INIT_10 => X"0000004700000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000005c00000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"000000000000000000000000000000000000001b000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000021000000000000000200000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000004d00000000",
            INIT_19 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000100000000000000000000000000000006700000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_20 => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"000000000000000000000000000000000000005c000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000006700000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000260000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000320000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000004200000000",
            INIT_30 => X"0000000000000000000000000000000000000012000000000000002900000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000002500000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_33 => X"0000000c00000000000000000000000000000048000000000000000000000000",
            INIT_34 => X"0000000300000000000000000000000000000000000000000000000100000000",
            INIT_35 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"000000000000000000000033000000000000000c000000000000005300000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000001200000000000000000000000000000012000000000000000000000000",
            INIT_3A => X"0000002e0000000000000004000000000000002d000000000000002700000000",
            INIT_3B => X"00000000000000000000008e000000000000006a000000000000001100000000",
            INIT_3C => X"000000330000000000000026000000000000002a000000000000000700000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_3E => X"0000000300000000000000000000000000000012000000000000001600000000",
            INIT_3F => X"00000019000000000000000000000000000000ad000000000000002200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000c000000000000002c0000000000000022000000000000002400000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000001700000000000000000000000000000000000000000000009c00000000",
            INIT_43 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000ac000000000000001d000000000000000c00000000",
            INIT_45 => X"0000004300000000000000000000000000000038000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000046000000000000006600000000",
            INIT_47 => X"0000003200000000000000000000000000000000000000000000000800000000",
            INIT_48 => X"000000150000000000000000000000000000005a000000000000000000000000",
            INIT_49 => X"0000003500000000000000000000000000000000000000000000006900000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000006800000000",
            INIT_4B => X"000000000000000000000062000000000000000a000000000000000000000000",
            INIT_4C => X"0000004c00000000000000220000000000000000000000000000001a00000000",
            INIT_4D => X"0000001800000000000000500000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_4F => X"00000019000000000000000b0000000000000087000000000000000a00000000",
            INIT_50 => X"0000000f000000000000002d000000000000002d000000000000000000000000",
            INIT_51 => X"000000240000000000000000000000000000004a000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"00000000000000000000002b000000000000002f000000000000003f00000000",
            INIT_54 => X"00000013000000000000001c000000000000000000000000000000ac00000000",
            INIT_55 => X"000000000000000000000000000000000000003e000000000000000000000000",
            INIT_56 => X"0000002600000000000000000000000000000000000000000000002800000000",
            INIT_57 => X"0000002900000000000000000000000000000076000000000000000000000000",
            INIT_58 => X"0000001d00000000000000110000000000000008000000000000000000000000",
            INIT_59 => X"0000002b00000000000000250000000000000000000000000000007900000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000007800000000",
            INIT_5B => X"0000000e00000000000000000000000000000000000000000000004400000000",
            INIT_5C => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"00000010000000000000002b0000000000000000000000000000007e00000000",
            INIT_5E => X"0000001000000000000000000000000000000022000000000000000700000000",
            INIT_5F => X"0000000100000000000000000000000000000000000000000000004200000000",
            INIT_60 => X"0000003300000000000000000000000000000000000000000000005000000000",
            INIT_61 => X"0000000a00000000000000000000000000000000000000000000004c00000000",
            INIT_62 => X"0000006900000000000000000000000000000010000000000000002800000000",
            INIT_63 => X"0000000c000000000000001d0000000000000000000000000000000000000000",
            INIT_64 => X"0000006800000000000000290000000000000000000000000000000000000000",
            INIT_65 => X"0000003800000000000000020000000000000001000000000000000000000000",
            INIT_66 => X"0000000000000000000000350000000000000016000000000000003a00000000",
            INIT_67 => X"0000000000000000000000000000000000000073000000000000000000000000",
            INIT_68 => X"000000000000000000000040000000000000002f000000000000000000000000",
            INIT_69 => X"0000002300000000000000030000000000000000000000000000000400000000",
            INIT_6A => X"000000000000000000000000000000000000004b000000000000002400000000",
            INIT_6B => X"0000001900000000000000140000000000000026000000000000004900000000",
            INIT_6C => X"0000000f00000000000000000000000000000001000000000000003000000000",
            INIT_6D => X"0000001300000000000000080000000000000000000000000000002f00000000",
            INIT_6E => X"0000001c00000000000000000000000000000000000000000000004400000000",
            INIT_6F => X"0000004f000000000000000f0000000000000036000000000000003c00000000",
            INIT_70 => X"00000027000000000000000e0000000000000000000000000000000000000000",
            INIT_71 => X"0000003b00000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000c00000000000000000000000000000000000000000000000900000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_75 => X"00000029000000000000000f0000000000000000000000000000000000000000",
            INIT_76 => X"0000004300000000000000000000000000000000000000000000000300000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_7A => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"000000000000000000000000000000000000001f000000000000004200000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE58;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE59 : if BRAM_NAME = "samplegold_layersamples_instance59" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000004200000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_0D => X"0000003c00000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000007400000000000000c80000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000003f00000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000004e00000000",
            INIT_14 => X"0000002a00000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"00000000000000000000000f0000000000000000000000000000000f00000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000003d00000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000100000000000000000000000000000000000000000000000d00000000",
            INIT_27 => X"0000001d00000000000000310000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_2D => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000200000000000000000000000000000000000000000",
            INIT_2F => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_32 => X"0000000000000000000000490000000000000019000000000000000000000000",
            INIT_33 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000004200000000",
            INIT_36 => X"0000001800000000000000260000000000000034000000000000000300000000",
            INIT_37 => X"00000000000000000000001b0000000000000000000000000000000000000000",
            INIT_38 => X"000000000000000000000000000000000000001a000000000000000d00000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"00000000000000000000001e0000000000000020000000000000001700000000",
            INIT_3B => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000270000000000000001000000000000002700000000",
            INIT_3F => X"00000013000000000000000b0000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000003500000000000000060000000000000019000000000000000000000000",
            INIT_42 => X"000000000000000000000015000000000000002b000000000000000000000000",
            INIT_43 => X"0000000000000000000000190000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"00000027000000000000001b0000000000000026000000000000001700000000",
            INIT_46 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_47 => X"0000000d00000000000000000000000000000010000000000000000000000000",
            INIT_48 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000430000000000000034000000000000003700000000",
            INIT_4A => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_4B => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_4C => X"0000000f00000000000000030000000000000008000000000000000300000000",
            INIT_4D => X"0000000000000000000000230000000000000027000000000000001d00000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000220000000000000007000000000000000600000000",
            INIT_51 => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000001100000000000000000000000000000014000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"00000034000000000000001f0000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000140000000000000019000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000080000000000000014000000000000001400000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000007400000000000000900000000000000038000000000000000d00000000",
            INIT_63 => X"0000007300000000000000840000000000000072000000000000005c00000000",
            INIT_64 => X"0000008b00000000000000320000000000000045000000000000006300000000",
            INIT_65 => X"0000000d000000000000009d000000000000009a000000000000009800000000",
            INIT_66 => X"000000310000000000000054000000000000008d000000000000002500000000",
            INIT_67 => X"0000006a00000000000000640000000000000049000000000000003a00000000",
            INIT_68 => X"0000007600000000000000650000000000000065000000000000003200000000",
            INIT_69 => X"0000001f00000000000000120000000000000088000000000000008000000000",
            INIT_6A => X"000000250000000000000031000000000000006a000000000000007100000000",
            INIT_6B => X"0000001c000000000000003c0000000000000042000000000000003a00000000",
            INIT_6C => X"0000004400000000000000410000000000000038000000000000005f00000000",
            INIT_6D => X"00000080000000000000002d0000000000000061000000000000005100000000",
            INIT_6E => X"000000360000000000000015000000000000003c000000000000004a00000000",
            INIT_6F => X"0000004000000000000000350000000000000037000000000000004800000000",
            INIT_70 => X"0000003600000000000000450000000000000037000000000000003800000000",
            INIT_71 => X"0000003b000000000000004e0000000000000060000000000000003300000000",
            INIT_72 => X"0000002e000000000000002b0000000000000022000000000000004a00000000",
            INIT_73 => X"0000005b000000000000002f000000000000002a000000000000002c00000000",
            INIT_74 => X"00000047000000000000004e000000000000003d000000000000003c00000000",
            INIT_75 => X"000000470000000000000033000000000000004c000000000000004400000000",
            INIT_76 => X"0000003700000000000000130000000000000031000000000000002500000000",
            INIT_77 => X"0000003300000000000000430000000000000033000000000000002900000000",
            INIT_78 => X"00000048000000000000004e000000000000004c000000000000003800000000",
            INIT_79 => X"000000160000000000000048000000000000005d000000000000005500000000",
            INIT_7A => X"0000003200000000000000330000000000000011000000000000002700000000",
            INIT_7B => X"0000003000000000000000380000000000000053000000000000002300000000",
            INIT_7C => X"0000006000000000000000480000000000000040000000000000003000000000",
            INIT_7D => X"0000000600000000000000360000000000000026000000000000006800000000",
            INIT_7E => X"00000044000000000000002b0000000000000033000000000000003f00000000",
            INIT_7F => X"0000002600000000000000450000000000000040000000000000003100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE59;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE60 : if BRAM_NAME = "samplegold_layersamples_instance60" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000061000000000000004c0000000000000042000000000000004500000000",
            INIT_01 => X"0000002f00000000000000270000000000000038000000000000001c00000000",
            INIT_02 => X"000000690000000000000059000000000000003a000000000000004200000000",
            INIT_03 => X"00000034000000000000003d0000000000000030000000000000005700000000",
            INIT_04 => X"0000003800000000000000430000000000000049000000000000003600000000",
            INIT_05 => X"00000051000000000000001c0000000000000016000000000000002500000000",
            INIT_06 => X"00000055000000000000005c000000000000005a000000000000004800000000",
            INIT_07 => X"0000003400000000000000340000000000000065000000000000006000000000",
            INIT_08 => X"000000400000000000000035000000000000003c000000000000003500000000",
            INIT_09 => X"000000630000000000000027000000000000002e000000000000004100000000",
            INIT_0A => X"00000046000000000000005b0000000000000059000000000000003b00000000",
            INIT_0B => X"0000004000000000000000390000000000000037000000000000004d00000000",
            INIT_0C => X"00000057000000000000002d000000000000003e000000000000002b00000000",
            INIT_0D => X"0000005d000000000000003b0000000000000049000000000000004400000000",
            INIT_0E => X"0000004c00000000000000480000000000000052000000000000004b00000000",
            INIT_0F => X"000000340000000000000043000000000000003a000000000000003900000000",
            INIT_10 => X"0000004e000000000000005d0000000000000031000000000000005300000000",
            INIT_11 => X"0000004300000000000000590000000000000041000000000000004b00000000",
            INIT_12 => X"0000003a00000000000000550000000000000040000000000000004d00000000",
            INIT_13 => X"0000002d000000000000002e000000000000003b000000000000004000000000",
            INIT_14 => X"0000004a00000000000000580000000000000068000000000000005b00000000",
            INIT_15 => X"0000004400000000000000490000000000000059000000000000003b00000000",
            INIT_16 => X"00000045000000000000002f000000000000004c000000000000005100000000",
            INIT_17 => X"00000045000000000000002a000000000000002e000000000000003000000000",
            INIT_18 => X"00000045000000000000004e0000000000000058000000000000004000000000",
            INIT_19 => X"000000570000000000000046000000000000004e000000000000004c00000000",
            INIT_1A => X"0000000000000000000000060000000000000000000000000000005000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000310000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_23 => X"0000000700000000000000100000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000028000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"000000000000000000000000000000000000001e000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_54 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_56 => X"000000500000000000000000000000000000000e000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_5A => X"0000000000000000000000480000000000000000000000000000000a00000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000001400000000000000380000000000000000000000000000000000000000",
            INIT_5D => X"0000002100000000000000000000000000000004000000000000000500000000",
            INIT_5E => X"0000000000000000000000000000000000000058000000000000000000000000",
            INIT_5F => X"0000000400000000000000020000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000029000000000000000000000000",
            INIT_61 => X"0000000a0000000000000029000000000000000a000000000000001400000000",
            INIT_62 => X"0000000000000000000000030000000000000000000000000000002e00000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000002c0000000000000011000000000000002e000000000000000f00000000",
            INIT_65 => X"0000003a000000000000000f0000000000000028000000000000003000000000",
            INIT_66 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_68 => X"0000005b000000000000004f0000000000000027000000000000003f00000000",
            INIT_69 => X"000000200000000000000000000000000000000c000000000000003400000000",
            INIT_6A => X"0000000000000000000000090000000000000000000000000000000200000000",
            INIT_6B => X"0000003000000000000000000000000000000006000000000000000c00000000",
            INIT_6C => X"0000003500000000000000200000000000000036000000000000002000000000",
            INIT_6D => X"0000000000000000000000160000000000000000000000000000000200000000",
            INIT_6E => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000f00000000000000000000000000000002000000000000000000000000",
            INIT_70 => X"0000001000000000000000590000000000000016000000000000004000000000",
            INIT_71 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000019000000000000000000000000",
            INIT_73 => X"0000002d00000000000000130000000000000000000000000000003a00000000",
            INIT_74 => X"0000000000000000000000070000000000000054000000000000001c00000000",
            INIT_75 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_76 => X"0000000100000000000000020000000000000000000000000000000000000000",
            INIT_77 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000130000000000000023000000000000003c00000000",
            INIT_79 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_7A => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_7B => X"0000003300000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000012000000000000005100000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"00000059000000000000003c0000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE60;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE61 : if BRAM_NAME = "samplegold_layersamples_instance61" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000210000000000000000000000000000001e00000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_03 => X"0000002600000000000000590000000000000036000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_05 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000001c0000000000000017000000000000006c000000000000002a00000000",
            INIT_08 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_09 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000007f00000000000000770000000000000091000000000000000000000000",
            INIT_0C => X"0000006e000000000000007b0000000000000083000000000000007c00000000",
            INIT_0D => X"000000a100000000000000a9000000000000001d000000000000003b00000000",
            INIT_0E => X"000000000000000000000000000000000000009e000000000000009f00000000",
            INIT_0F => X"0000008200000000000000850000000000000055000000000000008e00000000",
            INIT_10 => X"0000004300000000000000a60000000000000094000000000000008900000000",
            INIT_11 => X"000000b200000000000000b800000000000000bb000000000000006200000000",
            INIT_12 => X"000000500000000000000000000000000000000000000000000000ad00000000",
            INIT_13 => X"00000061000000000000009200000000000000a5000000000000006400000000",
            INIT_14 => X"000000b6000000000000003d0000000000000080000000000000008400000000",
            INIT_15 => X"000000bc00000000000000c400000000000000c400000000000000b900000000",
            INIT_16 => X"0000008b00000000000000980000000000000000000000000000000000000000",
            INIT_17 => X"0000005c0000000000000064000000000000009a00000000000000a100000000",
            INIT_18 => X"000000b500000000000000c20000000000000061000000000000004a00000000",
            INIT_19 => X"0000008800000000000000ba00000000000000e800000000000000dc00000000",
            INIT_1A => X"0000008f000000000000006900000000000000b5000000000000008a00000000",
            INIT_1B => X"00000053000000000000006c00000000000000aa00000000000000ad00000000",
            INIT_1C => X"000000ec00000000000000dc00000000000000a9000000000000005a00000000",
            INIT_1D => X"000000ab00000000000000b200000000000000af00000000000000c300000000",
            INIT_1E => X"000000ac000000000000009f000000000000006f00000000000000c000000000",
            INIT_1F => X"00000061000000000000006b0000000000000043000000000000009900000000",
            INIT_20 => X"000000cd00000000000000f200000000000000df000000000000009e00000000",
            INIT_21 => X"000000a500000000000000a500000000000000b700000000000000a600000000",
            INIT_22 => X"0000009b0000000000000076000000000000008d000000000000009700000000",
            INIT_23 => X"0000009000000000000000810000000000000090000000000000005500000000",
            INIT_24 => X"000000a600000000000000e400000000000000ef00000000000000de00000000",
            INIT_25 => X"000000a4000000000000008d00000000000000a500000000000000b900000000",
            INIT_26 => X"00000092000000000000008300000000000000a300000000000000b100000000",
            INIT_27 => X"000000bc00000000000000a9000000000000007c000000000000007e00000000",
            INIT_28 => X"000000ba00000000000000ba000000000000010200000000000000d300000000",
            INIT_29 => X"000000ad00000000000000aa0000000000000093000000000000008700000000",
            INIT_2A => X"000000670000000000000095000000000000009d00000000000000b800000000",
            INIT_2B => X"00000093000000000000005800000000000000a8000000000000006600000000",
            INIT_2C => X"0000009200000000000000bc00000000000000b500000000000000b400000000",
            INIT_2D => X"000000d100000000000000b900000000000000b300000000000000bb00000000",
            INIT_2E => X"000000870000000000000082000000000000009000000000000000b600000000",
            INIT_2F => X"00000091000000000000005b0000000000000073000000000000009600000000",
            INIT_30 => X"000000ac00000000000000b000000000000000c6000000000000009000000000",
            INIT_31 => X"000000a800000000000000ae00000000000000ba00000000000000ba00000000",
            INIT_32 => X"0000004f00000000000000ab00000000000000ae00000000000000af00000000",
            INIT_33 => X"0000007800000000000000760000000000000092000000000000007e00000000",
            INIT_34 => X"000000cf00000000000000ad00000000000000b500000000000000c800000000",
            INIT_35 => X"000000a800000000000000a9000000000000009700000000000000d800000000",
            INIT_36 => X"00000080000000000000006b000000000000006a00000000000000b400000000",
            INIT_37 => X"000000c2000000000000005a000000000000007e000000000000009700000000",
            INIT_38 => X"000000d300000000000000ca00000000000000a000000000000000b000000000",
            INIT_39 => X"0000009a00000000000000a700000000000000bb000000000000004600000000",
            INIT_3A => X"00000089000000000000006b0000000000000072000000000000006400000000",
            INIT_3B => X"000000a300000000000000ba000000000000006b000000000000006400000000",
            INIT_3C => X"0000008000000000000000ac00000000000000cb000000000000008500000000",
            INIT_3D => X"000000390000000000000075000000000000008700000000000000a700000000",
            INIT_3E => X"000000520000000000000056000000000000005f000000000000006900000000",
            INIT_3F => X"0000006e00000000000000980000000000000099000000000000007300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007d00000000000000b700000000000000b300000000000000c000000000",
            INIT_41 => X"0000005300000000000000380000000000000059000000000000006b00000000",
            INIT_42 => X"0000006800000000000000650000000000000049000000000000006400000000",
            INIT_43 => X"000000000000000000000031000000000000005f000000000000001200000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"00000011000000000000003b0000000000000000000000000000000000000000",
            INIT_46 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000054000000000000004a00000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"00000000000000000000000000000000000000dc000000000000000000000000",
            INIT_4A => X"0000002c00000000000000170000000000000000000000000000000000000000",
            INIT_4B => X"000000000000000000000013000000000000001b000000000000007100000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000006b00000000",
            INIT_4E => X"000001020000000000000094000000000000004c000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000330000000000000001000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_52 => X"000000000000000000000000000000000000005c000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000004900000000",
            INIT_54 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000003300000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000050000000000000000000000000000001c00000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000005200000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000700000000000000000000000000000000000000000000003000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_6C => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000003500000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000003700000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000003e000000000000004e0000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000005f00000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000200000000000000dc0000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE61;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE62 : if BRAM_NAME = "samplegold_layersamples_instance62" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000003f00000000000000000000000000000103000000000000000000000000",
            INIT_04 => X"0000002f00000000000000640000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000080000000000000000000000000000000600000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000760000000000000000000000000000000000000000",
            INIT_08 => X"0000001900000000000000120000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000011000000000000001900000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_0B => X"000000000000000000000000000000000000004f000000000000000000000000",
            INIT_0C => X"000000540000000000000000000000000000000b000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_10 => X"0000006100000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000340000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"00000000000000000000000000000000000000d2000000000000000000000000",
            INIT_17 => X"00000000000000000000005b0000000000000000000000000000001200000000",
            INIT_18 => X"00000000000000000000004500000000000000c2000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000003200000000000000000000000000000035000000000000000000000000",
            INIT_1C => X"00000068000000000000007a00000000000000b1000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"000000000000000000000004000000000000001e000000000000000000000000",
            INIT_1F => X"0000001800000000000000000000000000000005000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"000000000000000000000000000000000000002e000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000043000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000180000000000000000000000000000000200000000",
            INIT_28 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000005300000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"000000000000000000000014000000000000001e000000000000000000000000",
            INIT_2C => X"0000000e00000000000000010000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000180000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_30 => X"0000000000000000000000460000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"00000007000000000000000f000000000000002d000000000000001e00000000",
            INIT_6D => X"00000006000000000000002a0000000000000026000000000000003200000000",
            INIT_6E => X"00000027000000000000000f0000000000000035000000000000000000000000",
            INIT_6F => X"000000000000000000000000000000000000002f000000000000003000000000",
            INIT_70 => X"000000000000000000000000000000000000001c000000000000002000000000",
            INIT_71 => X"0000000000000000000000000000000000000014000000000000001500000000",
            INIT_72 => X"0000002400000000000000150000000000000009000000000000001400000000",
            INIT_73 => X"0000002300000000000000000000000000000000000000000000002300000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_75 => X"0000000000000000000000190000000000000000000000000000000200000000",
            INIT_76 => X"00000009000000000000000a0000000000000009000000000000001600000000",
            INIT_77 => X"0000000300000000000000000000000000000034000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000002f00000000000000170000000000000000000000000000000000000000",
            INIT_7B => X"000000000000000000000008000000000000000b000000000000000800000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000010000000000000002000000000000000000000000",
            INIT_7E => X"0000000e000000000000001a000000000000002d000000000000001400000000",
            INIT_7F => X"0000000000000000000000000000000000000022000000000000001200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE62;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE63 : if BRAM_NAME = "samplegold_layersamples_instance63" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000002200000000000000070000000000000015000000000000000000000000",
            INIT_02 => X"0000001200000000000000250000000000000025000000000000003e00000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000002600000000000000160000000000000013000000000000000800000000",
            INIT_06 => X"000000000000000000000000000000000000001e000000000000002800000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000002400000000000000000000000000000007000000000000000100000000",
            INIT_09 => X"0000001800000000000000380000000000000000000000000000001b00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_0B => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000001300000000000000000000000000000000000000000000000700000000",
            INIT_0D => X"0000001e000000000000002b0000000000000041000000000000002400000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000140000000000000016000000000000000000000000",
            INIT_11 => X"000000040000000000000007000000000000001f000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000040000000000000014000000000000001b00000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_18 => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"000000000000000000000000000000000000001b000000000000003100000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_1B => X"0000000000000000000000040000000000000007000000000000000500000000",
            INIT_1C => X"0000003500000000000000210000000000000000000000000000000800000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000003a00000000",
            INIT_1E => X"0000001200000000000000070000000000000003000000000000000000000000",
            INIT_1F => X"0000000800000000000000000000000000000004000000000000000200000000",
            INIT_20 => X"0000003e00000000000000350000000000000027000000000000000c00000000",
            INIT_21 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"00000004000000000000001e0000000000000000000000000000000400000000",
            INIT_23 => X"0000000000000000000000030000000000000006000000000000000600000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000001200000000000000150000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000060000000000000008000000000000001200000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000004c00000000000000540000000000000076000000000000000300000000",
            INIT_2D => X"0000000600000000000000450000000000000042000000000000003f00000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000002900000000000000090000000000000003000000000000008400000000",
            INIT_31 => X"00000000000000000000001e000000000000003f000000000000003c00000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000009100000000000000050000000000000000000000000000000000000000",
            INIT_34 => X"0000003c00000000000000600000000000000017000000000000002200000000",
            INIT_35 => X"00000000000000000000002d0000000000000021000000000000002d00000000",
            INIT_36 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_37 => X"000000480000000000000075000000000000004b000000000000000500000000",
            INIT_38 => X"00000059000000000000004e0000000000000059000000000000006100000000",
            INIT_39 => X"0000000000000000000000020000000000000035000000000000004900000000",
            INIT_3A => X"00000051000000000000000f0000000000000000000000000000000000000000",
            INIT_3B => X"0000003b000000000000000f000000000000008c000000000000004d00000000",
            INIT_3C => X"00000018000000000000002d000000000000004f000000000000005e00000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_3E => X"000000390000000000000064000000000000003d000000000000000000000000",
            INIT_3F => X"0000008e000000000000009b0000000000000075000000000000003e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006200000000000000730000000000000067000000000000007800000000",
            INIT_41 => X"00000000000000000000002c0000000000000041000000000000004000000000",
            INIT_42 => X"000000860000000000000006000000000000004d000000000000002600000000",
            INIT_43 => X"00000057000000000000002e0000000000000014000000000000004400000000",
            INIT_44 => X"0000001300000000000000220000000000000000000000000000002400000000",
            INIT_45 => X"0000003200000000000000000000000000000014000000000000000000000000",
            INIT_46 => X"0000003600000000000000570000000000000037000000000000005e00000000",
            INIT_47 => X"00000053000000000000001c0000000000000046000000000000005f00000000",
            INIT_48 => X"0000004300000000000000560000000000000059000000000000004a00000000",
            INIT_49 => X"0000007d00000000000000220000000000000000000000000000007000000000",
            INIT_4A => X"0000004f000000000000004c000000000000005b000000000000003500000000",
            INIT_4B => X"0000007800000000000000690000000000000045000000000000004000000000",
            INIT_4C => X"0000004800000000000000640000000000000064000000000000007800000000",
            INIT_4D => X"0000004600000000000000820000000000000029000000000000000000000000",
            INIT_4E => X"0000002500000000000000290000000000000049000000000000003c00000000",
            INIT_4F => X"0000002400000000000000340000000000000000000000000000009000000000",
            INIT_50 => X"0000000000000000000000490000000000000072000000000000000000000000",
            INIT_51 => X"0000005000000000000000000000000000000081000000000000004200000000",
            INIT_52 => X"0000003700000000000000380000000000000044000000000000006300000000",
            INIT_53 => X"0000004400000000000000000000000000000000000000000000003100000000",
            INIT_54 => X"000000240000000000000000000000000000003c000000000000004900000000",
            INIT_55 => X"0000004700000000000000510000000000000061000000000000004c00000000",
            INIT_56 => X"0000000b00000000000000280000000000000034000000000000006000000000",
            INIT_57 => X"0000005a000000000000008e0000000000000046000000000000000400000000",
            INIT_58 => X"0000004000000000000000410000000000000000000000000000001800000000",
            INIT_59 => X"0000005200000000000000470000000000000058000000000000005800000000",
            INIT_5A => X"0000004100000000000000390000000000000038000000000000003400000000",
            INIT_5B => X"0000002a0000000000000044000000000000008a000000000000003f00000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000003700000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"000000c700000000000000870000000000000054000000000000005700000000",
            INIT_62 => X"000000000000000000000019000000000000005d00000000000000a700000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"000000000000000000000000000000000000001e000000000000001200000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"000000000000000000000000000000000000001e000000000000000000000000",
            INIT_6B => X"0000006500000000000000000000000000000000000000000000001100000000",
            INIT_6C => X"0000001f000000000000003e0000000000000000000000000000001500000000",
            INIT_6D => X"0000000000000000000000000000000000000006000000000000000400000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000a00000000000000000000000000000012000000000000000300000000",
            INIT_70 => X"0000004b00000000000000030000000000000000000000000000007b00000000",
            INIT_71 => X"0000005a0000000000000079000000000000003b000000000000005d00000000",
            INIT_72 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000058000000000000005a00000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"000000a3000000000000003f000000000000001b000000000000000800000000",
            INIT_76 => X"0000008e000000000000002e0000000000000000000000000000007400000000",
            INIT_77 => X"0000002900000000000000480000000000000000000000000000000000000000",
            INIT_78 => X"000000b500000000000000c90000000000000055000000000000002700000000",
            INIT_79 => X"0000004400000000000000ad00000000000000d8000000000000008300000000",
            INIT_7A => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"000000000000000000000000000000000000000000000000000000b900000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000003200000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000640000000000000012000000000000000000000000",
            INIT_7F => X"0000003800000000000000730000000000000019000000000000006800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE63;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE64 : if BRAM_NAME = "samplegold_layersamples_instance64" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007000000000000000840000000000000064000000000000007400000000",
            INIT_01 => X"0000000000000000000000000000000000000059000000000000005300000000",
            INIT_02 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000003f00000000000000210000000000000000000000000000002600000000",
            INIT_04 => X"0000004600000000000000000000000000000005000000000000000f00000000",
            INIT_05 => X"0000004400000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000003000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"000000160000000000000057000000000000005200000000000000ec00000000",
            INIT_08 => X"000000c700000000000000450000000000000060000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000028000000000000000000000000",
            INIT_0D => X"0000001000000000000000000000000000000016000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"00000030000000000000006500000000000000b9000000000000000000000000",
            INIT_10 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000b000000000000002e0000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000210000000000000058000000000000000f00000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000003100000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"000000000000000000000026000000000000000e000000000000001600000000",
            INIT_1B => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_1E => X"0000000000000000000000710000000000000000000000000000000000000000",
            INIT_1F => X"00000000000000000000005a0000000000000000000000000000000000000000",
            INIT_20 => X"0000006c00000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000002c00000000",
            INIT_22 => X"0000000000000000000000420000000000000000000000000000000000000000",
            INIT_23 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_24 => X"0000002c00000000000000170000000000000000000000000000000000000000",
            INIT_25 => X"0000002300000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000100000000000000051000000000000000000000000",
            INIT_27 => X"000000000000000000000000000000000000002d000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000062000000000000000000000000",
            INIT_29 => X"0000000f000000000000000b0000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000059000000000000005a00000000",
            INIT_2B => X"0000000000000000000000080000000000000000000000000000001c00000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_2D => X"0000006000000000000000000000000000000000000000000000001700000000",
            INIT_2E => X"0000000000000000000000050000000000000064000000000000005700000000",
            INIT_2F => X"000000000000000000000000000000000000008d000000000000000000000000",
            INIT_30 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000008f000000000000003b0000000000000000000000000000002c00000000",
            INIT_32 => X"000000000000000000000000000000000000007c000000000000005b00000000",
            INIT_33 => X"0000003200000000000000330000000000000000000000000000004100000000",
            INIT_34 => X"0000002400000000000000000000000000000000000000000000002500000000",
            INIT_35 => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_36 => X"000000030000000000000000000000000000000000000000000000f500000000",
            INIT_37 => X"0000002c00000000000000000000000000000038000000000000000000000000",
            INIT_38 => X"000000000000000000000011000000000000000000000000000000b300000000",
            INIT_39 => X"0000014900000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"00000000000000000000003e0000000000000050000000000000000100000000",
            INIT_3C => X"0000001000000000000000000000000000000000000000000000007b00000000",
            INIT_3D => X"0000000000000000000001250000000000000008000000000000000000000000",
            INIT_3E => X"000000000000000000000000000000000000003c000000000000000000000000",
            INIT_3F => X"000000da00000000000000000000000000000083000000000000002500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_41 => X"0000000000000000000000000000000000000182000000000000000400000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000009a00000000000000650000000000000019000000000000000200000000",
            INIT_44 => X"0000005000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000013500000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000003b000000000000005c0000000000000043000000000000001e00000000",
            INIT_48 => X"00000113000000000000007a0000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"00000000000000000000003c000000000000001f000000000000001300000000",
            INIT_4C => X"0000000000000000000001110000000000000053000000000000000000000000",
            INIT_4D => X"0000000000000000000000080000000000000002000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000019000000000000001e00000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000001d00000000000000430000000000000054000000000000000c00000000",
            INIT_56 => X"0000000900000000000000a10000000000000081000000000000003500000000",
            INIT_57 => X"0000001a00000000000000020000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000300000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000002c00000000000000090000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_5C => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_60 => X"0000002d00000000000000590000000000000000000000000000000000000000",
            INIT_61 => X"0000003c000000000000001d0000000000000000000000000000002000000000",
            INIT_62 => X"00000000000000000000003f0000000000000049000000000000000b00000000",
            INIT_63 => X"0000003300000000000000230000000000000024000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"000000000000000000000000000000000000001d000000000000000000000000",
            INIT_67 => X"000000000000000000000008000000000000004a000000000000000000000000",
            INIT_68 => X"0000003900000000000000da00000000000000c5000000000000002f00000000",
            INIT_69 => X"0000000000000000000000190000000000000026000000000000000000000000",
            INIT_6A => X"0000000000000000000000320000000000000063000000000000003600000000",
            INIT_6B => X"00000000000000000000006a0000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"00000037000000000000000a0000000000000000000000000000000000000000",
            INIT_70 => X"0000009e00000000000000360000000000000000000000000000007900000000",
            INIT_71 => X"0000007000000000000000190000000000000093000000000000008000000000",
            INIT_72 => X"0000001600000000000000000000000000000002000000000000003e00000000",
            INIT_73 => X"0000000300000000000000220000000000000025000000000000000000000000",
            INIT_74 => X"000000a300000000000000a7000000000000009d000000000000001000000000",
            INIT_75 => X"000000000000000000000000000000000000009000000000000000a400000000",
            INIT_76 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_77 => X"0000001700000000000000390000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000e000000000000004c0000000000000068000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000002a00000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000004100000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE64;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE65 : if BRAM_NAME = "samplegold_layersamples_instance65" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000080000000000000029000000000000007e00000000",
            INIT_01 => X"0000000200000000000000060000000000000009000000000000000a00000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_03 => X"0000001e000000000000001c000000000000000e000000000000000100000000",
            INIT_04 => X"00000020000000000000000b0000000000000000000000000000001900000000",
            INIT_05 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000005900000000000000c70000000000000000000000000000000000000000",
            INIT_0A => X"0000004f00000000000000780000000000000036000000000000002000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_0D => X"0000000000000000000000000000000000000061000000000000001600000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000006f0000000000000018000000000000000000000000000000d500000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000005c00000000000000bc0000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000190000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"00000000000000000000009a0000000000000000000000000000002a00000000",
            INIT_19 => X"0000001700000000000000170000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_1B => X"0000006700000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000d00000000000000000000000000000000000000000000000a00000000",
            INIT_1D => X"0000006d00000000000000000000000000000007000000000000002e00000000",
            INIT_1E => X"0000000200000000000000190000000000000000000000000000003f00000000",
            INIT_1F => X"000000000000000000000099000000000000003d000000000000000000000000",
            INIT_20 => X"000000000000000000000000000000000000001b000000000000009200000000",
            INIT_21 => X"0000000e00000000000000450000000000000063000000000000000300000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000006000000000",
            INIT_23 => X"000000e80000000000000000000000000000005f000000000000000000000000",
            INIT_24 => X"0000000000000000000000020000000000000022000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_27 => X"0000004100000000000000000000000000000036000000000000009900000000",
            INIT_28 => X"0000006500000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"000000140000000000000000000000000000001a000000000000000000000000",
            INIT_2A => X"0000009800000000000000000000000000000000000000000000002600000000",
            INIT_2B => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000058000000000000000000000000",
            INIT_2D => X"0000000000000000000000430000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000dd0000000000000000000000000000000000000000",
            INIT_2F => X"0000001c000000000000000f0000000000000049000000000000000000000000",
            INIT_30 => X"00000000000000000000002c0000000000000000000000000000004000000000",
            INIT_31 => X"0000000000000000000000630000000000000066000000000000004700000000",
            INIT_32 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"00000000000000000000000d0000000000000024000000000000000000000000",
            INIT_34 => X"00000095000000000000002e0000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000006e00000000",
            INIT_36 => X"0000000000000000000000510000000000000000000000000000003700000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000002f00000000",
            INIT_38 => X"00000007000000000000007e0000000000000000000000000000004900000000",
            INIT_39 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_3A => X"0000001200000000000000000000000000000071000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000290000000000000046000000000000000000000000",
            INIT_3D => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_3F => X"0000000300000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003000000000000000000000000000000037000000000000000000000000",
            INIT_41 => X"0000004c00000000000000220000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000030000000000000000000000000",
            INIT_45 => X"0000000000000000000000ef0000000000000010000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000400000000000000000000000000000000000000000000005200000000",
            INIT_49 => X"00000000000000000000000000000000000000b9000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_4B => X"0000005100000000000000050000000000000000000000000000000000000000",
            INIT_4C => X"0000000200000000000000100000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000006500000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000001400000000000000480000000000000000000000000000000000000000",
            INIT_50 => X"0000008800000000000000400000000000000029000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"00000000000000000000003c0000000000000000000000000000002000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000003a00000000000000050000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000077000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"00000000000000000000006d0000000000000022000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_5D => X"0000007e0000000000000000000000000000001d000000000000001900000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000003400000000",
            INIT_5F => X"00000060000000000000000000000000000000af000000000000002500000000",
            INIT_60 => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"00000000000000000000002f000000000000001100000000000000be00000000",
            INIT_64 => X"0000000000000000000000390000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"000000da00000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"000000000000000000000063000000000000002d000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000056000000000000000000000000",
            INIT_69 => X"00000000000000000000008b0000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000c90000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000430000000000000058000000000000001500000000",
            INIT_6C => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"000000000000000000000000000000000000002800000000000000dc00000000",
            INIT_6E => X"00000013000000000000004a0000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000010000000000000071000000000000000000000000",
            INIT_70 => X"000000c500000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000003300000000",
            INIT_72 => X"000000000000000000000000000000000000003f000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000003000000000000002200000000",
            INIT_74 => X"0000003000000000000000330000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"00000007000000000000000d0000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"00000074000000000000006a0000000000000051000000000000003a00000000",
            INIT_7B => X"0000000b00000000000000a700000000000000c800000000000000a700000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000580000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE65;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE66 : if BRAM_NAME = "samplegold_layersamples_instance66" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000c0000000000000000000000000000000000000000",
            INIT_01 => X"0000004400000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"000000000000000000000009000000000000000000000000000000a500000000",
            INIT_03 => X"0000000000000000000000260000000000000000000000000000001500000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"000000000000000000000004000000000000002b000000000000002100000000",
            INIT_06 => X"000000190000000000000016000000000000000a000000000000004000000000",
            INIT_07 => X"000000000000000000000000000000000000002d000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_0A => X"000000390000000000000000000000000000000e000000000000001b00000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"00000015000000000000004f0000000000000002000000000000000000000000",
            INIT_0E => X"0000004c000000000000004b00000000000000a5000000000000005e00000000",
            INIT_0F => X"00000008000000000000000700000000000000b6000000000000005e00000000",
            INIT_10 => X"000000000000000000000000000000000000004a000000000000000000000000",
            INIT_11 => X"0000004d00000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"00000059000000000000007d0000000000000007000000000000003f00000000",
            INIT_13 => X"0000000c00000000000000000000000000000038000000000000000000000000",
            INIT_14 => X"00000077000000000000000c000000000000003d000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000007500000000",
            INIT_16 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000005f00000000000000000000000000000000000000000000007d00000000",
            INIT_18 => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000007f00000000",
            INIT_1A => X"0000003300000000000000000000000000000032000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000024000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000250000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000074000000000000000000000000",
            INIT_20 => X"0000006f0000000000000075000000000000002f000000000000000000000000",
            INIT_21 => X"000000620000000000000032000000000000000f00000000000000b200000000",
            INIT_22 => X"0000000000000000000000000000000000000052000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000005900000000000000000000000000000000000000000000000300000000",
            INIT_25 => X"0000001100000000000000000000000000000000000000000000001200000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000001000000000000000300000000",
            INIT_28 => X"0000002c00000000000000000000000000000033000000000000000000000000",
            INIT_29 => X"0000001600000000000000000000000000000006000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_2C => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000002f00000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000001d00000000000000150000000000000042000000000000002b00000000",
            INIT_2F => X"0000003000000000000000310000000000000021000000000000001a00000000",
            INIT_30 => X"000000310000000000000016000000000000001d000000000000002200000000",
            INIT_31 => X"000000370000000000000039000000000000001b000000000000000d00000000",
            INIT_32 => X"0000005b0000000000000058000000000000003f000000000000004900000000",
            INIT_33 => X"00000004000000000000002e000000000000002d000000000000003000000000",
            INIT_34 => X"000000090000000000000018000000000000001c000000000000000000000000",
            INIT_35 => X"00000045000000000000003a000000000000003a000000000000000000000000",
            INIT_36 => X"000000b100000000000000b90000000000000097000000000000009800000000",
            INIT_37 => X"00000000000000000000007600000000000000b100000000000000c800000000",
            INIT_38 => X"00000000000000000000000f0000000000000022000000000000002800000000",
            INIT_39 => X"000000ab000000000000002f000000000000004d000000000000003900000000",
            INIT_3A => X"000000c100000000000000bf0000000000000069000000000000007000000000",
            INIT_3B => X"00000000000000000000007900000000000000a100000000000000bf00000000",
            INIT_3C => X"0000003300000000000000000000000000000023000000000000001c00000000",
            INIT_3D => X"0000009800000000000000990000000000000049000000000000004c00000000",
            INIT_3E => X"000000a800000000000000b400000000000000a6000000000000009200000000",
            INIT_3F => X"00000028000000000000001b00000000000000be000000000000009e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004d0000000000000017000000000000002a000000000000004e00000000",
            INIT_41 => X"0000009e000000000000005100000000000000b8000000000000005000000000",
            INIT_42 => X"0000009e000000000000009b00000000000000a000000000000000a900000000",
            INIT_43 => X"0000003b0000000000000020000000000000004e000000000000007a00000000",
            INIT_44 => X"00000014000000000000002e000000000000001d000000000000003a00000000",
            INIT_45 => X"000000c50000000000000097000000000000009a000000000000006200000000",
            INIT_46 => X"0000006200000000000000950000000000000088000000000000009500000000",
            INIT_47 => X"000000380000000000000000000000000000001c000000000000003300000000",
            INIT_48 => X"0000007100000000000000000000000000000010000000000000001e00000000",
            INIT_49 => X"000000760000000000000075000000000000008c000000000000009000000000",
            INIT_4A => X"0000003a00000000000000530000000000000047000000000000004900000000",
            INIT_4B => X"0000002c00000000000000190000000000000055000000000000003d00000000",
            INIT_4C => X"000000660000000000000007000000000000001d000000000000002d00000000",
            INIT_4D => X"00000069000000000000006e000000000000005a000000000000002e00000000",
            INIT_4E => X"0000006c00000000000000700000000000000096000000000000004a00000000",
            INIT_4F => X"0000005800000000000000410000000000000000000000000000006700000000",
            INIT_50 => X"00000060000000000000003c0000000000000035000000000000001800000000",
            INIT_51 => X"0000005e00000000000000800000000000000010000000000000004500000000",
            INIT_52 => X"00000056000000000000006b0000000000000066000000000000006c00000000",
            INIT_53 => X"00000042000000000000005b0000000000000037000000000000000000000000",
            INIT_54 => X"00000055000000000000001c000000000000002c000000000000005000000000",
            INIT_55 => X"0000007700000000000000740000000000000035000000000000006c00000000",
            INIT_56 => X"000000000000000000000078000000000000003a000000000000006f00000000",
            INIT_57 => X"00000076000000000000000f0000000000000069000000000000005f00000000",
            INIT_58 => X"0000003e000000000000000a0000000000000023000000000000005000000000",
            INIT_59 => X"0000004500000000000000600000000000000031000000000000000000000000",
            INIT_5A => X"0000006e00000000000000000000000000000037000000000000003d00000000",
            INIT_5B => X"000000680000000000000081000000000000005500000000000000ab00000000",
            INIT_5C => X"0000000a0000000000000020000000000000001f000000000000003d00000000",
            INIT_5D => X"0000002b00000000000000b00000000000000066000000000000002600000000",
            INIT_5E => X"00000078000000000000006d000000000000000e000000000000001f00000000",
            INIT_5F => X"00000052000000000000005a000000000000006f000000000000008600000000",
            INIT_60 => X"0000002e0000000000000022000000000000001e000000000000002000000000",
            INIT_61 => X"0000001b000000000000002200000000000000ac000000000000003900000000",
            INIT_62 => X"0000009400000000000000860000000000000080000000000000001b00000000",
            INIT_63 => X"0000002e00000000000000400000000000000053000000000000004400000000",
            INIT_64 => X"0000003e000000000000003c0000000000000033000000000000003600000000",
            INIT_65 => X"000000300000000000000027000000000000002a000000000000006e00000000",
            INIT_66 => X"0000001200000000000000290000000000000029000000000000001b00000000",
            INIT_67 => X"0000002300000000000000120000000000000010000000000000001600000000",
            INIT_68 => X"00000020000000000000002a000000000000001f000000000000003300000000",
            INIT_69 => X"00000014000000000000001b0000000000000032000000000000001600000000",
            INIT_6A => X"0000000000000000000000000000000000000018000000000000001600000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000002a000000000000002e0000000000000016000000000000000000000000",
            INIT_6D => X"0000001300000000000000130000000000000034000000000000002b00000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000002900000000000000310000000000000038000000000000000000000000",
            INIT_71 => X"00000000000000000000001d0000000000000013000000000000002c00000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"00000042000000000000002d0000000000000017000000000000001000000000",
            INIT_75 => X"0000000000000000000000000000000000000015000000000000001600000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000001a0000000000000022000000000000001a000000000000001e00000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"00000013000000000000002f0000000000000015000000000000001400000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE66;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE67 : if BRAM_NAME = "samplegold_layersamples_instance67" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000050000000000000006000000000000004a000000000000001200000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000002c00000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"00000000000000000000004f0000000000000000000000000000002000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000001200000000000000110000000000000000000000000000000400000000",
            INIT_07 => X"0000001700000000000000020000000000000000000000000000001b00000000",
            INIT_08 => X"0000000000000000000000000000000000000017000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"00000000000000000000000a0000000000000000000000000000000a00000000",
            INIT_13 => X"0000000b000000000000000a0000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"000000130000000000000015000000000000000a000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_58 => X"0000000c000000000000000a0000000000000000000000000000000000000000",
            INIT_59 => X"0000001d00000000000000000000000000000003000000000000000900000000",
            INIT_5A => X"0000000400000000000000000000000000000000000000000000000800000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000003500000000000000230000000000000001000000000000000d00000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000001100000000000000100000000000000000000000000000000000000000",
            INIT_61 => X"00000000000000000000002f000000000000001b000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE67;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE68 : if BRAM_NAME = "samplegold_layersamples_instance68" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_04 => X"0000000000000000000000000000000000000019000000000000000000000000",
            INIT_05 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000029000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000002600000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"000000d300000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000009b00000000000000a500000000000000e000000000000000cd00000000",
            INIT_10 => X"000000e000000000000000b6000000000000009a000000000000009400000000",
            INIT_11 => X"000000bc00000000000000d700000000000000e000000000000000e400000000",
            INIT_12 => X"000000f100000000000000f2000000000000009900000000000000c500000000",
            INIT_13 => X"000000950000000000000090000000000000008a00000000000000ff00000000",
            INIT_14 => X"000000c500000000000000cb00000000000000a6000000000000008800000000",
            INIT_15 => X"000000d200000000000000e300000000000000e200000000000000bc00000000",
            INIT_16 => X"000000e800000000000000fb00000000000000f900000000000000c000000000",
            INIT_17 => X"0000004400000000000000560000000000000031000000000000006700000000",
            INIT_18 => X"0000009500000000000000740000000000000056000000000000004d00000000",
            INIT_19 => X"000000ac00000000000000b900000000000000ea00000000000000e700000000",
            INIT_1A => X"0000007f00000000000000c1000000000000010200000000000000f800000000",
            INIT_1B => X"0000007800000000000000920000000000000095000000000000007b00000000",
            INIT_1C => X"000000cd00000000000000a80000000000000067000000000000007300000000",
            INIT_1D => X"000000f4000000000000009a00000000000000c800000000000000c000000000",
            INIT_1E => X"0000006f000000000000004b00000000000000bd00000000000000fd00000000",
            INIT_1F => X"0000007d000000000000006a0000000000000067000000000000007700000000",
            INIT_20 => X"000000df00000000000000b70000000000000090000000000000006f00000000",
            INIT_21 => X"0000010000000000000000e000000000000000a600000000000000d200000000",
            INIT_22 => X"0000004100000000000000240000000000000053000000000000007200000000",
            INIT_23 => X"0000005b000000000000004c000000000000004e000000000000005400000000",
            INIT_24 => X"000000f800000000000000db0000000000000077000000000000007000000000",
            INIT_25 => X"0000008300000000000000b900000000000000d000000000000000fa00000000",
            INIT_26 => X"0000005200000000000000520000000000000035000000000000002600000000",
            INIT_27 => X"00000043000000000000006f0000000000000040000000000000003100000000",
            INIT_28 => X"000000f100000000000000c400000000000000ba000000000000006400000000",
            INIT_29 => X"0000009b000000000000004f000000000000005f00000000000000ce00000000",
            INIT_2A => X"0000002c000000000000001d000000000000001c000000000000003200000000",
            INIT_2B => X"0000001d00000000000000170000000000000000000000000000001600000000",
            INIT_2C => X"000000b000000000000000da000000000000005e000000000000001f00000000",
            INIT_2D => X"000000320000000000000018000000000000008a000000000000003c00000000",
            INIT_2E => X"000000190000000000000010000000000000002e000000000000004a00000000",
            INIT_2F => X"000000450000000000000018000000000000003e000000000000001800000000",
            INIT_30 => X"0000004e00000000000000b900000000000000a1000000000000007400000000",
            INIT_31 => X"0000001400000000000000210000000000000000000000000000006200000000",
            INIT_32 => X"0000006600000000000000720000000000000033000000000000002000000000",
            INIT_33 => X"00000028000000000000008f000000000000005f000000000000006900000000",
            INIT_34 => X"0000002c000000000000003900000000000000be000000000000005700000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_36 => X"0000002a0000000000000038000000000000000c000000000000003900000000",
            INIT_37 => X"000000490000000000000036000000000000002c000000000000003000000000",
            INIT_38 => X"000000360000000000000016000000000000003f00000000000000bb00000000",
            INIT_39 => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_3A => X"000000a500000000000000590000000000000039000000000000003000000000",
            INIT_3B => X"000000940000000000000010000000000000003c000000000000000000000000",
            INIT_3C => X"0000000a000000000000007a000000000000003f000000000000003b00000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000970000000000000098000000000000006400000000",
            INIT_3F => X"0000009800000000000000a4000000000000002e000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000000000000000000027000000000000006f000000000000005f00000000",
            INIT_41 => X"0000006300000000000000020000000000000000000000000000000000000000",
            INIT_42 => X"000000000000000000000000000000000000008a000000000000006500000000",
            INIT_43 => X"0000007400000000000000790000000000000089000000000000002800000000",
            INIT_44 => X"0000000000000000000000000000000000000021000000000000002500000000",
            INIT_45 => X"0000003c00000000000000160000000000000000000000000000000000000000",
            INIT_46 => X"0000003700000000000000000000000000000000000000000000004500000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000004000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"00000018000000000000000c0000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000082000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000003100000000",
            INIT_58 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"00000000000000000000001f0000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000480000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"00000000000000000000006a0000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000002900000000",
            INIT_67 => X"000000aa000000000000004000000000000000b600000000000000cd00000000",
            INIT_68 => X"000000000000000000000000000000000000000000000000000000ea00000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000039000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000002c00000000",
            INIT_6F => X"000000550000000000000000000000000000002b000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000150000000000000000000000000000005e00000000",
            INIT_72 => X"0000000000000000000000000000000000000083000000000000000000000000",
            INIT_73 => X"0000002900000000000000000000000000000000000000000000002200000000",
            INIT_74 => X"00000000000000000000007b0000000000000000000000000000000000000000",
            INIT_75 => X"00000011000000000000000c0000000000000000000000000000000000000000",
            INIT_76 => X"000000000000000000000008000000000000011c000000000000000700000000",
            INIT_77 => X"000000000000000000000093000000000000000e000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000005200000000000000390000000000000022000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000034000000000000006200000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000900000000000000140000000000000021000000000000001100000000",
            INIT_7E => X"0000004100000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"000000000000000000000000000000000000000000000000000000ab00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE68;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE69 : if BRAM_NAME = "samplegold_layersamples_instance69" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000008000000000000000360000000000000064000000000000002c00000000",
            INIT_05 => X"00000000000000000000000d000000000000006800000000000000b200000000",
            INIT_06 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_07 => X"0000004900000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"00000000000000000000000000000000000000a0000000000000000000000000",
            INIT_0A => X"000000000000000000000000000000000000004c000000000000000000000000",
            INIT_0B => X"0000002000000000000000930000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_0D => X"00000000000000000000000000000000000000ae000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000b00000000000000000000000000000083000000000000000000000000",
            INIT_10 => X"000000000000000000000000000000000000000f000000000000001100000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000005e00000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000003500000000",
            INIT_13 => X"000000180000000000000000000000000000001a000000000000008300000000",
            INIT_14 => X"000000130000000000000076000000000000001a000000000000002600000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000008600000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000009c00000000000000340000000000000000000000000000002c00000000",
            INIT_19 => X"000000000000000000000003000000000000000100000000000000a200000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000006d00000000",
            INIT_1B => X"0000006200000000000000610000000000000004000000000000001f00000000",
            INIT_1C => X"0000002c000000000000008f000000000000005d000000000000002e00000000",
            INIT_1D => X"0000000200000000000000000000000000000000000000000000010d00000000",
            INIT_1E => X"000000000000000000000020000000000000002d000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000009800000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000d00000000000000000000000000000000000000000",
            INIT_22 => X"0000007500000000000000260000000000000000000000000000007b00000000",
            INIT_23 => X"00000046000000000000002d0000000000000048000000000000000000000000",
            INIT_24 => X"000000000000000000000082000000000000000000000000000000ab00000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"000000a400000000000000000000000000000000000000000000006800000000",
            INIT_27 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"000000000000000000000000000000000000000000000000000000e600000000",
            INIT_2A => X"00000000000000000000009a0000000000000010000000000000007900000000",
            INIT_2B => X"000000b000000000000000000000000000000043000000000000000300000000",
            INIT_2C => X"0000000000000000000000000000000000000001000000000000005700000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000004200000000",
            INIT_2E => X"0000000000000000000000bf0000000000000000000000000000000800000000",
            INIT_2F => X"0000001400000000000000270000000000000000000000000000000000000000",
            INIT_30 => X"0000005c00000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"00000000000000000000008c0000000000000087000000000000000000000000",
            INIT_33 => X"000000000000000000000030000000000000002c000000000000000000000000",
            INIT_34 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"000000000000000000000078000000000000003c000000000000000e00000000",
            INIT_37 => X"0000000000000000000000000000000000000034000000000000002800000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000600000000000000000000000000000000000000000000000e00000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000002e00000000000000030000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE69;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE70 : if BRAM_NAME = "samplegold_layersamples_instance70" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE70;

MEM_EMPTY_36Kb : if BRAM_NAME(1 to 7) = "default" generate
    BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
    generic map (
        BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
        DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
        DO_REG => 0,                     -- Optional output register (0 or 1)
        INIT => X"000000000000000000",   -- Initial values on output port
        INIT_FILE => "NONE",
        WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        SRVAL => X"000000000000000000",  -- Set/Reset value for port output
        WRITE_MODE => "WRITE_FIRST"      -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
    )
    port map (
        DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
        ADDR => bram_addr,  -- Input address, width defined by read/write port depth
        CLK => CLK,    -- 1-bit input clock
        DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
        EN => EN,      -- 1-bit input RAM enable
        REGCE => '1', -- 1-bit input output register enable
        RST => RST,    -- 1-bit input reset
        WE => bram_wr_en       -- Input write enable, width defined by write port depth
    );
-- End of BRAM_SINGLE_MACRO_inst instantiation
end generate;


end a1;