-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;


-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity bram_single is
    generic (
        DEVICE: string := "7SERIES";
        N_BRAM: integer := 0
        );

    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic_vector(2-1 downto 0);;
        DI   : in std_logic_vector(16-1 downto 0);
        ADDR : in std_logic_vector(10-1 downto 0);
        DO   : out std_logic_vector(16-1 downto 0)
    );
 end bram_single;

  architecture a1 of bram is

    begin


    MEM_IWGHT_18K_LAYER2_ENTITY0 : if N_BRAM = 0 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"-2681-aba-dc2-468-7734a571017-5ea0ea50a32218541710277-25ad-d421a10",
            INIT_01 => X"41b444f2-c110d1f13052f1d0aed-12e5-4e52f06-2ff1-7bc-56e1b8c-da22a6e",
            INIT_02 => X"1aee4eda2657172922b71e3d-2a0b05d9-12c01361-17b8091d-2d56-ac81eef-f51",
            INIT_03 => X"0be82c7a227f-51117562c6e-139-6990ac318cc2da42571380e-1f001e3c2be4",
            INIT_04 => X"-013000a-00c0006-01500000019-0010010-00d-010001f-005000b001d-01a",
            INIT_05 => X"-006-0200027002a002d0028008f003400280064002300140038-002-00a000b",
            INIT_06 => X"-0070006-02a-02a0011003f00430054008d0045003a006000070000001a-01a",
            INIT_07 => X"0019000f00000024001f0011-0020000001b-02d-0040021-028-014-0020000",
            INIT_08 => X"-002-014-023-010-028-009-021-00e002000030018-0030012003b0002-012",
            INIT_09 => X"-00c-00c001a0009-004-0020004-008-0060005-01b00260011-004000d-004",
            INIT_0A => X"-018-028-0160008-005-0240007-006-024-03800090003000f001100020007",
            INIT_0B => X"-011-003000b000e00220010000f0025-01d-00900150000-00600040000-008",
            INIT_0C => X"-03500100015001000020024000a00100003-027-009-031-0100001-017-00f",
            INIT_0D => X"00110009000e-00b001100370001-010-021000700200013-003-00d000c-01b",
            INIT_0E => X"-0190000-043-02e-03a-001-049-029-02c-06f-021-0120008-007-00c0001",
            INIT_0F => X"-006002200000012-01b-009-028-00c-022-00e0002-010-0040009-00a-01c",
            INIT_10 => X"0011-001-00a001000010018-0080005-00b-010-01000020002-015-0110001",
            INIT_11 => X"-0090002000c0007002c-008-01d001a00070010-013000d0006-0390013-01a",
            INIT_12 => X"-068000d000e0030-00500120011-00a000800040003-0120022001d-002001a",
            INIT_13 => X"-001-01d-024000a-0040016-0180000001b0008-01200210019001900020010",
            INIT_14 => X"00150012-02b-013-025001c-0200014-00b-004-006-019000e-005-0150004",
            INIT_15 => X"0002-01700030016-00100140019-001-01500100006001d0004-003-034-018",
            INIT_16 => X"000000010012001e-010000200230000-003-023-03a-022-029000000050025",
            INIT_17 => X"006e002c0011-01e-03200240026-0150069002a0043-00a-00a-0510009-065",
            INIT_18 => X"0000-00d001c003b-009-00f000700140039003e003f00460022-00f0007-01b",
            INIT_19 => X"-00b0051-002-045-042-013000200210033-016-003-023-04e-04c-0160010",
            INIT_1A => X"00020003-030-03a-0410019000c0011-014-002-00e-0080012001400000020",
            INIT_1B => X"00140034002200040013002200080018-00b-029-0130009-00e001200290020",
            INIT_1C => X"001f0021-024-0010003-01e00540036-0260023-01f-0060011-004-0260006",
            INIT_1D => X"0003-030-046-031-03f00390043000e-027-023-01c001200250038-024-011",
            INIT_1E => X"-02b0025003e0018-034-033-03a0019001f001800050004-002-027-069-072",
            INIT_1F => X"003400310042-011000c-00c0005002a001700300033000d0023001e0005-01e",
            INIT_20 => X"-003000500040023-0190007004d0010-006001d-00900050004-004-0070022",
            INIT_21 => X"-003-00e-020-01b-002001a0003001d0008000d0000-009-020001b00040010",
            INIT_22 => X"0009001f0000-01a-02e-01d0007-002-010-009000d0007-02c-010-023-026",
            INIT_23 => X"-0020000003100490023-019-024-028-022-04a-00f0028-053-039004d-02d",
            INIT_24 => X"-034-016-022-00a-020-032-0110014002400310030003800160013002a0020",
            INIT_25 => X"0011-00d-03d-0120015-00a-032002400140000-045-012-0050004-045-00f",
            INIT_26 => X"-0130001000e0026003b-00100000005-049001a-03e-006-026-0270003-00d",
            INIT_27 => X"-01c0008-01c-012-01f-017001800320013-009-0110013-005-01a-01a-023",
            INIT_28 => X"001100220014-00e-0120007-0070000-0080002-00a0008-00b-021-04d001c",
            INIT_29 => X"0019-01b-017-012-003-039-027-011-004000f000b000d001f001d0059001f",
            INIT_2A => X"003c000e00350019-03b-02d-027-012-03c00010006-00d0025-004000a000d",
            INIT_2B => X"00060026000a-00c000c001e-003-001-00b-02700060004-023-024-0160035",
            INIT_2C => X"001a00180000-01c-036000f-00f-011-0190022-02e000d0000-00500370010",
            INIT_2D => X"-020-00100310038-02a0019002e-031-01e0028001c-004-005001f001e-01d",
            INIT_2E => X"-003-004-01d0019-008000f-00400260011-0170024002c-00d-0180013-016",
            INIT_2F => X"0002000f-019000c0016001d00070038-02a-028-028001b-0040002000f-003",
            INIT_30 => X"-02c0008-002-016-032-00c0005-02e-0140036-03100040038-038-032002c",
            INIT_31 => X"002d-010-00a0023-02c-03100310007-010000a0001003c-01b00080028-03a",
            INIT_32 => X"-01b00240006-037-023001f0000001f-00c-01a-0080001-001-01a00180011",
            INIT_33 => X"0000-00a-0050009001f-01a-017000f0010000d000b0004-0060024-002-018",
            INIT_34 => X"0023-00a0007-00e00000002-00d001d0031-028-0060022-037-034001f0000",
            INIT_35 => X"-00d-04900160014-012-0080003-035-0150032000d001b0027002200260036",
            INIT_36 => X"00300003-015-020-003-018-0490037001d-01d-024-0010023-03d-0270023",
            INIT_37 => X"-042-0130020-01c002e002d-017-0040030-01b-018002c00020017001f000f",
            INIT_38 => X"003e004900250044002c-0080013001c-024000f0035-028-01d-0040005-004",
            INIT_39 => X"-03600300013001a0012001b0006-015-00c0029-041-001000e-0400003003e",
            INIT_3A => X"-003000000000003-003-005000c-0120008-010-01c000a-016-008-00d-00a",
            INIT_3B => X"-016-00d0006-013000b-019-00c-00a-00a000e0000-0100008-00b-010-018",
            INIT_3C => X"000d-0150005-003-014000000050000-006-00a0003-012-013-00f0007-00c",
            INIT_3D => X"0000-005000200110006-00a-005-00c-00d-010-009-00d0006-003-003000d",
            INIT_3E => X"000a00050007-0120000-015-0230000000c-0190002000900040007-007-014",
            INIT_3F => X"-004-0130008-00100020002-009-007-004-001-015000f-00e000300000010",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY0;


    MEM_IWGHT_18K_LAYER2_ENTITY1 : if N_BRAM = 1 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"-016-006-021-015-0080011-00800070004-00e-00400080005-0080005-00c",
            INIT_01 => X"0000-0150002-00c-004-01f-003-01e000a000b-00e0000-00300000001-012",
            INIT_02 => X"-007-012000800120007000b-00b-008-014-00f00030005-00e-005-005-00b",
            INIT_03 => X"000b-0100000-009-018-001-0050000-013-0010006-014-015-011-017-019",
            INIT_04 => X"-003-006-00c0000-002-00a000a-00e-00b-00c-008-016000c-002-00f0000",
            INIT_05 => X"-010-019-00c-015-014000f-013-007-005-015-005-00d-013-00c00030004",
            INIT_06 => X"0001-0060007-012000b-00e-002000c0005-0170000-015-008-019-0040004",
            INIT_07 => X"0003-004-0160000-0080003-00e-013-0160005-001-016-0180005-0040000",
            INIT_08 => X"-020-012-0100001-00d0009-00a-0100009-013-00500020004001100000001",
            INIT_09 => X"00000005-014000b000b-01600100008-0140002-00a-018-016-00e-002-010",
            INIT_0A => X"-007-00f-00f-00b0009-00a00070007-013000b000b0001-006-00f0009-00a",
            INIT_0B => X"0006-0060008000d0009-005-00c-00d-011-01d00040012-00d-0090008-010",
            INIT_0C => X"0009001b0017-005-00a0001000c0001-004-01d-02b-01d0012003e-006-01a",
            INIT_0D => X"-012-00d-04a-02a-016000c-009-0270011001e0007-01a-0320032-01c-042",
            INIT_0E => X"-02b-021-01c-03e-030-032-033000a-02f-030-008-02a-01b-03d-03d-02d",
            INIT_0F => X"-041-016-017-00200160016002300250031001b000f-0050008001c0036-001",
            INIT_10 => X"00160018-01f-009-013000e001f-00e00070008-00a002b0011-00f0003000e",
            INIT_11 => X"0024-007-03d-010-04a-031-055-029-022000f0009000300000028003a000e",
            INIT_12 => X"-006000f001d-01700140001-00c0024-010-003-012-0240016001a-009-00c",
            INIT_13 => X"-0220000-00b-020-021-00d0038001c-04b-031-056-04e-015-01e-0160000",
            INIT_14 => X"0000-001-006-00e00160003000c000f-0060000-011-0200000-004-01b-038",
            INIT_15 => X"0027000d-018002a0041006000120035001d000f001a0017-013003f0022-007",
            INIT_16 => X"0046003700060000-0080006002c000c-01c0000-02c0016-003000a000d0001",
            INIT_17 => X"00020004-0020002002b0018001f000d001300160013-00500040002-01a000e",
            INIT_18 => X"0010-02100150014-006000d-026001b-010-032-012-01d-009-0140002-00b",
            INIT_19 => X"-00e-0010022003f0032001a001200110017-032-019002e-00b-02a0023-014",
            INIT_1A => X"-042-013-026-026-019002e-02a-00f00050008-034-020-01b-02c-017-012",
            INIT_1B => X"000800060028000b-008-02b0006-017-017001c-009-003-059-04a0015-027",
            INIT_1C => X"-039-02f-044-029-00d000d-004-02700240003-00f00140006001100290005",
            INIT_1D => X"0014000c-009-0170011000f-010-00a-015-014-01b000a-017-025-014-00a",
            INIT_1E => X"000f-014-003-001-010001c-008-00b-007003800260005000c-00f-017-00d",
            INIT_1F => X"000e002c-006-053-06e-035-061-0530036-019-02b-005-073-03c-030-01b",
            INIT_20 => X"-0350004-025-002-00e-049-014-010-062-03a-02f-009-015002300350022",
            INIT_21 => X"0012001a00310000-003-013-020-028-022-00d-003-0280008-00e-004001b",
            INIT_22 => X"000a00120007-011001c-01d-0120019-002-02c-00c-046-049-020-02d-00f",
            INIT_23 => X"000c-0060024000d002d0018-00f001500180000-006-029-021-011-01c-020",
            INIT_24 => X"000e00160058-018-024-02000070000-0430010-01e-042-004000d00100000",
            INIT_25 => X"-00300070001-0120006001000140000001900120016001a000b001000190008",
            INIT_26 => X"001a-01c-002-011-01d-012-007000400200012000f0011-008000e0000-02b",
            INIT_27 => X"-01b-02f-023-017-0440001-029-0130002-00300030016003e000f-0080014",
            INIT_28 => X"-003-02d-0070007-03c-002000a-00600150022-01e0000001200110002000d",
            INIT_29 => X"0023-0250007000a0014002500210023001c0034-0190005000d000c0005002f",
            INIT_2A => X"00090027003c-0030005-001-00c000b-01b00050016-017-0130006-038-013",
            INIT_2B => X"-01b-008-02e-006000a000f0013002b001c-04d-022-005-008-00f0033-007",
            INIT_2C => X"-01e001b-00e-0120007000e00050015001a003100220021-009002e000a-02e",
            INIT_2D => X"00440004-014-009-00f-007-03d00070005-00100000002-042-088-043-02c",
            INIT_2E => X"-048-033-010-02b-02d000f000b0015-00400210030001e-016-008000b001d",
            INIT_2F => X"001000040019001a-004-005002f00170019001e00370017-0080025000c-03a",
            INIT_30 => X"-028-01b-00f-00f-016-005-007-00e-0150026002a0029003200250015-009",
            INIT_31 => X"-045-0480000000e-003-01e-0160026-01b-00b001a-00a00120031-02a-026",
            INIT_32 => X"000d-018-0130023-026001c-016002e00350016-010001a0007000400080005",
            INIT_33 => X"00150036001c0027003100330038000200240019-007-013-00e-033-02d-00e",
            INIT_34 => X"-00f-00f-04b-05f-055-021-032-0350028002600220053003f0037000e0003",
            INIT_35 => X"-010-005-00e-00a000a0001000b0014-010000c0005-0020017001b000a000b",
            INIT_36 => X"-022-00f-023000b-0110021000200000040-004-0030030002100210020-01b",
            INIT_37 => X"00190013-018-00b-00e-022-03c-019-034-03f-036-012-023-02e000a0025",
            INIT_38 => X"002c0022003a00230006-00d00130018-010-009-001-002000e-01c001a002c",
            INIT_39 => X"00110002-00b-055-04d-013-052-06b-05d001a0005001300220016002f-00b",
            INIT_3A => X"00080006-02d000c0016-02b-0060031-0140034001100340032001d-00a0016",
            INIT_3B => X"-011-010-00b-00f0004-0120004-032-003-017-0040004001500250027001a",
            INIT_3C => X"000e0016-005001f001500110029002d001f00170002000f-01b-030-01d000b",
            INIT_3D => X"0012-001-017000a-002-01b-015-005002b-006-032-018-024-054-045-011",
            INIT_3E => X"-033000700020013-050-054-04a-03a-04a-055001900110003-014-0020024",
            INIT_3F => X"-020-0010003001a000a-014000b-008-046-04a-046-049-004-008-002-033",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY1;


    MEM_IWGHT_18K_LAYER2_ENTITY2 : if N_BRAM = 2 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0010002f-00c004e002e0009-01e-022-010-02d-04d-01c-03d-03d-00a0005",
            INIT_01 => X"0006-02d-01100000010-008-002-007-00b001f0013-0110016-0020010001e",
            INIT_02 => X"-003000f000c-00b000b000e000c0012-005-00e-002-014000c-005-00c-01b",
            INIT_03 => X"-006-01900090001-0040001-00d0000-0080002-006-01a0001-016-00b0000",
            INIT_04 => X"0005-001-00a0000-00c-0120003-01b-00a-006-012-01500060001-014-017",
            INIT_05 => X"000a00090000-00c-00c00010005-002-005-0010011-015-00b-013-007-011",
            INIT_06 => X"-00a00060004-01800050007-00b0004-020-00f-00a-00500050005-001-01d",
            INIT_07 => X"00050000-0100006-004000b-0110014-0130006-01d-00f-004-01b-01d0000",
            INIT_08 => X"-01b0000-0190003-004-00c000d-0030008-00e-006000c0006001300130007",
            INIT_09 => X"-012-015000d-0080013-006-00d-007-00800040000-00e0007000000030000",
            INIT_0A => X"-003-016-009000e-008000d-001-01c-00800040008-013000b-00e-010-003",
            INIT_0B => X"-010-01600010000-009-002000c-003-010-008-005-009-003-014-00e0005",
            INIT_0C => X"-0100004-0190003-005-002-012-01300070009-00c-0080000-017-0190009",
            INIT_0D => X"00060001-00d-017-00b-00e-001-016-01d-00f-007-0110008-004-011-008",
            INIT_0E => X"000a-0190002-004-00f0005-0070009-004000e0011-00f-012000e-00b-008",
            INIT_0F => X"-005-007-00a-01a-007-010-006-016-00b0001000b-009-003-01f0004-014",
            INIT_10 => X"-016-004-01a0003-00f-00f-00f-0260000-0140010-00b-00d001100020007",
            INIT_11 => X"00140007-011000f-006000a0003-01300040001-002-013-018-001000d-009",
            INIT_12 => X"-00f-00e0000000a0000-00400010002-003-001-0080001-00b000500040006",
            INIT_13 => X"0001-00200050006-00a0008-004-004-0170003-0100000-014-015000b0000",
            INIT_14 => X"0000-007000f-0150003-003-009-003000a-00f0004-00400020015-025-024",
            INIT_15 => X"-048-0270022-012-009001900100021002e00050005001c002f000a-00c0030",
            INIT_16 => X"002e000200480022-01a-0130028-00a0014001e003600420019-009001d0011",
            INIT_17 => X"002b0048-0130027003b0034-023000f000a-024-037-002-02b-00c00290024",
            INIT_18 => X"000d-00f-001-026-003-01a000c0016-018-0020003-01d-012001a001c-016",
            INIT_19 => X"0010-0240010002f-013-02f00000006-0100001-014-0150002-042-021-001",
            INIT_1A => X"-047-039-01e-006-0040006-011-006000f-018-00c0015-00b-015-022-005",
            INIT_1B => X"-0040017-027-011-00d-010000a-0320000-0120003-041-027-008-015-009",
            INIT_1C => X"0013-010000d000f-00700020000-003-02f-0190006-016-020-021-037-022",
            INIT_1D => X"0018-0070015-0430024-02a-056-022000a-0110013002e-03f-0270000-040",
            INIT_1E => X"-011-0100012-00c000700110031002e000e002e-005-016-0190000-0040004",
            INIT_1F => X"-00600020005-011000100040022-010-00b0002-002-006-00f-0210009-006",
            INIT_20 => X"000f-0050004-004-016-010-04d-00e0023-026-0090005-00c-024-005-035",
            INIT_21 => X"-0060018-04f-01a000f-05e-0200016-03c-02b004d001e000200240008-01b",
            INIT_22 => X"-010-001-014-027-02f-012-01d-044-0040012-0180009000c000c-01e0024",
            INIT_23 => X"-008-031000a-015-008001a-02200080005-021-033-01c0014002a001d002a",
            INIT_24 => X"0016002a005600690038-01700250004-035-005-00b-02a-065-00a001a0003",
            INIT_25 => X"0015-017-00a-002-02a00050028000a-0030007-00400060017001f0018000e",
            INIT_26 => X"0005-015-017-009001e00020001000f-010001e-002-010002c002f00220019",
            INIT_27 => X"00160000-01c-02c-01b-00700110012-008001a00100027-00d-01b00050037",
            INIT_28 => X"0006002500350006-011-030-01400100000-02600000046-016-00c-0030022",
            INIT_29 => X"0026-007000800060000001a-004-00b-021001d000d00050026000800180020",
            INIT_2A => X"0000-00d00280013-015-0050009-00d-011-019-03000110011-00e-014-00f",
            INIT_2B => X"-030-02700080022-03f-0150018-018-02f0020002d0014-0090031000d0014",
            INIT_2C => X"0013-003-016-029-01f0008-038-01c000d-031-021-005-008001a0011-003",
            INIT_2D => X"-004000e000d00000004000d001f-005-010-0090000-037-00f-011-001-00a",
            INIT_2E => X"0016-004-02e-0310019-007-031-040-0030012-017-01c0047-02700020049",
            INIT_2F => X"0002-004000d0018000800130014-0110004-01a-02e-01b-040-01d0030-027",
            INIT_30 => X"-0100010-02d0006-00c-021-0030035-005-013000f000c00170013001c0011",
            INIT_31 => X"-001002e00020016001b0012-0040016-01e000a0004-026-00d-00e00020012",
            INIT_32 => X"0019-00d000b-017-0090002-00f001b0000-017-00c002d000a-0120008-015",
            INIT_33 => X"-017-0110030000a-0340023-00c-02a0021001d-01300130048004600250053",
            INIT_34 => X"004f00380010-0170021003b000a00200018-01f-02b-0160021-068-035002d",
            INIT_35 => X"-022-005001e0002-01f0014002c-003-020003c001a-008-004-022-016-00e",
            INIT_36 => X"002b-00d0045004e0021-026-007002d0000-01f-0080009-030-02800170034",
            INIT_37 => X"000c00290001-023000a-02a-027-052-01b0024-065-0300017-0270011004f",
            INIT_38 => X"-004-002-007-002000300000008000a-0010002-049-0520013-050-0510017",
            INIT_39 => X"-001-00f-02300280043-024002a00500006-005001d-01a0001-005-00b0014",
            INIT_3A => X"002a-01b002d0030-017002c-006000d006e0045-01d-0070016-017-0130018",
            INIT_3B => X"-01b0009002c-01a-00400050000-020-02c-00f0006-0080027001e00030006",
            INIT_3C => X"-005-0250005-01700020005-01e-020-006-0250027-007-00e00040017-018",
            INIT_3D => X"000b-00e-01d-05b0021-030-0450004-02e-038-017-02e00160007-02a000a",
            INIT_3E => X"000a0009-005-00d000d0016-022-0120008-01f-005-023-01e001e001e0009",
            INIT_3F => X"0007000d0016002b00120012-029-04500640000-03d0033-018-043-030-01a",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY2;


    MEM_IWGHT_18K_LAYER2_ENTITY3 : if N_BRAM = 3 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0029-01a000c0003-021-027-021-00e0007000a000f0036002600130003000a",
            INIT_01 => X"002a-033-084-006-066-05e-00c-047-0310018-00e-01c0040-00f-0290027",
            INIT_02 => X"-010-023-010000b000d-0160019-012-008001b0000-00d002b00340001-002",
            INIT_03 => X"001d00050014000e001c001e000400110009-012-006001f-016001300000010",
            INIT_04 => X"0007001200260000-0040000-012-009-004-00d000f-0180000001c00180007",
            INIT_05 => X"00110027-0160003002a-011000e-00b-037002a0058-03500140053-00d-01d",
            INIT_06 => X"00280006-029-0260015-004-00f000b-003-00e000f0007-02a0033-007-005",
            INIT_07 => X"0009-01a-03d0000-01f-014-0120001-004-007-008001a001800260017-007",
            INIT_08 => X"0007-006-028-0080009-00d0013-0080018-014000a-01a-019-019-00c001f",
            INIT_09 => X"000a000d-002-01400090016-013-009-007000300260008000f00200007-017",
            INIT_0A => X"000400100007-00c0009-00a-001-026-008-067-042-058-076-08c-057-05c",
            INIT_0B => X"-060-034001200210022001000370015002b-005001a0024-01d-00200220000",
            INIT_0C => X"-01c-00a-004-01c00460029002c005f0015000400510029-00f000d0004-008",
            INIT_0D => X"0000001d00060002-01a-012-01e-001-015-004-00d000b0019-003-00a-00f",
            INIT_0E => X"0024001f0017000a000b0028003c-009-003-0030003-031-05f-029-03d-038",
            INIT_0F => X"0016-00b-017-001-013-010-013-007-0090025-02e-01e-01b-02e-060-031",
            INIT_10 => X"-010-037-007-024-028-02100180004-01b0009-016-015-018-01b-011000c",
            INIT_11 => X"0009-016001b001d0010000d001b0002-006-00b00130015000e-004-002-001",
            INIT_12 => X"-01c-01800070002-008-01f-00e-018-00b-0270014-018-018002b0018000c",
            INIT_13 => X"-050-02d-011-04f-029-010-020-012000f-007-027-02a-008-0140003000d",
            INIT_14 => X"-0020006-01000290019-00a000b-00a-00c-015-01c0005000a-00200050017",
            INIT_15 => X"-006000f001e0005-008-004000700140006-013001c-003-022-017-00e-004",
            INIT_16 => X"-017-00a-0140012-005000a-011-01b-00c-01c-0070008-00d-00a00140027",
            INIT_17 => X"00050012-015-00a0012-01000080004-002-001000f0000-00f002a-0300010",
            INIT_18 => X"0031001d001400200008001b00090008-013-00f-009-0020014001e00060006",
            INIT_19 => X"00000001003a-003-01600050003-019001f0014-00400000034002900110003",
            INIT_1A => X"0031000300090021000c-02500090015-01f0002002e-00b000c000000030011",
            INIT_1B => X"000f000d000d-0090002-00a-023001700000015001a0017001e002d0018000a",
            INIT_1C => X"00080001-021-009-015000a0007-00800000004000a-00d0023002d-0130005",
            INIT_1D => X"-032-052000b002e0056001e0006-00d-013-01c-011000400150000-03a000c",
            INIT_1E => X"002a-046-00e00130037001b0022-00d0006-028-00f-029-030-027-04d-01f",
            INIT_1F => X"000c-04f000f0029002900440019-00d0012-021-0160017-00c-01d-01f000b",
            INIT_20 => X"00050013-00f001f-0010002-011-016-0130011001a0028-0020021-01e-02b",
            INIT_21 => X"-01b-02b-018-010-012-01d-029-00b-020-00500110000-01c0033-002-013",
            INIT_22 => X"-007-011-0230017-00e-00e-009-022-017-005-018-008-006-028-02a0012",
            INIT_23 => X"000400080008001e0031000500050031001e00150009-0190003-0160003-053",
            INIT_24 => X"-0520044-03400090036001d003d0000000c0019000c001100150003-01b0018",
            INIT_25 => X"000d-017-0250003000c-041001e-024-02a-029-00a0002-03b-00a-007-01e",
            INIT_26 => X"-0260026-004003400250010004d004d001c-001-0130001-021-0150010-028",
            INIT_27 => X"00250026-00100180024-012000b-014-02400000000-014-003-013-0180016",
            INIT_28 => X"-00f-01e0020000c0007001f-036-002-00c-021-0060000-014-00b000c-00c",
            INIT_29 => X"-044-015000c0010001b002b001100280010006d00310026003b-007-024-01b",
            INIT_2A => X"-01b-00800130028-0050004-00f-010-014-041-00a-00100090017-00e001a",
            INIT_2B => X"-013-0070006000b-025-0200005000e-00d00100006-009001800130035-003",
            INIT_2C => X"000f000a-00f-007-0010002-026-02200080019-01e-014-009-0090006-022",
            INIT_2D => X"-0060006-01b0000000200050011-0060001000b-002001b001d001f00180028",
            INIT_2E => X"0008-0050001-009001d00000014-007-002-00f0010-008-006-009-008-012",
            INIT_2F => X"-00b0023-020-008-036-009002a0017005100600059001c000b0008-025-01a",
            INIT_30 => X"-00b0019-00e-025-008-027-04f0025000d-02c004f00270014000700150013",
            INIT_31 => X"-014-0230003000a-01a0001-012000a0019-01d-01f0008000b-00e-00c-007",
            INIT_32 => X"-028001f-01300020000000c0016001e0004-028-04500140016-027001c-013",
            INIT_33 => X"0000-014-006-0020027002f-00d000f000b-025-01e-00e-03c00060007-008",
            INIT_34 => X"-026-010-002-011-00f001d-012-00200320001002c-002-011000e0002-006",
            INIT_35 => X"-00b0014-02f-024-007000a0008002d000b0018-021000c001300060015000e",
            INIT_36 => X"00100001000200000012-01e0010-01c-02b000a-013-003-00a00120000-02d",
            INIT_37 => X"0025002f002d0071004a00600023-004001f-01b000d000500050015000c0012",
            INIT_38 => X"0007-013-0010001-00e0002-02a-00d-025-025-010-009-01e0024-007-039",
            INIT_39 => X"-030-009-00f-00500060013002a-00e-036-01f000100040004-00c-003001f",
            INIT_3A => X"-033-007-01d0017-005-002-00d-008-0100024000c-00d00150003-0110000",
            INIT_3B => X"-015001c0003-0090024-016-03f-01000090010-01d-00b-012-02300140002",
            INIT_3C => X"0000-001000000000008-0150003001300260015-004000f-01f000e002a-009",
            INIT_3D => X"0003-014-02d-028-0190007-00d-012-00e0014001d0027-03e-00b-004-007",
            INIT_3E => X"-00a-0050023-00d-01b-0020032002d-006-00d0042-017-005001400320000",
            INIT_3F => X"0027-006-029-00e-007-00d-00a-0110019-007-008001d0014000a-003-010",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY3;


    MEM_IWGHT_18K_LAYER2_ENTITY4 : if N_BRAM = 4 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"-011-014001e00090014000b002a001c001c00270013-003002c0006000c-02a",
            INIT_01 => X"-02c000d000e-0020011001400520034004100210027002c0038001f002b003d",
            INIT_02 => X"000e0002-004-022002d-004-02000340050-01d0005-009-019-00d000c0032",
            INIT_03 => X"-001-009000f002f000f001d0002-023-007-02a-02a-0460006000f-00c-004",
            INIT_04 => X"-0190002000b0026000a001c001e0003002c0024-010-0020002-00c-01c-020",
            INIT_05 => X"00040008001e0023-026-02100000000-00d-0030025-00d-01a0002-010-01b",
            INIT_06 => X"-008-02a-017000f-0210002-0230009-00d0018-024-016-02e00050007-038",
            INIT_07 => X"-01d-009-01a00070004-00a-032-00e002900010005001c0015001e-003001b",
            INIT_08 => X"0001-020000100170042003d001a-03b-00d000a-05d-0380010-01f000d-011",
            INIT_09 => X"0043-02f-00a000a-015-03e-015-0010026-01e-007001c0009-00900010022",
            INIT_0A => X"000c0002-02d-01f001e-042-01d-0210020-0070004-00b0005-00d-023-00d",
            INIT_0B => X"0011001c-018-00f0023-00f001f-029-0200018-016-00b00100001002a0023",
            INIT_0C => X"-01d-0030016000b00110006-008-009000a-034-00c001e-01000340024003a",
            INIT_0D => X"-008-0080001-02a-03b0001-019-023-00e0029004b002500320020-013-00b",
            INIT_0E => X"-005-004-01b-020001e0012-016-012-00b0000-002-0140032-004-0130028",
            INIT_0F => X"0014001d0005-021-00a000c-01a00040017000c-01600110017005800030015",
            INIT_10 => X"005c-0190019001c-030-040-067000d-019-01d-00a-0020015-00a0005-008",
            INIT_11 => X"000d-00c00000002000a000600290000000f0013-00e-00600200004-002-002",
            INIT_12 => X"-00c00090009000200130017000c000b000d002a001b0036-00c00000010000e",
            INIT_13 => X"0021001d0039000a002500420019-001001500180017-024-01f0013-030-033",
            INIT_14 => X"-01f-041-047-03b001b0021002c001000430040-018-0060005-00a000c000f",
            INIT_15 => X"-02500150000001e-00a-006-0030018003200020018-005-002-01a-0160000",
            INIT_16 => X"-001-016001300070000-018000a0018000d-030-00b001e000a-0100028-005",
            INIT_17 => X"00000005001a0000-0040003-015-011-010000c0015-010000c-0060015001b",
            INIT_18 => X"001b0017001a001f00130027-039000d-00e0003002d-01a-001000e002c0000",
            INIT_19 => X"-019000c-01f-01f-02f-009000d0006000f00190009-0230015001100170015",
            INIT_1A => X"0034-036-016-00d-0010011-007000c002200330005000d0009-00c0000-017",
            INIT_1B => X"00020034-01b-00c0006002f-001002200120025001b001c-00f001a-00a-02a",
            INIT_1C => X"0001-016-065-034-034-039-010-034-02d0015-02a0000-005000e-008-005",
            INIT_1D => X"0006000b0008-00e-0120000-026-026-02a-00f-014000c00080016001b-008",
            INIT_1E => X"-01b-013-01b001d-007000e001b00240035-003-015001f0005-022-015-025",
            INIT_1F => X"0012000e-024000d-01900100020-01f-00d-03e-02b0007-017-033001d-010",
            INIT_20 => X"0019-008-012-035001b000d-003-015000e-00a00190025-0070019-00c-019",
            INIT_21 => X"-00f000a-020-00b-00e-002-006-01f-00e0002-026-02b-026-0250010-040",
            INIT_22 => X"-045-016-023-02c-03c-01a-019-00d-00f-00e-02300030001-015-017-01b",
            INIT_23 => X"-03b-027-025-02f-00f000f-012002500390043000e00000000-014-024-02c",
            INIT_24 => X"-010000d0016-00f-00700150005-001-005-021-01e-017-00600010027001f",
            INIT_25 => X"00050014000e-039-01f-03a-04d-05a-01c-057-057001b-04a-04d-00e-03b",
            INIT_26 => X"-0590019001e-06c-026-058-03a-060-03b-065-03c-00c-058-03f-02c-016",
            INIT_27 => X"-026-0100015-005000b0010-00c-00e-025-00d000b-01f000a0000-0360029",
            INIT_28 => X"001d-00f00310026000c0027000a-025000100000022-01a00170015-0040017",
            INIT_29 => X"000a-017-0140036-002-02c0027-01000210047-00a00080016-00e0007-001",
            INIT_2A => X"-003-0080001-07a-064-043-02f-086-0420015-00b-018-01e-00e-02f0003",
            INIT_2B => X"0000-00c-00e-002-00b00070000-018-002-00e-0140017-01c0000-053-034",
            INIT_2C => X"-01d-02c-052-021-030-01d-02a-027-015-00b00110016002f000800130017",
            INIT_2D => X"00330026001000120002000c0002000c-022-00f-012-028-00c-01c-00a-006",
            INIT_2E => X"-017-0050011001c0010-012-028-026-050-046-040-0050034001a002e0024",
            INIT_2F => X"001e001d002d-006-019-015-010-0070015-0110000-006-004-01000000005",
            INIT_30 => X"-004-0080017000c0028000000060000-0120013000c002a000b0004001a0005",
            INIT_31 => X"0029-00c0011-0050003-009001e-00b0006001a0033004f006d002f007a0054",
            INIT_32 => X"0064002a0013-00500320003-00c000d0010-02b-008-0090023-013-007001e",
            INIT_33 => X"0003-001003a-008-00e0013001b000d-00f-003000b-00d-008-045-00a-04f",
            INIT_34 => X"-05d-047-016-02e-051001800150006-023-01800000015-008-00100270020",
            INIT_35 => X"-004001200210001-00b-00a-02d-021-00f0006-00b-012001a001400150037",
            INIT_36 => X"0000-007-007-002-006000f000a-0100006-04a-075-067-054-07a-031-00a",
            INIT_37 => X"-036-02a-02400470042000200070014-018-018-029-00500160044-00f0009",
            INIT_38 => X"-01d0001-020-031003000300021001c0006004d0011-002000f0019003e001e",
            INIT_39 => X"001f001f001f000700180013-024-029-03e-010-029-01b-02f-0150003-006",
            INIT_3A => X"001900100016001e0005002400190009-006-01c-008-023-035-011-027-02f",
            INIT_3B => X"0000-05e-01c-011-03f-0050004-01b0009-021-019-044-035-005-033-023",
            INIT_3C => X"000d-021-01a-037-0300013-015-01d-01f0012-02a-0230000-00c0011-00b",
            INIT_3D => X"0001000f-00700110018-031-02d-02c-00c-02e-01f-037-0120006-005-015",
            INIT_3E => X"0012-00d-002-015-00d0000-02a-03d-019-00a-02a000a0006-00c00390024",
            INIT_3F => X"-02b-016-059-05a-03b-042-039-041-049-022-041-0240001-011-01d001c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY4;


    MEM_IWGHT_18K_LAYER2_ENTITY5 : if N_BRAM = 5 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000-01a001e000e0027-018-0170007-0560000-0110008-0020006000f0027",
            INIT_01 => X"0022-0070017002f-015000f0020-01100100003-00700160019-008-004-001",
            INIT_02 => X"000a0008000c0001001a0016-03e-026-03b-034-00b-01c000c-015-0030018",
            INIT_03 => X"000a001100190015-011-00a000c-006-013002b-001-049-00e0005-05c-022",
            INIT_04 => X"00060010002a0025-001-00e0005-00b-01a0005-019-005000f-010-00d-006",
            INIT_05 => X"-00d0009-008-015-038-020-01b0008-00a-04200000004001c001300370008",
            INIT_06 => X"0000-00e-01d-0530012-0060005-027-02a-00e-021-01f0002-03500190032",
            INIT_07 => X"000c-008001f0011-008001a00170000-015000000120016-003002a-0030004",
            INIT_08 => X"-012-0120014000d0003000a0000-01700170016000f003e0005001c000a-00b",
            INIT_09 => X"00000003-01700000001-004001b000e-00c000a001c-032-01d000f00320006",
            INIT_0A => X"-019002f000b0000-012-0040002000b-00500080022-0040007-00900180003",
            INIT_0B => X"-013-0120009-011000400220000001b000f000300010018-012-001000f-016",
            INIT_0C => X"00000025-01b00170031004800180050001e-023-039001b0034-02400280001",
            INIT_0D => X"-00900110022-00e-013-002-028-057-01e-030001b00000011-007000d-01b",
            INIT_0E => X"-01a0009-00e000d-010002c-02d-036-038-03c-02c-015002300260024-019",
            INIT_0F => X"-01f0008-007-00700130014002b0020-009001b00190011-0090043-00e-023",
            INIT_10 => X"-022-014-01b-021002c003d003e004a00460021-01c-0080000-042-03e-03a",
            INIT_11 => X"-039-02f-04c-014001c000c-02f-011-02100210025000f-01e-002-00a-04a",
            INIT_12 => X"-0060003-01f-022-02d00020031-008-046-017-033000d-001-00b-017-006",
            INIT_13 => X"-016-010-01b001e0000000a000e00130011002e-005-01300040021001e0016",
            INIT_14 => X"-00b-00f0013000e-02400030052002d001a00000000-032-00a-00f-00a-034",
            INIT_15 => X"-054-030-017-01e-008-01600120012-028-05b-051-00c-011-01f-00b-02c",
            INIT_16 => X"-044-04e-029-009000e0034000c002a-009-003-002000e-004-030-00b-025",
            INIT_17 => X"-04e-015000f000f0000000f000000120014-01d-00e0037-010-00f-036001d",
            INIT_18 => X"-006-033000f0000-03400180007-00e-0020015003b0001-00e003c-02a-018",
            INIT_19 => X"-004001b00230022001b001e000b00100029001c-01d0000000b-034-012-018",
            INIT_1A => X"000c0006001a000e-00c-00400150002-0070033004b002a00430040003e0042",
            INIT_1B => X"0038003a-010-046-00b-044-076-044-042-06c-026-022-021-01d-022-040",
            INIT_1C => X"-011-05e-01c-01b-009-01e-01a-03c-045000c-07a-042-01f-006-017-027",
            INIT_1D => X"000c0000-0010037002f0042-00200420027-009-015000d-024-020-011000e",
            INIT_1E => X"0001-005001000210005002700150008000a00150022001e-00f000a000c0010",
            INIT_1F => X"00380014000b001b-02500050002-035-025000300210010000d0022-00b0029",
            INIT_20 => X"-012-0030017-008-010-028-010-009-019-01c001e000a000b-017-015-011",
            INIT_21 => X"-00d-00f-001000c-00e001300210016001400310032-01300070009000c-017",
            INIT_22 => X"-002-0130000-005001e00100006-01c-004-017-02600000003-00600100009",
            INIT_23 => X"0033005d005e-0070048003a002000130025000e001e-003000a00050000-009",
            INIT_24 => X"000e000d-0160000-018-01d000d-01a-018-008-01c001d000f001f0001-00a",
            INIT_25 => X"0008001400140019-02e-00b-016000f0018-019001a00020007001100190003",
            INIT_26 => X"-004000f-01a000b00070011001c0012002900030011001c-00c-00a00030003",
            INIT_27 => X"-00f0004-007000d0006-02d0004-00d-045-022-009-049-06c-03d-069-090",
            INIT_28 => X"-040000a002100240010000f0023000400110019000300130021-028002d0009",
            INIT_29 => X"-01a000a0006003200180009000a-005-01300250010-014-00a-02c-00c-02e",
            INIT_2A => X"-02b0009-038-0190008-011-017000100090008-0160004-016-021-00f-018",
            INIT_2B => X"-01a001800120003000d00150000-010000f-0040003000e0003-00500000009",
            INIT_2C => X"-015-0160000-016000b00030003000a000a00110004-004-011-039-01e-02c",
            INIT_2D => X"-028-022-03e-03f-034-055-066-013000b-00500150009-009-02a00290003",
            INIT_2E => X"-01b00360035-002-06a-03f-04d-04e-02a-017000500240005001a00420033",
            INIT_2F => X"000000160027-031-00f-02a-028-017-041-05d-022-01b0009-015002c001b",
            INIT_30 => X"000e000f-0090000001e001c000a0034-006-003-007-026-036-00a-035-019",
            INIT_31 => X"-01200100014-0040001-0130007-008000a-012-00e0007-00b-028-00d-013",
            INIT_32 => X"-00d002900240014001d00070008000c-00e-006001e-03a-004000300180002",
            INIT_33 => X"-007000500000001-026-025-02a-02d0003-007-00e004d0030003b000e0036",
            INIT_34 => X"0018-019000e-014-03c-013-01d-0170001-00f-003-003-015-028-0130000",
            INIT_35 => X"00040007-02b000b00100034001700360016-00c-00b0006001b-00f-0010008",
            INIT_36 => X"0014000b-02a-007-02e-0100005-001002a000a-01c-005000c001b-0130015",
            INIT_37 => X"-00a-01100050013000c000d-00c001f001c-00a-0090004-01500310010-001",
            INIT_38 => X"-006000e-019-02e-0120014-003001a000c000200150028-0150006-0090003",
            INIT_39 => X"000f00120006-00a-014000d001a0011-03c001d002d-03100340050-03a000e",
            INIT_3A => X"008d-037-033-035-01e0000-01a002a003a002e0001-00d0004-00c-011-00d",
            INIT_3B => X"003100200001-01c0008000a-01b-00f-007-04100150016-010-00c-027002a",
            INIT_3C => X"0009-01900370036-0150011002e0016-0160006000d-028-017001d0022000e",
            INIT_3D => X"-00d0025001e-003001b0010-00800250017002800360016-027001c0022-006",
            INIT_3E => X"-0020008000c0006000a001a00040017-00b-0090004-00d0003000600180005",
            INIT_3F => X"0030-013000f-006-00d-010-016-0170015-027-005-009-01e-02f0006-016",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY5;


    MEM_IWGHT_18K_LAYER2_ENTITY6 : if N_BRAM = 6 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"002c0002001a004d-01e-041-006-022-02e-001-002-05d-056-00c-014000f",
            INIT_01 => X"0000-00d-005-014-01e-00f00210025-00f-05e-058-02a-03b-03b0000-014",
            INIT_02 => X"001b0007-036-010000a-020000e002e00220015001100040006-016-005-00d",
            INIT_03 => X"-017000a-01b-03700160006-02b0011-00e-054000a0016001f001d0022-01c",
            INIT_04 => X"-016-014-02b0000-00a-00700070008-0110022000a0009-01f-017-01c-028",
            INIT_05 => X"-0070001-01f0002000600180023-00b-003001d000b00160006000e000b0005",
            INIT_06 => X"000100060015-012-03a-055-02f-008-003-0130028-004-00e-00b0003-00c",
            INIT_07 => X"0036002600210047003b0002000c000d0002-009000f000000050021-008-007",
            INIT_08 => X"-01e000600230027-005-0210026-00b-04b-00d-039000e000d0014-00f-013",
            INIT_09 => X"0007-045-02f-0010033002f001c-01f-0310015-03e-02200020033001d0021",
            INIT_0A => X"000e-008000d-020-0350023-014-027-00100060007-02700100009-001-003",
            INIT_0B => X"00240020000c0010000f-063-03d-0260036-018-0090028-04f00060024-03e",
            INIT_0C => X"-0280004000300050009-00c000f-0120001001900220026-00f000f002a-00e",
            INIT_0D => X"000b0024-034-019-01c-030-005-00a-013-016-02c-0070006-028-017-01f",
            INIT_0E => X"-0110012000700030034-012-005-00e-017-014-008000c-022-018001d000b",
            INIT_0F => X"0002-027-001-004-053-02c0027000a0013-0200022002c-00d0029001d-005",
            INIT_10 => X"0001001800040013-00a000d0016000a00010000-006001b0013002800350010",
            INIT_11 => X"0031-011003b0021-00c001f002d0012-0270001-0070013-008-011-037-01d",
            INIT_12 => X"-0130004-02a-00f0028000600130000002300040007000d-001-01a-02c-008",
            INIT_13 => X"-01e-042-027-00d-047-02b-01c-00a0009-008001f000c-01e00110009-003",
            INIT_14 => X"-00a000000040020000e-01c001f00290011-00a-00a-007-013000a-020-00d",
            INIT_15 => X"000e-002-004-001002d0006-015-002-00a-02900270020001a001900200010",
            INIT_16 => X"-006-009001e000500030018-03c-0020000-009-02c-0200006001c000e-01c",
            INIT_17 => X"-008-00a0006-00a-028-013-027-019-018001d000c-0030004-019-010-02e",
            INIT_18 => X"-010-018-043-017-00e-032-00c00110008000a0025-023-0100032-003-028",
            INIT_19 => X"-00d00300010-0350017-032-02600180001001d002c-008-0020012002f-028",
            INIT_1A => X"0017-0170012-01a001e0036002b-0070039-027-01f00120010000b-003-02f",
            INIT_1B => X"0000-004-01e-00600080010000e0012-019-00a-015-022-01a000b0011000a",
            INIT_1C => X"-00c-02c000d0005-017-00c-022-00f0015-006-008000d0008-00d-00c0020",
            INIT_1D => X"0000000c-002-010000d-00f-00500330011-02a-00900090004-008001a0001",
            INIT_1E => X"000300100022000c0011003c0029-0290029001d-00600020000000f00080000",
            INIT_1F => X"00450005-02a0003-00a001d-0380006-019-00f-004-02f-00e-0140001-02f",
            INIT_20 => X"-042-024-019-057-02b-008-01b0000-01f-033-03f0003002b-02800040000",
            INIT_21 => X"-006-009-0030001-012000200090005000e00050020-0050019001c-00f-020",
            INIT_22 => X"-00a-00a0010000a-002-00e000a-010-00b-022-037-0250025-015-03c0028",
            INIT_23 => X"0004-014-01d-039-02a-01a-010000d-025000a0029-00c-048-028-01a-005",
            INIT_24 => X"0028-018-0100033-016-049-038-012-0160010-00e0054004d-026-005-012",
            INIT_25 => X"-01e000e-01a00290029002f001b0017-001001e0031001a-027-039-03e0028",
            INIT_26 => X"00180013003f003a0018-010-0130011-031-00b-014-00f-006-012002e0049",
            INIT_27 => X"00100018001a002400280020003a-038-029-00b-031-023-027-00700070003",
            INIT_28 => X"000c00210000-024-024-00c00000028000a-01c000c00350009-005-0130006",
            INIT_29 => X"0015-008-007-00900120042000e0025006e00280019-012-03d-010-05e-01b",
            INIT_2A => X"-0440000003c00090023003f000d00050014-006-013-01b-00b000d-025-013",
            INIT_2B => X"002c0030003100510030004600150035000e0005-003-00e-0010000-004-024",
            INIT_2C => X"-033-012-00f0004000d-01f-0120001-0290006-02b-02e-014-0400000-001",
            INIT_2D => X"-021001900350002-024-020-0340017001a-009003b003b-007-015-007-042",
            INIT_2E => X"000f-006-0220042003500030024000700120013-0050001-024-035-012-035",
            INIT_2F => X"-02b-0140001002d-013000a000c-031-04700340000-02800400018-0340018",
            INIT_30 => X"004b0023-037-01e004500050004-004-01b-01f-008002d001a-00d-006003c",
            INIT_31 => X"-01f-042-006001e0044002d00140023001c-0110008-00f-011-02b000a000d",
            INIT_32 => X"-0260013-00f-003003a000c00430048000d001d002f-043-029-02b0002-018",
            INIT_33 => X"-0140022002a0010002a000d-00900030018002c-003-0190013-016-0110001",
            INIT_34 => X"0000-00600000008000a-00e-00900070012-0130013-00c0002-00a-00b-00b",
            INIT_35 => X"-00d-006-0040007000a-007-00d-0100010-007-0050000000e-00b0000-001",
            INIT_36 => X"00020007-00c000b-003-013-01a0000-0040000-012-001-007000500000003",
            INIT_37 => X"-009-00c-00c-015-004-00f-002-00a0010-003-014000000000004-00a-00d",
            INIT_38 => X"-00c000d0001-017000400100003-006-00f0009-011-003-010-005-0040000",
            INIT_39 => X"-005000a0000000a000a000300110003-00a-00b-0030013-0050002-0020004",
            INIT_3A => X"0017-00f-003-00700060007000c-00b-00d000000000007000f-0140002-009",
            INIT_3B => X"000300010000000d-0030006-015000b-0110002-010-00b-009-005-003000e",
            INIT_3C => X"00000000-007000b-00f-014-00c00030000-016-0160006-001-0140011-016",
            INIT_3D => X"00100011-012-010000c000f-00b0005000e-015-008-00a0000-00b00070004",
            INIT_3E => X"-00f000a001500110002-00d0007-005-006-007-0100003000e-013-00d000c",
            INIT_3F => X"-00d000e-0010002-007-001-0180004000d0002-00b0003-0030006000b-00c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY6;


    MEM_IWGHT_18K_LAYER2_ENTITY7 : if N_BRAM = 7 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"-017-00c000a0009-015000a-010000d-004-0060005-017-0120012-007-003",
            INIT_01 => X"-00f-00c-00e-0100004-00d-013-016-010-008-00a0003-002000a0005-002",
            INIT_02 => X"-018-00c-002-0180004-00d-0070003-0020000-002-00a000b0005000f-00a",
            INIT_03 => X"00110007000d-00a0009-00b-011-005-006-0150004-012-00a00000004-008",
            INIT_04 => X"0001-00b-00a0003-00b0000-008-00e-015-007-00400000007-014-0160009",
            INIT_05 => X"-00d-0120000-007-009-005000300060008-001-007-005-012-00d-00c-017",
            INIT_06 => X"-008-006-002-0080008-0190006-017-012-00300150002-003-017-02b-006",
            INIT_07 => X"-01c-00d-023-004-021-0040014001f002e00430028001d00480040003a0018",
            INIT_08 => X"001e000b0002-01a-007-00e-0260030000b-010002c00310033-005-020-009",
            INIT_09 => X"-020-003-012-0170017-01f-016000a-002-002-029-009-00c-00a-0170005",
            INIT_0A => X"001800040013002200260020002700000016001c0019001b-00c0001000d-017",
            INIT_0B => X"0006-04e-066-018-025-03d-01b0022000000240008002f0002-00e-025-011",
            INIT_0C => X"000c-018-020-037-03f-01a-02e-03c-02b-012-041-0310001-032-01b-004",
            INIT_0D => X"0003-00b001300210010-013000c000200020005-0020017000d002e0016-012",
            INIT_0E => X"-00a0010-00e00150001-007-011-016-02f-00e-023-00e-00700070009001e",
            INIT_0F => X"-031-03a-011-051-052-023-01b-020-033-039-009-0010000-03d0009-003",
            INIT_10 => X"-00800070001001b-00c-048-04f-04f-046-05d-03900280009-0140026002c",
            INIT_11 => X"000600250013001f00150001-00c0013-015-00f-022-014-00b0027000b-014",
            INIT_12 => X"002b001300040009-0060009-02b-015-00a-00e-02f00060016000a001c-002",
            INIT_13 => X"00070014-00d-0010004-0070007-001002000300019002c0029-0030000-005",
            INIT_14 => X"000b002400420020002300070024002300010017-049-043-009-039-0040007",
            INIT_15 => X"-003000b00200017-01e-005-0040028001f000a000600130041002e00240024",
            INIT_16 => X"00140014000b-012-010-024-036000c0004-0260003000d00080001000f0010",
            INIT_17 => X"00130028000b001d-00b-011-00e-013-0480002-042-0240010000b00140022",
            INIT_18 => X"0000-00700150007-00a-009-0030006-0170035001300280003-00700230003",
            INIT_19 => X"00000002002a-004003c002d002e0015002c00300016-038-00f-017-009-021",
            INIT_1A => X"-0120012000c-031-0110019-0340037003500140014001d0002-025-023-028",
            INIT_1B => X"000e00270023000e001e0007004d00380033000e001c0020-00b-039-03d001c",
            INIT_1C => X"00330016-017-009-02d-018-037-005002e-00800070001002c002a0012001b",
            INIT_1D => X"0017002c0011-002002b-021-01900260000-0110001-0150006-02300000033",
            INIT_1E => X"-017-00e-00d-00a002d000e-01e001f001e0007-024-020001b00040004000a",
            INIT_1F => X"0011-0210006-008-01d0030001200350002-01e-023-00e-01b-017000c000d",
            INIT_20 => X"-0130010003f00210010003e0018000600080003001d-006-01b-00a-0190001",
            INIT_21 => X"-01c-0050013000b-0110029-02f-02a-007001a001000280005-00c0027-00a",
            INIT_22 => X"-022-017-00a0006-00b00180004000900240007-00f000e-003-00c00080035",
            INIT_23 => X"0000-00e0008-00a-003-00e-00c000a0003-022-00a000e000600000001-017",
            INIT_24 => X"000f00130010001c000b000f004a002a00280015000b00170028-011-009-01d",
            INIT_25 => X"-00e-0290005000a-00b000d-005-0200001-03100000012-008003f-0240001",
            INIT_26 => X"0022-002000b-006-011-019-024-044-039-04b0013-003-0010011-01f0001",
            INIT_27 => X"0019-028-00200480013001e001900030011-002-00c-00d-00f-00a-00c0001",
            INIT_28 => X"0004001f001a003a-00f002000250019001b0002-008-005-0250013-01f-006",
            INIT_29 => X"-023-009-00b-00f-0170001-015001e0010-005-00b-029-00a00190001-013",
            INIT_2A => X"000a-012-0150014000300080015000a0000-019-010-0110001-016-0020008",
            INIT_2B => X"000200000002000a0005-013-00b0008-003-015-013-018000b-00c000d0004",
            INIT_2C => X"-00d00110002-0030002-003-00a00070015-00a000c000a0002-002-008-004",
            INIT_2D => X"-002000b-01a0005-0010003000b0007-0010000-00c-00c-00f-01b00060007",
            INIT_2E => X"-0150001-004-016-008-005-00a0001-00f00090005-011-010-019-00b-00e",
            INIT_2F => X"-013000c-00f-01500090000-019-018-01b-007-019000500090001000a-012",
            INIT_30 => X"-003-007-012000a-007-003000f-00b-00700000000-003-014-015-004-00f",
            INIT_31 => X"-01b000b0009-006-001-0110009-00c-00b0002-002-0040000-01a-01a-00b",
            INIT_32 => X"-01700010000-00f000400040002-01000040007000f000f-00f-00f-0070001",
            INIT_33 => X"-004-00d-00b0000000b0000-00f0007-0040003000b0001-0150002-007-016",
            INIT_34 => X"0009-012-00b000d0008-01400020000-014000f000f0007-004-00e-001-00d",
            INIT_35 => X"-00a-002-01d-00a-00e-007000b-014-008-013-01d-0100000-015000e0005",
            INIT_36 => X"0007000d-00a-012000e-0140000000d-0010004-011-008-00c-0130007-010",
            INIT_37 => X"00040000-010-016-0070007-012000500000002-019-00e0004-01c0007000b",
            INIT_38 => X"-013-01f00000003-01a-021-022-00c-020-011-00800060013-00a-00d-003",
            INIT_39 => X"-00a0000-010-017-00d0001-006-008-015-0140005-019-00c0007-01a-003",
            INIT_3A => X"0007-00e00130005-01d-001-014000b0010-00c0005-00d-01b-004-005-019",
            INIT_3B => X"0000-00b-00e-002-0150006-003-00c-00c-003-007-0140006000f-0180005",
            INIT_3C => X"-00a-0030012-0130014-002-0030006-0110004-003-01500090003000a0003",
            INIT_3D => X"-0010000-013-009-00300050004001100010005-0170000-015-014-011-009",
            INIT_3E => X"-0140009-009-00e-012-00d0003-00400090006-010-00c-012-017-01c0002",
            INIT_3F => X"-01c-011-01e0009000b-00c-00c-018-002-00b00020002-006-014-002-016",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY7;


    MEM_IWGHT_18K_LAYER2_ENTITY8 : if N_BRAM = 8 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"-00d-0070005-00a-00f-00b-019-0140007-011-01900000000-0020000000b",
            INIT_01 => X"00030006-010-00a-013-002000800080008000500000005-004-004-01d0005",
            INIT_02 => X"-00b-0090000-015-007000b-016-017000e-004-01700030008000f-0060005",
            INIT_03 => X"00090008000f000b000400020004000c-017-003-014000a-00a-001-017000a",
            INIT_04 => X"-002-00e0006000000080006-015-006000e-00a0000-0080001-00d-009-004",
            INIT_05 => X"000e0012000c-00a-002-00f0000-0130004-0080006-00c-003-016-0130008",
            INIT_06 => X"-004-009-0040005000a-00a0005-0050013-011-006000d-016-007-004-007",
            INIT_07 => X"-00f-017000a-01b0002-014000a-001-010-00b0003-00e-0110002-00c0007",
            INIT_08 => X"-0070005-00e-014-015-00e-011-005-0140000-002-00a-00f0000-0130006",
            INIT_09 => X"0005000b0004-001-006-019-007-006-00c0009000a-00a000f-01a-006-015",
            INIT_0A => X"000c-015-00e0003-015-017-008-0120004-00d-007000f0000-010-016-00b",
            INIT_0B => X"-008-01c-004-01700050010-014-016-00f-006-00b-012-016-0050007-00b",
            INIT_0C => X"-0110009-00b-007-006-012-01b-00b-01500030002000e-00f0003-014-006",
            INIT_0D => X"-0060005-00b0000-006-00d-012-0120006-001-002-001-007000d-012-009",
            INIT_0E => X"000000080011-0170008-009-006-01300000002002d001e-024-012-00a0016",
            INIT_0F => X"000c00000022002e000500320026-00c00350031-007-003-017-02c-00e-037",
            INIT_10 => X"-0570012-059-04d001e-005-027003e000b-0040038000a000a000b000b-00e",
            INIT_11 => X"001600290017-017-018-01e002a0022000f-0060003-016-01c-014-049-01f",
            INIT_12 => X"-0010018-0210010-00d003a0015002d0035001a-00e0007-01f-0100003000f",
            INIT_13 => X"000e000d-02b0022-017-00400260016-008002a0004002e0001-02d-042-01c",
            INIT_14 => X"0013-009000c-0050026000e0018-020-00b0012-03700060001-016-023-003",
            INIT_15 => X"00070018001500080013-02400000013-02a-0010006-0060015-00b0038000c",
            INIT_16 => X"0004-0010018-002-004-00d-019-01400030015-01c-00f002a-02f00050020",
            INIT_17 => X"-03a-00e0014-043-02e-027-00c000e-035-002000100230002-017001a0000",
            INIT_18 => X"000c0005-03a-0090012000a-004003f-032-024-01b0016002e001a001d0009",
            INIT_19 => X"000b-007000d-00f-01d001b002a-01000000013-013001c00190031002d000a",
            INIT_1A => X"0005000d0003-014000e-00900180026000a0017-001-003000c001c-0040034",
            INIT_1B => X"0014-01a00060008-004-011-00c-0120016002d001e-017-025-00c-056-01c",
            INIT_1C => X"-02d-00e00030013-002000d-0150005-008-01d-00a-01a0018-00700080035",
            INIT_1D => X"-007-0010019001f001d-00f00170010000d-017001d-013-008-008-051-008",
            INIT_1E => X"-010-033-026-031-041-00800060000-015000d002b0009-001-011-0310003",
            INIT_1F => X"-007-0180000-02600150008000c0001-029001c000e-00d0017-01f00010007",
            INIT_20 => X"000c-002-0070007000d-011000c-00c000e0002-01d-01c-024-002-013-01f",
            INIT_21 => X"000a-010-0110002-021-018-009-013000d-012-0070004-017-003-0070009",
            INIT_22 => X"-009-013-02c-015-01c-00c-010-00b000c-006-00200030000-013000f-007",
            INIT_23 => X"00010004-00c00000001-017-01300020003-01b-005-012-0150000-00e-009",
            INIT_24 => X"0002-010-0150006-00c-0170007-003-00a0000000a-015-003-014-0170008",
            INIT_25 => X"-00f00090003-00e0007-008-018000d-0010016-00b-00b000d-002-00f-00d",
            INIT_26 => X"-016-0180004000000120013-017-008-01a-003-01700050006000f-016-00a",
            INIT_27 => X"-01c-013-002-002-00f0005-01c-00f0002-01800000001-009000a000b0011",
            INIT_28 => X"-012-017-00d-015-00c-01b-003-012-0070003-013-009-007000c0000-008",
            INIT_29 => X"00160010-005-009-002000c000800200000-0030019001400110000-0030001",
            INIT_2A => X"-00a00040005-00b0011-003-007-006-00a00020000-0180000-015-00f-01a",
            INIT_2B => X"-001-018-0090002-020-014-011-011-020-00c0000-014-01d-00b-0200000",
            INIT_2C => X"-009-015-00e-00300020008-020-01a-009000f-007000c-0030020-00d000b",
            INIT_2D => X"-00600120009000000000006-0130008-00f-00c-024-017-018-01a0000000c",
            INIT_2E => X"-025000b-004-027-01a-010-016-015-013-013-00d-00600110012000f-004",
            INIT_2F => X"-01b000e-01a00040008-010-008-01d-006-008-002-010-0180002-00c-009",
            INIT_30 => X"-00600010003-014-00b-00a0000-00f-016-0010009-016-00f-010000a0007",
            INIT_31 => X"-010-0150008-006-00e-007-002-01d-006-007000e-004-007-015-017-001",
            INIT_32 => X"0019001a-01200040007000e0018001a0005001c003c0042004a0062003a0057",
            INIT_33 => X"0006-03a0000-011-009-040-04a-052-07d-048-08c-01b-00b0012-01b-00c",
            INIT_34 => X"001c001b000f0063-0030006-003-024-044-03c-015-09d-042001a0018-006",
            INIT_35 => X"0004-020-013002a00340054-00a000a-00c0012000800000000-01b00000009",
            INIT_36 => X"0011-006-004-00c00060016002d00070016001400300019003a0014002c0009",
            INIT_37 => X"-045-01b-00f-03d-00b-020-0500007-00b-00f0025002400020047002a-001",
            INIT_38 => X"0023-062-092-003-00b-04b-037-07c-035-002-03f-021-023-012000e0004",
            INIT_39 => X"-013-007001d00310065000f0023-0240031001f-007-003-005-0070012-02a",
            INIT_3A => X"-029-010-01c-058000a001f0031-004-01f-02a0014-022-019000300160022",
            INIT_3B => X"000a00490014002c0007-013-00a0002-0160028000f000b0022002100170001",
            INIT_3C => X"-00400150002-026000e-01f0016-018-00a0018-005001b000e0015-0070002",
            INIT_3D => X"0002000900130013000e-007-003-024-016-00a-008-00a0001001d0000-003",
            INIT_3E => X"-00f0000000a-008-0050009-018000c000f-003000f-012-00d000900000021",
            INIT_3F => X"0001-00d001e-01a-01c-015-033-039-01a-048-001-048-02a-065-00b-04b",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY8;


    MEM_IWGHT_18K_LAYER2_ENTITY9 : if N_BRAM = 9 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"-05e002f002400320020002a0007000c-00c-017002e-007-014-006-005-022",
            INIT_01 => X"-009-001000f-00d-002-016000e-008-010000c000f000e-010-030001d-01c",
            INIT_02 => X"-00d-006003b0019000e-020-02e-02d-045-040-0310013000b0014-00f000f",
            INIT_03 => X"0001-007-01a00170009000b001a000e-01b-00a0005-001-002-003001a001b",
            INIT_04 => X"-004001800140004-0040008000e0010000200120021-0030017-009-011-011",
            INIT_05 => X"-030000c-007-013-034-012-02e-03c0003-02b-035001a00000007002f0019",
            INIT_06 => X"002c003b0021-010-00d-06a-020-01b-06c-031-027-016-01a-036-00e-03c",
            INIT_07 => X"-0170009-00b-021004000310016000000130009-012001d-01e-013-012-025",
            INIT_08 => X"-02d0005-00a00130029000f-004001f004d0032000f004d0005-016-007-001",
            INIT_09 => X"-00a0002-016-00b000a-00c-026-017-00a-01d00250021-0010024-029-020",
            INIT_0A => X"-00b0000-01f0000-015-014-002001d0002-00e-005-002-00d-021-005-00d",
            INIT_0B => X"00160029001500180017-022-019-0220015000500370022-00700010011-011",
            INIT_0C => X"-028-01c-00a000b-00c001200080001-026-020-017001900190001000d0012",
            INIT_0D => X"005f00390026002e00280026-00c000600240009000b00110012-00400260008",
            INIT_0E => X"-015-018-00a-030-04c-014-008-010-016-01200190000-012-01b000e-01f",
            INIT_0F => X"-003-01b0022002e-019-019-028-041-01a-018-028001c002a-00a-011-022",
            INIT_10 => X"-03f-024-028-00800400042-002-016-02f-00e-0120004-02d-016-0090040",
            INIT_11 => X"0019000a0017-01b-003-002-00a-00a-006-025-041004c-002-02e0000001e",
            INIT_12 => X"00170005-01b-00f-010000d000800010005000a-001000e0013002200050005",
            INIT_13 => X"0007-008-00d-023-028-033-006-0120009-015-00c00040006001900210030",
            INIT_14 => X"0008000f001f0001-022-00d-004-00a-00c000d-01a-00a-0190012-025-012",
            INIT_15 => X"-02c-050-01b-00c-00c000c0018-01d00020017-0050011002f0018-0070012",
            INIT_16 => X"-0090001-013-021-00a000a-01d-018-018001a-00a-015-065-066-047-088",
            INIT_17 => X"-079-03a00180019-016-0200006-0040026001b000e0002-04d-024000a-03f",
            INIT_18 => X"-0340011-017-02a000a-012000000270014-011002b002c000a00290022-001",
            INIT_19 => X"00390027-00a000c0017-00a-0110008-015-007-00b-020-003-00e-00d000c",
            INIT_1A => X"00200001-00c001b00380026001a0019-00c-01c-00a-048-037-012-036-010",
            INIT_1B => X"0003000100110005-001-009-017000c-007-00200010009-003-024-03d-039",
            INIT_1C => X"-026-00f000e000a000b-013001e-030-023002f-028-01d-006-00c-01f0005",
            INIT_1D => X"-003-00f00200010-038000d00220028-01d-006-0010006000300020003-00e",
            INIT_1E => X"-017003f000e-00e00130012-010-010-00b000d000f001b-00f0019000e-006",
            INIT_1F => X"-034-01e-03c-04c-020-0450004-050-03e001e0014001100000011-01c0002",
            INIT_20 => X"-006-032002c004a004c0007-026-013-004-045-026-005-01900000017000d",
            INIT_21 => X"000b000f002300190004-008001c00220004-008-007-00e00000007-009-007",
            INIT_22 => X"0019000b000000070008001a0000-009-00400050007-00b00000022-0110020",
            INIT_23 => X"-009-0030013000d000800200019000b-00d0010-027-01500030030-00f0021",
            INIT_24 => X"004200000011000d-025-00b-01f0017-013000e-006002600290000000e-011",
            INIT_25 => X"0026-00a-01d-004-015-034-01800000009000600210005001d0000-01a0019",
            INIT_26 => X"0008-027-005003a-018-00c0021-0340007002c-0010029-005-014-001-01a",
            INIT_27 => X"0001000e-014000e00140006000c0021001b0032000e001b000200100023-032",
            INIT_28 => X"-013-00b-01d-0040010000e0001-006-010-0030015000e003600160032000e",
            INIT_29 => X"00200020002f0011001a-0230011000c0015001c0042-018001500070018003b",
            INIT_2A => X"0007-02a-016000b001c-02600150010000f0029-01800080027-033-028-015",
            INIT_2B => X"-019-01c-012-048-039-019-016-007-02b-051-047-04b-002-00e-0040022",
            INIT_2C => X"003a-00b0012-00f-01b0011-0070015-014-0050002-01800090011-0380001",
            INIT_2D => X"003e-012000b00180009-00900020006000b000d-017000d001a0009-002001a",
            INIT_2E => X"000300290013-01b-058000e-049-00f-019-040-01e-031-016-00c-005-037",
            INIT_2F => X"-00e000f-006-03e-045-022-006-02b-028-034-01d-0030012-014-021-041",
            INIT_30 => X"-010-040-066-005-069-05b-037-0100000001e-016-0160001-00e-029-041",
            INIT_31 => X"-034-016-019-045-055-057-036-07e-029-02f0000001a-010-055-01f-027",
            INIT_32 => X"-003-01a-001-0040024-01f00000000-023-031001c000e0018001b00020014",
            INIT_33 => X"00030013-021-029000f0045003000170036003e-006-01d-013000e00330033",
            INIT_34 => X"001100350014-020-013-013-01e-0110002-017000b0007-0150001000e-011",
            INIT_35 => X"-009001b-01e-01d0015-023-036-01b0008001d-0140024003200160031001a",
            INIT_36 => X"-00d002b0013-0190000001600060005-00d-010000000150039000000210043",
            INIT_37 => X"-008001a0038-025-02e-022-012-050-02f002f-04a-06200080000002c0030",
            INIT_38 => X"00040031000c000d0011-069-06b-03d-03b-070-08a00220004-03300080015",
            INIT_39 => X"003200150031000d0004-01d-031-00c000c00440011002b001a-005-00c001f",
            INIT_3A => X"00130013-011-01f0002-00d000100000000-01a-032-066-030-044-059-016",
            INIT_3B => X"-020-00a0004-016-036000b-02200030002-002-01f-012-005-00f-01c0011",
            INIT_3C => X"0016-01e0005-006-00f-028-0370004-010-01b-02a-026-01b000f002d002e",
            INIT_3D => X"001f001c00200025-004-0030014-023-036000e-01400050022-0050014-005",
            INIT_3E => X"0017-0210029000f00180012000e-01d0019-01c-0060000-021-009-017-012",
            INIT_3F => X"000c-013-020-00d-013-00100020011002400150013-017-035001c-00f-007",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY9;


    MEM_IWGHT_18K_LAYER2_ENTITY10 : if N_BRAM = 10 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0004000c001a0005-00700370017001c0026001f000a0004-01d0009002e-008",
            INIT_01 => X"0001001e-00700040009-002-00f-034-014-039-021-02a000a-00e0019002a",
            INIT_02 => X"00210021001c000800240007-026-016-02a0010-026-01a0000-01f-003000a",
            INIT_03 => X"-01a-036-029-005-02a-03c-01f-00d-026-002-016000d001900000013000d",
            INIT_04 => X"0038001700330004002c-02f00040004-00c00000047-005001d00120011001c",
            INIT_05 => X"00060029-004-014001e0011000400110012-00900110019000d000e00160015",
            INIT_06 => X"-00b0004000b-003-00e0009-009-00f-010000c0008001a0011001b00150009",
            INIT_07 => X"001e-00f0018-00b-0030021-01b-0250063003d0047002d004c0069005b0022",
            INIT_08 => X"0011-006-027-043-012-041-0240004-022-007-00a0005-00d00050016001c",
            INIT_09 => X"0014003c00240001-005-0020022-007-006002f0028000c0011000b00140002",
            INIT_0A => X"0001001a-022-00e002300070000-00700110026001500410021000300140014",
            INIT_0B => X"00110012000e-016000d-010-006-011-00b00060000-013000f00060027001a",
            INIT_0C => X"-0010008-010-00d000e-00d00140016-0020008-002-029-032-00a-015-023",
            INIT_0D => X"-040-040-001004b001900340047000c002000070000-004-00f001f0009-026",
            INIT_0E => X"-016002d00050026002c0024003d-002-00b-01a004a0005003c000c00000006",
            INIT_0F => X"0032001d-0160000-005-02f-02c-019-00d-02800020016-03d-00a-003-018",
            INIT_10 => X"0011000b-006-02f-0140002000d001f001b0014000a0001000000240002-006",
            INIT_11 => X"001a-021-00b-01c001f0037-002-027-006000a0011-014-009-0050006001e",
            INIT_12 => X"-00c001c001f-021-00e00070017-031000f-01e-037-01f-05e-03c-023-032",
            INIT_13 => X"-036-039-006-021-02b00020004-0100012-01a-00e-028-010-02a0000-029",
            INIT_14 => X"-001-017-005-014-007-018-016-06f-06b-029-041-03a-02600120003-001",
            INIT_15 => X"-023-047-063-01e000e001600160003-021-044-013-033-00e-0210013-01b",
            INIT_16 => X"0015000c0026001b002a0037-001000c0024-0080029-014-01b-001-001-006",
            INIT_17 => X"-004-00d-00e001700090005-00e000d-0060009000f0001001d-017-018-002",
            INIT_18 => X"0007000a000c-011-015-002-05b-03c-024-00d-021-027-005-018-004-00e",
            INIT_19 => X"-017-001001600110019000c00070029-01e001c-001-03a-016-02e-0250024",
            INIT_1A => X"001000290003000000140025003300200031001e-001-009-0140018-003-023",
            INIT_1B => X"-003-0170001-047-00c-02f-03a-019-00f-04e0017-0240027002e00250011",
            INIT_1C => X"-00e-007002f001c0004-017-02e-04f-018-0110013-01c000b001700110003",
            INIT_1D => X"000500190002001b000d00190015000c-012-01e-00d-056-033-024-00f-012",
            INIT_1E => X"-00b-00f-00c00020005-009-0040010000d000f0001-019-0170009-01a-01f",
            INIT_1F => X"-00e-01b000f001a00360005002d002a001100360016005f0012-01b00170015",
            INIT_20 => X"-018-01a000d0014002b00250005001e0031-00c0001-0070010-04f-0540002",
            INIT_21 => X"-030-018001a-037-019-00a-016-035-02f-01c-016000b0025000c0027-00b",
            INIT_22 => X"0019000000360009003a002c000a000d-0220008-02a-057-007-011-033-00a",
            INIT_23 => X"-00c-042-034-022-012-016-0250008-00f-01a-012-01d0011-02a-0060013",
            INIT_24 => X"-00a-021-009-00c-00b001d-00e-045-005-036-02d-030-02f-016-00d-009",
            INIT_25 => X"00160003-00600110020001c0011-0150059001f000d002f-005-00e-056-025",
            INIT_26 => X"-01a-039-00300020002-024-021-009000a0000-00f00070011000100230002",
            INIT_27 => X"0042-00b00030048-007-03b0016-041-006-02a-01c-00e-011-01400100007",
            INIT_28 => X"00110024-021-040-02f-00b-015-0390011-01d000b-013000c0015-0100002",
            INIT_29 => X"0010000100020021-00f-0020003-002-007-007-0030007-01a-00500230004",
            INIT_2A => X"-0020020001b-004-012-018-014-0050013-001-01a0013000700130036-012",
            INIT_2B => X"-0290018-00e0000-00b000e000e002d-0070034002c-02c0014002f-027-034",
            INIT_2C => X"-017003700200012002f00130006002e00060004-013-005-00d002e0025-004",
            INIT_2D => X"-007000c0007-03c-024-02f0004-01900160000001e00200012-020-02d000d",
            INIT_2E => X"-003-032-0200020-017-046-02d001a-019-019-0060004-00b0033-0150014",
            INIT_2F => X"0019001100070012000a00010004-010000c-004000c0016001300190023-004",
            INIT_30 => X"-014-00a-017-015-00a-021-00700100003-00c-00a0015-00a0003001d-04e",
            INIT_31 => X"00020010-021-013-0150017-0060009-00100370018-002001f002800010009",
            INIT_32 => X"-017000d-008-02e-02c-031-02c0009002c00060024004d00000000-002-003",
            INIT_33 => X"00230010-0230034001e-00c0003000f0023-0100012000900090000000e-01f",
            INIT_34 => X"00020020-00e-010000c001a0007000300130024-00d00350025000200120000",
            INIT_35 => X"-027-05200140016-04d00360031-052000a004600030013-00c00210006-013",
            INIT_36 => X"-006-00f-026-01d-0040000-037-005000b-00a001d000000000009-008-018",
            INIT_37 => X"-009-00a0015-02f-022-04500190015-03f00200006-0650005003900040007",
            INIT_38 => X"-0250036000b-006002b0039-0110000-00b001c-00e00090020000d-0040012",
            INIT_39 => X"-006004a004a001900450052-03e-0050016-03a-00c002d-0210026001d-026",
            INIT_3A => X"0017001700390005-017-001-03200140005000a00170027-01e-026002c-00e",
            INIT_3B => X"-02e002a0000-02c0037-011-025002c-00f-02f003f0000-027002f-031-030",
            INIT_3C => X"0010-00a-037002c-00b-01b-01200180006-034000e002d-01f-018002b0002",
            INIT_3D => X"-01e-03400300002-024001c0003-054003f003100010015001a00070019-00f",
            INIT_3E => X"000d-02c000d-003000a0015-00c-022-0050001-061-00e0033-0300023004b",
            INIT_3F => X"-04a000c003f-006-00d-009-017-00800050014-00b0012-017001c-002000f",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY10;


    MEM_IWGHT_18K_LAYER2_ENTITY11 : if N_BRAM = 11 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00160015-00d-008-01d-033-00a000b-035-004001c-018-011001a002b-00b",
            INIT_01 => X"-0150023-017-0230050000a-034-024-001003b-0380000002e-03f-00a0015",
            INIT_02 => X"00140002-00a-01c0001-0180005-00f-0160023000a0027002f-004-0130003",
            INIT_03 => X"-01c-036-017-010-009000d-03a-02e00330016-007-031-03300160020-037",
            INIT_04 => X"-045002d-035-012-00d-039-0520015-039-040005f0025-00d0033-005-018",
            INIT_05 => X"0010-00a-011-019-00d-02a00370008-00e000d0000-01600050007-014-018",
            INIT_06 => X"00110052-037-0100011-032-013001b000e001c-013001f-005-02d0004-001",
            INIT_07 => X"-02c000e-040-02a0028-004-00b0015-003-03f000f0001000a-004-0110000",
            INIT_08 => X"-015000b-002-013-015002a-01f-025-00d-017-042-0270031-01d0009000b",
            INIT_09 => X"-018-032-01c-01f-0330002-0170026004c00130008001f000a-01300030005",
            INIT_0A => X"00070004-020-020-02e-023-03a0031-00d-005002b0003-00900210027000d",
            INIT_0B => X"00080029000f00430051004b003d0014-0070010-01000090012000b-0230008",
            INIT_0C => X"-005-039-034-01f-01b000800050006000c0021-00f00010003000a-00a-004",
            INIT_0D => X"0002-00c000b0008-00a-0020018-0130017000f-00b00060015-00700110003",
            INIT_0E => X"-002-0180013000c003e001100220002-02e0036-005-024-00c-005-03c0014",
            INIT_0F => X"-027-03900000001-001000800040016004b0070004d000f004a003e-0120015",
            INIT_10 => X"0033-014000b00020026-004001900270007001e001b-02d-025002e0007-006",
            INIT_11 => X"002e-008-028000c002d-005000600000004-01a0000-02a-020-04f-00a-00e",
            INIT_12 => X"-028-04d0039-008-01e0017000e000e-021-008001d-02f-018-03c-00f-020",
            INIT_13 => X"000f-01a-0090016-041-0210001001e-01f-0190033-002-01900110031-014",
            INIT_14 => X"-0010019-005-0050014001f001c001c000f-043-0400039-037-01200290008",
            INIT_15 => X"0008-00a-058-05d-035-043-056-0610003-01e0008001100310041000f0020",
            INIT_16 => X"000c0015001f000e-026-083-050-064-042-012-00c-002-00100410033001b",
            INIT_17 => X"0018001f00100007-0180005-00c-017-007-00c-0070000-0030018001e-00a",
            INIT_18 => X"000300010009-027-01d-01d0009-015-023-022003d-01f00000020-021-007",
            INIT_19 => X"000d-00f-0060015-017-002000c-01500150022-031-029-008-007-0100012",
            INIT_1A => X"0011-005000800100009-0010004000b-03b0008-008-010002d000c00080017",
            INIT_1B => X"001f0021000b000d001d-041-01a001e-02f00030017-01d0013000b0033002c",
            INIT_1C => X"001500110028-00c0018-007000f0016000c000b-01b0024-00700030028000c",
            INIT_1D => X"-039002b0044000200340048001700550039-022-026-0040000-0110003001e",
            INIT_1E => X"00030024-004002d-00d-0060022-006-00e001b-00f001e0024-00a0014000e",
            INIT_1F => X"000c0019000b001c0003001a-021001c-005-01d-00f000f-02700040000-012",
            INIT_20 => X"002a0018-00b00070003-008000b-00c002d-01c00260003-010001e0007000b",
            INIT_21 => X"0004-025000c00110003001a-00c0015000a-04e000b-011-008-027-0140029",
            INIT_22 => X"0001-03a-02a0016-007-0110034003a00290009-02000120017-02b00060015",
            INIT_23 => X"-01900070025-00100110014000d001c0015-007-0080001-00f-018001a0006",
            INIT_24 => X"000c000c000f000b002b-01100090006-006-009000b-0120002-00300000016",
            INIT_25 => X"-02000170004-00c0014-008-014-00e-0100002-01b00100011-01a00000004",
            INIT_26 => X"000f-00a-0070006-019-017-017-011-007-021-0040032-00500120016001f",
            INIT_27 => X"003c-010-034-018-01f-01a-02f0009-020-043-006-0120035001200130052",
            INIT_28 => X"00530032001e0038-0270022-001-00b00020039-023-009-0180010001e-00b",
            INIT_29 => X"00150000-00b-026-00b-00c-017-011002000160021002c0005-0010045-007",
            INIT_2A => X"0015002a-019-011-012000f-0220007-040-0180015-05c00190028-03b0036",
            INIT_2B => X"-01f0022-012-0150013-01e-043-0010003-012-03b-0220033-05500090025",
            INIT_2C => X"-012-01f-02f-00d-023-029-044-04f-04e-010-052-069001c0001000b0000",
            INIT_2D => X"-00c-01e001e0018000c0001-009-00e001d0011-0210027-008-002-0130005",
            INIT_2E => X"-002-019-0230002-014-033-0070023-009-01d0020-019-011000d0009-012",
            INIT_2F => X"-01c-017-02c-00e000200340010000b0013-009-013-0040014000800170028",
            INIT_30 => X"0004000800250034000b002b003c0017002f0003-02d0025002000250012-004",
            INIT_31 => X"000e-0160012002700160013-021-007-013-004-02f-01d-01900020016001b",
            INIT_32 => X"0012000b000f0013000a000b0001000700210026001b0006001a002e000e-047",
            INIT_33 => X"-0090018-0290015000b-00d0003002e-02d-03c-00e-03d-010-011-052-055",
            INIT_34 => X"-039-039000900280003003000270010001d-0030025-016-028002d0007-036",
            INIT_35 => X"000f0000-0130010-00a-0030009-002-01f-0050008-0140003-003-0060016",
            INIT_36 => X"0060004800000015002b000b-029-0200004-048-044-01b-02a-01200080015",
            INIT_37 => X"-008-02c00060009-0160006-010000900120003001a0002-00500220007-00f",
            INIT_38 => X"-0010009-0180008-014-008000000130019-015002a0001-017-042-01c0036",
            INIT_39 => X"001e-01500170037004200130047004d0011004100280028000e-01800450018",
            INIT_3A => X"0008-007001700220038004b001a004a0037003e0017002e002e001f0026002c",
            INIT_3B => X"0021003e0035-019-004-001002f00160010-037-004-01a-00b0004000b-010",
            INIT_3C => X"000b000b-038-026-039-010-00d-010000a00090000-027-021000000120003",
            INIT_3D => X"00190023002e0018-00e0013-009-016-007000a00000026-02f-00f-010-016",
            INIT_3E => X"0008001b000e001d-01c-02b00210006-0170027-007-0050022-00a-005-010",
            INIT_3F => X"0000-014-021-01f-00f-028-008-00c-046-045-037-004002a0029-0040024",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY11;


    MEM_IWGHT_18K_LAYER2_ENTITY12 : if N_BRAM = 12 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"-00f00070023000b-025-039-01e00340011-00b0022000d0006-0110000-03d",
            INIT_01 => X"000000080029-00f000a-00c0017002b-0020019-00a-015-00b-0020000000a",
            INIT_02 => X"0007-026-00b-024-0090012-03c000e-003-0050004-0030007-0200011-013",
            INIT_03 => X"0000-02e-020-011-015-025-0100006-0120018-019-011-0240024-008-005",
            INIT_04 => X"000e0017000d-01c-023-03400330023000c-003-004-00f-035-00d-01f-007",
            INIT_05 => X"-02c-034000e-007-017-007000b002c003d00400012001200530049-01b-014",
            INIT_06 => X"002f-0240018-015-028-028-029-01d000c-0030003000c-00a-001-003-01e",
            INIT_07 => X"-021-015-00f00240031-023-026001a-016-00d-00f-0080039001a-0080039",
            INIT_08 => X"00570015-01c0029-019-020-036-03a-024-002-02b-01a-026-025-00a-02b",
            INIT_09 => X"-00f00050000-0120006-0010004001b-0060012-001000a-01200090000-012",
            INIT_0A => X"000400130024002200100009000d0013-007-008-02c-0020014001300220036",
            INIT_0B => X"0036003d00000021-00c0029004c0027005600650051-001-023-0090012-007",
            INIT_0C => X"-02a-03d-0030018-0040014-0070052006c0033004400400057002f00480042",
            INIT_0D => X"-02300110000-07d-068-0470008001600140000-036-051-03e-03b-020-005",
            INIT_0E => X"-01f-01b002c-02a-00d000c00100010000a0017000e-015-007001300030019",
            INIT_0F => X"0020-00a0005-0080001-008000c-005-008-026001b00090023000d000d001e",
            INIT_10 => X"001400040001001200200027-003-00c-021-03d0000-01d000e00290017-012",
            INIT_11 => X"001e-025-0350004-019-0010003-01d-010-03a-010-00f00160013001f0027",
            INIT_12 => X"0023-036-032-005-074-046-02c-009000d001a-0200013000b-011-016-00e",
            INIT_13 => X"003600470040000b00280009-0030000-0220032001c0006-006-002-019-01a",
            INIT_14 => X"0006000d00380042004b-0050006-00b-048-05f-01b001100300023-00a0018",
            INIT_15 => X"0013-017-041-03800100014001c-00e-005-004-02b-05f-022002a00390018",
            INIT_16 => X"-00b00120018-043-029-019-00100040014-004-00a-006-00a-002-0180027",
            INIT_17 => X"00330044-010000f0000-063-06a-03f-012-015-034-024-02a000000120006",
            INIT_18 => X"000f0000-010-003001a-015001b0003-012-00e000e000a-00a-0190001-00e",
            INIT_19 => X"0004-00c-01f0001-009000c-023-00c0012-007-019-012-016-024-039-00a",
            INIT_1A => X"0001-020-03a-01a002100010005-006-034-004-02d000b001b-00e000f0016",
            INIT_1B => X"0020-016-012-01d-039-036-033001c00250021-00e00110005-00f0014-014",
            INIT_1C => X"-01100030005-002000e00010012000e001a-01b-014-012-01b-025-016-009",
            INIT_1D => X"-01d-02d00000045003d001400510070-009-00d0015-0020011-002-01a0047",
            INIT_1E => X"0029-02700290013003e003b-004002000440045-0250021-001000700010002",
            INIT_1F => X"000c000300130029001e0012-01a000e-019-0090008-023-00f0005000c0001",
            INIT_20 => X"0000-008-015-007-00a000b000c0019001000310021000a-00a0001-006-025",
            INIT_21 => X"0008-010-01e-00b0010-00a00010025-012-006-015000a001a00070000000a",
            INIT_22 => X"-037-048-034000500020019001400250007-009001d-032-00c-00e-00c0017",
            INIT_23 => X"-006-0210020002a0007000b-01e-0150006000500110028-002-0050000000f",
            INIT_24 => X"0020002e001a0026000e0031-0030018-032-02b0019-029-029004f00360034",
            INIT_25 => X"-00e-006-029-01d-01a-027004c0024002b-024-024-02e-01a-01b-0090005",
            INIT_26 => X"00240003000c0016000b0028001a0016000900330016-018-00f-0150010-002",
            INIT_27 => X"-02200030000001a0009-0210004-01c-015-02f001e001f-00f-008-01c-009",
            INIT_28 => X"0008-003-01700000017-003-027-034-01a00080000001900280031002b000c",
            INIT_29 => X"0023-01400050005-0150001-0140003000b004300580012002f0047-01e-028",
            INIT_2A => X"0011000a-01c-009-0010004000d001500090010-004-01a-002-001-01b-001",
            INIT_2B => X"002a000d001d-01c-027-031-00b000400070029001b00220029002e-005-00b",
            INIT_2C => X"0051003e-026001e0017-00f-0050012-00f0004000a001a0009002a000d0000",
            INIT_2D => X"-014-01a-012-01c002300260016-019-023-0150003-01b0000001e00240005",
            INIT_2E => X"-005-0010008-014-00a-0050008-010000f-006-00500060000-010-0200000",
            INIT_2F => X"00040004-0180006-009-0110000-014-009-0010010-015-00e-0040012000d",
            INIT_30 => X"001a-00a-018-018000c00020006001e-003-005000c-011-007001a0000000b",
            INIT_31 => X"-00b0007-008-002-00f-013-00b-0170007-026-01b-014-01c-015-017-01c",
            INIT_32 => X"-01b000d00070000000c0008000b0000-013-00e-016-00a-018-001-005-021",
            INIT_33 => X"00140006-01d-01b-015-015000b-013-013-010-0120008-019-016-0050004",
            INIT_34 => X"-008-0140000-018-00d-013-006-018-00d-00e-00d-015-013-00b0004-01a",
            INIT_35 => X"000a-012-013-01e-012-011-01f-021000000060009-010-01400050001-01b",
            INIT_36 => X"0008-015-024000a-010-008-005-0150001000a-01d0004-01800000001-010",
            INIT_37 => X"-01a-005-012-006-00c-00a0005000d-003-023-027-00c-00200010000000c",
            INIT_38 => X"-01b-008-00b-0040003-00f-010-00f000b000c0000-01b-01f-001-0020000",
            INIT_39 => X"-014-0120003-010000f-0190008-00b0006-0140000-01c000d000a-0060007",
            INIT_3A => X"-01d-01f-017-016-018-012-006-01e0001-02100050005-010-004-00b-01c",
            INIT_3B => X"00030003-014-01b000a-001-019-016-00a-01a-001-017-017-00c-01a000d",
            INIT_3C => X"-008-019-013-00b00080000-017-011-0050007-014-017-0190004-012-004",
            INIT_3D => X"0001-013-004-001-017000a0007-004-01e00020002-009-00d-00b000e0002",
            INIT_3E => X"-019000200010008-01e-0050000-0080005-011-0090000-006-00e-016000a",
            INIT_3F => X"00020000-013-01400090009-005000a-00e-0040008-007-00f-00100160008",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY12;


    MEM_IWGHT_18K_LAYER2_ENTITY13 : if N_BRAM = 13 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"-00a-01400000008-0180007000a000b-015-011-00e-02d0014-008-0130015",
            INIT_01 => X"0001-0250018000a000a003c00310010002f0037002b-025000b-028-03f-01b",
            INIT_02 => X"-048-028-04a-039-004-007001c001a003b004d002300550030-00600220017",
            INIT_03 => X"-016000a-005-010-022-0030021001b0017-028-02e-00f-01e-035-01a-004",
            INIT_04 => X"-019-0130016-001-008000b000b0005002a000d0023-00d001a-00e-047-06b",
            INIT_05 => X"-050000200000014-03700170000-00c-0020003-00c-01e0008-00a-026-021",
            INIT_06 => X"-02f-035-032-00900100000-005000c-007-03c-016001d0013000f-00f-017",
            INIT_07 => X"0010000e-01d00020014-0340006-004-005000f000f001500160022001b0011",
            INIT_08 => X"0019-02700010000-058-055-030-00e000b-03000100030000c002100440035",
            INIT_09 => X"-0170001000d-0070007001a00020021001400060019001f-011-011-00c-049",
            INIT_0A => X"-021-017-02a-013-043-03f-04a-03f-02b0002-01e000e000e00050004-010",
            INIT_0B => X"000800050019000e-01d-012-02a0027-00b-024003b0019-008-004-010-01a",
            INIT_0C => X"00150015-015002300190006001000220015-0120005000a-02c-034-023001d",
            INIT_0D => X"00160027-026-0040007-063-043-01b-0140032-012-030-034-027-005-066",
            INIT_0E => X"-0320015000500180020001e-0030027001f0007-01900010023-00e-0030015",
            INIT_0F => X"-00800150017000a00090003-01d-012000c000e-020-005-01a-0010009-03f",
            INIT_10 => X"-048-034-03b-037-014-022-00e0017-015-0090001-042-02b-0050007000b",
            INIT_11 => X"000500190021-013003900350012-00d000b001a00040017002f-028-004-009",
            INIT_12 => X"-002000c000f000d000100120024-001-005-009-017-00b-037-068-030-047",
            INIT_13 => X"-076-022-0100009000c00330035004e00430055002600260059002600340043",
            INIT_14 => X"0031002c00180008-003-014-01e002a0026-01a00310018-006000a0008-01a",
            INIT_15 => X"001b001b000f002c00280022-011-01c-033-002-009-01300250000-001-021",
            INIT_16 => X"0000-020-012-003-013-039-027-0100039000a-001001a-00c-004-005-00a",
            INIT_17 => X"0000-018-022-0120023-00a-015001e-004-003001600060010001b-013-01f",
            INIT_18 => X"-014-00f-00f-010-0040020-0070023001b002c00060022-013-00900000018",
            INIT_19 => X"000b0013001500280003-004-034-019001a-031-01f-015-031-01f000e-003",
            INIT_1A => X"000a00040022000000170034-007-001-002-01b001200180012000b0006000a",
            INIT_1B => X"0006-01d-013002a-055-025-01e-02d-02e0018-00b-01d00510009-029001a",
            INIT_1C => X"-00d-02e-02f-034-045-01b-024-006-016-010-00b-024-00f0014-023-016",
            INIT_1D => X"0017-010-00b0016-020000d000c-01900090022-025-0180007-037-01f0006",
            INIT_1E => X"-017000a001d-01700000022-0120000000500340002-02000350005-00f0011",
            INIT_1F => X"-00f-007-0080016-00b001600030004003600450020003f006f001d005a0045",
            INIT_20 => X"00350001-01e-00e-01f-01b-005-02e-052-02d0008-004-00c0031-006-02b",
            INIT_21 => X"0034-007-020-026-0190014-025-020-002-01f-00e001b003500490017007b",
            INIT_22 => X"005b0038006900270036-02a-0240011-0020005-018-01b-01a000f-01a-011",
            INIT_23 => X"0012-019001c0022-014-00f0016-0090000-00f001e-01b-00f0035-005-038",
            INIT_24 => X"0014-00900040016-0070000-01f00000008003f001e-043-029-0070026-010",
            INIT_25 => X"-028-007001a0001-028000a000a0021-011-0140009-02c-0210001-02f-010",
            INIT_26 => X"0010-036-00a-010001a000c0028000f-0040028-0020006-028-0170019000b",
            INIT_27 => X"-009000e0014001800230015-050-02a0003-029-01a-02c-010-008-02b-034",
            INIT_28 => X"-035-03e-0280002-01e-016-02f0006003100330035-021-0090033-027-008",
            INIT_29 => X"0023-01b-007-02d-030-00e-03f-004-00c-007000f0016000d-03b-0230044",
            INIT_2A => X"-027-01d0020-025-015-00f-010-03e00010010-023-010-029-032-016-023",
            INIT_2B => X"-061-0020003-035-03b-01e-034-0070001-021-006-018-0060002-0420022",
            INIT_2C => X"0048-027-0210003-008-023-01c-02e-00c-029-006-026-06400170016-033",
            INIT_2D => X"00070036-008-03c00050030-030000b002b-00d000e000b-04c-00e0028-004",
            INIT_2E => X"-00f-0090006003800390069004e003c005500660023-020-0060000-026-03c",
            INIT_2F => X"-04f-025-036-056-021-02a-007-004-00e-04c-006-003-0300004000d-004",
            INIT_30 => X"-009-016-01c-0050018-025-00f-011-00e-01b-024-01500130047-01c0001",
            INIT_31 => X"002e003d-030-0120023-02b-025001c-010000b-00e-022000b00270007-02a",
            INIT_32 => X"00030021-017000c-017-007000a-021-01f0015-017-00e-005-009-00b-01a",
            INIT_33 => X"-01300070032-02f-019-004-02a-01d-005-024000e-029-02a00140028-008",
            INIT_34 => X"000e003a000300110029-028-035-014-016-00c0007-01100170043-024-034",
            INIT_35 => X"00050004-01f-01e000c-011-02e001400240012000a-00700110021001a0023",
            INIT_36 => X"0012-004-004000c0014-010-010-00e001900360037-00f000300130009-00e",
            INIT_37 => X"-004000f-0320015000a-0040041-005-01a-0050009-02a-008-02e0010002c",
            INIT_38 => X"0011000c0023003a-02b-0020031001e-024-0040034-037-00a00060019000c",
            INIT_39 => X"00000008-007-00d0001-026-0060010-03c0000000e0006-006-001-020-015",
            INIT_3A => X"-0200000-00b0007001f-00c000d0013000a002a0007-00f0015-009-0070006",
            INIT_3B => X"0036000a-010-014-001-03c-049-010-01b-013-00f001c-015001d00070017",
            INIT_3C => X"001c-00a0024-004-02e-00f-003-023-019-03c-025-0580000-0160010-008",
            INIT_3D => X"-01b-015-030-027-02d-00d0007-023000b-00c0000000100060019-005-02c",
            INIT_3E => X"-0110007-010-023-034-033-0490007-026-027-01f-01d-03c-01c-015-00f",
            INIT_3F => X"-033-05c-043-06d-038-020-0210006-025001f0011-019002d0004-0060010",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY13;


    MEM_IWGHT_18K_LAYER2_ENTITY14 : if N_BRAM = 14 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000a000a0010004a0048000d0066005b005300900038-012-00d0007-027-020",
            INIT_01 => X"-004-022-036-00d-025-00f-003-019-0100010-00c-005-011-007-005-013",
            INIT_02 => X"-0300009-002-014-013-023001d0000-01e0023-007-002-00a-002-0130008",
            INIT_03 => X"-036-033000f-02e-031-026-038-0010009003e00120018003b-005-002-017",
            INIT_04 => X"000d-00400000007-0150006000b-013000f0045003b0000-01e000b0001-03a",
            INIT_05 => X"-019-026-027-009003a-001-01a-001-036-023-032-021-00c0012-00f0025",
            INIT_06 => X"004e0018002a0034003e0002-00b0013-0090006-041-01d-00d-01d-03a-006",
            INIT_07 => X"0008-026-00a0010-010001200070037000e-014001e000d-026-004000a-00e",
            INIT_08 => X"-008-003002400120004001b-020-002-00b0011000a0000-003-0100022000c",
            INIT_09 => X"00170016-03c-044-026-02a-031-034-008-023-012-03b0012001c-05f0025",
            INIT_0A => X"0000-01000160010-08a-060-01f-05b-085000b0003-03f0001000f000d001f",
            INIT_0B => X"00000028001600010022002c000400210011-01e-0180025-056-042-0090039",
            INIT_0C => X"0006-00e00280029-00e0020001a001e0037-01b-007-018-022-012-025-031",
            INIT_0D => X"-02a0027001c0028-01300210010-018-007-0050012001a-0070000-008000f",
            INIT_0E => X"001a-01b-028000d002c002d-02a00170015-0190013000d0010000f0019-016",
            INIT_0F => X"002000110000000b0020001b00100002-0010023-004-02100060025-008002a",
            INIT_10 => X"002e-018-0020020-01d-014000b-020-00e000f-020000600030012000c0023",
            INIT_11 => X"-04a-022-00a-037-03d-026-03c00390003-00400280038-003-00d0023-03f",
            INIT_12 => X"-0010005001c-010-019-009-02a0019-0090011-012-020-03d-0140016-01f",
            INIT_13 => X"-0190033-0050005-007-039-0260035-006-0490059001c-014-012-01d-01f",
            INIT_14 => X"0022-021-018003b0001-01d-00500020027-003000d-006-02d-00c0019-021",
            INIT_15 => X"-00d001b-020-0150016-018-017-00e-040-021-02b0016002a-0310023002a",
            INIT_16 => X"0000-01c0003-01d000600120004003a00170016-015000c0016-03b000c0013",
            INIT_17 => X"-048-00c0008-00c-00c000a-00e-00f000e-008-0390025-002-01e-002-058",
            INIT_18 => X"-00d-014-03f-002001b-01b00200027000c00250009-006000d00000002-009",
            INIT_19 => X"-013002d-010-024004d0016-011-01000130026-053000e000d-02c-003001c",
            INIT_1A => X"0000-008000400120006-005-0020012-009-00e0007-007-007-007-0160005",
            INIT_1B => X"-0120003-00f-008-00a-0020001-0100006000b-00a-00c0000-00100060000",
            INIT_1C => X"0000-0180005-00d0006-001000d-002-00e000e-00a-017-0030006-00e-00a",
            INIT_1D => X"0007-016-016-011-0010006-004000a-00f000c000c-006-00b-017-005-006",
            INIT_1E => X"0004-019-00e0006-00c000600000000-002-007000b-0110002-0090009-019",
            INIT_1F => X"-00e-00500020012-014-00c000a0008-0070000-013-00e0001-00f00000000",
            INIT_20 => X"000e-019000d-0140000-014000a000a-014-0050010-013000f-00b-00d000f",
            INIT_21 => X"000a-00c000d-0100011-005-001-00e-004-01200000001-01a0000-0080001",
            INIT_22 => X"-010-00f-016-009-0030007-0080006-003-007-005-015-013-011-011-012",
            INIT_23 => X"-0030002-008-004-00c-012-00f-0110009000b-016000f-00e000e-005-014",
            INIT_24 => X"-015-00d00120007000f000d-00c0009000d0001-007-018-015-01700060000",
            INIT_25 => X"-019-01b0008000c-013000e-00d-010-00d-014-019000a-01700060005-008",
            INIT_26 => X"0003000b-007000400010006-007-014-013-00a-009-012000d-01000010005",
            INIT_27 => X"-014-00c-0110000-00d-017-0040006-0140005-004000a-011-014-003-016",
            INIT_28 => X"-002-003-017-003-00d000a-0080009-01e00000001-0190007-0020001-016",
            INIT_29 => X"-00c-00b-005-0120008-0100003000d000f-002-01100070005-010000c000e",
            INIT_2A => X"0015-013-00d-005-01c-010000c000b-00f00050012000d-017-00c-005-013",
            INIT_2B => X"-010000b-018-015000f000d000a-01000070002000c0007-004-00d0004000d",
            INIT_2C => X"-0100000-016001000110004000c0015-009-003-01c-00b-004-01a000a-001",
            INIT_2D => X"-0020019001d0032000b00050026-005001a00240002-021-02b-0060000-007",
            INIT_2E => X"001100140008-006-00d0015-007-004002d00130003000f000a-01a-002000f",
            INIT_2F => X"-0320001-003-00f-039-00c-009-01f-01300040002-0040000-02d-033-003",
            INIT_30 => X"-00b-01a002b0013000500250018-01900000006000b-014000f002500050007",
            INIT_31 => X"-005-01a-041-0030009-03e-05e-006-00d-00900070018001c000d-0080014",
            INIT_32 => X"-00a0014002d001f000a-00e-00e-0010003-022-00c000000010016001a0004",
            INIT_33 => X"0001000b000f000c000f000d-03d-03a000f-040-03e-00c-00d0004-0170008",
            INIT_34 => X"0005-028-0050006-03b-017000e000f00060000000b0005-0060033-00c-036",
            INIT_35 => X"0013-020-0040000-03b-051-019-04c-010-00f-006-0100020-01d-03a-002",
            INIT_36 => X"-036-0310025003b0000-00d-01c-02e-009-038-038-010000b001d-0240009",
            INIT_37 => X"-002-01100000008-02a00000011-006-006-01b-029-017-00c-0100010000c",
            INIT_38 => X"-01c-0040006-00d-00c-001-0110004-01b000b-024-0120029-044-018000a",
            INIT_39 => X"-00600260004000b0017-001000d-008-00a00170019004d0012000100340053",
            INIT_3A => X"-0010010-0190000000e-0010000000b-00b002b-00d-019-009003b-023-017",
            INIT_3B => X"000e-019-01c-00a-015-01a0006-006000c-011-013-02c-01c-030-014-001",
            INIT_3C => X"-025-0100012-003-00a0009002000310018-01d-01e-018000c-010-02e0012",
            INIT_3D => X"0023-00f00030018-010001e002400290000-01d0028-00b-048001c-00b-03a",
            INIT_3E => X"-0010000000600080001-00d0000-0020007002300060013000e00380029-024",
            INIT_3F => X"00070010-008-0030019-003-02f-027-00e-042-051-047-030-028-049-067",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY14;


    MEM_IWGHT_18K_LAYER2_ENTITY15 : if N_BRAM = 15 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"-03b-051-07a-063-01900460026-049-011-005-00b-0400001003d00280013",
            INIT_01 => X"000000000023003400100023-004-00a-002000300050000-0080000-003-008",
            INIT_02 => X"0014000f001e001f00220022000f001c-024-015-004-0210012-030-010000a",
            INIT_03 => X"-011000a-015-013-00d-004000a-013-00b-007-016-00f-01e000a-014-00e",
            INIT_04 => X"000c00080001-008-0040001-0030001000400140002-00d000b00000012-005",
            INIT_05 => X"-0110015001b00140012000a0002000900120047003700000012001800250014",
            INIT_06 => X"003300070015001600210027002a0010000c-007-01b0003-004-01300050014",
            INIT_07 => X"-02d000c0018-01400280010-01a0024-00b-002-00200050009000e0005-004",
            INIT_08 => X"0016-0060018-016-0190014-032-014-007001d-007-009000d0001-00d-014",
            INIT_09 => X"-005002600130008-01c-001-008-00e-013-00a0000-0080014-00700090008",
            INIT_0A => X"-00f-00e-005-001-001001f-007-002-018000e001b-01a000f0005-004-004",
            INIT_0B => X"-01f-003-00f-024000500190008-00f-07c-01f-06b-093-092-06c-022-05d",
            INIT_0C => X"-07c000f0031001d000800320034000e-008-00e-006001d0001-00800110012",
            INIT_0D => X"000c0002-00f-006-012-010001a00080024002b002d0029-02d-01c-024-04b",
            INIT_0E => X"-05b-059-056-05f-0570000-005000d00060017001100300027002e-017-019",
            INIT_0F => X"-014-00d-00f-0030023-001001c001c001b0014-015000c-002-010-006-00d",
            INIT_10 => X"00090018-00100000017001500030015000e001500220009000a-0130015-017",
            INIT_11 => X"0002000e0019001800080027005700480035000b004900220001000e0015-01a",
            INIT_12 => X"0008-015-01c-0390018-00f-013002300290040001a000c002c-01e-01c-00e",
            INIT_13 => X"-00a00130004003c0026-007000a0032001f-00f0008-00e-02d-037-02f-007",
            INIT_14 => X"-001000f-01c0004-015-018-00d001b0033002b000a00370021000600170002",
            INIT_15 => X"000600080027-003-005001d-02100010004-02b001400360009000600150009",
            INIT_16 => X"0017-0090018-01f-00f0021000a000400240007000b-01a-025-0020016-029",
            INIT_17 => X"-01e-024-016-00f-037-0040038002c-02f0006-01d-01d00120012-01a-020",
            INIT_18 => X"-007001e-00a0007004300060016-026000d0032-042-01b0014-03200040007",
            INIT_19 => X"0013003a-02f-003-010-07f-039-00c-02600180037003c0003-00f-0100008",
            INIT_1A => X"-021-040-01c-009-00d-041-013-009-02c0003-037-00f-0100008-01e-015",
            INIT_1B => X"-00d000f-019-003-00100000011-02700060021-0200009002c-008-009002d",
            INIT_1C => X"-0130018002f-00d00020024-00a00190023-01800090009-009-018-03b0017",
            INIT_1D => X"000b-01b0008000f000800180006-00f-009-04b-030-030-04d0014-00b-030",
            INIT_1E => X"-02000110015-01a-016-018-01d-00d0011000c0003002e000b-016-004-00f",
            INIT_1F => X"000400130007-009-010001b-030-008-03f0013-02f-00e-002001d002d-009",
            INIT_20 => X"00150016-005-0180011-024-01e-004-058-016-046-01b-00c-00d0001-005",
            INIT_21 => X"-012-015-00a0021-00800090013000800060020-02900030002-031-00e-006",
            INIT_22 => X"-009-00e000000000010-003-00a0002-00800260014000f00490023-00c0018",
            INIT_23 => X"00330059000e000400200000-013-0060006-041-0170013-005001700280032",
            INIT_24 => X"003f001100360034-010002a002d-037-00d-002-01e-01a-01b-00400200013",
            INIT_25 => X"-028-025001a-02f-0160000-007001e0018-0300006003e-006-00f0013-007",
            INIT_26 => X"002e003b000300380024-007-016-01e0004-02c-008-0090013-014000a001f",
            INIT_27 => X"002a000a-01d-001-027-039-01e0005-025-013-011-004-011-028-0060010",
            INIT_28 => X"-0200012003b0018002d0020-036000c001b-042-01b001900260028001a-011",
            INIT_29 => X"000b0004-001000c0002000d000100020009-018-02e0026-00e-010-0100025",
            INIT_2A => X"0021-07c-0130006-078-01000190031001d-0030016-019-024001a-007-01d",
            INIT_2B => X"0003-012-0240008005000280022001b003e0029001700050004000f0030-01a",
            INIT_2C => X"0013001b-01f-005001a0013002e00170014001b0010-0040026000c-024-001",
            INIT_2D => X"0038-029000f-00b-027-001-00a-00e002e0016-02a-005-00a002a001c000f",
            INIT_2E => X"001a00250018-020-013-0020017-00e0008-021-0290017-01a-00f-011-023",
            INIT_2F => X"-00a0004-03d001a001f-0220024000e-018-0220012-01b-02b00020029-014",
            INIT_30 => X"-01e-017-016-001-01d-003-00a-01d-014-002-002-030-0110004-028-037",
            INIT_31 => X"002f0000-005000700160022-04d-03400200006-01b-0090002-00f0005-001",
            INIT_32 => X"000800260009001900190009-0070018-033-01c00110026-026-02a-0270000",
            INIT_33 => X"0016-024001c0006-03d000a000b0012-00900170029-008-029003300060013",
            INIT_34 => X"001400030010000c0022000e-007000e0002001700000002-00c001f-024-01c",
            INIT_35 => X"-01e0022003d002e-00500170038-004-004-010000a0037001d-00c003d0006",
            INIT_36 => X"-02000400007-02a-00f-01c-01c003c-017-0450043-031-003-02800000017",
            INIT_37 => X"0010000b001300380004002900000004002c-013-00a001f001a-0230009-02f",
            INIT_38 => X"-01a-036-045-00d-031-011-032-005000f-008-017-014000a-00a0002-027",
            INIT_39 => X"-017-00f00000006000b001a00150001001c0013000c0007000a-0170016000d",
            INIT_3A => X"-033-0200009-00d0009001a0000000300370017000a0001-015-0050012-025",
            INIT_3B => X"-01500060015000a002a001f0003-006-01a000f-00700220008-00d-03a-01c",
            INIT_3C => X"0018-00900050004-0170017-00a-027-01a-004-01d0006-006001300200009",
            INIT_3D => X"00000006-00c000b0020-007-004-015-011-01f000e002e0001001b002b000c",
            INIT_3E => X"000d-0020047002a0010005000060028004b006b0054-022-025-017-038-028",
            INIT_3F => X"-01a-039-00e-00f-0070012-034-0130009-02d-03d-00900090008-029-032",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY15;


    MEM_IWGHT_18K_LAYER2_ENTITY16 : if N_BRAM = 16 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"-011-010-030-020-018-0060007-0020016-008-0140017001f0006-00d-01c",
            INIT_01 => X"000c00090018-00500100015-017-01d-015-01d-01f001c0030-01b-0290005",
            INIT_02 => X"000b000e0002-00a-0020024-023-00d-02f-007-014-0120003000d0016-002",
            INIT_03 => X"00310027000b-01e-0140013-0180005-017-009001b001d000e0023-0030033",
            INIT_04 => X"-010-025000a001c0003-0160000-01700010022002200230037003c-006-02e",
            INIT_05 => X"-03e-0320002-020-03f-02a-009001800000009-00200000004004100160020",
            INIT_06 => X"-007000d-014-0090010000a-009001d0018000d001b00260019001a00170013",
            INIT_07 => X"001100210042-012-03e002d0028-05c0028-001-0030004-01e-030-011-040",
            INIT_08 => X"-071-00b-01a-052003f-04a-0410036-049-04200550009-054-009-014001d",
            INIT_09 => X"000600220009-016-00e0000000a0020-00e0006-001000a0007000e00130024",
            INIT_0A => X"0040003500230009000d0019001e0005-00e-012-044-0130000-0330002-01c",
            INIT_0B => X"-024-0180008-018-02c0027-004-0080003-0050002-012-019001e0030-005",
            INIT_0C => X"000b000e0012-019-007-01d-001-01f0000-032000100110000-005000f-014",
            INIT_0D => X"-00b002c-03f-0160013-0200036000e0001003b002c-0020012000c-00b000c",
            INIT_0E => X"-005-01f-0040028-01f0003-004000d000e000a-014001a000b-03e-016-009",
            INIT_0F => X"-03200280032001e0042001e000300040015-0330010000e-00800290014-009",
            INIT_10 => X"0018-00f-012-030-069-008000b000b-01b0009000a001b00030014-018001b",
            INIT_11 => X"001c-01c00000015000f0013000400000025003a-0090000001e001300210013",
            INIT_12 => X"000200060014-01b-01d000600220009-015-002-026-010-024000b0002-013",
            INIT_13 => X"-02e-025-00c-0020002-01f000100160028-067-0520003-063-0740038-03c",
            INIT_14 => X"-089001200260002001c0002000e-0030015001f-0130000000a-0010016000e",
            INIT_15 => X"001a0019000e-004-0070025-02d-0160003001b-00e0000-025-06f-044-03a",
            INIT_16 => X"-064-04f0006-033-049-031-01e-013-038000a-004-014-002000300100000",
            INIT_17 => X"00110002002b0016-012-00200180004-016-01b00060010001c000e00070001",
            INIT_18 => X"000c001f000e-00d0005-0010009-012-00700180031-00e00470025-008-00f",
            INIT_19 => X"001f0012-00f-03e-01e-00d-05a-0110017-02a-0270017003b002800410031",
            INIT_1A => X"003d00380028-001-037-059-024-027-04d-027-010-00e-019-043-033-00e",
            INIT_1B => X"-00d-04f-026002c-002-026-00c001a0045003a003e002f00000004-0230012",
            INIT_1C => X"000c00070011-0050015-028-0140015-0030048-009005200220013002d0018",
            INIT_1D => X"-00d0001-024-00a-00b0001-008-00500150003000f0016001e0021000c0011",
            INIT_1E => X"000d00140018-02a-06a-041-045-0450000-006-008000f0014-009-0010014",
            INIT_1F => X"00040010-011-013-00f00060012-02e00230015-01b-055-025-02d-01d-045",
            INIT_20 => X"-022-029-020002200120013-0010041-00e0004001a-010-00f0024-01a-01a",
            INIT_21 => X"00090005002c-0060004-025-01a001b0010001700220010000700110002000c",
            INIT_22 => X"0009000f00230017-02900460011-003001e-009-00f-00c000a002600090012",
            INIT_23 => X"000b0007-0060010000a-00f-009-01b-018-0170002002e0030-00400030020",
            INIT_24 => X"0004001000110025000d001a-00300110015000c0001000a00010003-00a-002",
            INIT_25 => X"00020018001f001e0029000b001b-020001d001600270029001f-00b00350045",
            INIT_26 => X"001c-0150017-01b-007-011-011-028-0010023000f0006-0150010000a-018",
            INIT_27 => X"001a-00800040000-0070009-01c00070024-00d-017-004001d000a003c0024",
            INIT_28 => X"-00f-00400140011-01f-013-03e-032-029-049-008-029-037-023-0100006",
            INIT_29 => X"-012-025000300250005002a-007001d-00900150026001a-0070049001d002d",
            INIT_2A => X"000b000800170003-00f000f00180010-00800140006-01e0025001c000e002d",
            INIT_2B => X"002a00190003000c-027-01600090000-01c000c-01a-017-03d-051-01c-014",
            INIT_2C => X"-042-03a-045-043004f002a000a0002003e000a-01b00120006-00a-00d-001",
            INIT_2D => X"-00700210014-0100008-01200180014000d-005-00e-00f-03a-032-0070017",
            INIT_2E => X"00010011000c-00e00000004000b00290003000500050005-006001c00080000",
            INIT_2F => X"00110028002c001c0016001c0002-06e-049-03a0015001b000800200008002a",
            INIT_30 => X"00040006-0110001-02c-0360009-00e-037-011-028-047-00c-00a-00b0013",
            INIT_31 => X"-002-003-013-01d0003000f0016001000050000-01b-005-002-01c-019-004",
            INIT_32 => X"00000008000d-009-005-01b-016000c0016-02b001f0015-001-002-00b-02b",
            INIT_33 => X"-02c-020-002-041-045-055-03e-072-05500190022001d000f-0100000-04a",
            INIT_34 => X"-048-03d0031003f-0110040-005-012001c002e000a-00a-002000100130016",
            INIT_35 => X"0001-0040029001000010002-00c002e002200010038000d00240007000a0005",
            INIT_36 => X"0012001f0018001e0005002a-017003d0019-013-001-020-080-035-064-00b",
            INIT_37 => X"-0010010-015-0050012-028-02f001a-01f-02f-015-032-045-047-066-030",
            INIT_38 => X"-03e0019002700230023001200170018-003000e00440046001e001e-00d-004",
            INIT_39 => X"-034-017-029-006-01d-002-02d-02d-006-015-029-02f001a-034-02a-013",
            INIT_3A => X"-013-011-013-045-015-026-0340021-05b-085-05a-02d-070-04f000a0017",
            INIT_3B => X"00000023000d00080018002500090016003d0004-00b00040029-041-01a-047",
            INIT_3C => X"000d0004-00c00100014-011-0030006000c0010000b000000090003-01c0006",
            INIT_3D => X"0018002400030011-002000f001000100011001d0020-03b-020-011-04e-016",
            INIT_3E => X"-022-031-01e-0160006-00a-00c0022002b001800010048002d0004-024000f",
            INIT_3F => X"0013-006-00800080018-01b001d-00c-006-002-00c-020-00a-00e-011-014",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY16;


    MEM_IWGHT_18K_LAYER2_ENTITY17 : if N_BRAM = 17 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"-00d-0130004-001000b0007002b002d000c001a00080047001e-0230015-004",
            INIT_01 => X"000c0016-0050008-021-0110021-024-028001c-0020018-007000f-013-013",
            INIT_02 => X"002b-013-006-019-018-01f-02b-031-010-02f-01f-0330004-00c0009-007",
            INIT_03 => X"-0020009000d-006-0160007001500000002001e0034-01500200019-009-012",
            INIT_04 => X"-01a000c-006-011001a0000-0340004001e0000001b002b0013-0130004001d",
            INIT_05 => X"-051-02d-042-020-036-00d-047-069-058-00c00010006-01b-025-026-010",
            INIT_06 => X"-028-022-00400060023-03a-030-026-073-021-015001a001b0013001d001d",
            INIT_07 => X"-0040010002e0023000b000a-006001a001200220004-0120021001d0000-008",
            INIT_08 => X"00080010000000190008000a-032-01b-014-035-01d-04e-038-03d-0300006",
            INIT_09 => X"001300220016-00c-0160006-00d-008-031-00b-026-032-029-0520006-023",
            INIT_0A => X"-027000d0010002c001b0016000f001d0014001b0007-004001b-009000f0009",
            INIT_0B => X"-02a-01b00120008-0180009001500000003000100000006-00700020013-01c",
            INIT_0C => X"-00f-003-0080000-0280000001b002b-022-03b-026-01e-032-0230002-002",
            INIT_0D => X"001600030004000a0001-013-0050012000f0001-0170009-002-036-022-014",
            INIT_0E => X"0008000e0005-009-014-00700000000-011001b-015-021-0210021001f-041",
            INIT_0F => X"-031-0150019-0050000000c00100019-02a-008-045-01a-01d-0010002-005",
            INIT_10 => X"0020-01b-0050012-00c-010-00d-008-006-01f000d-02a-00c-026-031-006",
            INIT_11 => X"0006-033-0030029000b-00e-0120002000b000d001f-03a0007-006-00f0000",
            INIT_12 => X"001f001f-01c0010002a-009-0050037-02700110008-00d-0020000-02b-01e",
            INIT_13 => X"-0130016-00f-0400015-017-039002a-010-009-0080044002c-0270003004e",
            INIT_14 => X"-04a-008-024000e0005000f00270007004700290012-015001c-025-0110023",
            INIT_15 => X"-00d-02500360025000c000f0019-01a-02c000b0005-005-00a0013-031-009",
            INIT_16 => X"0016-001-026-007002f00270003003a-030-024003c-019-0280040-0040006",
            INIT_17 => X"-00c001c-020-030002a-007-042-0140023-00b-011-012-019001a-02a0015",
            INIT_18 => X"0032000800310006-002-0030007-034002a-0080002-00c-029000b-010-012",
            INIT_19 => X"-002-00e0001-013-023-0080016001500020004-01500030027-01e-0110020",
            INIT_1A => X"-011-020001d0010-008-003-006-01e-0420006-018-04000220019-009-01d",
            INIT_1B => X"00190040-03f-0130055-012-00b00110042002e001b00500052005e0006001e",
            INIT_1C => X"0023-01e001b-01f-02600130016-03800030028001a0001-022000d-013-032",
            INIT_1D => X"002d001c-0090000-01d-003-00b-016-01d000a001c001d001700270005001e",
            INIT_1E => X"001f002100180012001d00050008-01a0029003e00320017003b0050-036-03d",
            INIT_1F => X"0008-024-02d-006-011-008-0020008-026-0360036-011-02a005400220011",
            INIT_20 => X"0006-002-00e-001-002-01b0004-010-00d00040029002e00250005001d001d",
            INIT_21 => X"00290007-04c-059-04b-045-077-071-06d-042-05f-0080037002f00280037",
            INIT_22 => X"-001002700290015-053-049-052-04d-06a-031-057-051-036000000270018",
            INIT_23 => X"0002002b0034-02900120010000e00280032-014-013-00d-03b-024-00a0026",
            INIT_24 => X"001c-011000d-00b000700020002-004-019-026-00c0004-00b001a-01c-00b",
            INIT_25 => X"-039-010-0110017-009-02e-009000000090000-007-017-002-0070000001e",
            INIT_26 => X"-023-012-036-014-00f-01b0004001c0009-009-0260014001d-002001e0002",
            INIT_27 => X"0028002a-0140000000a000f00060007000e-015-00f000f000e001a00110019",
            INIT_28 => X"00070007001a0019-01e-023-016-00100060000-0020012000a000e000f0011",
            INIT_29 => X"-01c-01c000700160000-0060021000e0019002600160027000c0005000f000b",
            INIT_2A => X"-009-00d0015-012-02e001e-028-054000d-01d-02a-00a001e002b00020017",
            INIT_2B => X"0027-009-007000b-002000b-008-003-003-015-01200050000001e0028000f",
            INIT_2C => X"000f-00300170013001a001f0010002300290007-003000c-007-00500000017",
            INIT_2D => X"0009001b000a00290016-03c-039-00e-089-03b-067-060-01d-02b-04e-01d",
            INIT_2E => X"000b-00e00070009-007-01b-006001e00050008-002000a0008-00f-00b-00d",
            INIT_2F => X"-005-00f001300130003000a-00e00230029-02200060002-0150017-0040018",
            INIT_30 => X"-00c-03a-00f000b-036-00b0007-006-002-01d-007-013-022-01400020008",
            INIT_31 => X"0007000d00080000-019-01c-0030011001300070019001b001d002000240005",
            INIT_32 => X"-003-00d-01b-014-0050012000900030005000f00180000001c002600180046",
            INIT_33 => X"0047002300220007-001000d-039-003-015-0290002-002-004000f-01a-01b",
            INIT_34 => X"-004-069-039000b-001-0190000-06a-044-030-060-031-019000e00230013",
            INIT_35 => X"000e000a-00f004100250023002700080027-0190013-011-036-016-00b0006",
            INIT_36 => X"00040005-008-00e-006-014000a-010-0010004-013-001001500240009-012",
            INIT_37 => X"001d000a001b0004000500130017-0070020-00d00000006-004000b000b0023",
            INIT_38 => X"000b00160005-027-01e-004-009-02e-01200060004-00c-011-00d000c-01d",
            INIT_39 => X"-018-01c000c-012-009-0260021-004-00c002c000f0000003a001b0003-013",
            INIT_3A => X"-003-016-021-003-0020004-0010009-004-00b-014-007-0110015000a000c",
            INIT_3B => X"0009001e0039001b00460045-008000e003f000b002300170006000b0001-01c",
            INIT_3C => X"-007000f00460026-01d-004-02c-050-02c-029-0360039000800120008-00c",
            INIT_3D => X"0003-012-013-013000c-00a0004-003-032-03f-018-048-039001b0027000c",
            INIT_3E => X"-00c-01b-01e-017-007-0240004001e0014-018000e-001-01a000d-02a000b",
            INIT_3F => X"00100012-00a00180010-013-006-016-00c-03c-03a-035-054-022000b-036",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY17;


    MEM_IWGHT_18K_LAYER2_ENTITY18 : if N_BRAM = 18 generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"-063001f0006001500120022001b-01300140012-0080008000c-00e00280016",
            INIT_01 => X"-0110016002d0006-0060005-007-003-00d0025-015-01b-00f0002-014-029",
            INIT_02 => X"-02b-01c-053-03c0016-020-02b-01d-011-013-02d001f-0020013002d0004",
            INIT_03 => X"-0090000-01d-02f-00c-02c-02b0002000b0000-02a000c-007-010000f001f",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => ADDR,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => REGCE, -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => WE       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_18K_LAYER2_ENTITY18;



end a1;