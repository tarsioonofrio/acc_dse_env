-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;


-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity gold_36k_layer2_entity1 is
    generic (
        DEVICE: string := "7SERIES"
        );

    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic_vector(2-1 downto 0);;
        DI   : in std_logic_vector(INPUT_SIZE-1 downto 0);
        ADDR : in std_logic_vector(11-1 downto 0);
        DO   : out std_logic_vector(INPUT_SIZE-1 downto 0)
    );
 end gold_36k_layer2_entity1;

  architecture a1 of bram is

    begin

    BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
    generic map (
       BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
       DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
       DO_REG => 0,                     -- Optional output register (0 or 1)
       INIT => X"000000000000000000",   -- Initial values on output port
       INIT_FILE => "NONE",
       WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       SRVAL => X"000000000000000000",  -- Set/Reset value for port output
       WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
       -- The following INIT_xx declarations specify the initial contents of the RAM
       INIT_00 => X"009c0000000000000000000000000000000000000000000000000000000f0071",
       INIT_01 => X"00000000000000000000002d00000000000a002b000000000072004f003200c7",
       INIT_02 => X"003a000000530000000001db01760128008300cc009e002c003f0104008c0000",
       INIT_03 => X"0000012900640000007b0000008a007e005c000a000000000000004300000051",
       INIT_04 => X"0000000000000021002b00000000017800f100010024008d0079004200580060",
       INIT_05 => X"0000000000000000000000000000000000000000000000000000000000030044",
       INIT_06 => X"000e00000096002b000000100008000000000000001f00000000000000000000",
       INIT_07 => X"000000000000000000000000000000000000000000000000000000000000003b",
       INIT_08 => X"00000000000000000050005a00f800620000000000e200000000000000000000",
       INIT_09 => X"00000000000000000000000000000000000000000000000000000051008700ae",
       INIT_0A => X"0000009000cf011a00e3010d00000000000000000091000000000052013800ae",
       INIT_0B => X"0047005000000197007c006a007f00f9002b00bc010100ef0000000000000098",
       INIT_0C => X"00e30000003d00210000017b010a003301c30162013b00890059013b00e70030",
       INIT_0D => X"01150113017f0000000000000000000000000063009b01320000000000000000",
       INIT_0E => X"00a50000000f0027000801aa00ca000001620000000000000000000001380164",
       INIT_0F => X"01580000009501920032002d015400420114007c0049015e00da012e0212026d",
       INIT_10 => X"003f000000000014000000000000007600000000000000000000000000000000",
       INIT_11 => X"0000000b00000009005500000036004900000000009c00000000000000000000",
       INIT_12 => X"00000000000000000000000000000000002b001c00000000000000aa010d0000",
       INIT_13 => X"00e000cf0074010e00b1004e0000000000000000000000000000000000710000",
       INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_15 => X"00000034006100590000006e017c00320000010000c500a001d300ee009c00e8",
       INIT_16 => X"0190014e007500ed006900ff00fc00e6002e005500de000000d4006501260084",
       INIT_17 => X"0094007b00520000000000000000000000000000000000000000000000540000",
       INIT_18 => X"000000000000003e0000000000080083004f000300000000004c007300000000",
       INIT_19 => X"0000001600000000008300800032000000000069000000f5007700bf00ad0078",
       INIT_1A => X"005a0079000000fb0011000000a900760037000000000000001a000000000000",
       INIT_1B => X"00000008000000000000000000000000000000000000005a002a000800070000",
       INIT_1C => X"001a00000000001b000000000044008d0000003e000000000000006000000000",
       INIT_1D => X"001000000000001f001b00660010004800000000000000000000000000000000",
       INIT_1E => X"000000970037003d0059014a00be0086007300e100000000000000000000001c",
       INIT_1F => X"00000000002e0000000000000000000000000000000000000000000000000000",
       INIT_20 => X"00000000000000000000002c002a00890048003700810039000100f800000000",
       INIT_21 => X"00000000000000000000000000000000003700000000003e0000003000000000",
       INIT_22 => X"00000000000000000000000000000000000000ee00d100b2015200d900ec001b",
       INIT_23 => X"008e009b00a600de006f0068000000420000000000000000000000000000000d",
       INIT_24 => X"00be0000003b00d300000000000000000000000000000000000000dd0151015c",
       INIT_25 => X"015600e600a90115009c0000000000000000000000000042000000000012010e",
       INIT_26 => X"00520078010f0000000000af0008002b00070000000000000000001700000055",
       INIT_27 => X"00b800000037000000000047000000390054000000000000000e003f00000000",
       INIT_28 => X"0000000000190000000000000000000000000000000000390047000000ad0075",
       INIT_29 => X"0000000c003f00f0000000000000000000000000000000000000000000f4010e",
       INIT_2A => X"019101530000000001a20166000000d100000017003b00000000000400150039",
       INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_2C => X"0000000000000000000000000000000000290000000000000000000000000000",
       INIT_2D => X"00000000000000000066000000000085003f0000000500a30000000000450000",
       INIT_2E => X"000000000060003c0000000000280005000000000000009200000000006d0000",
       INIT_2F => X"000000220095003e0000004a00a2000000000000000000000000000000000000",
       INIT_30 => X"0000000001110000003c00ab001600ce0000000000c7007f002b009600a50043",
       INIT_31 => X"00ba00dd001e0026015b00ab00d7003f000000f400da00000161015a013900f2",
       INIT_32 => X"00b2011b0190007b011400000000000000980000000000000044000000000000",
       INIT_33 => X"0000000000370000002300a60000000000000000000000000000000000000000",
       INIT_34 => X"007000a5010e00c6000000e000de0089008300190086007800a0005100540000",
       INIT_35 => X"0000000000000000000000000000003100000000000000000000000000000000",
       INIT_36 => X"000000000000000000e4011800cd002d00c40000003b00910096007d00000000",
       INIT_37 => X"0076002600000000000000000000000000560000000000d4003d0000002c0000",
       INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_39 => X"000000000048008a00be005d009700000056004e004d0003005c0000000100dd",
       INIT_3A => X"001a0000002a0020000000000055000000000000000000000000000000410000",
       INIT_3B => X"0000000000be002f002b000000000000001c0000000000000000000000000000",
       INIT_3C => X"00000026000000550000004900b00000000000000000001e0022003e00930025",
       INIT_3D => X"00340054003d004c00be0000000000290000006d000000000000000000000000",
       INIT_3E => X"000000000000000000000000000000000000000000000000002b0000000000df",
       INIT_3F => X"00000000005a000000cf00860000006d001e0000000000320000000000000000",

       -- The next set of INIT_xx are valid when configured as 36Kb
       INIT_40 => X"00000000000000000000000000000022004100000082002d004400ea010e0000",
       INIT_41 => X"000000000027002f000000000000000000000000000000000000000000000000",
       INIT_42 => X"000000cf008700a400de00c200bf00c300cc00e4000000000000000000030000",
       INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_44 => X"0000000000000000000000820070000000e4009d000000ae0073001000000000",
       INIT_45 => X"000000000000000000000000000000000000000000000000001b000000540000",
       INIT_46 => X"00000000000000000000000000000031007d00ed007e007201090000000000d3",
       INIT_47 => X"0023000000000000000000000000000000000000000000ca00b8009e00a60000",
       INIT_48 => X"003a00660000004e0092008f0083004e0006007c00db00b50136000000000000",
       INIT_49 => X"00000000000000000000004d0000000000000000000000000000000000000000",
       INIT_4A => X"0000000000000000000000000040000000bc00f8001500e40031000000000000",
       INIT_4B => X"00000000000000000000000000000000000000000000000000000000004900a5",
       INIT_4C => X"006500000000000000000000005c003400c4000000000000002d006900700000",
       INIT_4D => X"0000006400b50084006f00000000000000000000000000000000000000000000",
       INIT_4E => X"0000000000000000000000000000003b0000005c00c3000000bc00ae002a0078",
       INIT_4F => X"00000000000000000000000000000000004b0000000000000000000000000000",
       INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_51 => X"00000000000000000094006e00ae00b90077012c006e00bc0077000000000000",
       INIT_52 => X"00000000000000470000000000190000005d0082007e0070008200aa00e30000",
       INIT_53 => X"0000000000000000000000000000007000000000000000000000000000000000",
       INIT_54 => X"0000000000000000000000000000000000000000011500ae00e000fe01450116",
       INIT_55 => X"0059011c00f5000000000000000000000000000000000000005a0057003400bc",
       INIT_56 => X"00ac0096006400660034003200000000000000000000004e008000a7005e000b",
       INIT_57 => X"0000000000000000000000000000000000250000000000c10000000000400060",
       INIT_58 => X"004b004001080120000900e200d300570169016d0215000401b9000000000000",
       INIT_59 => X"01b701da000000000000007300410000008f00af000000000000000000000000",
       INIT_5A => X"0000000000000000037c02790120014900000000000000000000000000000000",
       INIT_5B => X"000000000000000000000000016000000000004b000000000000000000000000",
       INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_5D => X"000000000008009e013b01bf00eb003b000000be000000000000000000000134",
       INIT_5E => X"001e014200000000000000000000000000000000000000000000000000000000",
       INIT_5F => X"0000000000e3000000000000006900d100fe00eb000e00000000000000000000",
       INIT_60 => X"00000000016300cc016c00d000ca00b400730000000000000065002600940156",
       INIT_61 => X"00000000006c0000000000860000000000000000000000000000000000000000",
       INIT_62 => X"0000000000000000000000000000000000000000000001ec022f004200db0262",
       INIT_63 => X"005f009e008c000000c6017a00310027000d00000000006a0000001101b70000",
       INIT_64 => X"0170012000000000000000000051008c0148008200c400a400a1009701390000",
       INIT_65 => X"0000000000000000010000000000000000000000000000000000000000000000",
       INIT_66 => X"0000000000000062002900e6011c0109009f0000000000000000000000000000",
       INIT_67 => X"0000000002360000000000000000000000000000000000000000000000000000",
       INIT_68 => X"00000000000000000000008400aa00330040000000000000004600f500000000",
       INIT_69 => X"0000000000000000000000000000000000c80000019401f9008a000000000000",
       INIT_6A => X"028f026b016a01d2035600000127000000260000000000000000000000000000",
       INIT_6B => X"00000000000000000000000000000000008e020000d80135002a000000000000",
       INIT_6C => X"00000008000000000000000000fb000000000000000000000000000000000000",
       INIT_6D => X"0000008701cf003f0124000000110000000000f401120000012d000000590000",
       INIT_6E => X"004f00880084000000bc0000000000c7011501c9008201bf009a000000000046",
       INIT_6F => X"0000000000000000000000000089000001790000000000000000000000000028",
       INIT_70 => X"00d701ba019b00a602a201a8037400b301c70026027b02310064005e007a0053",
       INIT_71 => X"005a00d700ca0000000000000000000000000000000000000000000000000000",
       INIT_72 => X"000000000000000000000000001a009c00000000002b00780051000000b1009d",
       INIT_73 => X"00bb000000000000000000000000000000000000000000000000000000000078",
       INIT_74 => X"0000005000000000000000000000000000000000000000000000000000000000",
       INIT_75 => X"000000000000000000ce005901270017000000b3000000000037000000000000",
       INIT_76 => X"0000000000000000000000000224007f004000f3007200000175016801980000",
       INIT_77 => X"001100000000011e0000004501030000000000000000000000b5000000000078",
       INIT_78 => X"000000000000000000000000000000000000000002c801de0134012c02670182",
       INIT_79 => X"0154013801650000000000000000000000000000000000ad0000000000000010",
       INIT_7A => X"0000000000590000000000c3000000000000000000c1000000000010001a0153",
       INIT_7B => X"000000200000000000000000000001a501d1008901a00096000400af01340000",
       INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_7D => X"000000000033007500000000006f00000000002e000000000000000000000000",
       INIT_7E => X"000000000000000000000000000000000000001e00000029002a017e01b50155",
       INIT_7F => X"00bd016801ea0081018f01e80000006f000000000016009100f100d3003d0000",

       -- The next set of INITP_xx are for the parity bits
       INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

       -- The next set of INIT_xx are valid when configured as 36Kb
       INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000")
    port map (
       DO => DO,      -- Output data, width defined by READ_WIDTH parameter
       ADDR => ADDR,  -- Input address, width defined by read/write port depth
       CLK => CLK,    -- 1-bit input clock
       DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
       EN => EN,      -- 1-bit input RAM enable
       REGCE => REGCE, -- 1-bit input output register enable
       RST => RST,    -- 1-bit input reset
       WE => WE       -- Input write enable, width defined by write port depth
    );


-- End of BRAM_SINGLE_MACRO_inst instantiation
