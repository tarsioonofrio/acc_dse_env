library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    0, 0, 0, 108, 141, 68, 56, 
    59, 36, 110, 20, 0, 14, 48, 
    27, 93, 79, 0, 0, 38, 0, 
    50, 65, 0, 126, 26, 34, 0, 
    10, 18, 95, 0, 85, 134, 0, 
    29, 0, 212, 145, 8, 0, 0, 
    76, 130, 32, 0, 0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 0, 0, 11, 0, 
    0, 0, 0, 78, 0, 0, 166, 
    0, 99, 0, 45, 0, 134, 0, 
    0, 63, 0, 0, 0, 161, 0, 
    0, 0, 100, 0, 0, 38, 0, 
    0, 0, 181, 0, 48, 0, 0, 
    199, 0, 59, 4, 0, 0, 0, 
    
    -- channel=2
    72, 84, 56, 53, 0, 43, 49, 
    64, 86, 57, 64, 31, 58, 57, 
    48, 98, 0, 43, 26, 53, 13, 
    26, 35, 0, 0, 58, 37, 48, 
    8, 71, 109, 35, 0, 0, 28, 
    0, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    56, 81, 5, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 57, 0, 0, 0, 0, 0, 
    0, 0, 36, 3, 38, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    31, 0, 0, 0, 0, 0, 0, 
    0, 105, 0, 0, 0, 0, 0, 
    
    -- channel=4
    6, 1, 11, 32, 3, 0, 0, 
    67, 17, 0, 57, 71, 40, 5, 
    52, 19, 0, 45, 159, 50, 17, 
    29, 0, 1, 34, 42, 4, 16, 
    0, 125, 6, 0, 1, 0, 0, 
    0, 54, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    5, 0, 0, 0, 13, 0, 9, 
    39, 23, 0, 0, 0, 0, 66, 
    0, 110, 0, 0, 0, 0, 0, 
    0, 82, 0, 0, 0, 0, 0, 
    0, 0, 48, 0, 0, 104, 0, 
    0, 0, 0, 0, 56, 41, 0, 
    45, 0, 19, 0, 0, 0, 0, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 20, 
    113, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 0, 0, 0, 
    33, 0, 0, 92, 285, 345, 351, 
    204, 0, 227, 327, 367, 390, 383, 
    
    -- channel=7
    114, 0, 138, 79, 0, 0, 26, 
    0, 0, 0, 0, 32, 0, 0, 
    0, 0, 0, 0, 43, 0, 0, 
    0, 0, 75, 0, 31, 68, 3, 
    0, 0, 0, 0, 0, 0, 39, 
    0, 40, 76, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=8
    221, 221, 205, 297, 177, 123, 183, 
    95, 288, 121, 0, 0, 0, 0, 
    0, 135, 0, 0, 0, 0, 0, 
    0, 136, 8, 0, 0, 0, 0, 
    0, 0, 3, 0, 63, 92, 209, 
    0, 0, 0, 27, 37, 57, 17, 
    58, 0, 0, 13, 33, 20, 17, 
    
    -- channel=9
    0, 0, 12, 0, 0, 21, 0, 
    0, 0, 0, 47, 0, 62, 0, 
    203, 0, 104, 256, 0, 86, 179, 
    327, 26, 0, 56, 0, 62, 0, 
    224, 109, 0, 187, 0, 0, 0, 
    0, 0, 0, 0, 77, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 
    
    -- channel=10
    52, 27, 94, 62, 134, 116, 85, 
    115, 84, 165, 84, 34, 16, 54, 
    94, 47, 211, 92, 49, 59, 94, 
    95, 106, 25, 17, 0, 22, 0, 
    10, 52, 136, 153, 92, 116, 133, 
    93, 33, 253, 87, 92, 126, 63, 
    0, 142, 0, 0, 0, 0, 0, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 
    14, 0, 74, 0, 0, 24, 0, 
    0, 0, 0, 71, 0, 0, 56, 
    0, 0, 0, 0, 0, 0, 9, 
    0, 60, 121, 0, 0, 80, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 
    
    -- channel=12
    208, 213, 198, 120, 54, 46, 117, 
    118, 173, 120, 75, 67, 49, 44, 
    0, 120, 54, 66, 100, 45, 20, 
    0, 58, 62, 13, 45, 29, 60, 
    0, 42, 22, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=13
    0, 0, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 97, 0, 0, 
    0, 42, 0, 0, 194, 0, 0, 
    0, 0, 197, 0, 88, 0, 10, 
    0, 0, 0, 84, 0, 0, 141, 
    1, 294, 0, 0, 0, 97, 8, 
    0, 0, 23, 0, 57, 18, 105, 
    
    -- channel=14
    0, 0, 0, 0, 0, 26, 0, 
    71, 0, 70, 34, 0, 72, 0, 
    0, 0, 0, 189, 0, 75, 0, 
    72, 0, 0, 42, 0, 1, 0, 
    72, 109, 126, 0, 0, 0, 0, 
    0, 0, 107, 0, 0, 0, 0, 
    0, 0, 0, 50, 31, 10, 53, 
    
    -- channel=15
    0, 0, 0, 0, 5, 12, 27, 
    47, 0, 0, 0, 11, 0, 0, 
    0, 0, 0, 0, 36, 0, 0, 
    0, 0, 59, 0, 0, 0, 0, 
    0, 0, 0, 0, 31, 89, 67, 
    205, 0, 86, 113, 11, 17, 34, 
    80, 147, 80, 33, 13, 40, 30, 
    
    -- channel=16
    22, 90, 0, 0, 0, 0, 10, 
    0, 29, 0, 0, 20, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 82, 
    27, 0, 0, 0, 0, 0, 90, 
    0, 0, 0, 0, 53, 135, 76, 
    0, 0, 0, 91, 129, 104, 57, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 
    0, 36, 38, 0, 2, 0, 0, 
    0, 0, 0, 0, 20, 0, 5, 
    10, 39, 18, 0, 0, 0, 0, 
    0, 48, 46, 0, 0, 40, 2, 
    0, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 5, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=19
    177, 162, 188, 215, 121, 92, 114, 
    75, 185, 141, 71, 0, 0, 12, 
    0, 0, 0, 19, 0, 9, 0, 
    0, 49, 0, 0, 0, 6, 0, 
    0, 0, 18, 0, 30, 22, 5, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=20
    90, 123, 85, 16, 0, 0, 0, 
    0, 57, 0, 0, 50, 0, 0, 
    0, 5, 0, 0, 74, 0, 0, 
    0, 0, 13, 0, 55, 0, 12, 
    0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 52, 0, 0, 
    0, 0, 0, 0, 82, 0, 0, 
    0, 0, 67, 0, 81, 0, 24, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    155, 0, 51, 81, 85, 122, 106, 
    
    -- channel=22
    37, 22, 6, 118, 22, 51, 26, 
    49, 88, 85, 89, 0, 85, 0, 
    139, 26, 34, 145, 4, 147, 0, 
    164, 133, 70, 122, 0, 49, 0, 
    104, 84, 108, 18, 103, 0, 0, 
    0, 46, 120, 0, 17, 0, 12, 
    0, 18, 54, 29, 5, 16, 0, 
    
    -- channel=23
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 14, 17, 20, 
    65, 0, 0, 0, 9, 0, 16, 
    51, 0, 0, 0, 66, 0, 14, 
    87, 37, 123, 48, 38, 45, 27, 
    186, 138, 28, 154, 182, 265, 273, 
    345, 103, 155, 232, 264, 282, 314, 
    
    -- channel=24
    64, 80, 53, 29, 22, 54, 40, 
    10, 36, 0, 0, 14, 0, 33, 
    0, 11, 0, 0, 0, 0, 0, 
    4, 21, 49, 0, 19, 0, 47, 
    0, 0, 0, 23, 0, 0, 54, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 14, 
    54, 0, 0, 0, 147, 96, 86, 
    0, 0, 113, 0, 0, 0, 0, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=28
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=29
    196, 234, 131, 69, 0, 0, 62, 
    18, 126, 37, 13, 22, 78, 20, 
    0, 167, 116, 70, 0, 52, 5, 
    0, 16, 7, 27, 6, 30, 100, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=30
    89, 207, 84, 91, 0, 0, 5, 
    0, 104, 0, 0, 0, 39, 0, 
    0, 0, 0, 83, 0, 28, 5, 
    49, 0, 0, 0, 0, 0, 7, 
    111, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    0, 0, 41, 86, 0, 91, 0, 
    100, 4, 138, 103, 0, 35, 87, 
    0, 96, 0, 141, 41, 59, 6, 
    111, 109, 0, 0, 0, 26, 0, 
    0, 98, 137, 21, 103, 0, 0, 
    0, 0, 30, 0, 0, 0, 0, 
    39, 0, 0, 0, 0, 0, 0, 
    
    -- channel=32
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 50, 0, 0, 
    0, 0, 0, 0, 29, 0, 0, 
    0, 0, 58, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 166, 78, 
    48, 0, 0, 55, 120, 123, 101, 
    
    -- channel=33
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 42, 0, 3, 68, 56, 
    154, 0, 81, 143, 160, 213, 208, 
    316, 88, 172, 177, 195, 208, 212, 
    
    -- channel=34
    97, 37, 97, 137, 74, 55, 101, 
    42, 53, 43, 1, 4, 0, 50, 
    33, 150, 156, 0, 0, 14, 7, 
    5, 98, 111, 64, 37, 81, 15, 
    0, 0, 0, 0, 91, 65, 19, 
    162, 21, 186, 89, 0, 0, 0, 
    34, 239, 14, 0, 0, 0, 0, 
    
    -- channel=35
    0, 0, 0, 12, 0, 45, 0, 
    312, 0, 100, 100, 129, 112, 208, 
    75, 393, 0, 9, 301, 99, 0, 
    0, 0, 0, 11, 342, 3, 0, 
    0, 259, 421, 0, 17, 0, 0, 
    0, 118, 64, 0, 0, 0, 0, 
    193, 0, 41, 0, 0, 0, 0, 
    
    -- channel=36
    136, 154, 128, 130, 52, 27, 80, 
    50, 134, 41, 52, 0, 41, 51, 
    40, 191, 56, 61, 0, 59, 6, 
    4, 65, 14, 76, 51, 99, 26, 
    0, 4, 0, 0, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=37
    0, 0, 0, 82, 0, 0, 60, 
    0, 0, 0, 0, 44, 0, 0, 
    63, 101, 42, 0, 10, 22, 0, 
    0, 0, 121, 50, 26, 0, 0, 
    0, 0, 0, 0, 106, 0, 69, 
    155, 16, 174, 85, 0, 0, 0, 
    0, 112, 0, 0, 0, 0, 0, 
    
    -- channel=38
    0, 0, 0, 40, 0, 58, 0, 
    38, 0, 0, 142, 0, 122, 92, 
    104, 0, 0, 206, 0, 261, 45, 
    134, 107, 0, 138, 0, 172, 0, 
    0, 0, 139, 4, 36, 45, 0, 
    0, 0, 253, 0, 72, 0, 1, 
    8, 0, 36, 43, 11, 9, 0, 
    
    -- channel=39
    0, 0, 0, 63, 92, 0, 23, 
    0, 27, 93, 69, 0, 31, 57, 
    0, 72, 0, 52, 0, 151, 36, 
    49, 80, 0, 140, 0, 98, 0, 
    0, 54, 204, 0, 79, 133, 0, 
    0, 0, 129, 43, 0, 0, 0, 
    0, 143, 0, 0, 0, 0, 0, 
    
    -- channel=40
    6, 58, 0, 115, 0, 12, 12, 
    17, 12, 36, 115, 0, 155, 3, 
    223, 0, 0, 174, 0, 193, 8, 
    197, 34, 0, 179, 0, 97, 0, 
    127, 80, 92, 0, 39, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=41
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    61, 0, 0, 0, 30, 6, 0, 
    93, 81, 62, 32, 0, 23, 0, 
    112, 136, 146, 152, 179, 169, 193, 
    203, 167, 239, 155, 173, 194, 208, 
    
    -- channel=42
    31, 34, 0, 0, 0, 0, 21, 
    0, 48, 0, 0, 69, 34, 57, 
    207, 126, 61, 9, 34, 89, 41, 
    147, 139, 25, 34, 52, 81, 104, 
    63, 80, 20, 77, 0, 0, 17, 
    47, 30, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=43
    0, 64, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 74, 46, 
    0, 0, 0, 50, 66, 43, 0, 
    
    -- channel=44
    21, 27, 7, 21, 21, 60, 31, 
    33, 0, 31, 55, 12, 74, 73, 
    16, 22, 0, 40, 0, 71, 63, 
    10, 6, 0, 68, 0, 32, 54, 
    0, 20, 77, 0, 51, 59, 31, 
    0, 0, 118, 58, 38, 37, 38, 
    19, 0, 16, 16, 2, 4, 0, 
    
    -- channel=45
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 104, 13, 101, 129, 
    187, 0, 0, 175, 169, 199, 188, 
    
    -- channel=46
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 67, 
    0, 0, 0, 0, 0, 96, 130, 
    133, 230, 0, 0, 0, 117, 0, 
    0, 0, 0, 204, 17, 79, 0, 
    0, 0, 0, 0, 13, 7, 0, 
    118, 150, 0, 10, 5, 0, 0, 
    
    -- channel=47
    48, 27, 0, 0, 0, 6, 30, 
    7, 12, 0, 0, 27, 24, 6, 
    0, 0, 0, 0, 3, 0, 7, 
    0, 0, 0, 40, 33, 47, 58, 
    63, 58, 0, 0, 50, 58, 101, 
    126, 13, 44, 90, 88, 83, 118, 
    154, 174, 152, 137, 125, 150, 160, 
    
    -- channel=48
    104, 92, 106, 105, 75, 45, 80, 
    53, 129, 84, 66, 35, 29, 33, 
    20, 107, 36, 69, 52, 49, 10, 
    19, 95, 11, 26, 29, 40, 8, 
    0, 40, 17, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=49
    0, 0, 0, 21, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 54, 0, 
    0, 0, 0, 68, 0, 56, 0, 
    0, 0, 0, 0, 86, 153, 0, 
    195, 0, 277, 327, 163, 122, 189, 
    114, 426, 156, 172, 120, 218, 55, 
    
    -- channel=50
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 19, 0, 0, 
    0, 0, 30, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    34, 0, 0, 0, 0, 0, 0, 
    272, 87, 74, 193, 0, 47, 79, 
    95, 269, 56, 76, 67, 109, 96, 
    
    -- channel=51
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 78, 0, 0, 0, 0, 
    
    -- channel=52
    0, 0, 45, 0, 0, 24, 0, 
    30, 24, 53, 61, 0, 41, 0, 
    0, 0, 56, 129, 0, 0, 22, 
    0, 0, 0, 0, 0, 37, 0, 
    0, 85, 92, 104, 0, 28, 50, 
    0, 80, 71, 0, 31, 63, 31, 
    0, 0, 29, 20, 20, 0, 53, 
    
    -- channel=53
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 32, 0, 65, 11, 39, 
    87, 0, 164, 123, 105, 136, 117, 
    166, 114, 107, 91, 118, 139, 161, 
    
    -- channel=54
    0, 27, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 
    
    -- channel=55
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 61, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=56
    0, 0, 37, 69, 3, 32, 0, 
    0, 4, 46, 121, 34, 103, 63, 
    212, 143, 103, 132, 68, 155, 68, 
    255, 115, 132, 84, 83, 115, 8, 
    167, 137, 177, 153, 127, 0, 24, 
    95, 266, 105, 33, 52, 18, 40, 
    18, 225, 43, 0, 1, 0, 25, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 63, 32, 
    108, 0, 0, 33, 51, 37, 71, 
    
    -- channel=58
    0, 0, 0, 0, 164, 0, 24, 
    361, 210, 98, 0, 215, 0, 0, 
    0, 0, 125, 28, 440, 0, 13, 
    0, 0, 0, 0, 0, 0, 27, 
    41, 552, 157, 0, 0, 126, 0, 
    0, 0, 71, 0, 66, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=59
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 
    180, 0, 190, 31, 0, 43, 22, 
    98, 0, 0, 41, 0, 16, 4, 
    74, 0, 0, 9, 10, 0, 0, 
    140, 22, 312, 102, 116, 132, 108, 
    63, 146, 122, 88, 90, 122, 89, 
    
    -- channel=60
    38, 0, 120, 1, 113, 0, 51, 
    106, 163, 44, 0, 215, 0, 0, 
    231, 0, 128, 0, 339, 0, 89, 
    325, 147, 335, 0, 0, 0, 109, 
    289, 308, 0, 103, 101, 0, 166, 
    208, 308, 0, 81, 0, 0, 26, 
    0, 263, 0, 1, 23, 15, 76, 
    
    -- channel=61
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 81, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=62
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=63
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 156, 8, 0, 0, 0, 
    81, 0, 0, 0, 0, 0, 0, 
    128, 157, 0, 54, 0, 0, 0, 
    0, 219, 0, 38, 47, 61, 94, 
    
    
    others => 0);
end ifmap_package;
