library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    517, 513, 519, 522, 520, 524, 525, 532, 531, 513, 504, 510, 529, 552, 559, 562, 548, 524, 502, 487, 478, 476, 480, 489, 494, 512, 529, 546, 553, 550, 
    537, 530, 535, 530, 523, 523, 526, 532, 523, 479, 469, 496, 522, 541, 540, 529, 521, 489, 453, 428, 425, 434, 446, 461, 468, 485, 510, 534, 545, 545, 
    534, 530, 540, 537, 528, 525, 530, 532, 513, 404, 393, 448, 489, 499, 500, 500, 485, 430, 377, 340, 336, 352, 389, 411, 432, 455, 478, 502, 525, 537, 
    504, 493, 510, 528, 531, 532, 539, 540, 521, 394, 373, 413, 462, 482, 475, 470, 449, 362, 294, 248, 248, 279, 316, 350, 397, 430, 446, 460, 494, 521, 
    483, 470, 473, 504, 530, 541, 544, 548, 536, 434, 423, 417, 435, 456, 445, 443, 398, 298, 226, 206, 225, 251, 274, 304, 364, 411, 430, 430, 467, 505, 
    453, 444, 438, 473, 524, 546, 543, 540, 535, 500, 461, 403, 395, 414, 386, 374, 350, 270, 196, 198, 248, 278, 278, 307, 362, 405, 422, 417, 445, 488, 
    412, 374, 367, 429, 506, 536, 522, 493, 496, 473, 403, 328, 319, 348, 336, 330, 330, 290, 219, 210, 265, 305, 315, 332, 359, 397, 432, 428, 430, 468, 
    305, 257, 266, 369, 479, 515, 442, 344, 334, 346, 293, 245, 258, 309, 322, 328, 346, 334, 253, 226, 253, 296, 334, 343, 355, 373, 425, 449, 435, 446, 
    195, 123, 171, 318, 448, 502, 351, 170, 140, 190, 181, 190, 231, 285, 325, 336, 372, 366, 249, 206, 210, 273, 324, 324, 333, 350, 401, 448, 442, 441, 
    124, 54, 98, 279, 423, 505, 351, 116, 28, 107, 130, 155, 213, 271, 313, 333, 399, 343, 184, 158, 164, 251, 310, 310, 306, 321, 363, 420, 430, 441, 
    97, 32, 69, 251, 401, 508, 428, 202, 96, 145, 144, 120, 181, 244, 297, 299, 391, 287, 118, 114, 146, 255, 307, 307, 301, 310, 329, 369, 392, 438, 
    95, 22, 86, 246, 379, 486, 520, 312, 209, 190, 161, 81, 127, 205, 258, 270, 358, 225, 83, 102, 165, 271, 313, 323, 311, 304, 297, 325, 349, 429, 
    83, 14, 108, 251, 358, 449, 536, 387, 289, 197, 137, 65, 100, 157, 204, 246, 333, 189, 83, 107, 175, 255, 302, 316, 310, 290, 269, 295, 337, 418, 
    54, 10, 111, 241, 311, 385, 491, 404, 314, 137, 47, 46, 105, 154, 199, 249, 318, 206, 116, 126, 188, 260, 307, 310, 295, 265, 257, 305, 361, 426, 
    26, 0, 66, 211, 244, 294, 390, 402, 310, 126, 42, 85, 159, 206, 233, 274, 325, 243, 194, 184, 200, 252, 314, 313, 286, 266, 282, 349, 404, 452, 
    0, 0, 5, 166, 201, 212, 269, 351, 306, 187, 120, 180, 236, 266, 286, 284, 296, 288, 317, 260, 235, 284, 345, 349, 321, 297, 321, 382, 422, 463, 
    0, 0, 0, 111, 176, 166, 179, 283, 285, 296, 247, 258, 293, 272, 294, 281, 258, 281, 351, 316, 297, 328, 381, 385, 371, 351, 378, 414, 449, 481, 
    0, 0, 0, 66, 175, 151, 152, 193, 227, 331, 299, 297, 277, 209, 245, 269, 232, 270, 319, 315, 345, 388, 415, 381, 375, 362, 402, 433, 467, 493, 
    0, 0, 0, 43, 162, 141, 105, 141, 210, 319, 290, 283, 198, 120, 165, 233, 250, 289, 307, 336, 379, 408, 408, 344, 340, 334, 392, 438, 461, 473, 
    3, 0, 0, 50, 168, 128, 26, 26, 121, 237, 211, 183, 83, 18, 61, 163, 221, 300, 342, 362, 360, 351, 326, 271, 251, 246, 286, 325, 340, 345, 
    0, 0, 0, 55, 160, 77, 0, 0, 0, 99, 125, 75, 7, 0, 18, 109, 184, 263, 314, 312, 280, 256, 213, 188, 165, 149, 156, 186, 193, 197, 
    0, 0, 0, 29, 111, 0, 0, 0, 0, 36, 73, 65, 47, 48, 62, 106, 141, 199, 217, 200, 169, 147, 123, 104, 86, 73, 66, 84, 89, 89, 
    0, 0, 0, 10, 43, 0, 0, 0, 0, 71, 106, 118, 121, 124, 128, 140, 141, 151, 143, 123, 107, 98, 82, 63, 51, 42, 40, 50, 50, 47, 
    0, 0, 0, 4, 0, 0, 0, 0, 66, 116, 127, 132, 135, 144, 143, 141, 138, 134, 120, 99, 85, 74, 56, 34, 30, 31, 32, 30, 15, 0, 
    24, 19, 3, 25, 0, 0, 0, 46, 112, 117, 103, 108, 115, 123, 129, 134, 131, 123, 107, 85, 62, 41, 28, 19, 21, 27, 12, 0, 0, 0, 
    15, 38, 42, 37, 0, 0, 0, 93, 122, 115, 91, 100, 115, 122, 124, 124, 116, 103, 84, 66, 44, 18, 6, 14, 27, 21, 0, 0, 0, 0, 
    5, 29, 48, 38, 0, 0, 0, 96, 118, 104, 81, 90, 101, 114, 120, 117, 101, 84, 67, 54, 36, 20, 19, 27, 28, 0, 0, 0, 0, 0, 
    4, 17, 32, 44, 0, 0, 49, 107, 131, 114, 84, 79, 81, 96, 104, 101, 87, 73, 59, 54, 50, 46, 43, 30, 5, 0, 0, 0, 36, 53, 
    7, 20, 28, 43, 51, 34, 110, 135, 151, 134, 112, 100, 90, 96, 96, 91, 72, 51, 43, 52, 61, 69, 57, 18, 0, 0, 0, 0, 61, 78, 
    17, 35, 45, 46, 74, 94, 126, 154, 165, 152, 143, 131, 128, 134, 123, 103, 73, 40, 31, 50, 69, 86, 60, 3, 0, 0, 0, 12, 59, 92, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 76, 80, 63, 48, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 35, 0, 0, 0, 0, 0, 0, 0, 76, 148, 165, 134, 89, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    159, 126, 76, 55, 34, 0, 0, 0, 0, 19, 66, 73, 34, 0, 0, 0, 0, 0, 0, 0, 0, 25, 40, 37, 20, 7, 5, 0, 0, 0, 
    203, 88, 55, 97, 107, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 48, 61, 62, 56, 31, 1, 0, 0, 0, 0, 
    159, 0, 0, 29, 49, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 31, 45, 51, 52, 49, 39, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 33, 33, 41, 61, 90, 99, 98, 100, 95, 81, 68, 54, 
    189, 170, 154, 137, 123, 109, 101, 90, 79, 62, 38, 13, 11, 18, 29, 28, 40, 66, 86, 100, 114, 126, 138, 135, 120, 115, 114, 104, 91, 70, 
    378, 351, 317, 306, 309, 309, 306, 299, 290, 271, 232, 187, 156, 143, 135, 129, 137, 154, 170, 183, 187, 187, 181, 162, 136, 129, 135, 129, 113, 81, 
    471, 447, 384, 366, 392, 422, 443, 456, 463, 455, 410, 329, 286, 274, 266, 254, 253, 256, 257, 250, 235, 212, 179, 150, 138, 148, 155, 146, 124, 76, 
    502, 481, 405, 374, 397, 442, 481, 514, 533, 538, 502, 359, 256, 240, 256, 262, 263, 257, 251, 236, 215, 193, 174, 170, 170, 176, 175, 152, 110, 42, 
    532, 523, 458, 427, 436, 471, 505, 533, 549, 555, 534, 372, 213, 163, 188, 215, 222, 227, 231, 232, 234, 232, 228, 231, 227, 214, 183, 132, 72, 1, 
    544, 556, 526, 507, 509, 524, 542, 556, 562, 564, 559, 431, 270, 226, 258, 286, 291, 302, 315, 324, 327, 322, 309, 290, 253, 208, 157, 94, 31, 0, 
    524, 560, 562, 554, 554, 560, 567, 569, 570, 569, 571, 517, 395, 379, 428, 458, 463, 461, 451, 435, 412, 372, 319, 268, 223, 182, 133, 64, 4, 0, 
    500, 554, 570, 567, 563, 566, 568, 571, 572, 571, 571, 558, 483, 485, 558, 597, 588, 539, 484, 429, 375, 313, 257, 222, 196, 164, 116, 50, 0, 0, 
    483, 546, 570, 569, 565, 565, 566, 569, 571, 570, 567, 561, 512, 511, 568, 584, 551, 479, 403, 337, 285, 247, 221, 200, 176, 144, 98, 37, 0, 0, 
    471, 531, 556, 557, 555, 553, 554, 557, 558, 557, 550, 543, 510, 496, 513, 494, 445, 381, 321, 277, 248, 226, 207, 184, 156, 122, 78, 22, 0, 0, 
    447, 499, 519, 523, 522, 517, 516, 516, 513, 509, 502, 495, 473, 449, 430, 389, 346, 316, 285, 264, 244, 220, 196, 169, 141, 106, 63, 11, 0, 0, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 95, 95, 50, 29, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 55, 84, 140, 145, 130, 159, 137, 64, 0, 0, 0, 0, 0, 0, 
    54, 107, 74, 60, 56, 44, 27, 18, 29, 22, 7, 3, 3, 0, 22, 69, 108, 126, 146, 155, 161, 210, 189, 135, 71, 27, 62, 104, 70, 80, 
    149, 178, 158, 146, 154, 137, 126, 113, 117, 109, 91, 83, 54, 29, 64, 96, 109, 114, 131, 143, 136, 167, 156, 163, 115, 69, 134, 187, 163, 161, 
    201, 210, 183, 169, 181, 194, 186, 155, 155, 151, 128, 101, 63, 48, 70, 97, 110, 120, 140, 157, 124, 98, 71, 127, 144, 82, 142, 201, 212, 201, 
    184, 198, 162, 145, 168, 190, 165, 115, 106, 111, 99, 66, 39, 46, 73, 100, 115, 120, 132, 143, 77, 25, 4, 56, 140, 83, 122, 197, 230, 211, 
    144, 167, 144, 155, 172, 179, 137, 78, 52, 52, 48, 24, 16, 34, 60, 83, 94, 87, 90, 86, 16, 0, 0, 0, 110, 104, 117, 218, 256, 242, 
    120, 154, 155, 175, 183, 156, 95, 45, 11, 4, 0, 0, 0, 1, 10, 17, 23, 19, 31, 28, 0, 0, 0, 5, 78, 140, 162, 269, 291, 283, 
    92, 117, 124, 126, 109, 76, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 30, 25, 30, 27, 38, 58, 158, 211, 291, 311, 304, 
    44, 48, 52, 38, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 82, 81, 71, 54, 54, 47, 137, 196, 205, 233, 263, 
    0, 0, 14, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 105, 97, 78, 56, 51, 39, 93, 127, 112, 136, 176, 
    11, 23, 35, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 53, 61, 49, 44, 35, 37, 33, 65, 80, 82, 110, 126, 
    56, 53, 38, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 8, 5, 9, 19, 34, 53, 88, 121, 162, 172, 128, 
    61, 42, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 14, 0, 0, 0, 0, 5, 38, 73, 107, 149, 198, 235, 237, 196, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 94, 132, 79, 19, 2, 10, 27, 52, 95, 134, 177, 222, 257, 273, 287, 287, 
    0, 0, 0, 0, 0, 0, 16, 16, 16, 0, 0, 0, 33, 119, 172, 197, 129, 71, 55, 67, 92, 122, 167, 205, 238, 271, 291, 299, 333, 373, 
    0, 0, 0, 0, 12, 57, 89, 95, 99, 51, 0, 0, 53, 133, 178, 202, 158, 127, 126, 140, 167, 198, 232, 254, 281, 306, 319, 335, 379, 419, 
    31, 6, 0, 0, 55, 112, 139, 139, 129, 76, 41, 44, 95, 145, 168, 184, 176, 177, 189, 212, 232, 246, 264, 285, 316, 334, 348, 375, 408, 429, 
    58, 35, 24, 27, 82, 128, 148, 153, 152, 130, 123, 136, 161, 183, 193, 205, 210, 219, 234, 255, 273, 291, 293, 305, 337, 357, 373, 391, 407, 418, 
    112, 98, 97, 106, 143, 167, 177, 187, 194, 203, 216, 226, 233, 233, 235, 246, 252, 255, 270, 294, 312, 322, 312, 328, 358, 375, 386, 394, 399, 404, 
    216, 215, 217, 227, 242, 249, 248, 255, 265, 275, 279, 278, 271, 268, 275, 287, 280, 283, 302, 319, 333, 345, 346, 361, 380, 388, 390, 392, 392, 403, 
    334, 339, 338, 335, 335, 330, 319, 312, 310, 311, 310, 308, 302, 304, 319, 323, 286, 284, 312, 337, 354, 367, 374, 385, 390, 391, 391, 389, 397, 427, 
    402, 404, 397, 386, 377, 369, 357, 346, 339, 336, 334, 332, 326, 328, 347, 338, 279, 290, 330, 358, 374, 383, 392, 396, 394, 391, 388, 388, 424, 471, 
    418, 417, 410, 396, 387, 379, 372, 363, 353, 347, 341, 338, 334, 343, 372, 365, 302, 315, 350, 374, 387, 396, 402, 402, 398, 392, 385, 403, 465, 513, 
    412, 407, 399, 389, 381, 375, 369, 363, 356, 356, 358, 365, 376, 395, 429, 418, 346, 345, 367, 389, 402, 405, 409, 407, 405, 393, 394, 439, 504, 539, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 46, 51, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 85, 117, 93, 72, 65, 68, 83, 78, 66, 61, 59, 55, 46, 37, 44, 57, 12, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 78, 112, 116, 123, 119, 121, 136, 132, 111, 92, 87, 75, 68, 68, 68, 77, 23, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 84, 100, 93, 102, 104, 115, 138, 139, 107, 79, 59, 47, 53, 55, 53, 51, 20, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 81, 147, 145, 97, 85, 79, 101, 126, 130, 96, 78, 57, 45, 70, 74, 68, 40, 42, 25, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 70, 128, 123, 77, 63, 57, 73, 84, 86, 71, 71, 51, 49, 82, 83, 82, 41, 48, 41, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 25, 32, 18, 15, 9, 18, 12, 10, 7, 10, 0, 5, 37, 40, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 71, 117, 106, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 91, 165, 177, 111, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 76, 195, 218, 155, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 117, 238, 252, 210, 147, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 49, 220, 287, 304, 279, 227, 164, 102, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 30, 231, 312, 345, 340, 319, 286, 250, 214, 174, 134, 103, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 68, 260, 354, 382, 359, 344, 332, 323, 314, 296, 280, 275, 243, 173, 113, 71, 26, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 93, 224, 320, 381, 376, 366, 327, 272, 249, 264, 318, 333, 314, 287, 271, 247, 163, 69, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 16, 73, 149, 230, 260, 273, 227, 144, 91, 94, 174, 202, 195, 187, 216, 229, 156, 64, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 90, 111, 70, 0, 0, 0, 23, 28, 22, 23, 44, 56, 12, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 17, 50, 56, 57, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    97, 66, 73, 84, 88, 95, 104, 110, 111, 119, 122, 121, 113, 94, 70, 60, 56, 49, 48, 49, 48, 40, 29, 27, 25, 26, 30, 38, 40, 70, 
    183, 156, 157, 166, 172, 183, 198, 208, 215, 221, 224, 223, 215, 199, 179, 175, 185, 192, 195, 195, 198, 196, 191, 186, 181, 180, 190, 207, 211, 211, 
    261, 233, 234, 235, 237, 249, 260, 270, 286, 296, 297, 295, 292, 292, 285, 287, 299, 312, 320, 323, 324, 321, 320, 319, 318, 318, 332, 340, 307, 270, 
    337, 320, 323, 328, 334, 344, 349, 359, 372, 376, 375, 371, 370, 373, 371, 372, 379, 390, 399, 402, 401, 399, 398, 397, 397, 396, 386, 352, 291, 264, 
    395, 384, 385, 384, 389, 394, 393, 401, 410, 413, 405, 398, 401, 404, 401, 397, 400, 406, 410, 410, 408, 407, 409, 410, 404, 372, 319, 273, 245, 268, 
    401, 391, 388, 387, 388, 389, 391, 397, 401, 391, 379, 376, 381, 385, 379, 378, 381, 384, 387, 395, 399, 405, 411, 402, 358, 293, 247, 237, 270, 331, 
    413, 405, 400, 397, 393, 393, 398, 404, 408, 391, 374, 369, 375, 380, 375, 374, 372, 372, 372, 388, 399, 406, 399, 357, 296, 248, 244, 291, 352, 388, 
    
    -- channel=4
    362, 418, 441, 408, 388, 365, 345, 373, 464, 478, 430, 388, 393, 409, 369, 339, 338, 345, 321, 311, 361, 369, 269, 250, 409, 433, 407, 397, 372, 366, 
    324, 392, 395, 368, 364, 342, 331, 383, 471, 473, 429, 387, 401, 423, 369, 336, 346, 359, 329, 310, 369, 366, 254, 236, 399, 422, 381, 347, 336, 373, 
    286, 362, 352, 348, 346, 324, 319, 394, 476, 483, 455, 418, 417, 419, 367, 334, 336, 343, 323, 311, 375, 360, 239, 209, 347, 365, 323, 285, 304, 351, 
    283, 341, 333, 346, 334, 321, 322, 410, 479, 495, 469, 428, 406, 387, 344, 318, 318, 332, 347, 332, 370, 347, 223, 169, 274, 294, 272, 245, 269, 308, 
    324, 360, 348, 346, 326, 335, 343, 433, 480, 482, 434, 396, 361, 349, 358, 346, 310, 345, 396, 350, 357, 331, 202, 127, 213, 243, 242, 211, 248, 295, 
    387, 378, 362, 341, 324, 352, 375, 463, 470, 428, 372, 341, 329, 370, 418, 404, 332, 358, 414, 344, 338, 315, 196, 110, 177, 203, 213, 177, 251, 343, 
    409, 353, 310, 299, 324, 357, 388, 472, 441, 368, 321, 306, 343, 428, 469, 420, 350, 370, 381, 315, 315, 288, 200, 124, 169, 175, 186, 162, 294, 408, 
    389, 299, 234, 228, 299, 354, 388, 436, 380, 313, 288, 308, 395, 475, 452, 376, 338, 344, 330, 281, 282, 273, 215, 150, 179, 164, 170, 175, 343, 442, 
    364, 265, 182, 166, 250, 333, 395, 399, 323, 278, 259, 305, 413, 447, 381, 315, 310, 302, 279, 250, 266, 302, 232, 179, 189, 163, 159, 189, 380, 465, 
    370, 267, 180, 132, 187, 296, 379, 360, 300, 271, 257, 318, 365, 334, 278, 264, 272, 267, 258, 248, 285, 323, 226, 192, 197, 160, 149, 201, 406, 489, 
    391, 291, 206, 139, 139, 227, 306, 297, 285, 277, 279, 336, 336, 269, 223, 230, 246, 259, 265, 273, 310, 321, 218, 193, 210, 178, 153, 208, 415, 486, 
    390, 310, 238, 172, 131, 162, 208, 238, 270, 289, 304, 343, 320, 273, 251, 255, 258, 261, 269, 287, 293, 292, 227, 207, 221, 193, 160, 218, 391, 434, 
    361, 305, 254, 214, 155, 133, 148, 218, 280, 306, 309, 331, 321, 299, 288, 293, 295, 290, 278, 283, 259, 256, 229, 234, 239, 208, 165, 222, 358, 375, 
    335, 296, 253, 238, 177, 142, 137, 184, 265, 340, 326, 305, 296, 289, 276, 282, 297, 301, 293, 295, 255, 217, 195, 222, 245, 217, 174, 244, 366, 355, 
    323, 294, 243, 225, 178, 151, 154, 156, 210, 332, 336, 293, 263, 255, 252, 254, 260, 266, 265, 273, 259, 220, 166, 170, 220, 226, 200, 279, 392, 350, 
    302, 279, 231, 214, 181, 166, 169, 150, 163, 265, 287, 274, 245, 227, 224, 233, 240, 238, 236, 248, 243, 226, 180, 166, 200, 228, 229, 305, 406, 341, 
    259, 238, 209, 231, 212, 209, 200, 194, 172, 189, 209, 242, 231, 220, 212, 206, 211, 207, 205, 223, 236, 237, 201, 197, 237, 276, 270, 312, 368, 298, 
    210, 220, 219, 272, 264, 259, 224, 220, 216, 172, 164, 206, 213, 202, 183, 186, 190, 181, 200, 225, 222, 225, 222, 240, 285, 327, 318, 326, 323, 244, 
    201, 236, 252, 304, 310, 282, 258, 241, 246, 223, 206, 194, 182, 171, 148, 160, 164, 147, 173, 212, 211, 213, 233, 251, 317, 330, 333, 312, 268, 193, 
    242, 275, 277, 313, 329, 281, 273, 270, 259, 261, 247, 205, 149, 124, 130, 135, 145, 151, 180, 205, 218, 220, 242, 257, 315, 312, 301, 257, 206, 171, 
    296, 301, 287, 309, 334, 287, 262, 264, 248, 263, 248, 198, 147, 110, 117, 122, 135, 156, 196, 209, 219, 225, 248, 269, 303, 309, 265, 197, 181, 180, 
    288, 240, 246, 285, 327, 308, 246, 226, 227, 247, 234, 176, 145, 122, 128, 127, 141, 164, 199, 210, 226, 223, 245, 279, 310, 313, 246, 184, 182, 194, 
    202, 144, 157, 215, 291, 303, 248, 216, 234, 231, 215, 166, 151, 138, 153, 153, 141, 163, 200, 183, 200, 214, 244, 282, 320, 322, 253, 210, 191, 198, 
    152, 86, 86, 126, 213, 264, 250, 246, 263, 230, 172, 146, 158, 164, 197, 196, 159, 161, 188, 163, 177, 209, 255, 285, 325, 351, 290, 234, 198, 221, 
    203, 159, 108, 99, 138, 195, 232, 262, 274, 241, 191, 157, 173, 215, 273, 266, 198, 169, 177, 161, 176, 208, 252, 282, 338, 401, 322, 251, 230, 261, 
    304, 298, 224, 146, 128, 142, 175, 227, 264, 252, 235, 219, 216, 260, 318, 317, 232, 180, 175, 166, 176, 222, 248, 283, 376, 424, 320, 270, 268, 306, 
    364, 408, 370, 260, 176, 134, 127, 159, 222, 262, 264, 261, 262, 276, 298, 295, 231, 191, 188, 185, 178, 220, 265, 339, 417, 402, 331, 282, 248, 292, 
    373, 444, 465, 383, 270, 167, 114, 110, 149, 204, 235, 245, 260, 259, 271, 273, 231, 212, 211, 184, 190, 242, 294, 379, 432, 379, 357, 291, 219, 257, 
    386, 428, 475, 451, 367, 249, 157, 112, 103, 123, 156, 191, 224, 218, 239, 281, 291, 262, 258, 243, 247, 277, 295, 341, 362, 328, 332, 248, 176, 242, 
    424, 405, 436, 462, 439, 356, 245, 166, 127, 107, 95, 119, 165, 169, 183, 244, 318, 323, 324, 304, 296, 276, 230, 239, 246, 251, 233, 180, 143, 209, 
    
    -- channel=5
    446, 439, 421, 438, 453, 445, 443, 444, 469, 474, 485, 495, 506, 504, 473, 471, 492, 502, 483, 471, 469, 477, 480, 482, 475, 459, 434, 453, 463, 465, 
    378, 383, 403, 446, 451, 433, 435, 433, 458, 466, 478, 494, 508, 505, 494, 501, 528, 540, 507, 478, 468, 465, 466, 460, 453, 446, 447, 462, 459, 454, 
    349, 361, 395, 443, 443, 433, 434, 430, 446, 449, 463, 486, 503, 500, 494, 508, 541, 557, 525, 487, 468, 469, 463, 442, 437, 441, 457, 471, 463, 449, 
    357, 357, 385, 427, 427, 429, 429, 423, 433, 435, 446, 469, 493, 497, 491, 495, 517, 534, 516, 480, 461, 474, 468, 453, 448, 447, 458, 464, 452, 440, 
    369, 350, 372, 403, 412, 420, 418, 415, 412, 424, 441, 455, 477, 495, 482, 481, 476, 484, 483, 464, 455, 480, 480, 468, 465, 464, 459, 453, 444, 434, 
    368, 343, 361, 387, 404, 409, 405, 402, 397, 418, 438, 448, 458, 482, 471, 463, 448, 447, 454, 461, 460, 483, 488, 481, 484, 484, 466, 451, 441, 430, 
    355, 347, 360, 382, 399, 404, 395, 394, 397, 424, 434, 444, 447, 470, 466, 456, 437, 431, 436, 466, 459, 481, 496, 490, 490, 482, 466, 453, 442, 433, 
    348, 353, 358, 378, 393, 405, 400, 396, 399, 423, 430, 432, 428, 441, 440, 443, 439, 434, 429, 460, 435, 449, 484, 485, 479, 465, 456, 446, 442, 435, 
    358, 351, 355, 367, 382, 402, 398, 397, 404, 423, 414, 395, 378, 368, 373, 407, 436, 439, 426, 436, 405, 422, 475, 474, 463, 459, 455, 442, 440, 433, 
    374, 359, 372, 368, 373, 390, 389, 398, 407, 409, 360, 317, 308, 289, 293, 348, 417, 425, 413, 415, 403, 438, 487, 467, 460, 466, 466, 451, 445, 434, 
    361, 350, 361, 344, 349, 358, 362, 391, 402, 375, 289, 246, 259, 277, 310, 340, 397, 401, 383, 385, 404, 457, 497, 474, 467, 475, 476, 460, 447, 440, 
    348, 343, 330, 307, 306, 318, 341, 389, 375, 319, 235, 226, 261, 297, 351, 349, 368, 363, 340, 360, 405, 471, 493, 480, 470, 477, 481, 466, 455, 450, 
    365, 344, 288, 269, 280, 289, 318, 354, 319, 269, 241, 277, 299, 310, 339, 295, 303, 292, 287, 339, 395, 460, 481, 479, 469, 470, 480, 470, 465, 461, 
    412, 365, 281, 260, 274, 289, 305, 305, 258, 230, 244, 305, 319, 281, 268, 216, 220, 220, 241, 304, 376, 445, 468, 474, 459, 440, 452, 468, 472, 465, 
    452, 387, 289, 260, 278, 307, 301, 260, 209, 207, 233, 294, 310, 260, 221, 190, 195, 189, 214, 265, 357, 434, 468, 479, 446, 404, 401, 444, 473, 465, 
    446, 380, 288, 256, 268, 325, 310, 234, 207, 233, 228, 266, 292, 281, 257, 231, 230, 230, 248, 284, 384, 457, 498, 503, 445, 379, 353, 410, 464, 467, 
    437, 375, 279, 243, 247, 325, 336, 231, 230, 270, 244, 265, 320, 331, 341, 314, 313, 323, 336, 377, 458, 502, 532, 515, 446, 370, 322, 369, 449, 468, 
    441, 380, 277, 216, 203, 294, 377, 269, 253, 277, 252, 277, 347, 339, 361, 368, 401, 426, 438, 470, 505, 518, 535, 508, 447, 363, 296, 313, 426, 472, 
    438, 382, 280, 203, 181, 265, 425, 372, 312, 272, 250, 303, 382, 332, 335, 368, 452, 506, 494, 499, 496, 492, 521, 504, 455, 353, 269, 252, 387, 466, 
    423, 383, 289, 210, 193, 273, 469, 474, 411, 366, 332, 361, 410, 355, 345, 388, 466, 532, 517, 499, 478, 467, 504, 502, 468, 362, 250, 211, 348, 455, 
    401, 386, 313, 245, 238, 325, 488, 513, 483, 468, 445, 440, 455, 420, 416, 458, 497, 536, 525, 512, 502, 486, 497, 495, 469, 387, 271, 212, 327, 447, 
    398, 391, 343, 289, 285, 359, 454, 485, 502, 500, 488, 475, 472, 462, 493, 528, 534, 546, 537, 528, 533, 519, 507, 495, 469, 425, 328, 255, 324, 448, 
    405, 379, 363, 334, 305, 327, 381, 449, 486, 486, 476, 469, 465, 470, 515, 550, 548, 549, 542, 536, 544, 533, 520, 503, 468, 468, 405, 329, 332, 427, 
    406, 383, 380, 371, 336, 300, 310, 405, 433, 439, 443, 448, 444, 471, 509, 534, 539, 544, 544, 542, 550, 540, 534, 509, 472, 497, 468, 407, 365, 393, 
    400, 384, 381, 380, 357, 336, 311, 370, 393, 414, 431, 426, 420, 448, 476, 499, 505, 517, 518, 527, 539, 528, 524, 502, 486, 513, 489, 433, 406, 400, 
    401, 397, 368, 367, 373, 391, 352, 349, 371, 408, 437, 408, 390, 412, 453, 478, 473, 475, 479, 494, 511, 497, 490, 486, 490, 506, 475, 427, 433, 420, 
    408, 404, 359, 362, 391, 428, 389, 386, 409, 404, 427, 398, 383, 399, 441, 455, 443, 441, 448, 464, 475, 459, 454, 464, 472, 474, 458, 433, 456, 426, 
    417, 398, 366, 379, 399, 424, 402, 397, 414, 393, 409, 402, 399, 402, 432, 438, 431, 439, 445, 452, 453, 436, 430, 438, 443, 445, 458, 458, 453, 409, 
    414, 384, 374, 389, 402, 406, 393, 403, 390, 371, 399, 414, 425, 423, 429, 434, 438, 455, 453, 445, 439, 426, 415, 419, 422, 429, 456, 469, 434, 388, 
    390, 368, 390, 405, 403, 395, 382, 400, 390, 383, 405, 420, 439, 447, 444, 443, 445, 454, 444, 430, 426, 417, 401, 407, 414, 418, 433, 437, 413, 394, 
    
    -- channel=6
    757, 778, 779, 769, 779, 798, 796, 792, 793, 787, 774, 758, 754, 762, 759, 750, 710, 659, 646, 648, 673, 669, 639, 597, 548, 523, 522, 580, 644, 660, 
    786, 788, 773, 766, 775, 789, 784, 777, 771, 764, 751, 737, 735, 740, 737, 729, 706, 697, 681, 674, 680, 666, 622, 573, 540, 517, 523, 591, 656, 668, 
    761, 747, 735, 742, 752, 766, 761, 750, 742, 734, 722, 711, 713, 717, 713, 707, 693, 692, 685, 661, 628, 610, 589, 563, 551, 534, 540, 605, 656, 666, 
    705, 697, 699, 717, 724, 737, 735, 726, 716, 709, 698, 692, 698, 699, 695, 689, 682, 684, 678, 616, 538, 508, 517, 541, 560, 540, 551, 603, 644, 655, 
    666, 672, 686, 700, 701, 710, 711, 705, 699, 691, 683, 680, 688, 687, 685, 679, 678, 678, 659, 566, 468, 433, 442, 496, 538, 539, 569, 605, 642, 654, 
    669, 679, 685, 689, 684, 691, 693, 692, 688, 682, 675, 673, 680, 677, 676, 669, 663, 660, 627, 535, 468, 435, 429, 483, 533, 566, 603, 625, 657, 663, 
    674, 682, 680, 681, 674, 681, 680, 681, 679, 676, 672, 659, 652, 641, 646, 640, 635, 633, 594, 536, 504, 482, 465, 512, 573, 622, 645, 654, 673, 671, 
    668, 678, 677, 681, 672, 677, 674, 673, 669, 660, 649, 621, 607, 600, 615, 615, 605, 594, 558, 521, 493, 480, 478, 535, 613, 654, 667, 666, 670, 667, 
    663, 677, 679, 683, 674, 676, 674, 668, 657, 636, 620, 575, 551, 541, 539, 511, 463, 422, 422, 416, 405, 428, 444, 504, 576, 619, 649, 658, 659, 659, 
    667, 679, 677, 681, 673, 676, 674, 665, 650, 614, 566, 467, 398, 359, 329, 287, 223, 177, 198, 181, 216, 349, 430, 480, 487, 530, 604, 642, 651, 654, 
    674, 679, 672, 675, 671, 673, 672, 657, 618, 542, 453, 326, 243, 196, 168, 146, 113, 99, 102, 0, 21, 234, 410, 489, 447, 443, 529, 604, 636, 649, 
    677, 675, 667, 668, 671, 670, 663, 621, 544, 453, 351, 235, 190, 197, 211, 225, 249, 270, 171, 0, 0, 86, 342, 486, 456, 414, 467, 545, 604, 638, 
    671, 671, 666, 665, 672, 662, 632, 558, 472, 395, 325, 271, 289, 342, 394, 408, 437, 421, 212, 0, 0, 0, 204, 419, 474, 435, 458, 501, 562, 614, 
    664, 667, 667, 658, 638, 609, 560, 492, 424, 395, 366, 344, 379, 425, 465, 443, 419, 314, 90, 0, 0, 0, 87, 313, 445, 472, 475, 456, 480, 561, 
    659, 664, 662, 635, 562, 501, 452, 406, 395, 396, 368, 357, 359, 324, 304, 246, 185, 61, 0, 0, 0, 0, 109, 282, 423, 505, 471, 363, 342, 469, 
    658, 660, 647, 604, 497, 412, 354, 338, 365, 386, 375, 383, 299, 142, 57, 0, 0, 0, 0, 0, 0, 30, 248, 351, 442, 473, 383, 226, 180, 363, 
    660, 647, 589, 536, 443, 371, 321, 313, 377, 407, 394, 395, 224, 0, 0, 0, 0, 0, 0, 0, 0, 146, 347, 382, 384, 338, 224, 108, 71, 286, 
    658, 573, 436, 411, 393, 366, 321, 359, 430, 458, 413, 380, 145, 0, 0, 0, 0, 0, 0, 0, 0, 87, 231, 257, 213, 146, 74, 45, 48, 268, 
    614, 405, 219, 236, 305, 348, 340, 415, 471, 495, 434, 360, 103, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 38, 20, 0, 4, 35, 104, 315, 
    532, 254, 75, 111, 246, 328, 367, 457, 501, 510, 444, 349, 88, 0, 0, 0, 0, 32, 143, 173, 101, 0, 0, 0, 0, 0, 8, 94, 232, 400, 
    481, 271, 127, 98, 223, 306, 392, 486, 516, 477, 386, 288, 57, 0, 0, 0, 13, 215, 329, 364, 317, 157, 0, 0, 0, 2, 86, 224, 378, 478, 
    497, 393, 257, 149, 219, 302, 424, 496, 503, 409, 300, 200, 0, 0, 0, 0, 148, 331, 410, 434, 429, 319, 131, 20, 13, 66, 203, 367, 475, 507, 
    544, 468, 331, 177, 208, 303, 434, 478, 452, 331, 239, 128, 0, 0, 0, 0, 227, 345, 398, 415, 445, 422, 261, 118, 58, 128, 311, 446, 503, 510, 
    555, 448, 333, 175, 195, 313, 426, 436, 371, 259, 205, 90, 0, 0, 0, 0, 248, 333, 369, 382, 415, 456, 358, 193, 110, 203, 380, 478, 515, 518, 
    541, 428, 332, 182, 181, 287, 361, 330, 230, 131, 92, 3, 0, 0, 0, 6, 242, 317, 310, 306, 362, 439, 420, 274, 208, 303, 434, 502, 528, 527, 
    538, 432, 342, 208, 196, 276, 307, 265, 172, 93, 59, 11, 0, 0, 0, 60, 256, 309, 297, 285, 342, 422, 461, 380, 353, 416, 488, 527, 537, 524, 
    537, 463, 387, 288, 285, 339, 349, 321, 264, 222, 203, 185, 172, 170, 171, 231, 353, 339, 308, 300, 347, 426, 496, 473, 476, 507, 531, 541, 536, 513, 
    525, 485, 445, 392, 394, 416, 430, 431, 413, 402, 396, 390, 385, 388, 394, 418, 469, 418, 365, 331, 371, 452, 518, 535, 545, 549, 550, 545, 529, 502, 
    501, 484, 448, 416, 401, 400, 429, 450, 447, 442, 440, 445, 454, 466, 477, 494, 513, 471, 420, 385, 398, 476, 527, 549, 552, 550, 546, 536, 515, 492, 
    460, 424, 361, 314, 285, 287, 336, 364, 366, 359, 354, 362, 378, 396, 413, 436, 461, 462, 422, 394, 430, 487, 520, 529, 528, 528, 522, 510, 488, 479, 
    
    -- channel=7
    293, 303, 310, 308, 295, 293, 297, 314, 336, 349, 357, 362, 362, 357, 356, 358, 366, 371, 384, 396, 405, 417, 430, 444, 453, 458, 456, 464, 470, 473, 
    295, 304, 315, 311, 306, 332, 331, 339, 366, 377, 375, 376, 391, 397, 395, 388, 383, 381, 398, 415, 425, 433, 439, 445, 445, 442, 436, 439, 441, 441, 
    298, 304, 319, 314, 320, 369, 362, 369, 400, 418, 418, 415, 426, 436, 437, 432, 412, 396, 399, 409, 418, 420, 419, 420, 412, 405, 398, 400, 405, 411, 
    306, 306, 321, 323, 341, 387, 383, 402, 437, 462, 469, 468, 477, 488, 482, 467, 422, 386, 370, 374, 381, 380, 379, 380, 372, 368, 369, 379, 393, 409, 
    320, 318, 327, 342, 378, 412, 411, 441, 475, 499, 512, 516, 522, 525, 516, 494, 431, 371, 340, 336, 339, 340, 349, 358, 356, 358, 365, 383, 405, 426, 
    335, 333, 338, 366, 415, 448, 457, 480, 504, 523, 534, 543, 546, 541, 528, 513, 462, 395, 349, 327, 327, 340, 356, 361, 359, 360, 373, 395, 421, 444, 
    343, 336, 334, 349, 402, 466, 487, 509, 514, 518, 523, 530, 529, 530, 529, 527, 505, 458, 410, 373, 357, 367, 383, 377, 368, 369, 385, 408, 429, 445, 
    317, 297, 280, 269, 331, 442, 489, 521, 513, 491, 480, 474, 478, 501, 517, 536, 535, 512, 479, 442, 415, 410, 409, 390, 377, 376, 391, 409, 423, 433, 
    246, 216, 191, 164, 260, 411, 474, 515, 507, 464, 431, 413, 420, 467, 499, 524, 536, 536, 527, 509, 484, 454, 433, 399, 380, 379, 392, 404, 410, 416, 
    161, 134, 114, 97, 229, 397, 458, 494, 499, 456, 413, 397, 399, 441, 480, 505, 520, 532, 542, 539, 529, 493, 461, 420, 388, 380, 383, 389, 392, 399, 
    106, 96, 92, 88, 211, 378, 438, 460, 466, 438, 403, 401, 408, 439, 468, 479, 491, 508, 527, 537, 545, 520, 480, 441, 404, 383, 375, 376, 380, 389, 
    100, 100, 104, 104, 182, 337, 421, 440, 427, 404, 381, 395, 417, 447, 469, 460, 461, 476, 497, 516, 541, 532, 489, 456, 422, 392, 372, 368, 375, 390, 
    114, 119, 123, 124, 155, 267, 367, 416, 430, 414, 389, 400, 434, 457, 474, 450, 438, 444, 467, 494, 530, 538, 497, 465, 438, 404, 380, 374, 385, 401, 
    137, 138, 135, 130, 140, 203, 281, 349, 428, 446, 410, 409, 446, 466, 470, 437, 415, 412, 439, 478, 519, 539, 513, 475, 455, 428, 409, 397, 399, 408, 
    146, 138, 129, 122, 143, 190, 216, 271, 365, 414, 394, 395, 432, 461, 462, 428, 396, 391, 420, 466, 508, 530, 526, 486, 468, 448, 425, 410, 408, 418, 
    139, 127, 112, 99, 121, 191, 173, 186, 262, 314, 333, 339, 379, 435, 452, 426, 394, 383, 410, 453, 491, 514, 527, 495, 474, 454, 426, 415, 427, 454, 
    108, 83, 51, 19, 22, 111, 135, 123, 159, 198, 285, 292, 335, 406, 445, 434, 401, 386, 404, 437, 469, 495, 518, 502, 473, 457, 434, 441, 470, 504, 
    24, 0, 0, 0, 0, 0, 52, 84, 133, 130, 265, 281, 315, 389, 438, 438, 406, 389, 396, 417, 445, 475, 506, 507, 478, 473, 468, 487, 517, 538, 
    0, 0, 0, 0, 0, 0, 49, 112, 161, 145, 270, 305, 332, 392, 435, 437, 413, 394, 393, 405, 428, 465, 498, 511, 486, 490, 502, 520, 534, 537, 
    0, 0, 0, 0, 13, 46, 152, 206, 232, 233, 320, 361, 372, 413, 433, 431, 418, 404, 397, 406, 433, 471, 502, 516, 495, 487, 501, 518, 529, 531, 
    0, 0, 0, 26, 145, 195, 268, 307, 330, 356, 401, 420, 419, 441, 436, 426, 423, 417, 413, 420, 442, 470, 496, 512, 499, 474, 476, 500, 522, 530, 
    0, 0, 0, 93, 190, 243, 302, 360, 413, 456, 479, 460, 433, 452, 457, 449, 448, 443, 433, 430, 437, 452, 478, 504, 501, 470, 456, 481, 513, 529, 
    0, 2, 58, 141, 191, 228, 282, 353, 437, 493, 505, 460, 422, 443, 462, 466, 466, 459, 441, 420, 408, 410, 443, 493, 510, 487, 455, 463, 496, 522, 
    109, 149, 177, 200, 222, 240, 273, 325, 388, 443, 462, 432, 410, 434, 466, 470, 467, 455, 417, 379, 369, 381, 417, 472, 508, 506, 476, 457, 473, 508, 
    227, 238, 243, 255, 267, 280, 287, 312, 357, 395, 424, 427, 426, 429, 455, 465, 458, 441, 387, 340, 340, 366, 408, 457, 493, 511, 502, 469, 461, 490, 
    285, 288, 289, 295, 301, 315, 333, 358, 381, 393, 419, 449, 456, 438, 451, 471, 466, 449, 393, 343, 343, 375, 415, 449, 485, 509, 519, 493, 469, 479, 
    321, 322, 322, 332, 351, 382, 412, 442, 448, 430, 441, 466, 461, 450, 466, 492, 490, 476, 439, 401, 388, 401, 427, 454, 485, 515, 529, 518, 495, 482, 
    340, 354, 374, 397, 426, 459, 486, 507, 492, 450, 442, 458, 458, 470, 494, 521, 522, 511, 495, 474, 454, 446, 453, 472, 502, 531, 541, 537, 523, 499, 
    387, 417, 447, 470, 491, 514, 525, 533, 506, 465, 450, 452, 463, 495, 520, 546, 547, 536, 532, 525, 507, 496, 496, 507, 530, 549, 554, 550, 544, 525, 
    457, 488, 509, 521, 529, 536, 537, 542, 515, 479, 471, 458, 478, 512, 536, 559, 561, 550, 548, 548, 536, 531, 533, 537, 549, 562, 566, 559, 553, 543, 
    
    -- channel=8
    496, 479, 340, 246, 240, 252, 242, 223, 227, 243, 248, 248, 253, 247, 229, 211, 236, 314, 363, 340, 216, 147, 153, 171, 192, 197, 197, 204, 214, 225, 
    493, 494, 370, 250, 242, 253, 217, 167, 161, 192, 202, 194, 192, 188, 171, 149, 163, 248, 338, 308, 168, 106, 109, 131, 153, 162, 167, 176, 187, 198, 
    493, 499, 403, 271, 264, 273, 205, 115, 86, 132, 166, 170, 162, 148, 135, 122, 137, 218, 308, 248, 114, 60, 60, 85, 107, 122, 133, 146, 157, 171, 
    491, 495, 434, 304, 290, 294, 209, 89, 20, 70, 138, 176, 186, 167, 148, 139, 164, 216, 254, 171, 74, 34, 30, 43, 59, 69, 78, 92, 104, 119, 
    494, 493, 460, 332, 281, 274, 204, 77, 0, 21, 120, 201, 233, 217, 205, 191, 209, 220, 184, 87, 41, 18, 6, 3, 5, 5, 10, 24, 37, 48, 
    501, 501, 444, 295, 219, 221, 186, 71, 0, 0, 81, 180, 230, 238, 253, 240, 247, 220, 131, 32, 23, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    420, 438, 353, 209, 136, 167, 187, 93, 1, 0, 32, 109, 161, 203, 250, 249, 252, 216, 110, 17, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    274, 288, 205, 110, 80, 151, 210, 131, 36, 0, 0, 38, 88, 152, 228, 234, 231, 207, 113, 30, 20, 0, 0, 0, 0, 0, 21, 44, 15, 0, 
    142, 140, 89, 56, 61, 158, 222, 149, 58, 1, 0, 10, 61, 135, 210, 220, 216, 202, 124, 52, 24, 0, 0, 0, 0, 0, 63, 90, 58, 0, 
    75, 72, 51, 33, 54, 156, 200, 130, 53, 8, 0, 19, 81, 161, 220, 205, 203, 196, 123, 67, 29, 0, 0, 0, 0, 0, 67, 108, 96, 42, 
    61, 64, 49, 37, 62, 144, 164, 110, 47, 19, 13, 40, 105, 184, 208, 171, 171, 166, 107, 71, 37, 0, 0, 0, 0, 0, 41, 98, 115, 85, 
    64, 74, 62, 73, 103, 130, 140, 115, 84, 70, 48, 63, 120, 167, 156, 119, 132, 121, 92, 74, 39, 0, 0, 0, 0, 0, 0, 61, 96, 80, 
    68, 83, 73, 115, 160, 128, 120, 103, 99, 98, 64, 59, 114, 152, 110, 75, 104, 96, 78, 68, 37, 0, 0, 0, 0, 0, 0, 11, 44, 29, 
    69, 85, 70, 137, 205, 131, 94, 67, 71, 73, 51, 48, 87, 122, 98, 74, 94, 104, 79, 65, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    76, 93, 75, 131, 216, 135, 65, 18, 28, 29, 30, 45, 68, 93, 117, 110, 104, 132, 103, 78, 84, 95, 60, 0, 0, 0, 0, 0, 0, 0, 
    92, 119, 100, 114, 178, 124, 48, 0, 0, 0, 16, 40, 44, 60, 141, 158, 131, 163, 136, 98, 117, 184, 197, 128, 28, 0, 1, 2, 0, 0, 
    97, 137, 119, 93, 118, 94, 40, 0, 0, 0, 0, 0, 9, 32, 141, 200, 165, 190, 163, 112, 139, 217, 262, 235, 152, 90, 96, 68, 1, 0, 
    80, 124, 104, 63, 52, 48, 31, 0, 0, 0, 0, 0, 0, 6, 92, 183, 184, 194, 154, 113, 157, 202, 255, 267, 213, 164, 161, 139, 82, 22, 
    46, 92, 73, 34, 16, 18, 23, 11, 0, 0, 0, 0, 0, 0, 19, 100, 150, 160, 138, 136, 190, 203, 224, 234, 198, 172, 187, 187, 157, 107, 
    13, 60, 58, 25, 3, 3, 15, 12, 3, 11, 32, 9, 0, 0, 0, 19, 87, 109, 141, 180, 216, 208, 202, 185, 159, 162, 193, 206, 201, 182, 
    0, 39, 65, 32, 0, 0, 0, 0, 0, 16, 75, 63, 34, 20, 0, 0, 47, 92, 178, 225, 223, 195, 175, 146, 137, 165, 199, 214, 225, 239, 
    0, 25, 76, 45, 0, 0, 0, 0, 0, 12, 74, 74, 53, 42, 25, 19, 47, 119, 219, 245, 211, 179, 158, 124, 129, 164, 192, 217, 242, 266, 
    0, 25, 83, 56, 0, 0, 0, 0, 0, 37, 77, 63, 47, 45, 40, 40, 69, 154, 238, 238, 198, 178, 166, 126, 126, 154, 185, 220, 246, 265, 
    12, 37, 90, 69, 8, 0, 0, 0, 18, 119, 124, 73, 47, 51, 56, 66, 105, 182, 239, 227, 196, 189, 181, 146, 145, 162, 191, 219, 241, 257, 
    26, 59, 107, 96, 29, 0, 0, 0, 67, 204, 184, 104, 71, 76, 91, 110, 151, 209, 247, 228, 207, 210, 201, 184, 193, 200, 209, 214, 229, 246, 
    40, 82, 129, 131, 58, 0, 0, 0, 83, 203, 177, 123, 107, 118, 141, 167, 197, 248, 270, 241, 224, 227, 219, 226, 241, 247, 230, 212, 215, 230, 
    57, 99, 152, 165, 83, 0, 0, 0, 55, 130, 124, 124, 143, 163, 186, 213, 241, 293, 288, 255, 238, 239, 232, 253, 276, 273, 240, 209, 200, 212, 
    85, 113, 167, 195, 110, 3, 0, 0, 21, 62, 85, 132, 176, 198, 221, 245, 282, 325, 296, 269, 252, 242, 237, 262, 282, 273, 242, 213, 203, 216, 
    122, 127, 171, 217, 145, 28, 0, 0, 6, 35, 94, 168, 221, 236, 248, 269, 314, 329, 294, 279, 260, 243, 240, 259, 268, 260, 245, 229, 221, 227, 
    171, 160, 184, 240, 192, 73, 0, 0, 16, 54, 135, 229, 292, 301, 293, 301, 327, 317, 295, 287, 267, 246, 245, 255, 263, 263, 258, 243, 228, 227, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 30, 32, 23, 15, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 13, 8, 
    0, 0, 0, 0, 0, 0, 24, 13, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 50, 31, 34, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 104, 77, 54, 2, 3, 13, 0, 13, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 22, 0, 0, 
    0, 0, 0, 0, 0, 5, 119, 87, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 64, 12, 0, 
    0, 0, 0, 0, 0, 0, 97, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 84, 52, 0, 
    0, 0, 0, 0, 0, 0, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 86, 82, 7, 
    0, 0, 0, 0, 0, 0, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 52, 0, 
    0, 0, 0, 0, 0, 6, 72, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 40, 102, 50, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 49, 133, 130, 98, 45, 0, 0, 0, 5, 2, 1, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 75, 131, 134, 94, 45, 0, 0, 0, 19, 38, 32, 13, 0, 0, 19, 44, 53, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 56, 66, 112, 125, 99, 37, 4, 0, 0, 0, 33, 62, 54, 25, 0, 0, 59, 98, 101, 43, 0, 0, 0, 0, 0, 0, 0, 
    0, 40, 98, 119, 90, 97, 104, 79, 35, 46, 82, 87, 101, 113, 127, 114, 94, 77, 100, 145, 161, 156, 120, 80, 31, 0, 0, 0, 0, 0, 
    0, 124, 181, 161, 88, 70, 107, 109, 79, 91, 143, 165, 172, 178, 219, 242, 255, 261, 250, 253, 266, 267, 254, 206, 121, 68, 0, 0, 0, 0, 
    12, 154, 205, 161, 85, 116, 172, 145, 125, 128, 133, 151, 142, 169, 235, 273, 284, 295, 245, 222, 260, 286, 299, 250, 146, 62, 0, 0, 0, 0, 
    0, 137, 187, 137, 106, 227, 258, 185, 130, 125, 118, 110, 74, 116, 159, 168, 174, 179, 110, 92, 139, 166, 198, 144, 72, 42, 12, 0, 0, 0, 
    0, 115, 182, 136, 146, 302, 308, 228, 160, 157, 167, 171, 125, 133, 72, 49, 63, 68, 7, 0, 39, 52, 72, 11, 0, 52, 68, 31, 0, 0, 
    0, 113, 214, 184, 201, 313, 318, 270, 224, 216, 231, 239, 204, 193, 79, 29, 38, 45, 27, 28, 39, 46, 53, 2, 20, 104, 139, 100, 0, 0, 
    0, 93, 214, 235, 252, 297, 312, 323, 304, 286, 262, 254, 227, 223, 166, 141, 127, 120, 119, 124, 135, 120, 121, 102, 113, 143, 136, 108, 0, 0, 
    0, 82, 202, 236, 265, 285, 301, 348, 353, 349, 288, 234, 159, 206, 255, 225, 156, 144, 163, 160, 170, 122, 93, 173, 200, 146, 107, 107, 0, 0, 
    0, 81, 210, 233, 244, 241, 255, 324, 368, 392, 338, 272, 169, 217, 308, 285, 173, 147, 158, 141, 153, 85, 56, 201, 250, 187, 150, 149, 0, 0, 
    0, 91, 244, 264, 245, 171, 177, 267, 343, 399, 376, 343, 267, 302, 355, 321, 212, 165, 137, 102, 106, 55, 69, 227, 275, 251, 247, 221, 7, 0, 
    0, 56, 214, 249, 218, 117, 121, 214, 306, 381, 411, 412, 385, 391, 395, 371, 281, 165, 74, 23, 36, 15, 112, 273, 327, 331, 317, 246, 15, 0, 
    0, 0, 91, 157, 153, 74, 116, 185, 258, 342, 409, 438, 442, 431, 411, 407, 344, 161, 27, 0, 0, 0, 136, 295, 369, 372, 315, 222, 2, 0, 
    0, 0, 0, 45, 95, 57, 133, 176, 219, 300, 387, 434, 444, 431, 403, 381, 311, 141, 28, 0, 0, 0, 142, 314, 398, 385, 294, 196, 0, 0, 
    0, 0, 0, 9, 82, 73, 155, 180, 201, 273, 365, 420, 432, 418, 388, 354, 295, 187, 120, 64, 16, 0, 173, 334, 412, 381, 287, 193, 0, 0, 
    0, 0, 0, 2, 79, 113, 189, 198, 215, 270, 344, 394, 405, 394, 369, 336, 300, 253, 209, 152, 89, 52, 195, 336, 410, 376, 297, 198, 0, 0, 
    0, 0, 0, 0, 58, 154, 221, 228, 239, 283, 329, 364, 369, 360, 348, 336, 310, 279, 244, 200, 154, 118, 217, 333, 399, 374, 302, 173, 0, 0, 
    0, 0, 0, 0, 21, 165, 244, 267, 272, 291, 313, 330, 322, 311, 305, 298, 275, 249, 227, 202, 179, 159, 210, 300, 348, 336, 257, 102, 0, 0, 
    
    
    others => 0);
end gold_package;
