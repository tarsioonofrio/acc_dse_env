-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use IEEE.std_logic_arith.all;

-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity bram_single is
    generic (
        DEVICE     : string := "7SERIES";
        BRAM_NAME  : string := "default"
        );

    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic;
        DI   : in std_logic_vector(36-1 downto 0);
        ADDR : in std_logic_vector(9-1 downto 0);
        DO   : out std_logic_vector(36-1 downto 0)
    );
    attribute dont_touch : string;
    attribute dont_touch of bram_single : entity is "true";
   end bram_single;

  architecture a1 of bram_single is
    signal bram_wr_en    : std_logic_vector(8-1 downto 0);
    signal bram_addr     : std_logic_vector(9-1 downto 0);
    signal bram_di     : std_logic_vector(44-1 downto 0);
    signal bram_do     : std_logic_vector(44-1 downto 0);
    constant bram_par     : std_logic_vector(8-1 downto 0) := "00000000";

    begin
    bram_wr_en <= (others => '1') when WE = '1' else (others => '0');
    bram_addr <= ADDR(9-1 downto 0);
    bram_di <= bram_par & DI;
    DO <= bram_do(36-1 downto 0);


    MEM_IWGHT_LAYER0_INSTANCE0 : if BRAM_NAME = "iwght_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000151600000000ffffb971ffffffffffffabcbffffffff0000012600000000",
            INIT_01 => X"0000198d00000000fffffa62ffffffff000022be0000000000000f5d00000000",
            INIT_02 => X"fffff1b0fffffffffffff3a4ffffffff0000053100000000000003bc00000000",
            INIT_03 => X"fffffa2bffffffff00000f3500000000ffffeab4fffffffffffff10bffffffff",
            INIT_04 => X"ffffffaeffffffff0000000a00000000ffffffe6ffffffffffffffe1ffffffff",
            INIT_05 => X"0000004700000000ffffffd0ffffffff00000025000000000000002600000000",
            INIT_06 => X"0000000c000000000000002100000000ffffffc9ffffffff0000001600000000",
            INIT_07 => X"ffffffd7ffffffff0000004800000000fffffffdffffffffffffffc1ffffffff",
            INIT_08 => X"ffffffddffffffffffffffe0fffffffffffffff5ffffffff0000003f00000000",
            INIT_09 => X"00000001000000000000000700000000ffffffb1ffffffff0000001300000000",
            INIT_0A => X"ffffffbdffffffff00000043000000000000003b00000000ffffffe4ffffffff",
            INIT_0B => X"0000001000000000000000010000000000000020000000000000001c00000000",
            INIT_0C => X"00000026000000000000001f00000000ffffffe7ffffffff0000001200000000",
            INIT_0D => X"0000001d000000000000001d0000000000000039000000000000001500000000",
            INIT_0E => X"0000003900000000000000190000000000000034000000000000003d00000000",
            INIT_0F => X"00000003000000000000003400000000fffffffcffffffff0000003c00000000",
            INIT_10 => X"00000009000000000000001500000000ffffffffffffffff0000001900000000",
            INIT_11 => X"0000003000000000fffffffbffffffff0000003e000000000000002800000000",
            INIT_12 => X"00000002000000000000002300000000ffffffefffffffff0000003700000000",
            INIT_13 => X"fffffff7ffffffff0000001800000000fffffffbffffffffffffffd8ffffffff",
            INIT_14 => X"ffffffe0ffffffffffffffd0fffffffffffffff4fffffffffffffff4ffffffff",
            INIT_15 => X"0000000600000000ffffffd1fffffffffffffffaffffffff0000001c00000000",
            INIT_16 => X"ffffffffffffffff0000003d0000000000000048000000000000001500000000",
            INIT_17 => X"0000002800000000ffffffedffffffff0000004c000000000000001800000000",
            INIT_18 => X"ffffffe8ffffffff00000008000000000000000600000000ffffffe6ffffffff",
            INIT_19 => X"ffffffe5fffffffffffffffeffffffffffffffc9fffffffffffffff0ffffffff",
            INIT_1A => X"ffffffceffffffff000000050000000000000017000000000000000e00000000",
            INIT_1B => X"ffffffdeffffffff0000000d000000000000000100000000ffffffe5ffffffff",
            INIT_1C => X"0000002b00000000ffffffcfffffffffffffffd9ffffffffffffffcfffffffff",
            INIT_1D => X"fffffff8ffffffff000000180000000000000010000000000000001a00000000",
            INIT_1E => X"0000004200000000000000070000000000000048000000000000003700000000",
            INIT_1F => X"0000000d000000000000002d0000000000000027000000000000000c00000000",
            INIT_20 => X"0000002200000000000000270000000000000040000000000000002500000000",
            INIT_21 => X"ffffffd1ffffffff0000002200000000ffffffc6ffffffff0000000000000000",
            INIT_22 => X"fffffffdffffffff0000001f00000000ffffffdcffffffff0000000a00000000",
            INIT_23 => X"0000000600000000ffffffd5ffffffff0000000b00000000fffffffdffffffff",
            INIT_24 => X"fffffffcffffffffffffffecfffffffffffffffbffffffff0000000000000000",
            INIT_25 => X"ffffffccffffffffffffffe9ffffffffffffffdaffffffffffffffc0ffffffff",
            INIT_26 => X"fffffff2ffffffffffffffd1ffffffff0000001100000000ffffffe8ffffffff",
            INIT_27 => X"ffffffeaffffffff0000001200000000ffffffc5ffffffff0000002700000000",
            INIT_28 => X"000000270000000000000048000000000000003b00000000ffffffefffffffff",
            INIT_29 => X"00000017000000000000001b000000000000002f000000000000000700000000",
            INIT_2A => X"ffffffdbffffffff0000002600000000ffffffedffffffff0000001e00000000",
            INIT_2B => X"0000000100000000ffffffe2ffffffffffffffd3ffffffffffffffd3ffffffff",
            INIT_2C => X"0000000000000000ffffffcbffffffffffffffc8ffffffff0000000400000000",
            INIT_2D => X"fffffff3ffffffffffffffd9ffffffffffffffbcffffffffffffffe7ffffffff",
            INIT_2E => X"0000000800000000ffffffd6ffffffff0000000900000000ffffffb8ffffffff",
            INIT_2F => X"fffffff9ffffffff000000110000000000000022000000000000003c00000000",
            INIT_30 => X"0000000f00000000000000080000000000000037000000000000001600000000",
            INIT_31 => X"000000260000000000000033000000000000002f000000000000002000000000",
            INIT_32 => X"0000002700000000fffffffaffffffff0000000b000000000000002600000000",
            INIT_33 => X"fffffff3ffffffffffffffe2ffffffff0000001d000000000000000700000000",
            INIT_34 => X"0000002c00000000fffffff3ffffffff0000002a00000000fffffff6ffffffff",
            INIT_35 => X"fffffff3ffffffff00000035000000000000002b000000000000002c00000000",
            INIT_36 => X"0000002f00000000ffffffe2ffffffff00000038000000000000001100000000",
            INIT_37 => X"ffffffd1fffffffffffffff5fffffffffffffff0ffffffff0000002c00000000",
            INIT_38 => X"ffffffcfffffffffffffffd7ffffffffffffffe5ffffffff0000001d00000000",
            INIT_39 => X"ffffffefffffffffffffffc7ffffffffffffffc8ffffffffffffffdfffffffff",
            INIT_3A => X"ffffffbaffffffff0000004700000000fffffff4ffffffffffffffebffffffff",
            INIT_3B => X"0000000f00000000ffffffb8ffffffff0000002700000000fffffffaffffffff",
            INIT_3C => X"0000004f000000000000001a00000000ffffffdbffffffff0000003300000000",
            INIT_3D => X"ffffffbbffffffff00000007000000000000002d00000000ffffffdfffffffff",
            INIT_3E => X"fffffff3ffffffffffffffffffffffff0000001200000000ffffffd3ffffffff",
            INIT_3F => X"0000003b00000000ffffffeaffffffffffffffd8ffffffff0000002600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000042000000000000003600000000ffffffe6ffffffffffffffddffffffff",
            INIT_41 => X"fffffff3ffffffff000000220000000000000039000000000000003000000000",
            INIT_42 => X"ffffffd8ffffffffffffffc2ffffffffffffffbaffffffffffffffccffffffff",
            INIT_43 => X"ffffffe3ffffffff000000190000000000000018000000000000003800000000",
            INIT_44 => X"ffffffd9ffffffffffffffedffffffff00000025000000000000001200000000",
            INIT_45 => X"0000001a000000000000002b00000000ffffffeeffffffffffffffd8ffffffff",
            INIT_46 => X"ffffffcfffffffff0000001e00000000fffffff0ffffffff0000000400000000",
            INIT_47 => X"0000002000000000ffffffdfffffffff0000001200000000ffffffc1ffffffff",
            INIT_48 => X"00000036000000000000002700000000ffffffeaffffffff0000003700000000",
            INIT_49 => X"fffffff0ffffffff0000001d000000000000003f000000000000001600000000",
            INIT_4A => X"000000160000000000000017000000000000001e000000000000000a00000000",
            INIT_4B => X"00000021000000000000002300000000fffffff2ffffffff0000002c00000000",
            INIT_4C => X"0000000a00000000ffffffcfffffffffffffffbfffffffffffffffb8ffffffff",
            INIT_4D => X"ffffffd6ffffffff00000021000000000000001600000000ffffffd3ffffffff",
            INIT_4E => X"ffffffc3fffffffffffffff2ffffffff0000002700000000ffffffeeffffffff",
            INIT_4F => X"0000003300000000ffffffdcffffffff00000023000000000000003200000000",
            INIT_50 => X"ffffffd5ffffffff0000002f00000000fffffff8ffffffff0000000900000000",
            INIT_51 => X"ffffffcfffffffff00000002000000000000003800000000ffffffeeffffffff",
            INIT_52 => X"0000002500000000ffffffd8ffffffffffffffd5ffffffff0000001800000000",
            INIT_53 => X"0000000700000000000000500000000000000005000000000000003400000000",
            INIT_54 => X"ffffffeaffffffffffffffe1ffffffff0000000100000000ffffffd7ffffffff",
            INIT_55 => X"0000003b00000000ffffffe3ffffffff00000000000000000000001d00000000",
            INIT_56 => X"0000000b00000000ffffffefffffffffffffffe7ffffffff0000003800000000",
            INIT_57 => X"ffffffdaffffffff00000016000000000000004b00000000fffffffbffffffff",
            INIT_58 => X"0000003700000000ffffffc2fffffffffffffff3ffffffff0000001a00000000",
            INIT_59 => X"ffffffeeffffffff0000005200000000fffffffaffffffff0000001b00000000",
            INIT_5A => X"ffffffd8ffffffff00000024000000000000002100000000ffffffebffffffff",
            INIT_5B => X"0000003300000000ffffffc5ffffffffffffffe5ffffffff0000003700000000",
            INIT_5C => X"0000000d00000000ffffffefffffffff00000018000000000000002e00000000",
            INIT_5D => X"0000001500000000ffffffdefffffffffffffffbffffffff0000004300000000",
            INIT_5E => X"ffffffe9ffffffff0000001c00000000ffffffeaffffffff0000002900000000",
            INIT_5F => X"fffffffeffffffffffffffe5ffffffff00000001000000000000000800000000",
            INIT_60 => X"ffffffc9ffffffffffffffd0ffffffffffffffeeffffffff0000001d00000000",
            INIT_61 => X"0000000a00000000ffffffb7ffffffffffffffceffffffff0000001f00000000",
            INIT_62 => X"00000045000000000000001400000000ffffffd7ffffffff0000000e00000000",
            INIT_63 => X"0000003200000000ffffffefffffffff00000042000000000000002600000000",
            INIT_64 => X"ffffffe3fffffffffffffffbffffffffffffffdcffffffff0000002e00000000",
            INIT_65 => X"ffffffeaffffffffffffffefffffffff00000004000000000000000800000000",
            INIT_66 => X"ffffffb6ffffffffffffffdcffffffffffffffb8ffffffffffffffc9ffffffff",
            INIT_67 => X"0000000c000000000000003600000000fffffff1ffffffff0000004400000000",
            INIT_68 => X"fffffff5ffffffffffffffefffffffffffffffcaffffffff0000000800000000",
            INIT_69 => X"0000002c000000000000001a000000000000002a00000000ffffffddffffffff",
            INIT_6A => X"ffffffceffffffff0000003c000000000000001f000000000000000900000000",
            INIT_6B => X"ffffffcdffffffff0000001800000000ffffffccffffffffffffffbdffffffff",
            INIT_6C => X"0000002700000000fffffff3ffffffff0000000100000000ffffffdaffffffff",
            INIT_6D => X"ffffffceffffffffffffffe6ffffffff0000000e00000000ffffffd5ffffffff",
            INIT_6E => X"000000390000000000000032000000000000002500000000ffffffebffffffff",
            INIT_6F => X"ffffffe2ffffffff00000000000000000000000d00000000fffffff0ffffffff",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER0_INSTANCE0;


    MEM_IWGHT_LAYER1_INSTANCE0 : if BRAM_NAME = "iwght_layer1_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000249000000000000010d200000000000001b6000000000000069600000000",
            INIT_01 => X"000004be00000000ffffde10ffffffffffffeae6fffffffffffffbbdffffffff",
            INIT_02 => X"ffffe556ffffffffffffeb0dffffffff0000098b00000000ffffe494ffffffff",
            INIT_03 => X"000046b600000000000018a60000000000004b7c00000000fffff7d6ffffffff",
            INIT_04 => X"00001e8200000000000016270000000000003f8a000000000000130400000000",
            INIT_05 => X"ffffe587ffffffff0000227900000000fffffbafffffffff0000289b00000000",
            INIT_06 => X"00002dc400000000000002f500000000ffffe951ffffffff00000b3700000000",
            INIT_07 => X"fffff522fffffffffffffa4dffffffff00002cfe0000000000002d4700000000",
            INIT_08 => X"0000002c000000000000004a000000000000004a00000000ffffffd0ffffffff",
            INIT_09 => X"0000007e00000000000000170000000000000027000000000000006600000000",
            INIT_0A => X"0000000500000000ffffffdafffffffffffffff3ffffffff0000001e00000000",
            INIT_0B => X"0000000c00000000fffffff6ffffffff0000000400000000ffffffe8ffffffff",
            INIT_0C => X"fffffff4ffffffff00000017000000000000001d00000000ffffffe7ffffffff",
            INIT_0D => X"0000000e00000000ffffffe7ffffffffffffffdeffffffffffffffecffffffff",
            INIT_0E => X"000000250000000000000009000000000000000000000000ffffffe1ffffffff",
            INIT_0F => X"000000270000000000000036000000000000001b000000000000004700000000",
            INIT_10 => X"0000000200000000000000040000000000000025000000000000002c00000000",
            INIT_11 => X"fffffffaffffffff0000002c00000000fffffff0fffffffffffffff5ffffffff",
            INIT_12 => X"0000002200000000000000030000000000000027000000000000002200000000",
            INIT_13 => X"ffffffdaffffffffffffffe7ffffffffffffffd8ffffffff0000000200000000",
            INIT_14 => X"ffffffddffffffffffffffe0fffffffffffffff6ffffffffffffffd9ffffffff",
            INIT_15 => X"ffffffceffffffff0000002600000000ffffffe8fffffffffffffffbffffffff",
            INIT_16 => X"0000000a00000000ffffffdcffffffffffffffeeffffffffffffffd6ffffffff",
            INIT_17 => X"ffffffe9ffffffffffffffebffffffff0000001000000000fffffff8ffffffff",
            INIT_18 => X"fffffff5ffffffff0000000d00000000ffffffe7fffffffffffffff2ffffffff",
            INIT_19 => X"0000002900000000fffffff3ffffffff0000000a000000000000002300000000",
            INIT_1A => X"ffffffeaffffffff00000003000000000000000900000000ffffffcaffffffff",
            INIT_1B => X"0000005d000000000000001c0000000000000012000000000000003b00000000",
            INIT_1C => X"ffffffc8ffffffffffffffceffffffffffffffefffffffff0000000b00000000",
            INIT_1D => X"ffffffb6ffffffffffffffa4ffffffffffffffe2fffffffffffffff9ffffffff",
            INIT_1E => X"fffffff6ffffffffffffffdaffffffffffffff94ffffffffffffff7bffffffff",
            INIT_1F => X"0000002200000000ffffffe5ffffffffffffffdfffffffff0000000700000000",
            INIT_20 => X"0000004b0000000000000002000000000000001100000000ffffffdbffffffff",
            INIT_21 => X"fffffff6ffffffff0000003b00000000fffffffaffffffff0000001b00000000",
            INIT_22 => X"0000000200000000fffffffdffffffff00000017000000000000000c00000000",
            INIT_23 => X"0000002a000000000000000600000000fffffff9ffffffff0000000a00000000",
            INIT_24 => X"00000003000000000000002300000000ffffffe8ffffffffffffffe4ffffffff",
            INIT_25 => X"ffffffd4fffffffffffffff1ffffffffffffffe2fffffffffffffff3ffffffff",
            INIT_26 => X"0000002b00000000ffffffc3ffffffffffffffe4fffffffffffffffaffffffff",
            INIT_27 => X"0000006900000000000000650000000000000010000000000000000d00000000",
            INIT_28 => X"0000003c000000000000003e0000000000000062000000000000001f00000000",
            INIT_29 => X"0000001500000000000000370000000000000047000000000000004200000000",
            INIT_2A => X"ffffffeaffffffffffffffe6ffffffff0000000f000000000000003a00000000",
            INIT_2B => X"ffffff8fffffffffffffffcfffffffffffffffcbffffffffffffffb2ffffffff",
            INIT_2C => X"0000000c000000000000001f000000000000003000000000fffffffaffffffff",
            INIT_2D => X"000000f10000000000000044000000000000007200000000000000ec00000000",
            INIT_2E => X"ffffffe0ffffffffffffffeaffffffff0000003600000000000000a700000000",
            INIT_2F => X"ffffffeffffffffffffffff0ffffffffffffffd0ffffffff0000002000000000",
            INIT_30 => X"0000000d00000000fffffffcffffffffffffffebffffffffffffffc7ffffffff",
            INIT_31 => X"fffffff9ffffffffffffffc9ffffffffffffffe6fffffffffffffff0ffffffff",
            INIT_32 => X"fffffff8ffffffffffffffd5ffffffffffffffd9ffffffffffffffc3ffffffff",
            INIT_33 => X"00000008000000000000001c00000000ffffffeeffffffff0000001200000000",
            INIT_34 => X"ffffffe4ffffffff0000000b000000000000002900000000ffffffe4ffffffff",
            INIT_35 => X"00000000000000000000000000000000ffffffe8ffffffff0000001d00000000",
            INIT_36 => X"ffffffa1ffffffffffffffc3ffffffffffffffeaffffffffffffffc2ffffffff",
            INIT_37 => X"000000110000000000000015000000000000001400000000ffffffcaffffffff",
            INIT_38 => X"ffffffc4ffffffff0000002f0000000000000002000000000000000600000000",
            INIT_39 => X"000000030000000000000012000000000000002a00000000ffffffc9ffffffff",
            INIT_3A => X"0000000900000000000000020000000000000021000000000000001600000000",
            INIT_3B => X"00000038000000000000000d00000000ffffffebfffffffffffffff3ffffffff",
            INIT_3C => X"00000000000000000000003f00000000fffffffbfffffffffffffff6ffffffff",
            INIT_3D => X"ffffffb2fffffffffffffff7fffffffffffffffaffffffffffffffbbffffffff",
            INIT_3E => X"ffffffd4ffffffff0000002a000000000000001300000000ffffffb6ffffffff",
            INIT_3F => X"0000004900000000ffffffecffffffff0000002d000000000000001000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003b000000000000000f00000000ffffffc1ffffffff0000000e00000000",
            INIT_41 => X"00000080000000000000000d0000000000000029000000000000002500000000",
            INIT_42 => X"0000001a00000000000000020000000000000051000000000000006500000000",
            INIT_43 => X"ffffffedffffffffffffffdeffffffff00000023000000000000000f00000000",
            INIT_44 => X"0000003d00000000ffffffe7ffffffffffffffbfffffffffffffffe1ffffffff",
            INIT_45 => X"0000000c000000000000005300000000fffffff6ffffffff0000001200000000",
            INIT_46 => X"ffffffefffffffff0000001d000000000000002e00000000fffffffdffffffff",
            INIT_47 => X"000000170000000000000013000000000000002e000000000000004600000000",
            INIT_48 => X"00000005000000000000000e000000000000000100000000fffffffeffffffff",
            INIT_49 => X"000000600000000000000053000000000000007100000000ffffffdbffffffff",
            INIT_4A => X"0000005d00000000000000280000000000000011000000000000001900000000",
            INIT_4B => X"0000002300000000ffffffe3ffffffff0000002400000000ffffffd8ffffffff",
            INIT_4C => X"ffffffdaffffffff0000000b0000000000000013000000000000001300000000",
            INIT_4D => X"ffffffbcffffffffffffffd7ffffffff00000010000000000000000e00000000",
            INIT_4E => X"ffffffffffffffff000000150000000000000027000000000000000800000000",
            INIT_4F => X"00000043000000000000006e0000000000000066000000000000002800000000",
            INIT_50 => X"0000001e000000000000002b00000000fffffff3ffffffff0000000a00000000",
            INIT_51 => X"000000060000000000000007000000000000000e00000000fffffff3ffffffff",
            INIT_52 => X"fffffffcffffffff0000001e00000000fffffff1ffffffff0000005100000000",
            INIT_53 => X"0000001200000000ffffffe2ffffffff0000001b000000000000000c00000000",
            INIT_54 => X"ffffffcbffffffffffffffe2ffffffff0000000f00000000fffffff9ffffffff",
            INIT_55 => X"ffffffd4ffffffffffffffaafffffffffffffff1ffffffffffffffc7ffffffff",
            INIT_56 => X"ffffffdaffffffffffffffbdffffffffffffffa0ffffffffffffffd5ffffffff",
            INIT_57 => X"ffffff96ffffffffffffff9dffffffffffffffb9ffffffffffffffbcffffffff",
            INIT_58 => X"ffffffb4ffffffffffffffbfffffffffffffff91ffffffffffffffa8ffffffff",
            INIT_59 => X"0000000500000000ffffffedffffffff00000002000000000000000300000000",
            INIT_5A => X"ffffffefffffffffffffffecfffffffffffffff8ffffffffffffffdbffffffff",
            INIT_5B => X"0000001e00000000000000500000000000000030000000000000000800000000",
            INIT_5C => X"0000006b0000000000000036000000000000004e000000000000006400000000",
            INIT_5D => X"fffffffdffffffff000000340000000000000044000000000000005d00000000",
            INIT_5E => X"00000029000000000000001000000000ffffffffffffffff0000000600000000",
            INIT_5F => X"0000002a00000000fffffffbffffffff00000001000000000000001c00000000",
            INIT_60 => X"00000020000000000000002e0000000000000031000000000000000f00000000",
            INIT_61 => X"000000340000000000000020000000000000002d000000000000002d00000000",
            INIT_62 => X"0000002300000000ffffffcfffffffffffffffd5ffffffffffffffdfffffffff",
            INIT_63 => X"fffffff5fffffffffffffff8fffffffffffffff9ffffffffffffffcfffffffff",
            INIT_64 => X"000000320000000000000046000000000000005900000000ffffffedffffffff",
            INIT_65 => X"0000005700000000000000700000000000000055000000000000005800000000",
            INIT_66 => X"fffffff4ffffffffffffffebffffffff0000004d000000000000005b00000000",
            INIT_67 => X"00000016000000000000000b00000000fffffff3fffffffffffffffbffffffff",
            INIT_68 => X"0000001c000000000000001a00000000ffffffe6ffffffff0000000200000000",
            INIT_69 => X"ffffffe6fffffffffffffffdfffffffffffffff6ffffffff0000000700000000",
            INIT_6A => X"fffffffbfffffffffffffff8fffffffffffffffcffffffffffffffe9ffffffff",
            INIT_6B => X"0000001b000000000000000800000000ffffffeeffffffff0000001a00000000",
            INIT_6C => X"fffffff7ffffffff0000001400000000fffffff2fffffffffffffffaffffffff",
            INIT_6D => X"ffffffceffffffffffffffe0ffffffffffffffeffffffffffffffffaffffffff",
            INIT_6E => X"ffffffa9fffffffffffffff4ffffffffffffffc9ffffffffffffffd8ffffffff",
            INIT_6F => X"ffffffb2ffffffffffffff93ffffffffffffffd5ffffffffffffffa7ffffffff",
            INIT_70 => X"ffffff80ffffffffffffff73ffffffffffffff9bffffffffffffffceffffffff",
            INIT_71 => X"0000000300000000ffffff97ffffffffffffffa9ffffffffffffff83ffffffff",
            INIT_72 => X"0000000b000000000000000100000000ffffffdbfffffffffffffffcffffffff",
            INIT_73 => X"ffffffe1ffffffff0000000a0000000000000009000000000000001e00000000",
            INIT_74 => X"ffffffc3fffffffffffffff2ffffffffffffffadffffffffffffff8affffffff",
            INIT_75 => X"ffffffb1ffffffffffffff98ffffffffffffffc9ffffffffffffffacffffffff",
            INIT_76 => X"000000170000000000000000000000000000001d00000000ffffff9cffffffff",
            INIT_77 => X"ffffffdaffffffff0000001800000000fffffff5ffffffff0000000600000000",
            INIT_78 => X"0000001c000000000000002300000000ffffffe3fffffffffffffff4ffffffff",
            INIT_79 => X"ffffffe7fffffffffffffff0ffffffffffffffe3ffffffff0000000800000000",
            INIT_7A => X"0000001e00000000fffffff5ffffffff0000000200000000ffffffe8ffffffff",
            INIT_7B => X"ffffffe7fffffffffffffffdffffffff00000037000000000000002800000000",
            INIT_7C => X"ffffffacffffffffffffffb9ffffffffffffffbeffffffffffffffe2ffffffff",
            INIT_7D => X"0000001700000000000000060000000000000011000000000000001800000000",
            INIT_7E => X"0000002500000000000000550000000000000027000000000000001100000000",
            INIT_7F => X"fffffff0ffffffff0000000200000000ffffffd7ffffffff0000002800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE0;


    MEM_IWGHT_LAYER1_INSTANCE1 : if BRAM_NAME = "iwght_layer1_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff8ffffffffffffffd5ffffffffffffffe9ffffffffffffffd5ffffffff",
            INIT_01 => X"000000270000000000000019000000000000001a000000000000000700000000",
            INIT_02 => X"ffffffdbffffffff0000000000000000ffffffe8ffffffff0000001900000000",
            INIT_03 => X"0000001700000000ffffffeaffffffffffffffe6ffffffffffffffdbffffffff",
            INIT_04 => X"00000004000000000000002500000000ffffffffffffffffffffffd8ffffffff",
            INIT_05 => X"0000003f00000000000000410000000000000032000000000000001200000000",
            INIT_06 => X"ffffffdcffffffff0000003700000000fffffffbffffffff0000002700000000",
            INIT_07 => X"ffffffc6ffffffffffffffdbffffffffffffffe9ffffffffffffffc5ffffffff",
            INIT_08 => X"0000000000000000fffffff9ffffffff0000002000000000ffffffb8ffffffff",
            INIT_09 => X"fffffffaffffffffffffffd6ffffffffffffffe0ffffffffffffffdcffffffff",
            INIT_0A => X"ffffffd2ffffffff0000000c000000000000000f00000000ffffffdcffffffff",
            INIT_0B => X"fffffffaffffffff00000009000000000000001200000000ffffffecffffffff",
            INIT_0C => X"ffffffffffffffff00000028000000000000001c000000000000000e00000000",
            INIT_0D => X"fffffff0ffffffffffffffcaffffffff00000006000000000000002d00000000",
            INIT_0E => X"ffffffedfffffffffffffffbffffffffffffffd3ffffffffffffffe4ffffffff",
            INIT_0F => X"ffffffe1ffffffff0000001300000000fffffff6ffffffffffffffe8ffffffff",
            INIT_10 => X"0000001a00000000fffffffcfffffffffffffff0ffffffff0000001300000000",
            INIT_11 => X"ffffffb2ffffffffffffffa8ffffffffffffffa9fffffffffffffff8ffffffff",
            INIT_12 => X"ffffff8bffffffffffffffb8ffffffffffffff55ffffffffffffff87ffffffff",
            INIT_13 => X"0000001800000000fffffffbffffffffffffff8fffffffffffffff92ffffffff",
            INIT_14 => X"fffffff9ffffffff000000070000000000000007000000000000003000000000",
            INIT_15 => X"fffffffbffffffff00000048000000000000004a000000000000003e00000000",
            INIT_16 => X"ffffffb3ffffffffffffffe2ffffffffffffffe9ffffffffffffffdaffffffff",
            INIT_17 => X"ffffffedffffffff0000001e00000000fffffffeffffffffffffffe3ffffffff",
            INIT_18 => X"ffffffd9ffffffffffffffe5ffffffff0000003d00000000fffffff0ffffffff",
            INIT_19 => X"ffffffc3ffffffffffffffdeffffffff0000000400000000ffffffffffffffff",
            INIT_1A => X"0000001f00000000fffffff0fffffffffffffffbffffffffffffffdaffffffff",
            INIT_1B => X"0000002d00000000ffffffeaffffffffffffffcffffffffffffffffbffffffff",
            INIT_1C => X"0000003f00000000ffffffddfffffffffffffff4fffffffffffffffbffffffff",
            INIT_1D => X"00000039000000000000001400000000ffffffb2ffffffff0000000300000000",
            INIT_1E => X"fffffffaffffffffffffffd9ffffffffffffffcbffffffff0000002c00000000",
            INIT_1F => X"fffffff1fffffffffffffffdffffffff0000002300000000fffffff6ffffffff",
            INIT_20 => X"ffffffc7fffffffffffffffaffffffff0000004c00000000ffffffe2ffffffff",
            INIT_21 => X"ffffffcaffffffff0000001f000000000000003900000000fffffffaffffffff",
            INIT_22 => X"ffffffeeffffffffffffffe6ffffffff0000001a00000000ffffffeeffffffff",
            INIT_23 => X"0000000e000000000000004600000000fffffff1fffffffffffffffbffffffff",
            INIT_24 => X"ffffffcfffffffff00000043000000000000000200000000ffffffbaffffffff",
            INIT_25 => X"0000001f0000000000000001000000000000001500000000ffffffc1ffffffff",
            INIT_26 => X"fffffffeffffffffffffffdeffffffffffffffe9ffffffff0000002300000000",
            INIT_27 => X"ffffffefffffffffffffffcfffffffffffffffd0ffffffff0000002b00000000",
            INIT_28 => X"ffffffe6ffffffffffffffebfffffffffffffffcfffffffffffffff4ffffffff",
            INIT_29 => X"00000000000000000000001700000000fffffff6ffffffff0000000300000000",
            INIT_2A => X"ffffffb8ffffffff0000004e00000000000000ba000000000000005900000000",
            INIT_2B => X"fffffff2ffffffff00000034000000000000009f000000000000009800000000",
            INIT_2C => X"0000001e000000000000005800000000ffffffddffffffff0000002300000000",
            INIT_2D => X"00000003000000000000005a000000000000004800000000ffffffc4ffffffff",
            INIT_2E => X"fffffff0ffffffffffffffe6ffffffff0000005a00000000ffffff92ffffffff",
            INIT_2F => X"0000001600000000ffffffe3ffffffff00000015000000000000000300000000",
            INIT_30 => X"0000000b00000000ffffffe6ffffffff00000008000000000000003100000000",
            INIT_31 => X"00000012000000000000004a00000000ffffffffffffffffffffffadffffffff",
            INIT_32 => X"ffffffe9ffffffff0000003e000000000000000e00000000ffffffabffffffff",
            INIT_33 => X"00000029000000000000003900000000ffffffd5fffffffffffffff1ffffffff",
            INIT_34 => X"00000044000000000000003e00000000ffffffe4ffffffffffffffe0ffffffff",
            INIT_35 => X"00000054000000000000003c000000000000002a00000000fffffffdffffffff",
            INIT_36 => X"ffffffd8ffffffff00000051000000000000000000000000ffffffd5ffffffff",
            INIT_37 => X"0000000800000000ffffffe6ffffffffffffffeefffffffffffffff7ffffffff",
            INIT_38 => X"0000003b000000000000003100000000ffffffd0fffffffffffffff9ffffffff",
            INIT_39 => X"00000001000000000000001800000000ffffffb3ffffffffffffff8bffffffff",
            INIT_3A => X"0000006300000000ffffffddffffffff0000000b000000000000001e00000000",
            INIT_3B => X"0000005e00000000ffffffd7ffffffffffffffdfffffffff0000009200000000",
            INIT_3C => X"ffffffddffffffffffffff9affffffffffffffceffffffff0000000500000000",
            INIT_3D => X"ffffff74ffffffffffffffacffffffffffffff3fffffffffffffff7affffffff",
            INIT_3E => X"fffffff3ffffffff0000000a000000000000001200000000ffffff72ffffffff",
            INIT_3F => X"ffffffe3ffffffff000000240000000000000016000000000000001f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffffdffffffff0000002200000000ffffffecffffffff0000000500000000",
            INIT_41 => X"0000001000000000000000130000000000000026000000000000000f00000000",
            INIT_42 => X"0000000f000000000000000f000000000000000100000000ffffffdbffffffff",
            INIT_43 => X"ffffffeeffffffffffffffe3ffffffff0000000f00000000fffffffaffffffff",
            INIT_44 => X"fffffffdffffffffffffffb6ffffffffffffffcaffffffffffffffe4ffffffff",
            INIT_45 => X"fffffffefffffffffffffffbfffffffffffffffbffffffff0000001600000000",
            INIT_46 => X"0000003600000000000000130000000000000000000000000000000000000000",
            INIT_47 => X"ffffffacffffffffffffffd2ffffffffffffffb9ffffffff0000000d00000000",
            INIT_48 => X"00000004000000000000000c00000000ffffffbfffffffffffffffc8ffffffff",
            INIT_49 => X"fffffff7fffffffffffffff3ffffffff0000002f000000000000000800000000",
            INIT_4A => X"00000005000000000000000600000000fffffffaffffffff0000000500000000",
            INIT_4B => X"fffffff8ffffffffffffffe8ffffffffffffffe4ffffffffffffffdcffffffff",
            INIT_4C => X"00000000000000000000000900000000ffffffd9fffffffffffffff3ffffffff",
            INIT_4D => X"00000014000000000000002d0000000000000038000000000000002400000000",
            INIT_4E => X"ffffffcdffffffffffffffbcffffffffffffffbaffffffffffffffdeffffffff",
            INIT_4F => X"ffffffb5ffffffffffffffe8ffffffffffffffcdffffffffffffff97ffffffff",
            INIT_50 => X"ffffffb5ffffffffffffffd0ffffffffffffffcaffffffffffffffc6ffffffff",
            INIT_51 => X"ffffffecffffffffffffffc0ffffffffffffffaaffffffffffffffccffffffff",
            INIT_52 => X"00000017000000000000000f0000000000000000000000000000000200000000",
            INIT_53 => X"0000001200000000fffffff8ffffffff00000007000000000000001c00000000",
            INIT_54 => X"0000002000000000fffffff4ffffffff0000000d000000000000000300000000",
            INIT_55 => X"0000001b00000000000000000000000000000013000000000000002800000000",
            INIT_56 => X"ffffffd4ffffffffffffffe2ffffffffffffffecfffffffffffffffaffffffff",
            INIT_57 => X"00000027000000000000000b000000000000001e00000000fffffff0ffffffff",
            INIT_58 => X"000000050000000000000012000000000000000900000000fffffffbffffffff",
            INIT_59 => X"ffffffd4ffffffffffffffe2ffffffff00000003000000000000000900000000",
            INIT_5A => X"fffffff4fffffffffffffff4fffffffffffffffeffffffffffffffdfffffffff",
            INIT_5B => X"ffffffeaffffffff0000000c00000000ffffffe5ffffffff0000001800000000",
            INIT_5C => X"ffffffb9ffffffffffffffe3ffffffff0000000500000000ffffffbeffffffff",
            INIT_5D => X"ffffff8efffffffffffffffcffffffff0000001b000000000000001200000000",
            INIT_5E => X"ffffffaaffffffffffffffe5ffffffffffffffa5ffffffffffffff99ffffffff",
            INIT_5F => X"ffffffcfffffffffffffffd0ffffffffffffffbbffffffffffffffa4ffffffff",
            INIT_60 => X"ffffffbdffffffffffffffc9ffffffffffffff73ffffffffffffffd3ffffffff",
            INIT_61 => X"ffffffc1ffffffffffffffd7ffffffffffffffecffffffffffffffb9ffffffff",
            INIT_62 => X"0000000d00000000ffffffd9fffffffffffffffaffffffffffffff8bffffffff",
            INIT_63 => X"0000001d0000000000000005000000000000001a000000000000001500000000",
            INIT_64 => X"0000000f00000000fffffffcffffffffffffffeaffffffff0000001700000000",
            INIT_65 => X"0000001700000000ffffffe9ffffffff0000002c000000000000000100000000",
            INIT_66 => X"0000001a00000000000000090000000000000018000000000000000c00000000",
            INIT_67 => X"fffffff4ffffffff0000000c0000000000000003000000000000000700000000",
            INIT_68 => X"ffffffe2fffffffffffffff2ffffffff00000020000000000000000800000000",
            INIT_69 => X"0000000900000000ffffffd7fffffffffffffff8fffffffffffffff0ffffffff",
            INIT_6A => X"0000000400000000fffffffdffffffffffffffeffffffffffffffffaffffffff",
            INIT_6B => X"ffffffbdffffffffffffff9effffffffffffff91ffffffff0000001400000000",
            INIT_6C => X"ffffffb9ffffffffffffffb6ffffffffffffffa7ffffffffffffffa7ffffffff",
            INIT_6D => X"0000000c000000000000002b00000000ffffffd8ffffffffffffffe3ffffffff",
            INIT_6E => X"fffffffcfffffffffffffff9ffffffff0000001400000000fffffff6ffffffff",
            INIT_6F => X"ffffffd0ffffffff000000050000000000000009000000000000001400000000",
            INIT_70 => X"ffffffcdffffffffffffffeeffffffffffffffeafffffffffffffffcffffffff",
            INIT_71 => X"fffffff7ffffffff0000001000000000ffffffe3ffffffffffffffc0ffffffff",
            INIT_72 => X"ffffff9bffffffff0000004a00000000ffffffe4ffffffffffffffdfffffffff",
            INIT_73 => X"ffffffddffffffff00000016000000000000002b00000000ffffffdfffffffff",
            INIT_74 => X"0000002c000000000000000d000000000000000c00000000ffffffe3ffffffff",
            INIT_75 => X"ffffffe8ffffffff0000001b0000000000000027000000000000000400000000",
            INIT_76 => X"ffffffdfffffffffffffffe4ffffffff0000000700000000fffffff6ffffffff",
            INIT_77 => X"0000001a00000000fffffff4ffffffffffffffedffffffffffffffd6ffffffff",
            INIT_78 => X"0000002200000000fffffff6ffffffff0000001e000000000000000a00000000",
            INIT_79 => X"fffffff9ffffffff000000440000000000000005000000000000002900000000",
            INIT_7A => X"fffffffdfffffffffffffffaffffffff0000001a00000000fffffff1ffffffff",
            INIT_7B => X"0000003100000000fffffffbffffffff0000001a000000000000001500000000",
            INIT_7C => X"0000001d000000000000001500000000ffffffdfffffffffffffffefffffffff",
            INIT_7D => X"ffffffbbffffffff0000000500000000ffffffedffffffffffffffe6ffffffff",
            INIT_7E => X"ffffffabffffffffffffffe6fffffffffffffff2fffffffffffffff1ffffffff",
            INIT_7F => X"00000040000000000000000f00000000ffffffe3ffffffffffffff9dffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE1;


    MEM_IWGHT_LAYER1_INSTANCE2 : if BRAM_NAME = "iwght_layer1_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff2ffffffff00000012000000000000002200000000fffffff3ffffffff",
            INIT_01 => X"0000000f00000000fffffff9ffffffff0000002600000000fffffff4ffffffff",
            INIT_02 => X"fffffff5fffffffffffffffbffffffff00000020000000000000000200000000",
            INIT_03 => X"0000000500000000ffffffe2ffffffffffffffd6ffffffff0000000400000000",
            INIT_04 => X"ffffffe7ffffffffffffffc5fffffffffffffff1ffffffff0000001800000000",
            INIT_05 => X"00000042000000000000003c00000000ffffffc7ffffffffffffffc0ffffffff",
            INIT_06 => X"ffffffccffffffffffffffd7ffffffffffffffcbffffffff0000001e00000000",
            INIT_07 => X"0000002a00000000ffffffe1ffffffff0000001f000000000000001300000000",
            INIT_08 => X"ffffff96ffffffffffffffc4ffffffff00000018000000000000003b00000000",
            INIT_09 => X"ffffffdbffffffff00000009000000000000002f00000000ffffffb6ffffffff",
            INIT_0A => X"ffffffeffffffffffffffff7ffffffff00000028000000000000003300000000",
            INIT_0B => X"0000001400000000ffffffd3ffffffffffffffe2fffffffffffffff9ffffffff",
            INIT_0C => X"0000004c00000000000000360000000000000017000000000000001000000000",
            INIT_0D => X"00000000000000000000002b0000000000000000000000000000001400000000",
            INIT_0E => X"fffffff3ffffffff0000001c000000000000000a00000000fffffff2ffffffff",
            INIT_0F => X"fffffff7fffffffffffffffcfffffffffffffffcffffffffffffffefffffffff",
            INIT_10 => X"ffffffe7ffffffffffffffd7ffffffffffffffe2fffffffffffffff4ffffffff",
            INIT_11 => X"ffffffc6ffffffffffffffc9ffffffffffffffacffffffffffffffe7ffffffff",
            INIT_12 => X"00000004000000000000001f00000000ffffffeeffffffffffffffddffffffff",
            INIT_13 => X"0000000a00000000000000390000000000000020000000000000002500000000",
            INIT_14 => X"fffffffeffffffff000000170000000000000008000000000000000000000000",
            INIT_15 => X"ffffffedffffffffffffffdaffffffff0000000800000000fffffff2ffffffff",
            INIT_16 => X"ffffffbdffffffffffffffc6ffffffffffffffb7ffffffffffffffdcffffffff",
            INIT_17 => X"0000001600000000ffffffeefffffffffffffffeffffffffffffffb8ffffffff",
            INIT_18 => X"ffffffeaffffffffffffffb7ffffffffffffffc9fffffffffffffff0ffffffff",
            INIT_19 => X"0000000600000000ffffffd2ffffffffffffffe4ffffffffffffffddffffffff",
            INIT_1A => X"0000000a000000000000000200000000ffffffa0ffffffff0000000100000000",
            INIT_1B => X"ffffffefffffffff00000009000000000000001a00000000fffffff4ffffffff",
            INIT_1C => X"ffffffbcffffffff0000000a000000000000001e000000000000003a00000000",
            INIT_1D => X"0000002100000000fffffffbfffffffffffffff0ffffffffffffffd8ffffffff",
            INIT_1E => X"0000003300000000000000000000000000000002000000000000000900000000",
            INIT_1F => X"ffffffefffffffffffffffe6ffffffffffffffcaffffffffffffffdeffffffff",
            INIT_20 => X"0000002f000000000000000a000000000000000b000000000000001500000000",
            INIT_21 => X"00000011000000000000000900000000ffffffffffffffff0000000700000000",
            INIT_22 => X"ffffffdeffffffff0000000b000000000000000c00000000ffffffefffffffff",
            INIT_23 => X"0000001400000000ffffffcaffffffff0000000000000000ffffffa9ffffffff",
            INIT_24 => X"0000003000000000ffffffd3ffffffffffffffd8ffffffff0000000100000000",
            INIT_25 => X"0000002800000000ffffffb6ffffffffffffffb7fffffffffffffff9ffffffff",
            INIT_26 => X"0000002d00000000ffffffd1ffffffff00000067000000000000002300000000",
            INIT_27 => X"ffffffddffffffffffffffc4ffffffffffffffc2ffffffff0000003200000000",
            INIT_28 => X"0000002b00000000ffffffa4ffffffff00000039000000000000003e00000000",
            INIT_29 => X"ffffffc0ffffffffffffffe7ffffffffffffff87ffffffffffffffa5ffffffff",
            INIT_2A => X"0000002c0000000000000013000000000000001400000000fffffff6ffffffff",
            INIT_2B => X"0000001700000000ffffffffffffffff0000001b000000000000000600000000",
            INIT_2C => X"0000002b00000000fffffff9ffffffffffffffd9ffffffffffffffefffffffff",
            INIT_2D => X"ffffffe1fffffffffffffff3ffffffff00000027000000000000002c00000000",
            INIT_2E => X"0000001800000000ffffffe6ffffffffffffffd2ffffffff0000002500000000",
            INIT_2F => X"fffffff2ffffffffffffffdcffffffffffffffeaffffffffffffffe5ffffffff",
            INIT_30 => X"fffffffafffffffffffffff9ffffffff0000000500000000ffffffe1ffffffff",
            INIT_31 => X"0000000000000000000000220000000000000006000000000000001c00000000",
            INIT_32 => X"ffffffe3fffffffffffffff8fffffffffffffff3ffffffff0000001900000000",
            INIT_33 => X"ffffff9affffffffffffffe7ffffffffffffffceffffffffffffffd0ffffffff",
            INIT_34 => X"ffffffe0ffffffffffffffccffffffffffffffa1fffffffffffffff2ffffffff",
            INIT_35 => X"fffffffeffffffffffffffeaffffffffffffffeaffffffffffffffcdffffffff",
            INIT_36 => X"ffffffdbfffffffffffffffffffffffffffffffbffffffff0000001700000000",
            INIT_37 => X"0000001800000000ffffffecffffffffffffffdafffffffffffffff1ffffffff",
            INIT_38 => X"0000000f000000000000000800000000fffffffcfffffffffffffffcffffffff",
            INIT_39 => X"ffffffcefffffffffffffffbffffffffffffffe9ffffffffffffffe0ffffffff",
            INIT_3A => X"ffffffd5ffffffffffffff5effffffffffffffd6ffffffff0000002700000000",
            INIT_3B => X"ffffffa7ffffffffffffffb8ffffffffffffff76ffffffffffffff7bffffffff",
            INIT_3C => X"ffffffdbffffffffffffffd2ffffffffffffffefffffffffffffffd7ffffffff",
            INIT_3D => X"ffffffd9ffffffffffffffdbffffffffffffffe5ffffffffffffff90ffffffff",
            INIT_3E => X"0000002e000000000000001e00000000ffffffdefffffffffffffffdffffffff",
            INIT_3F => X"0000000100000000ffffffedffffffff00000029000000000000000b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff4ffffffffffffffe3ffffffffffffffd9ffffffff0000000700000000",
            INIT_41 => X"00000033000000000000001c000000000000001e000000000000001800000000",
            INIT_42 => X"ffffffddfffffffffffffffdffffffff0000000a000000000000002200000000",
            INIT_43 => X"000000250000000000000012000000000000002900000000ffffffddffffffff",
            INIT_44 => X"0000001000000000fffffffeffffffff00000005000000000000002000000000",
            INIT_45 => X"ffffffcbffffffffffffffe1ffffffffffffffeefffffffffffffffbffffffff",
            INIT_46 => X"0000000d00000000fffffff1fffffffffffffff1ffffffff0000001d00000000",
            INIT_47 => X"00000020000000000000001200000000ffffffedffffffff0000000400000000",
            INIT_48 => X"00000049000000000000004a0000000000000029000000000000001300000000",
            INIT_49 => X"ffffffc3fffffffffffffff1ffffffff00000044000000000000002200000000",
            INIT_4A => X"ffffffd8ffffffffffffffe9ffffffffffffffccffffffffffffffa2ffffffff",
            INIT_4B => X"ffffffbdffffffffffffffd9fffffffffffffff1ffffffffffffffd9ffffffff",
            INIT_4C => X"0000007f000000000000003200000000ffffffa9ffffffff0000006a00000000",
            INIT_4D => X"ffffff8cffffffff0000005a000000000000006e00000000ffffff8cffffffff",
            INIT_4E => X"ffffffdfffffffff00000022000000000000000d000000000000007000000000",
            INIT_4F => X"0000000200000000fffffff5fffffffffffffff1ffffffff0000001d00000000",
            INIT_50 => X"ffffffebffffffff0000002d00000000ffffffdcffffffff0000000700000000",
            INIT_51 => X"ffffffeaffffffffffffffe5ffffffff0000000b00000000ffffffecffffffff",
            INIT_52 => X"fffffffdffffffffffffffe3ffffffffffffffceffffffff0000002100000000",
            INIT_53 => X"0000002e00000000ffffffddffffffff0000000100000000fffffff7ffffffff",
            INIT_54 => X"ffffffecffffffff000000150000000000000009000000000000001800000000",
            INIT_55 => X"00000025000000000000000900000000ffffffeeffffffff0000002c00000000",
            INIT_56 => X"ffffffe6ffffffff0000002900000000ffffffddffffffffffffffd3ffffffff",
            INIT_57 => X"fffffff7ffffffffffffffd3ffffffff00000011000000000000000200000000",
            INIT_58 => X"00000044000000000000001600000000ffffffa3ffffffff0000005000000000",
            INIT_59 => X"0000000c000000000000001e00000000ffffffe9ffffffffffffffe4ffffffff",
            INIT_5A => X"ffffffdcfffffffffffffff5ffffffff0000002f00000000ffffffe4ffffffff",
            INIT_5B => X"fffffffdfffffffffffffffefffffffffffffffbfffffffffffffffbffffffff",
            INIT_5C => X"00000000000000000000001600000000fffffffcffffffff0000002100000000",
            INIT_5D => X"fffffff8ffffffff0000002200000000ffffffe6fffffffffffffff0ffffffff",
            INIT_5E => X"00000052000000000000006000000000ffffffb7ffffffff0000007600000000",
            INIT_5F => X"ffffffb8ffffffff00000023000000000000005200000000ffffff78ffffffff",
            INIT_60 => X"0000001400000000ffffffb4ffffffff00000004000000000000006f00000000",
            INIT_61 => X"ffffff90ffffffffffffffebffffffffffffff8cffffffffffffffaaffffffff",
            INIT_62 => X"00000000000000000000001e00000000ffffffcbffffffffffffff9fffffffff",
            INIT_63 => X"fffffff0ffffffffffffffedffffffff0000000200000000fffffffaffffffff",
            INIT_64 => X"fffffffdffffffffffffffddffffffffffffffddffffffff0000002500000000",
            INIT_65 => X"0000000f00000000ffffffc9ffffffffffffffddffffffff0000002700000000",
            INIT_66 => X"ffffffd9ffffffff0000002900000000ffffffd3ffffffffffffffdaffffffff",
            INIT_67 => X"ffffffe5ffffffffffffffd9ffffffff0000002600000000ffffffe4ffffffff",
            INIT_68 => X"00000005000000000000001000000000fffffff1ffffffff0000003300000000",
            INIT_69 => X"fffffff2ffffffffffffffe2ffffffff0000000500000000fffffffaffffffff",
            INIT_6A => X"0000000700000000ffffffeefffffffffffffff9fffffffffffffff7ffffffff",
            INIT_6B => X"0000002000000000fffffffbffffffff00000009000000000000002900000000",
            INIT_6C => X"0000000b000000000000000200000000ffffffdaffffffff0000001500000000",
            INIT_6D => X"fffffff2fffffffffffffff5ffffffff0000000200000000ffffffffffffffff",
            INIT_6E => X"ffffffa9ffffffffffffff9bffffffffffffffe1fffffffffffffff5ffffffff",
            INIT_6F => X"ffffffd3ffffffffffffffb9ffffffffffffff9effffffffffffffcaffffffff",
            INIT_70 => X"0000002900000000fffffff9ffffffff0000001e00000000ffffffe6ffffffff",
            INIT_71 => X"000000600000000000000011000000000000000d000000000000002b00000000",
            INIT_72 => X"fffffff9ffffffffffffffd9ffffffffffffffe0ffffffff0000004b00000000",
            INIT_73 => X"0000002400000000ffffffecffffffffffffffeeffffffffffffffffffffffff",
            INIT_74 => X"0000002e00000000000000170000000000000032000000000000000a00000000",
            INIT_75 => X"fffffffaffffffff00000004000000000000001d000000000000001300000000",
            INIT_76 => X"0000001400000000000000200000000000000023000000000000002300000000",
            INIT_77 => X"0000001c000000000000000800000000fffffffafffffffffffffff7ffffffff",
            INIT_78 => X"00000026000000000000002f000000000000002a000000000000000b00000000",
            INIT_79 => X"ffffffe7ffffffffffffffdbffffffffffffffe0ffffffffffffffd2ffffffff",
            INIT_7A => X"ffffffeaffffffff00000008000000000000001200000000ffffffd3ffffffff",
            INIT_7B => X"ffffffc9ffffffff0000000300000000ffffffadfffffffffffffff0ffffffff",
            INIT_7C => X"ffffff8affffffffffffffa4ffffffffffffffd1ffffffffffffffadffffffff",
            INIT_7D => X"0000001300000000ffffffd6ffffffffffffffbbffffffffffffffabffffffff",
            INIT_7E => X"00000006000000000000000a000000000000000400000000ffffffe0ffffffff",
            INIT_7F => X"ffffffeaffffffff0000001c000000000000001300000000fffffffeffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE2;


    MEM_IWGHT_LAYER1_INSTANCE3 : if BRAM_NAME = "iwght_layer1_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000006000000000000000200000000ffffffd5ffffffffffffffecffffffff",
            INIT_01 => X"00000011000000000000001600000000ffffffefffffffffffffffd8ffffffff",
            INIT_02 => X"fffffffafffffffffffffffeffffffff0000003600000000ffffffd6ffffffff",
            INIT_03 => X"0000002500000000ffffffe5fffffffffffffff9ffffffff0000003e00000000",
            INIT_04 => X"ffffffeeffffffffffffffa3ffffffffffffff98ffffffff0000003800000000",
            INIT_05 => X"ffffff82ffffffffffffff99ffffffffffffff9effffffffffffffaaffffffff",
            INIT_06 => X"fffffff1ffffffffffffffffffffffffffffffabffffffffffffffb0ffffffff",
            INIT_07 => X"00000007000000000000000700000000fffffffcffffffffffffffceffffffff",
            INIT_08 => X"0000003a00000000000000090000000000000027000000000000001f00000000",
            INIT_09 => X"0000000d00000000000000320000000000000006000000000000000c00000000",
            INIT_0A => X"000000040000000000000025000000000000003b00000000ffffffe6ffffffff",
            INIT_0B => X"ffffffffffffffffffffffe6fffffffffffffff5fffffffffffffff7ffffffff",
            INIT_0C => X"000000130000000000000031000000000000000a00000000ffffffe5ffffffff",
            INIT_0D => X"0000001e000000000000000300000000fffffffbfffffffffffffffdffffffff",
            INIT_0E => X"ffffffdeffffffff0000002e0000000000000001000000000000004100000000",
            INIT_0F => X"ffffffcaffffffffffffffdeffffffffffffffcdffffffffffffffcbffffffff",
            INIT_10 => X"0000000b00000000ffffffd3fffffffffffffffeffffffff0000001100000000",
            INIT_11 => X"ffffffcfffffffffffffffbdfffffffffffffff3fffffffffffffff7ffffffff",
            INIT_12 => X"ffffffa9ffffffffffffffbcffffffffffffffeaffffffffffffffdbffffffff",
            INIT_13 => X"ffffffb2ffffffffffffff88ffffffffffffffc2ffffffffffffffa9ffffffff",
            INIT_14 => X"ffffffbdffffffff0000003d0000000000000044000000000000001200000000",
            INIT_15 => X"0000003600000000ffffff9effffffff00000042000000000000004f00000000",
            INIT_16 => X"0000001d000000000000001300000000fffffff4ffffffff0000007400000000",
            INIT_17 => X"ffffffddffffffff0000001e00000000ffffffefffffffff0000000200000000",
            INIT_18 => X"00000028000000000000000a000000000000001c00000000ffffffd6ffffffff",
            INIT_19 => X"00000027000000000000003200000000ffffffebffffffff0000004b00000000",
            INIT_1A => X"ffffffc3ffffffff0000002200000000fffffff5ffffffffffffffcaffffffff",
            INIT_1B => X"ffffffe2fffffffffffffff8ffffffff0000000400000000fffffff5ffffffff",
            INIT_1C => X"0000000a00000000fffffffbffffffffffffffe3ffffffff0000000700000000",
            INIT_1D => X"ffffffffffffffffffffffebffffffff0000001c00000000fffffff6ffffffff",
            INIT_1E => X"ffffffedfffffffffffffffbffffffffffffffe1ffffffffffffffedffffffff",
            INIT_1F => X"ffffffdafffffffffffffff2fffffffffffffff5ffffffffffffffe5ffffffff",
            INIT_20 => X"ffffffefffffffffffffffe6ffffffff0000001300000000ffffffe1ffffffff",
            INIT_21 => X"0000000700000000000000090000000000000010000000000000001c00000000",
            INIT_22 => X"0000001700000000fffffffdffffffffffffffffffffffff0000002e00000000",
            INIT_23 => X"ffffffe7ffffffff00000000000000000000001e000000000000000700000000",
            INIT_24 => X"00000007000000000000001400000000ffffffdfffffffffffffffc9ffffffff",
            INIT_25 => X"fffffff0fffffffffffffffaffffffff0000001500000000ffffffd3ffffffff",
            INIT_26 => X"ffffffbfffffffff000000580000000000000070000000000000001b00000000",
            INIT_27 => X"0000004700000000fffffffeffffffff00000042000000000000004800000000",
            INIT_28 => X"00000010000000000000001900000000ffffff97ffffffff0000009c00000000",
            INIT_29 => X"ffffffdffffffffffffffffdffffffffffffffd9ffffffffffffffe7ffffffff",
            INIT_2A => X"ffffffdfffffffff00000003000000000000002100000000ffffffecffffffff",
            INIT_2B => X"0000000c00000000ffffffeeffffffff00000008000000000000001c00000000",
            INIT_2C => X"ffffffdfffffffff0000001300000000ffffffceffffffffffffffc3ffffffff",
            INIT_2D => X"ffffffdeffffffff000000150000000000000035000000000000000400000000",
            INIT_2E => X"ffffffebffffffff00000004000000000000001e000000000000002000000000",
            INIT_2F => X"0000000d000000000000000e00000000ffffffe0ffffffff0000000c00000000",
            INIT_30 => X"000000040000000000000017000000000000001e00000000ffffffd8ffffffff",
            INIT_31 => X"ffffffd0ffffffffffffffc2ffffffffffffffc9ffffffffffffffceffffffff",
            INIT_32 => X"0000000000000000ffffff82ffffffffffffffd1fffffffffffffff3ffffffff",
            INIT_33 => X"ffffff98ffffffffffffff7effffffffffffffbaffffffffffffffe4ffffffff",
            INIT_34 => X"ffffff94ffffffffffffffa3ffffffffffffff9bffffffffffffffa6ffffffff",
            INIT_35 => X"ffffffb9ffffffffffffffb1ffffffffffffffaaffffffffffffffcfffffffff",
            INIT_36 => X"ffffffdcffffffffffffffc1ffffffffffffffeaffffffffffffffddffffffff",
            INIT_37 => X"0000000c00000000ffffffbdffffffffffffffd6ffffffffffffffb5ffffffff",
            INIT_38 => X"00000009000000000000005f000000000000004600000000fffffffdffffffff",
            INIT_39 => X"ffffffa3fffffffffffffffcffffffffffffffe8ffffffff0000001d00000000",
            INIT_3A => X"fffffff1ffffffffffffffccffffffffffffffd1ffffffffffffffc3ffffffff",
            INIT_3B => X"000000280000000000000018000000000000000900000000fffffff0ffffffff",
            INIT_3C => X"ffffffecffffffff0000000f0000000000000020000000000000000700000000",
            INIT_3D => X"0000000200000000ffffffe3fffffffffffffff2ffffffffffffffd0ffffffff",
            INIT_3E => X"0000003000000000fffffff4ffffffff0000000d000000000000000700000000",
            INIT_3F => X"fffffff0ffffffff00000015000000000000000b000000000000003800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002200000000ffffffedffffffff0000000a000000000000000900000000",
            INIT_41 => X"ffffffeeffffffffffffffc9ffffffffffffffa0ffffffffffffffd0ffffffff",
            INIT_42 => X"0000003100000000000000340000000000000000000000000000000000000000",
            INIT_43 => X"0000000900000000fffffff5ffffffffffffffebffffffff0000002700000000",
            INIT_44 => X"0000002100000000ffffffebffffffff0000001500000000ffffffe7ffffffff",
            INIT_45 => X"0000001700000000fffffff0ffffffff00000010000000000000001d00000000",
            INIT_46 => X"0000001c00000000fffffffbffffffffffffffeeffffffff0000000c00000000",
            INIT_47 => X"ffffffecffffffffffffffdeffffffff00000009000000000000000000000000",
            INIT_48 => X"00000019000000000000000a00000000ffffffccffffffffffffffc3ffffffff",
            INIT_49 => X"000000280000000000000024000000000000001e000000000000002000000000",
            INIT_4A => X"ffffffd3ffffffff0000001a000000000000001f00000000fffffff3ffffffff",
            INIT_4B => X"ffffffbdffffffffffffffe3ffffffffffffff72ffffffffffffff96ffffffff",
            INIT_4C => X"00000000000000000000005a000000000000006800000000ffffffa3ffffffff",
            INIT_4D => X"000000540000000000000017000000000000004000000000000000a300000000",
            INIT_4E => X"ffffffbeffffffffffffffd4ffffffff00000055000000000000005100000000",
            INIT_4F => X"fffffffbffffffff0000002e000000000000001800000000ffffffd8ffffffff",
            INIT_50 => X"fffffff1fffffffffffffffdffffffff00000023000000000000004200000000",
            INIT_51 => X"00000029000000000000000000000000ffffffbffffffffffffffff2ffffffff",
            INIT_52 => X"0000001200000000000000250000000000000025000000000000003600000000",
            INIT_53 => X"0000000c00000000ffffffcefffffffffffffffbffffffffffffffecffffffff",
            INIT_54 => X"0000002e000000000000001f0000000000000000000000000000000000000000",
            INIT_55 => X"ffffffcaffffffffffffffe0ffffffffffffffc3ffffffff0000000000000000",
            INIT_56 => X"00000040000000000000001700000000ffffffeaffffffff0000001200000000",
            INIT_57 => X"ffffffcaffffffffffffffe8ffffffff00000034000000000000005e00000000",
            INIT_58 => X"0000000a00000000ffffffe5ffffffffffffffd3ffffffffffffffb9ffffffff",
            INIT_59 => X"0000003200000000fffffff6ffffffff00000039000000000000001c00000000",
            INIT_5A => X"000000a000000000000000b300000000ffffffe7ffffffff0000003a00000000",
            INIT_5B => X"ffffffffffffffff000000410000000000000002000000000000006300000000",
            INIT_5C => X"ffffffabffffffff00000028000000000000001900000000ffffffacffffffff",
            INIT_5D => X"ffffffc9ffffffffffffffbffffffffffffffff7ffffffff0000000400000000",
            INIT_5E => X"fffffff2ffffffffffffffccfffffffffffffff3fffffffffffffffaffffffff",
            INIT_5F => X"0000000b00000000fffffff7ffffffffffffffd7ffffffffffffffe4ffffffff",
            INIT_60 => X"ffffffdfffffffffffffffc6ffffffffffffffd8ffffffffffffffecffffffff",
            INIT_61 => X"0000003100000000ffffffd1ffffffffffffffc4ffffffff0000004400000000",
            INIT_62 => X"00000016000000000000000400000000ffffffe3ffffffff0000003b00000000",
            INIT_63 => X"00000001000000000000000d000000000000004a000000000000002500000000",
            INIT_64 => X"0000001c000000000000000a000000000000001e000000000000003c00000000",
            INIT_65 => X"0000000c000000000000001800000000fffffffcffffffffffffffedffffffff",
            INIT_66 => X"fffffffeffffffff0000001400000000fffffff7fffffffffffffff7ffffffff",
            INIT_67 => X"0000000b00000000000000260000000000000017000000000000001800000000",
            INIT_68 => X"ffffffd5ffffffff0000001a000000000000001800000000ffffffdcffffffff",
            INIT_69 => X"ffffffe4ffffffffffffffd2ffffffff0000001900000000ffffffe0ffffffff",
            INIT_6A => X"0000001a00000000ffffffd5ffffffffffffffe2ffffffff0000001d00000000",
            INIT_6B => X"fffffffaffffffffffffffdaffffffffffffffaaffffffff0000000200000000",
            INIT_6C => X"00000004000000000000001d00000000ffffffe5fffffffffffffff3ffffffff",
            INIT_6D => X"0000001f000000000000002d000000000000002d000000000000000b00000000",
            INIT_6E => X"ffffffd8ffffffff00000058000000000000005a000000000000002900000000",
            INIT_6F => X"0000002c0000000000000011000000000000005c000000000000006300000000",
            INIT_70 => X"0000005600000000fffffff9ffffffffffffffddffffffff0000004300000000",
            INIT_71 => X"fffffff3ffffffff0000005d000000000000000000000000ffffffa5ffffffff",
            INIT_72 => X"ffffffdaffffffffffffffc6ffffffff0000001600000000ffffffc7ffffffff",
            INIT_73 => X"fffffff0ffffffffffffffdbfffffffffffffff8fffffffffffffff2ffffffff",
            INIT_74 => X"ffffffeaffffffffffffffe9ffffffff0000001d000000000000002f00000000",
            INIT_75 => X"fffffffaffffffff0000002e00000000ffffffbeffffffffffffffb6ffffffff",
            INIT_76 => X"ffffffecffffffff00000014000000000000005100000000ffffffd0ffffffff",
            INIT_77 => X"0000003e00000000ffffffcbffffffffffffffd4ffffffffffffffeaffffffff",
            INIT_78 => X"00000006000000000000004e00000000ffffffefffffffffffffffe7ffffffff",
            INIT_79 => X"ffffffc0fffffffffffffff9ffffffff0000002500000000fffffff9ffffffff",
            INIT_7A => X"0000001200000000ffffffb8fffffffffffffff1ffffffffffffffd6ffffffff",
            INIT_7B => X"0000002500000000fffffffeffffffffffffffc1ffffffff0000001000000000",
            INIT_7C => X"0000001200000000ffffffecffffffffffffffe7ffffffff0000001100000000",
            INIT_7D => X"ffffffefffffffff00000017000000000000000e00000000fffffffdffffffff",
            INIT_7E => X"ffffffacffffffffffffff9effffffff00000029000000000000001400000000",
            INIT_7F => X"ffffffc9ffffffffffffffbeffffffffffffffbeffffffffffffffedffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE3;


    MEM_IWGHT_LAYER1_INSTANCE4 : if BRAM_NAME = "iwght_layer1_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffff6bffffffffffffffbcffffffffffffff8effffffffffffffb5ffffffff",
            INIT_01 => X"ffffff63ffffffffffffff7fffffffffffffff5dffffffffffffff13ffffffff",
            INIT_02 => X"00000011000000000000000d000000000000000100000000ffffff7fffffffff",
            INIT_03 => X"fffffff2ffffffff000000090000000000000004000000000000000200000000",
            INIT_04 => X"000000200000000000000014000000000000001200000000ffffffe0ffffffff",
            INIT_05 => X"fffffff4fffffffffffffffffffffffffffffffafffffffffffffff0ffffffff",
            INIT_06 => X"0000001d00000000ffffffe8ffffffffffffffcbffffffffffffffdaffffffff",
            INIT_07 => X"0000001500000000000000290000000000000018000000000000001600000000",
            INIT_08 => X"ffffffd7fffffffffffffff3ffffffff00000008000000000000001500000000",
            INIT_09 => X"ffffffebffffffffffffffe1ffffffffffffffedffffffffffffffd8ffffffff",
            INIT_0A => X"0000000600000000fffffff5ffffffff0000001d000000000000000300000000",
            INIT_0B => X"ffffffdeffffffffffffffb7ffffffffffffffc8ffffffff0000002600000000",
            INIT_0C => X"fffffff4ffffffffffffffe7ffffffffffffffdeffffffffffffffb4ffffffff",
            INIT_0D => X"0000002a000000000000000700000000fffffff2ffffffffffffffffffffffff",
            INIT_0E => X"0000000900000000000000270000000000000011000000000000001d00000000",
            INIT_0F => X"ffffffe5ffffffffffffffe8fffffffffffffff8fffffffffffffff2ffffffff",
            INIT_10 => X"ffffffe0ffffffffffffffcdffffffffffffffc3ffffffffffffffcfffffffff",
            INIT_11 => X"0000001d0000000000000004000000000000000f00000000ffffffffffffffff",
            INIT_12 => X"0000000200000000ffffffdcffffffffffffffe3ffffffff0000000700000000",
            INIT_13 => X"ffffffa1ffffffffffffffdbffffffffffffffefffffffffffffffdaffffffff",
            INIT_14 => X"0000000e000000000000002d000000000000005800000000ffffffddffffffff",
            INIT_15 => X"0000000600000000000000510000000000000043000000000000002d00000000",
            INIT_16 => X"ffffffdcffffffffffffffdfffffffff0000001f000000000000000300000000",
            INIT_17 => X"ffffffedffffffffffffffdbffffffff0000000f00000000fffffffcffffffff",
            INIT_18 => X"000000020000000000000013000000000000000600000000ffffffeeffffffff",
            INIT_19 => X"0000000e00000000ffffffebffffffff00000016000000000000000000000000",
            INIT_1A => X"ffffffd7fffffffffffffff3ffffffff0000000f000000000000000200000000",
            INIT_1B => X"0000001700000000fffffffefffffffffffffff7fffffffffffffffbffffffff",
            INIT_1C => X"ffffffe7fffffffffffffffaffffffffffffffefffffffff0000001500000000",
            INIT_1D => X"0000002f00000000ffffffd8ffffffffffffffe0ffffffff0000000d00000000",
            INIT_1E => X"0000003b000000000000003b000000000000000300000000ffffffd9ffffffff",
            INIT_1F => X"00000013000000000000003e000000000000003f000000000000003100000000",
            INIT_20 => X"0000004100000000000000450000000000000049000000000000003000000000",
            INIT_21 => X"0000005a00000000000000630000000000000064000000000000004f00000000",
            INIT_22 => X"0000004b0000000000000036000000000000001d000000000000004300000000",
            INIT_23 => X"00000054000000000000002b0000000000000021000000000000006d00000000",
            INIT_24 => X"ffffffd2ffffffffffffffe8ffffffffffffffd6ffffffffffffff9affffffff",
            INIT_25 => X"fffffffcffffffffffffff90ffffffff00000048000000000000000700000000",
            INIT_26 => X"ffffffdaffffffffffffff96ffffffffffffff98ffffffff0000001a00000000",
            INIT_27 => X"ffffff82ffffffff0000002a00000000ffffffabffffffffffffff61ffffffff",
            INIT_28 => X"ffffffedffffffffffffffd1ffffffffffffffd6ffffffffffffff9affffffff",
            INIT_29 => X"0000004800000000fffffffbffffffff0000002300000000ffffffabffffffff",
            INIT_2A => X"000000430000000000000047000000000000002e000000000000000c00000000",
            INIT_2B => X"0000002600000000000000320000000000000030000000000000003f00000000",
            INIT_2C => X"0000002a00000000000000390000000000000035000000000000005d00000000",
            INIT_2D => X"0000001900000000ffffffffffffffff00000006000000000000001f00000000",
            INIT_2E => X"fffffff0fffffffffffffffdffffffff0000002100000000fffffff5ffffffff",
            INIT_2F => X"00000019000000000000002d000000000000002a00000000fffffff3ffffffff",
            INIT_30 => X"00000037000000000000001f000000000000002b000000000000005a00000000",
            INIT_31 => X"ffffffc0ffffffffffffff8effffffff0000001d000000000000003300000000",
            INIT_32 => X"0000001c00000000ffffffbbffffffffffffff7effffffffffffffadffffffff",
            INIT_33 => X"0000003f000000000000002200000000ffffffe0ffffffffffffff9bffffffff",
            INIT_34 => X"0000002f0000000000000021000000000000001c000000000000003400000000",
            INIT_35 => X"0000000200000000fffffffdffffffff00000022000000000000003200000000",
            INIT_36 => X"ffffffecffffffff0000000100000000ffffffe0ffffffffffffffb2ffffffff",
            INIT_37 => X"000000240000000000000011000000000000005b000000000000000600000000",
            INIT_38 => X"ffffffc2ffffffffffffffffffffffff00000011000000000000002f00000000",
            INIT_39 => X"ffffffffffffffffffffffb0ffffffffffffffe2ffffffff0000002900000000",
            INIT_3A => X"ffffffa1ffffffffffffff9bffffffff0000008c000000000000003000000000",
            INIT_3B => X"0000000500000000ffffffa0ffffffffffffff7fffffffffffffffb4ffffffff",
            INIT_3C => X"ffffffc3ffffffffffffffe6ffffffffffffff82ffffffffffffff95ffffffff",
            INIT_3D => X"ffffff8dffffffffffffff7cffffffffffffffb1ffffffffffffffd8ffffffff",
            INIT_3E => X"ffffffe8ffffffffffffffccffffffffffffffeaffffffffffffffaaffffffff",
            INIT_3F => X"ffffff7bffffffffffffff99ffffffffffffffc0ffffffffffffffacffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffff75ffffffffffffffb5ffffffffffffffacffffffffffffff5dffffffff",
            INIT_41 => X"ffffffa4ffffffffffffffcbffffffffffffffecffffffffffffffb3ffffffff",
            INIT_42 => X"ffffffb0ffffffffffffffbdffffffffffffffafffffffffffffffa5ffffffff",
            INIT_43 => X"00000014000000000000000c00000000ffffffc6ffffffffffffffe0ffffffff",
            INIT_44 => X"ffffffd9fffffffffffffff2ffffffff0000001000000000ffffffecffffffff",
            INIT_45 => X"00000006000000000000007b000000000000002d00000000fffffff8ffffffff",
            INIT_46 => X"ffffffceffffffffffffffffffffffffffffffbaffffffffffffffedffffffff",
            INIT_47 => X"000000820000000000000067000000000000000400000000ffffffeaffffffff",
            INIT_48 => X"000000450000000000000042000000000000004200000000fffffff5ffffffff",
            INIT_49 => X"00000053000000000000006a000000000000002e000000000000000a00000000",
            INIT_4A => X"fffffff7ffffffffffffffd5ffffffffffffffbcffffffff0000000100000000",
            INIT_4B => X"00000034000000000000002e000000000000000f00000000ffffffcfffffffff",
            INIT_4C => X"ffffffb3ffffffffffffffc3ffffffff00000044000000000000002e00000000",
            INIT_4D => X"0000001a00000000fffffffeffffffffffffffe8ffffffffffffffd7ffffffff",
            INIT_4E => X"fffffff0ffffffff000000240000000000000016000000000000000300000000",
            INIT_4F => X"0000000200000000ffffffd9fffffffffffffffeffffffff0000000f00000000",
            INIT_50 => X"0000001b0000000000000004000000000000001c000000000000000900000000",
            INIT_51 => X"ffffffe0ffffffffffffffd7ffffffffffffffffffffffff0000000800000000",
            INIT_52 => X"0000000c00000000ffffffe3ffffffff0000000700000000ffffffe6ffffffff",
            INIT_53 => X"0000000200000000ffffffc6ffffffffffffffd9fffffffffffffffaffffffff",
            INIT_54 => X"fffffff1ffffffff0000000a0000000000000008000000000000000300000000",
            INIT_55 => X"ffffffeaffffffffffffffe0ffffffff0000003b00000000ffffffffffffffff",
            INIT_56 => X"0000001b00000000ffffffeeffffffffffffffd3ffffffffffffffefffffffff",
            INIT_57 => X"ffffffd9ffffffff000000220000000000000012000000000000002a00000000",
            INIT_58 => X"ffffffd8fffffffffffffff3ffffffffffffffedffffffffffffffdbffffffff",
            INIT_59 => X"fffffffaffffffff000000110000000000000004000000000000000200000000",
            INIT_5A => X"ffffff94ffffffffffffffffffffffffffffffc0ffffffffffffffb6ffffffff",
            INIT_5B => X"ffffffbbffffffffffffffb7ffffffff0000000000000000ffffffa2ffffffff",
            INIT_5C => X"fffffff6ffffffff0000000c000000000000004200000000ffffffacffffffff",
            INIT_5D => X"ffffffefffffffff0000001200000000fffffffaffffffff0000002d00000000",
            INIT_5E => X"ffffffdfffffffffffffffe5ffffffff0000000300000000fffffffbffffffff",
            INIT_5F => X"fffffffcffffffff0000001c00000000fffffff4fffffffffffffff9ffffffff",
            INIT_60 => X"ffffffeaffffffff000000380000000000000018000000000000001c00000000",
            INIT_61 => X"ffffffbcffffffffffffffbeffffffffffffffbbffffffffffffffa0ffffffff",
            INIT_62 => X"0000000000000000ffffffe4fffffffffffffff2ffffffffffffffd9ffffffff",
            INIT_63 => X"ffffffc3ffffffffffffffd8ffffffffffffffd7ffffffffffffffbfffffffff",
            INIT_64 => X"fffffff4fffffffffffffff6fffffffffffffffcffffffffffffffc8ffffffff",
            INIT_65 => X"ffffffc5ffffffffffffffd0ffffffff00000017000000000000001d00000000",
            INIT_66 => X"0000000700000000ffffffc1ffffffff00000003000000000000000a00000000",
            INIT_67 => X"00000023000000000000005a000000000000002400000000fffffff8ffffffff",
            INIT_68 => X"00000020000000000000001d000000000000007000000000fffffffdffffffff",
            INIT_69 => X"0000007300000000ffffffe1fffffffffffffff6ffffffff0000001100000000",
            INIT_6A => X"0000001a0000000000000069000000000000002c000000000000004500000000",
            INIT_6B => X"ffffffe8ffffffff000000000000000000000006000000000000002800000000",
            INIT_6C => X"ffffff31ffffffffffffff62ffffffffffffff22ffffffffffffff64ffffffff",
            INIT_6D => X"ffffff20ffffffffffffff67ffffffffffffff41fffffffffffffedcffffffff",
            INIT_6E => X"0000000100000000fffffff4ffffffff0000000300000000ffffff8affffffff",
            INIT_6F => X"0000001600000000fffffffeffffffff0000000d000000000000000b00000000",
            INIT_70 => X"ffffffcaffffffffffffffcdffffffff00000003000000000000000e00000000",
            INIT_71 => X"ffffffc9ffffffffffffffccffffffffffffffe0ffffffffffffffe9ffffffff",
            INIT_72 => X"0000001200000000ffffffbdffffffffffffffaeffffffffffffffcfffffffff",
            INIT_73 => X"0000002000000000fffffff4ffffffff00000006000000000000001e00000000",
            INIT_74 => X"00000001000000000000000a0000000000000019000000000000003200000000",
            INIT_75 => X"0000002800000000000000200000000000000031000000000000000800000000",
            INIT_76 => X"00000029000000000000002b00000000fffffffbffffffff0000000e00000000",
            INIT_77 => X"0000002f000000000000004e0000000000000033000000000000000600000000",
            INIT_78 => X"0000002900000000000000050000000000000014000000000000002600000000",
            INIT_79 => X"0000001d00000000fffffffbffffffff0000000d000000000000004500000000",
            INIT_7A => X"0000000c00000000fffffff5ffffffffffffffe8ffffffff0000001100000000",
            INIT_7B => X"0000000c000000000000001a0000000000000007000000000000001800000000",
            INIT_7C => X"0000000d0000000000000006000000000000001f000000000000000c00000000",
            INIT_7D => X"00000025000000000000000e0000000000000011000000000000002100000000",
            INIT_7E => X"ffffff5bffffffffffffff9affffffffffffff49ffffffffffffff78ffffffff",
            INIT_7F => X"ffffff33ffffffffffffff4bffffffffffffff61ffffffffffffff1fffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE4;


    MEM_IWGHT_LAYER1_INSTANCE5 : if BRAM_NAME = "iwght_layer1_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffd1ffffffffffffffa7ffffffffffffffe3ffffffffffffff72ffffffff",
            INIT_01 => X"ffffffa5ffffffffffffff63ffffffffffffff6dffffffffffffff7effffffff",
            INIT_02 => X"fffffffdffffffff0000001b00000000ffffff9dffffffffffffffc5ffffffff",
            INIT_03 => X"fffffff7ffffffff0000000a000000000000000b00000000ffffffeeffffffff",
            INIT_04 => X"ffffffdcfffffffffffffff0ffffffff00000012000000000000000500000000",
            INIT_05 => X"0000001000000000000000000000000000000008000000000000000400000000",
            INIT_06 => X"ffffffd8ffffffffffffffdbffffffffffffffeaffffffff0000000700000000",
            INIT_07 => X"0000001d00000000fffffffeffffffff00000020000000000000002600000000",
            INIT_08 => X"fffffff8ffffffff0000000100000000fffffff2ffffffff0000000600000000",
            INIT_09 => X"ffffffdaffffffffffffffbcffffffffffffffb1ffffffffffffffecffffffff",
            INIT_0A => X"ffffffa4ffffffffffffffb6ffffffffffffffbeffffffffffffffd1ffffffff",
            INIT_0B => X"ffffff99ffffffffffffffb2ffffffffffffff94ffffffffffffffe5ffffffff",
            INIT_0C => X"ffffff86ffffffffffffff87ffffffffffffff75ffffffffffffffafffffffff",
            INIT_0D => X"fffffff7ffffffffffffffcfffffffffffffffc7ffffffffffffffb3ffffffff",
            INIT_0E => X"ffffffccffffffffffffffb6fffffffffffffff4ffffffffffffffafffffffff",
            INIT_0F => X"ffffff86ffffffffffffff9affffffffffffffc7ffffffffffffff97ffffffff",
            INIT_10 => X"ffffff83ffffffff0000001600000000ffffffe7ffffffffffffffd4ffffffff",
            INIT_11 => X"ffffff62ffffffffffffffaeffffffffffffffb5ffffffffffffff78ffffffff",
            INIT_12 => X"ffffffedffffffffffffffebffffffff0000000000000000ffffffd9ffffffff",
            INIT_13 => X"fffffff4ffffffff00000025000000000000001700000000ffffffedffffffff",
            INIT_14 => X"ffffffd4ffffffffffffffe1ffffffff00000002000000000000000000000000",
            INIT_15 => X"0000001d000000000000000600000000ffffffeaffffffffffffffffffffffff",
            INIT_16 => X"ffffffdfffffffff0000001800000000fffffff2ffffffffffffffe7ffffffff",
            INIT_17 => X"00000023000000000000001400000000ffffffe6ffffffffffffffdaffffffff",
            INIT_18 => X"fffffff3ffffffff000000080000000000000012000000000000001a00000000",
            INIT_19 => X"ffffffe3ffffffff0000000b000000000000002e00000000ffffffddffffffff",
            INIT_1A => X"ffffffc6ffffffffffffffe0fffffffffffffffcffffffffffffffe0ffffffff",
            INIT_1B => X"00000049000000000000003b000000000000003700000000ffffffc8ffffffff",
            INIT_1C => X"0000002f0000000000000056000000000000002e000000000000002000000000",
            INIT_1D => X"0000001800000000000000050000000000000025000000000000003d00000000",
            INIT_1E => X"0000000b0000000000000027000000000000002900000000fffffffdffffffff",
            INIT_1F => X"00000004000000000000002d0000000000000004000000000000000000000000",
            INIT_20 => X"ffffffc7ffffffffffffffeaffffffff00000013000000000000002300000000",
            INIT_21 => X"fffffff7fffffffffffffffcffffffffffffffdcfffffffffffffff4ffffffff",
            INIT_22 => X"0000000e00000000000000450000000000000013000000000000001a00000000",
            INIT_23 => X"0000001400000000000000160000000000000036000000000000002200000000",
            INIT_24 => X"0000001f0000000000000002000000000000004e000000000000003400000000",
            INIT_25 => X"0000004a000000000000002f0000000000000053000000000000004700000000",
            INIT_26 => X"0000001c00000000000000090000000000000061000000000000004600000000",
            INIT_27 => X"0000000c00000000fffffff9ffffffffffffffebffffffff0000002c00000000",
            INIT_28 => X"ffffffbaffffffffffffffe2ffffffffffffffe8ffffffffffffffe7ffffffff",
            INIT_29 => X"ffffffbbffffffffffffffe7ffffffffffffffe5ffffffffffffffdeffffffff",
            INIT_2A => X"ffffffcbffffffffffffffe9ffffffffffffffebffffffff0000000d00000000",
            INIT_2B => X"fffffff4ffffffff00000014000000000000000b00000000fffffff4ffffffff",
            INIT_2C => X"ffffffd6ffffffffffffffccfffffffffffffffcffffffff0000000000000000",
            INIT_2D => X"00000088000000000000005b000000000000005f000000000000000e00000000",
            INIT_2E => X"ffffffe8ffffffff0000002f000000000000005000000000ffffffd9ffffffff",
            INIT_2F => X"ffffffa6ffffffffffffffacffffffff0000002d000000000000000200000000",
            INIT_30 => X"ffffffccffffffffffffffc8ffffffffffffffc6ffffffffffffffecffffffff",
            INIT_31 => X"0000001700000000fffffff5ffffffffffffffdbffffffffffffffffffffffff",
            INIT_32 => X"0000003900000000000000150000000000000029000000000000003b00000000",
            INIT_33 => X"0000003500000000000000370000000000000029000000000000003300000000",
            INIT_34 => X"ffffffc5ffffffff0000005a000000000000002d000000000000003700000000",
            INIT_35 => X"fffffff2ffffffff000000140000000000000021000000000000000300000000",
            INIT_36 => X"ffffffe3ffffffff0000000000000000ffffffffffffffffffffffd2ffffffff",
            INIT_37 => X"0000001d00000000ffffffffffffffffffffffdfffffffffffffffedffffffff",
            INIT_38 => X"ffffffe1ffffffffffffffd4ffffffff0000002c000000000000002b00000000",
            INIT_39 => X"ffffffdbffffffffffffffeaffffffff0000000700000000fffffffeffffffff",
            INIT_3A => X"fffffff6ffffffff0000000600000000fffffff4ffffffffffffffe8ffffffff",
            INIT_3B => X"0000001200000000000000150000000000000012000000000000001b00000000",
            INIT_3C => X"000000200000000000000016000000000000000e00000000fffffff7ffffffff",
            INIT_3D => X"fffffffaffffffffffffffc8ffffffffffffffd2ffffffffffffffd3ffffffff",
            INIT_3E => X"0000000a000000000000002600000000ffffffe2ffffffffffffffebffffffff",
            INIT_3F => X"0000000700000000000000110000000000000028000000000000002b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffe0ffffffff00000007000000000000001500000000ffffffe2ffffffff",
            INIT_41 => X"0000000200000000fffffffcffffffffffffffdeffffffffffffffe0ffffffff",
            INIT_42 => X"0000000c00000000ffffffe3ffffffffffffffebfffffffffffffff2ffffffff",
            INIT_43 => X"ffffffedffffffffffffffe0fffffffffffffff8ffffffff0000000b00000000",
            INIT_44 => X"fffffff6ffffffff00000005000000000000000100000000ffffffe4ffffffff",
            INIT_45 => X"0000000c000000000000002a000000000000001e00000000ffffffe4ffffffff",
            INIT_46 => X"ffffffd3fffffffffffffffeffffffff0000001a000000000000002900000000",
            INIT_47 => X"ffffff0cffffffffffffff9bfffffffffffffff4fffffffffffffffeffffffff",
            INIT_48 => X"0000004d000000000000005d000000000000006500000000ffffff0cffffffff",
            INIT_49 => X"ffffffbcffffffff0000004c000000000000009500000000000000a900000000",
            INIT_4A => X"0000000400000000ffffffdefffffffffffffffaffffffffffffffb7ffffffff",
            INIT_4B => X"ffffffefffffffffffffffefffffffff0000000000000000fffffff8ffffffff",
            INIT_4C => X"000000060000000000000011000000000000002a000000000000001200000000",
            INIT_4D => X"ffffffdaffffffff0000000900000000fffffffafffffffffffffffaffffffff",
            INIT_4E => X"0000000300000000fffffff4fffffffffffffff9ffffffffffffffebffffffff",
            INIT_4F => X"ffffffebffffffffffffffdcffffffffffffffe6fffffffffffffff4ffffffff",
            INIT_50 => X"0000002100000000fffffff8ffffffffffffffefffffffff0000000000000000",
            INIT_51 => X"fffffffdffffffff000000500000000000000010000000000000000e00000000",
            INIT_52 => X"ffffffe9ffffffff000000150000000000000005000000000000000b00000000",
            INIT_53 => X"0000003000000000ffffffe8ffffffffffffffffffffffffffffffbeffffffff",
            INIT_54 => X"ffffffe9ffffffff000000120000000000000027000000000000000000000000",
            INIT_55 => X"0000004800000000ffffffe5ffffffffffffffa7ffffffffffffffb8ffffffff",
            INIT_56 => X"0000005600000000000000670000000000000030000000000000007200000000",
            INIT_57 => X"0000001f000000000000002600000000ffffffd8ffffffff0000005100000000",
            INIT_58 => X"0000000d00000000fffffff5ffffffff0000002f000000000000000600000000",
            INIT_59 => X"0000002b000000000000000d0000000000000001000000000000006e00000000",
            INIT_5A => X"0000000800000000fffffff2fffffffffffffffbffffffff0000005200000000",
            INIT_5B => X"fffffffeffffffffffffffedffffffff00000017000000000000000300000000",
            INIT_5C => X"ffffffdcffffffffffffffcfffffffffffffffedffffffff0000000800000000",
            INIT_5D => X"ffffffe6ffffffff0000000600000000ffffffd4fffffffffffffff4ffffffff",
            INIT_5E => X"ffffffbdffffffffffffffcefffffffffffffffbfffffffffffffffcffffffff",
            INIT_5F => X"ffffffd1ffffffffffffffeafffffffffffffffafffffffffffffff4ffffffff",
            INIT_60 => X"ffffffe3fffffffffffffffeffffffffffffffd2fffffffffffffff9ffffffff",
            INIT_61 => X"0000001d00000000fffffff4ffffffff00000029000000000000001100000000",
            INIT_62 => X"000000030000000000000024000000000000000e000000000000001400000000",
            INIT_63 => X"ffffffdeffffffffffffffe9ffffffffffffffebffffffffffffffffffffffff",
            INIT_64 => X"ffffffe0ffffffff00000016000000000000000000000000ffffffc6ffffffff",
            INIT_65 => X"fffffff0fffffffffffffffaffffffff00000025000000000000001200000000",
            INIT_66 => X"00000003000000000000000700000000ffffffe1ffffffffffffffc9ffffffff",
            INIT_67 => X"0000002800000000fffffff9ffffffff0000000300000000fffffff8ffffffff",
            INIT_68 => X"fffffff5fffffffffffffff8fffffffffffffff8ffffffff0000000b00000000",
            INIT_69 => X"000000230000000000000022000000000000000d000000000000000c00000000",
            INIT_6A => X"ffffffeaffffffffffffffeaffffffff0000004800000000ffffffe8ffffffff",
            INIT_6B => X"000000310000000000000005000000000000000d000000000000004600000000",
            INIT_6C => X"ffffffd4ffffffffffffffcfffffffffffffffceffffffffffffffefffffffff",
            INIT_6D => X"0000001500000000ffffffecffffffffffffffeaffffffffffffffd5ffffffff",
            INIT_6E => X"0000000c00000000000000240000000000000016000000000000001500000000",
            INIT_6F => X"fffffffbffffffff0000002100000000ffffffe6fffffffffffffff8ffffffff",
            INIT_70 => X"0000001100000000000000140000000000000008000000000000001700000000",
            INIT_71 => X"fffffff0ffffffff0000002b000000000000000000000000fffffff5ffffffff",
            INIT_72 => X"fffffff5ffffffff000000210000000000000022000000000000001100000000",
            INIT_73 => X"00000016000000000000001600000000fffffffdfffffffffffffffbffffffff",
            INIT_74 => X"0000001f000000000000002a000000000000001900000000ffffffe4ffffffff",
            INIT_75 => X"ffffffbfffffffffffffffdcffffffffffffffb8fffffffffffffffbffffffff",
            INIT_76 => X"ffffffb8ffffffffffffffefffffffffffffff7cffffffffffffff7affffffff",
            INIT_77 => X"ffffffecffffffff0000000300000000ffffffc5ffffffffffffffbcffffffff",
            INIT_78 => X"0000000400000000ffffffedffffffffffffffddffffffffffffffe2ffffffff",
            INIT_79 => X"ffffffdcffffffff0000002200000000fffffffcfffffffffffffff8ffffffff",
            INIT_7A => X"ffffffcaffffffffffffffadffffffffffffffe0fffffffffffffff2ffffffff",
            INIT_7B => X"0000002600000000ffffffe7ffffffff0000000300000000ffffffe1ffffffff",
            INIT_7C => X"000000630000000000000040000000000000009e000000000000007f00000000",
            INIT_7D => X"0000007d00000000000000680000000000000036000000000000007000000000",
            INIT_7E => X"ffffffdfffffffff000000020000000000000006000000000000001e00000000",
            INIT_7F => X"ffffffe7ffffffff000000020000000000000016000000000000000b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE5;


    MEM_IWGHT_LAYER1_INSTANCE6 : if BRAM_NAME = "iwght_layer1_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffffaffffffffffffffedfffffffffffffffeffffffff0000000b00000000",
            INIT_01 => X"fffffffdfffffffffffffffaffffffff0000000e00000000ffffffe3ffffffff",
            INIT_02 => X"0000002d000000000000000300000000fffffffdfffffffffffffffdffffffff",
            INIT_03 => X"00000013000000000000004e000000000000002c00000000fffffff6ffffffff",
            INIT_04 => X"0000001c00000000000000110000000000000026000000000000002e00000000",
            INIT_05 => X"ffffffd6ffffffff0000000300000000ffffffdeffffffffffffffdcffffffff",
            INIT_06 => X"000000040000000000000003000000000000001e00000000ffffffe4ffffffff",
            INIT_07 => X"ffffffeaffffffff0000002c0000000000000020000000000000002f00000000",
            INIT_08 => X"0000001c00000000000000140000000000000000000000000000000500000000",
            INIT_09 => X"00000022000000000000000100000000fffffff2ffffffffffffffedffffffff",
            INIT_0A => X"fffffff6fffffffffffffffefffffffffffffffeffffffff0000000000000000",
            INIT_0B => X"0000000d00000000ffffffcdffffffff0000000c000000000000000100000000",
            INIT_0C => X"ffffffe8fffffffffffffff0ffffffff00000009000000000000000e00000000",
            INIT_0D => X"0000000600000000000000190000000000000018000000000000001300000000",
            INIT_0E => X"ffffffb3ffffffffffffffd6ffffffffffffffedffffffffffffff9effffffff",
            INIT_0F => X"ffffffc3ffffffff0000001c00000000ffffffb9ffffffffffffffb1ffffffff",
            INIT_10 => X"00000011000000000000001500000000ffffffcaffffffffffffffd0ffffffff",
            INIT_11 => X"0000001f00000000000000010000000000000025000000000000000a00000000",
            INIT_12 => X"0000000d00000000ffffffe5ffffffffffffffcbfffffffffffffff4ffffffff",
            INIT_13 => X"0000001300000000ffffffdefffffffffffffffefffffffffffffffdffffffff",
            INIT_14 => X"000000060000000000000005000000000000000f00000000ffffffe0ffffffff",
            INIT_15 => X"00000018000000000000001600000000ffffffe9ffffffffffffffe4ffffffff",
            INIT_16 => X"fffffff2ffffffff00000015000000000000001000000000fffffff7ffffffff",
            INIT_17 => X"0000001a0000000000000000000000000000000f00000000ffffffe2ffffffff",
            INIT_18 => X"0000000200000000fffffffffffffffffffffff8ffffffff0000000300000000",
            INIT_19 => X"0000000800000000ffffffebffffffff0000001300000000ffffffe1ffffffff",
            INIT_1A => X"00000033000000000000002200000000fffffffbffffffff0000001300000000",
            INIT_1B => X"00000023000000000000002300000000ffffffd7fffffffffffffffeffffffff",
            INIT_1C => X"0000003b00000000000000260000000000000036000000000000002c00000000",
            INIT_1D => X"0000003200000000000000460000000000000049000000000000005c00000000",
            INIT_1E => X"000000550000000000000042000000000000004c000000000000001200000000",
            INIT_1F => X"ffffffeeffffffff00000019000000000000004b000000000000003f00000000",
            INIT_20 => X"0000002e0000000000000006000000000000002b000000000000000b00000000",
            INIT_21 => X"00000067000000000000002e0000000000000048000000000000001200000000",
            INIT_22 => X"fffffff0ffffffff0000001c00000000fffffffbffffffff0000004000000000",
            INIT_23 => X"0000001800000000fffffffaffffffff0000001500000000fffffff7ffffffff",
            INIT_24 => X"ffffffceffffffffffffffcaffffffff0000001b00000000fffffff8ffffffff",
            INIT_25 => X"0000000000000000fffffff4ffffffffffffffe7ffffffffffffffe8ffffffff",
            INIT_26 => X"fffffffdfffffffffffffff9ffffffffffffffeeffffffffffffffeeffffffff",
            INIT_27 => X"ffffffedfffffffffffffffbffffffff00000014000000000000001300000000",
            INIT_28 => X"ffffffe0ffffffffffffffe8ffffffffffffffd6ffffffffffffffe3ffffffff",
            INIT_29 => X"0000000700000000000000300000000000000006000000000000000100000000",
            INIT_2A => X"fffffffdfffffffffffffff3ffffffffffffffffffffffff0000000800000000",
            INIT_2B => X"00000021000000000000000d00000000fffffff6ffffffff0000000700000000",
            INIT_2C => X"0000002b000000000000002f00000000fffffff7fffffffffffffffaffffffff",
            INIT_2D => X"fffffff9fffffffffffffffdfffffffffffffffeffffffff0000000d00000000",
            INIT_2E => X"0000001200000000fffffff1ffffffff0000000f00000000ffffffdeffffffff",
            INIT_2F => X"0000002000000000fffffffdffffffffffffffe7ffffffffffffffe5ffffffff",
            INIT_30 => X"00000019000000000000000100000000fffffffcffffffff0000001200000000",
            INIT_31 => X"0000001500000000000000290000000000000006000000000000003100000000",
            INIT_32 => X"ffffffe8fffffffffffffff7ffffffffffffffddffffffff0000000d00000000",
            INIT_33 => X"0000002b00000000fffffffbffffffff0000000800000000fffffff8ffffffff",
            INIT_34 => X"ffffffbcffffffffffffffdaffffffffffffffc6ffffffffffffffd2ffffffff",
            INIT_35 => X"0000000400000000ffffffa5ffffffffffffffb3ffffffffffffffa0ffffffff",
            INIT_36 => X"0000001d0000000000000008000000000000000600000000fffffff9ffffffff",
            INIT_37 => X"fffffffbffffffff000000080000000000000014000000000000000400000000",
            INIT_38 => X"0000000c000000000000001b000000000000001b000000000000000800000000",
            INIT_39 => X"fffffff4ffffffff0000000000000000ffffffddffffffffffffffd9ffffffff",
            INIT_3A => X"fffffff2fffffffffffffffcffffffff0000000d00000000ffffffe3ffffffff",
            INIT_3B => X"0000000700000000ffffffe6ffffffffffffffe2ffffffff0000001b00000000",
            INIT_3C => X"0000000d00000000ffffffeefffffffffffffff3ffffffff0000000e00000000",
            INIT_3D => X"ffffffdbffffffffffffffd3ffffffffffffffeffffffffffffffff4ffffffff",
            INIT_3E => X"ffffffd4ffffffffffffffe5ffffffffffffffb2ffffffffffffff96ffffffff",
            INIT_3F => X"fffffffeffffffffffffffc8ffffffffffffffe6ffffffffffffffa1ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffe9ffffffffffffffdcffffffffffffffbbffffffffffffffe1ffffffff",
            INIT_41 => X"ffffffb6ffffffff0000001600000000ffffffedffffffffffffffdcffffffff",
            INIT_42 => X"ffffffdcffffffffffffffd8ffffffffffffffd2ffffffffffffff9bffffffff",
            INIT_43 => X"000000190000000000000015000000000000001f00000000ffffffdcffffffff",
            INIT_44 => X"00000057000000000000003a0000000000000068000000000000001c00000000",
            INIT_45 => X"000000410000000000000068000000000000001400000000000000af00000000",
            INIT_46 => X"00000004000000000000000600000000ffffffd9ffffffff0000000000000000",
            INIT_47 => X"ffffffeffffffffffffffffcffffffff0000000b00000000ffffffe6ffffffff",
            INIT_48 => X"0000002000000000000000010000000000000016000000000000001900000000",
            INIT_49 => X"00000012000000000000000d00000000fffffffcffffffff0000000600000000",
            INIT_4A => X"0000001f00000000ffffffefffffffff0000002a00000000ffffffeeffffffff",
            INIT_4B => X"ffffffe4ffffffff00000010000000000000000a000000000000001800000000",
            INIT_4C => X"fffffffcfffffffffffffff4ffffffffffffffedffffffff0000000000000000",
            INIT_4D => X"00000012000000000000002700000000fffffff8fffffffffffffffbffffffff",
            INIT_4E => X"0000001b00000000000000090000000000000004000000000000001900000000",
            INIT_4F => X"fffffff9ffffffff0000001800000000ffffffecffffffffffffffe0ffffffff",
            INIT_50 => X"0000002000000000000000240000000000000021000000000000000000000000",
            INIT_51 => X"0000002500000000000000000000000000000015000000000000002a00000000",
            INIT_52 => X"00000032000000000000001d00000000fffffff5ffffffff0000000900000000",
            INIT_53 => X"0000000c0000000000000034000000000000003500000000ffffffe0ffffffff",
            INIT_54 => X"0000000e00000000fffffff9fffffffffffffff8ffffffff0000000000000000",
            INIT_55 => X"00000007000000000000000500000000fffffff6fffffffffffffff7ffffffff",
            INIT_56 => X"0000000f000000000000001c0000000000000010000000000000002f00000000",
            INIT_57 => X"00000039000000000000002100000000ffffffffffffffff0000005200000000",
            INIT_58 => X"ffffffdeffffffffffffffd1ffffffffffffffe8ffffffff0000001c00000000",
            INIT_59 => X"fffffff6ffffffffffffffe3ffffffffffffffddffffffff0000001200000000",
            INIT_5A => X"0000000000000000fffffff3ffffffffffffffeaffffffffffffffb2ffffffff",
            INIT_5B => X"00000017000000000000000c00000000ffffffd9ffffffff0000001e00000000",
            INIT_5C => X"fffffff8ffffffffffffffe9ffffffff00000007000000000000000f00000000",
            INIT_5D => X"ffffffbcffffffffffffffe1ffffffff0000000200000000ffffffbbffffffff",
            INIT_5E => X"0000001000000000ffffffe1ffffffffffffffe8ffffffff0000000400000000",
            INIT_5F => X"ffffffd6ffffffff0000001600000000ffffffdafffffffffffffff5ffffffff",
            INIT_60 => X"ffffffe1ffffffffffffffe4ffffffff0000001200000000ffffffd6ffffffff",
            INIT_61 => X"ffffffe9ffffffff00000019000000000000000e00000000fffffffdffffffff",
            INIT_62 => X"00000025000000000000001000000000ffffffe0ffffffff0000003d00000000",
            INIT_63 => X"fffffff5ffffffff0000001a000000000000001d00000000ffffffedffffffff",
            INIT_64 => X"0000001e00000000ffffffbeffffffff00000022000000000000002000000000",
            INIT_65 => X"ffffffe6ffffffffffffffe4ffffffffffffffe0ffffffff0000000400000000",
            INIT_66 => X"ffffffb5ffffffffffffff9dfffffffffffffff3ffffffffffffffd8ffffffff",
            INIT_67 => X"ffffffb4ffffffffffffffbbffffffffffffff92fffffffffffffff4ffffffff",
            INIT_68 => X"ffffffe0ffffffffffffffbdffffffffffffff9effffffff0000001900000000",
            INIT_69 => X"ffffffc0ffffffff0000000700000000ffffffa4ffffffffffffff55ffffffff",
            INIT_6A => X"ffffffdefffffffffffffff6ffffffff0000002000000000ffffffb3ffffffff",
            INIT_6B => X"0000003200000000ffffffd3ffffffffffffffffffffffff0000002800000000",
            INIT_6C => X"fffffffcfffffffffffffffbffffffffffffffd1ffffffffffffffecffffffff",
            INIT_6D => X"ffffff93ffffffffffffffd5ffffffff0000000400000000ffffffe1ffffffff",
            INIT_6E => X"0000002500000000ffffffa4fffffffffffffff6ffffffff0000002a00000000",
            INIT_6F => X"00000026000000000000003c00000000ffffffe8fffffffffffffff0ffffffff",
            INIT_70 => X"ffffffebffffffff00000024000000000000004300000000ffffffd4ffffffff",
            INIT_71 => X"0000000700000000fffffff4ffffffffffffffdafffffffffffffff2ffffffff",
            INIT_72 => X"ffffffe9fffffffffffffff9fffffffffffffff8ffffffffffffffdfffffffff",
            INIT_73 => X"0000001900000000fffffff8ffffffffffffffe3fffffffffffffffcffffffff",
            INIT_74 => X"ffffffbcffffffff0000001200000000ffffffe1ffffffffffffffbcffffffff",
            INIT_75 => X"00000004000000000000003800000000fffffffdffffffffffffffceffffffff",
            INIT_76 => X"ffffffcdffffffffffffffe9ffffffff0000003b00000000ffffffd5ffffffff",
            INIT_77 => X"ffffffebffffffffffffffc1ffffffff00000010000000000000001a00000000",
            INIT_78 => X"0000001a000000000000000e000000000000002e00000000fffffffaffffffff",
            INIT_79 => X"0000001400000000000000110000000000000017000000000000002700000000",
            INIT_7A => X"ffffffd4ffffffff0000000700000000ffffffafffffffffffffffd9ffffffff",
            INIT_7B => X"ffffffd6ffffffff0000002d00000000fffffff7ffffffffffffff83ffffffff",
            INIT_7C => X"00000016000000000000000200000000ffffffcdffffffffffffffc2ffffffff",
            INIT_7D => X"0000000f000000000000000b00000000ffffffadfffffffffffffff3ffffffff",
            INIT_7E => X"0000000200000000ffffffffffffffffffffffd0ffffffffffffffe3ffffffff",
            INIT_7F => X"ffffffd3fffffffffffffffbffffffff0000001f00000000fffffff7ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE6;


    MEM_IWGHT_LAYER1_INSTANCE7 : if BRAM_NAME = "iwght_layer1_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003b00000000ffffffdfffffffff00000013000000000000001800000000",
            INIT_01 => X"00000004000000000000002e000000000000000000000000fffffff6ffffffff",
            INIT_02 => X"0000000000000000000000250000000000000034000000000000001a00000000",
            INIT_03 => X"0000003200000000ffffffdfffffffff00000019000000000000003400000000",
            INIT_04 => X"0000002b000000000000004900000000ffffffe6ffffffff0000000a00000000",
            INIT_05 => X"0000002e000000000000000200000000ffffffbdfffffffffffffff6ffffffff",
            INIT_06 => X"ffffffcdffffffff0000001f00000000fffffff0ffffffffffffffd8ffffffff",
            INIT_07 => X"0000001c00000000fffffff1ffffffff0000001d000000000000002200000000",
            INIT_08 => X"00000039000000000000000c00000000ffffffdfffffffff0000005100000000",
            INIT_09 => X"ffffffbcffffffff0000002900000000fffffffefffffffffffffffbffffffff",
            INIT_0A => X"ffffffeaffffffffffffffe2ffffffff00000004000000000000001400000000",
            INIT_0B => X"ffffffc1ffffffffffffffd2ffffffffffffffd0ffffffffffffffddffffffff",
            INIT_0C => X"00000036000000000000000e00000000ffffffd3ffffffff0000000700000000",
            INIT_0D => X"0000006400000000000000570000000000000067000000000000003a00000000",
            INIT_0E => X"ffffffe9fffffffffffffff6ffffffff00000022000000000000006000000000",
            INIT_0F => X"fffffff3ffffffff0000001800000000ffffffe1ffffffffffffffdcffffffff",
            INIT_10 => X"00000006000000000000002c000000000000000d00000000fffffff7ffffffff",
            INIT_11 => X"ffffffeeffffffff0000002000000000ffffffeffffffffffffffffdffffffff",
            INIT_12 => X"00000039000000000000003500000000ffffffd0ffffffffffffffc4ffffffff",
            INIT_13 => X"ffffffe9ffffffff0000000c0000000000000011000000000000002900000000",
            INIT_14 => X"fffffff1ffffffffffffffd5ffffffffffffffedffffffffffffffe9ffffffff",
            INIT_15 => X"ffffffefffffffffffffffdaffffffffffffffd6ffffffff0000000000000000",
            INIT_16 => X"0000002d00000000000000040000000000000015000000000000000800000000",
            INIT_17 => X"0000001500000000ffffffd1ffffffff00000010000000000000001500000000",
            INIT_18 => X"0000000b00000000000000370000000000000002000000000000001900000000",
            INIT_19 => X"0000000f0000000000000037000000000000002c000000000000002e00000000",
            INIT_1A => X"fffffffbfffffffffffffff0ffffffff00000013000000000000000a00000000",
            INIT_1B => X"ffffffd8fffffffffffffffeffffffffffffffd8ffffffffffffffe4ffffffff",
            INIT_1C => X"0000000f000000000000001e00000000ffffffe4ffffffffffffffdcffffffff",
            INIT_1D => X"000000200000000000000024000000000000000c000000000000002400000000",
            INIT_1E => X"fffffff2fffffffffffffff3ffffffffffffffb5ffffffff0000000500000000",
            INIT_1F => X"ffffffedfffffffffffffffdffffffff0000000c000000000000002900000000",
            INIT_20 => X"ffffffc6ffffffff000000440000000000000016000000000000003300000000",
            INIT_21 => X"ffffffd4ffffffff0000000d000000000000004d000000000000002b00000000",
            INIT_22 => X"ffffffd2ffffffffffffffecffffffff00000052000000000000001e00000000",
            INIT_23 => X"0000002100000000ffffffe0fffffffffffffffdffffffffffffffe3ffffffff",
            INIT_24 => X"000000280000000000000029000000000000001f00000000ffffffffffffffff",
            INIT_25 => X"0000000200000000fffffffdffffffff00000026000000000000004700000000",
            INIT_26 => X"ffffffdaffffffffffffffd0ffffffffffffffe0ffffffff0000001400000000",
            INIT_27 => X"ffffffeeffffffff0000000f000000000000000a000000000000001000000000",
            INIT_28 => X"ffffffe7ffffffffffffffceffffffffffffffebffffffffffffffe8ffffffff",
            INIT_29 => X"ffffffcaffffffffffffffcfffffffffffffffbfffffffffffffffe0ffffffff",
            INIT_2A => X"0000001300000000fffffff6ffffffff00000026000000000000003300000000",
            INIT_2B => X"fffffff9ffffffff000000260000000000000031000000000000001c00000000",
            INIT_2C => X"ffffffe6ffffffff00000039000000000000004100000000ffffffc3ffffffff",
            INIT_2D => X"000000050000000000000031000000000000004400000000ffffffedffffffff",
            INIT_2E => X"0000001b000000000000005c00000000ffffffd7ffffffff0000000d00000000",
            INIT_2F => X"0000004c000000000000003e0000000000000010000000000000000400000000",
            INIT_30 => X"0000001500000000000000270000000000000011000000000000001b00000000",
            INIT_31 => X"ffffffebfffffffffffffff5ffffffffffffffe7fffffffffffffff0ffffffff",
            INIT_32 => X"00000001000000000000000a000000000000001b000000000000001c00000000",
            INIT_33 => X"fffffffeffffffff0000001900000000ffffffeafffffffffffffff3ffffffff",
            INIT_34 => X"ffffffecffffffffffffffedffffffffffffffddfffffffffffffff2ffffffff",
            INIT_35 => X"0000001700000000fffffff5ffffffff0000001b00000000fffffff3ffffffff",
            INIT_36 => X"0000001c000000000000001500000000fffffff3ffffffff0000001200000000",
            INIT_37 => X"00000008000000000000000500000000ffffffecffffffffffffffefffffffff",
            INIT_38 => X"0000001d00000000fffffff0ffffffffffffffe8ffffffffffffffe8ffffffff",
            INIT_39 => X"0000001e0000000000000026000000000000001f000000000000000500000000",
            INIT_3A => X"fffffff6ffffffffffffffd4ffffffff0000000400000000fffffff0ffffffff",
            INIT_3B => X"000000020000000000000000000000000000000e00000000ffffffedffffffff",
            INIT_3C => X"0000000100000000ffffffd4fffffffffffffff3ffffffff0000000400000000",
            INIT_3D => X"ffffffffffffffffffffffe4ffffffffffffffc5ffffffffffffffcfffffffff",
            INIT_3E => X"0000000a00000000fffffff0ffffffff0000001c00000000fffffff5ffffffff",
            INIT_3F => X"0000000c00000000fffffff6ffffffff0000000700000000ffffffedffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffffbffffffffffffffdefffffffffffffff9ffffffff0000002700000000",
            INIT_41 => X"ffffffc7ffffffffffffffc5ffffffffffffffdcffffffffffffffeeffffffff",
            INIT_42 => X"0000003100000000fffffffcffffffffffffffeaffffffff0000001e00000000",
            INIT_43 => X"0000002b000000000000000800000000ffffffe6fffffffffffffffcffffffff",
            INIT_44 => X"00000033000000000000002e0000000000000044000000000000000b00000000",
            INIT_45 => X"0000002f00000000000000220000000000000050000000000000005800000000",
            INIT_46 => X"0000002f00000000000000240000000000000041000000000000006500000000",
            INIT_47 => X"fffffff5ffffffff0000000400000000fffffff2fffffffffffffff7ffffffff",
            INIT_48 => X"ffffffe7ffffffffffffffd3ffffffffffffffe4ffffffff0000000100000000",
            INIT_49 => X"fffffffcffffffff0000001b000000000000000000000000fffffffbffffffff",
            INIT_4A => X"ffffffe6ffffffff0000000e00000000ffffffe2ffffffff0000001600000000",
            INIT_4B => X"00000009000000000000000800000000fffffff7ffffffff0000002900000000",
            INIT_4C => X"ffffffe9ffffffff0000000d00000000fffffffcffffffff0000000600000000",
            INIT_4D => X"ffffffeaffffffff00000001000000000000001e00000000fffffff4ffffffff",
            INIT_4E => X"ffffffd2ffffffff000000130000000000000019000000000000000800000000",
            INIT_4F => X"00000037000000000000003a00000000fffffff9ffffffffffffffc1ffffffff",
            INIT_50 => X"0000003f000000000000002b0000000000000042000000000000002f00000000",
            INIT_51 => X"0000003700000000000000330000000000000026000000000000003800000000",
            INIT_52 => X"000000910000000000000083000000000000002e000000000000004100000000",
            INIT_53 => X"0000003200000000000000660000000000000050000000000000004500000000",
            INIT_54 => X"ffffffe7ffffffffffffffcbffffffffffffffcfffffffffffffffd0ffffffff",
            INIT_55 => X"0000002600000000fffffff4ffffffffffffffebffffffffffffffeeffffffff",
            INIT_56 => X"0000000900000000fffffff7ffffffffffffffe8ffffffff0000000900000000",
            INIT_57 => X"0000000f00000000fffffff6ffffffff0000001200000000fffffff0ffffffff",
            INIT_58 => X"ffffffe9ffffffffffffffe5fffffffffffffffcffffffff0000002200000000",
            INIT_59 => X"fffffffdffffffffffffffefffffffff0000000900000000ffffffdbffffffff",
            INIT_5A => X"0000001f00000000ffffffddffffffffffffffe5ffffffffffffffebffffffff",
            INIT_5B => X"0000001900000000ffffffefffffffff0000000300000000fffffff0ffffffff",
            INIT_5C => X"00000016000000000000001300000000fffffffeffffffff0000001200000000",
            INIT_5D => X"ffffffbdffffffffffffffb4ffffffffffffffc6ffffffffffffffeeffffffff",
            INIT_5E => X"ffffffbdffffffffffffffe4ffffffffffffffb6ffffffffffffffd0ffffffff",
            INIT_5F => X"00000027000000000000001c000000000000002700000000ffffffd5ffffffff",
            INIT_60 => X"0000005600000000000000100000000000000025000000000000001700000000",
            INIT_61 => X"000000000000000000000022000000000000002d000000000000005000000000",
            INIT_62 => X"0000002b00000000000000280000000000000020000000000000000400000000",
            INIT_63 => X"ffffffc8ffffffff0000002e0000000000000036000000000000003400000000",
            INIT_64 => X"ffffffd6ffffffffffffffdbffffffffffffffc8ffffffffffffffbeffffffff",
            INIT_65 => X"ffffffeeffffffff0000000800000000ffffffeaffffffffffffffc2ffffffff",
            INIT_66 => X"0000002d000000000000000500000000fffffff4ffffffff0000001100000000",
            INIT_67 => X"0000000d000000000000000d0000000000000002000000000000000c00000000",
            INIT_68 => X"00000051000000000000003c000000000000003a000000000000002200000000",
            INIT_69 => X"0000004b0000000000000041000000000000003a000000000000001600000000",
            INIT_6A => X"fffffff0ffffffff0000000b0000000000000028000000000000002500000000",
            INIT_6B => X"0000000b00000000ffffffedffffffffffffffeaffffffff0000001100000000",
            INIT_6C => X"fffffffdfffffffffffffff2ffffffffffffffebffffffff0000000000000000",
            INIT_6D => X"ffffffedfffffffffffffffefffffffffffffffefffffffffffffff7ffffffff",
            INIT_6E => X"00000011000000000000001a00000000fffffffcffffffffffffffe9ffffffff",
            INIT_6F => X"fffffffbffffffff0000000d000000000000001800000000fffffffdffffffff",
            INIT_70 => X"0000001f00000000000000010000000000000017000000000000000000000000",
            INIT_71 => X"0000001500000000ffffffe2ffffffffffffffdbffffffff0000001100000000",
            INIT_72 => X"ffffffb2ffffffffffffffb5ffffffffffffff80ffffffffffffffdbffffffff",
            INIT_73 => X"ffffffb2ffffffffffffffcbffffffff0000000400000000ffffffa0ffffffff",
            INIT_74 => X"ffffffc4ffffffffffffffb5ffffffffffffffa9ffffffffffffffd6ffffffff",
            INIT_75 => X"fffffff1ffffffffffffffb7ffffffffffffffbdffffffffffffffbdffffffff",
            INIT_76 => X"ffffffe0ffffffff00000008000000000000002000000000ffffffebffffffff",
            INIT_77 => X"fffffff8ffffffffffffffc9ffffffffffffffe2ffffffffffffffe9ffffffff",
            INIT_78 => X"ffffffd9ffffffff00000031000000000000001b00000000ffffffadffffffff",
            INIT_79 => X"ffffffc7ffffffffffffffc7ffffffff00000034000000000000002700000000",
            INIT_7A => X"0000001700000000ffffffecffffffff0000000400000000ffffffe9ffffffff",
            INIT_7B => X"ffffffffffffffff0000000a000000000000000700000000fffffffeffffffff",
            INIT_7C => X"000000180000000000000003000000000000000a000000000000000c00000000",
            INIT_7D => X"fffffffefffffffffffffff9ffffffffffffffd6fffffffffffffff3ffffffff",
            INIT_7E => X"00000035000000000000000700000000fffffffeffffffffffffffdeffffffff",
            INIT_7F => X"0000003c00000000000000220000000000000003000000000000003c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE7;


    MEM_IWGHT_LAYER1_INSTANCE8 : if BRAM_NAME = "iwght_layer1_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000002e000000000000002c000000000000000000000000",
            INIT_01 => X"000000050000000000000007000000000000000a00000000ffffffe6ffffffff",
            INIT_02 => X"0000001800000000fffffff6ffffffff0000001c000000000000000d00000000",
            INIT_03 => X"00000028000000000000002f00000000ffffffe9ffffffff0000000700000000",
            INIT_04 => X"00000010000000000000001f00000000fffffff9ffffffff0000000900000000",
            INIT_05 => X"0000001b000000000000001f00000000ffffffffffffffff0000000b00000000",
            INIT_06 => X"0000001e00000000fffffffbffffffffffffffeaffffffffffffffebffffffff",
            INIT_07 => X"fffffffafffffffffffffff9ffffffff0000001a000000000000001100000000",
            INIT_08 => X"fffffffeffffffffffffffddffffffff00000014000000000000000d00000000",
            INIT_09 => X"0000000600000000ffffffe4ffffffff0000000d000000000000001900000000",
            INIT_0A => X"fffffff2ffffffff00000033000000000000003600000000ffffffdaffffffff",
            INIT_0B => X"00000005000000000000000c0000000000000035000000000000001500000000",
            INIT_0C => X"ffffff72ffffffffffffff81ffffffffffffff84fffffffffffffff2ffffffff",
            INIT_0D => X"ffffff8affffffffffffff8effffffffffffff2cffffffffffffff3fffffffff",
            INIT_0E => X"0000001100000000ffffffe8ffffffffffffff7fffffffffffffff6dffffffff",
            INIT_0F => X"00000019000000000000000400000000fffffffbffffffff0000001600000000",
            INIT_10 => X"0000002b00000000ffffffe8ffffffffffffffe1ffffffff0000000500000000",
            INIT_11 => X"0000000100000000fffffff1ffffffff0000002e000000000000001800000000",
            INIT_12 => X"ffffffecfffffffffffffffeffffffffffffffecffffffff0000000d00000000",
            INIT_13 => X"ffffffd7fffffffffffffff0fffffffffffffff9ffffffff0000001f00000000",
            INIT_14 => X"0000000d00000000ffffffe8ffffffff0000001a00000000ffffffe1ffffffff",
            INIT_15 => X"0000000700000000ffffffe0ffffffffffffffceffffffffffffffe9ffffffff",
            INIT_16 => X"ffffffadffffffffffffffd4ffffffffffffffb4ffffffffffffffb9ffffffff",
            INIT_17 => X"ffffff88ffffffffffffff9bffffffffffffffcaffffffffffffff87ffffffff",
            INIT_18 => X"ffffffe6ffffffffffffffeeffffffffffffffd2ffffffffffffffbbffffffff",
            INIT_19 => X"ffffff88ffffffffffffffd7ffffffffffffff98ffffffffffffffa0ffffffff",
            INIT_1A => X"ffffff77ffffffffffffff6affffffffffffff74ffffffffffffff3dffffffff",
            INIT_1B => X"ffffff92ffffffffffffff8fffffffffffffff95ffffffffffffff80ffffffff",
            INIT_1C => X"000000600000000000000060000000000000004b000000000000006200000000",
            INIT_1D => X"00000010000000000000001d000000000000002a000000000000003200000000",
            INIT_1E => X"fffffff8ffffffff0000000000000000ffffffe6ffffffff0000002100000000",
            INIT_1F => X"000000040000000000000000000000000000001300000000fffffff1ffffffff",
            INIT_20 => X"ffffffddffffffffffffffe1ffffffff0000000900000000ffffffeaffffffff",
            INIT_21 => X"fffffff5ffffffffffffffdbffffffffffffffc3ffffffffffffffe4ffffffff",
            INIT_22 => X"ffffffebfffffffffffffffeffffffffffffffd7ffffffffffffffd8ffffffff",
            INIT_23 => X"ffffffdaffffffffffffffceffffffff0000000a00000000ffffffe6ffffffff",
            INIT_24 => X"ffffffdefffffffffffffffeffffffffffffffeeffffffff0000000200000000",
            INIT_25 => X"0000001e00000000000000290000000000000020000000000000000500000000",
            INIT_26 => X"00000025000000000000001d000000000000000e000000000000002500000000",
            INIT_27 => X"ffffffe9ffffffff0000000000000000fffffff1ffffffff0000001f00000000",
            INIT_28 => X"0000000000000000fffffff2ffffffff0000000600000000ffffffe6ffffffff",
            INIT_29 => X"ffffffd4fffffffffffffff1ffffffff0000000c00000000fffffffcffffffff",
            INIT_2A => X"00000000000000000000000600000000ffffffcfffffffffffffffefffffffff",
            INIT_2B => X"fffffff8ffffffff0000000400000000ffffffccffffffffffffffecffffffff",
            INIT_2C => X"0000002100000000fffffff6ffffffff00000017000000000000002400000000",
            INIT_2D => X"0000001200000000000000110000000000000016000000000000000000000000",
            INIT_2E => X"ffffffdeffffffff0000001200000000fffffff3ffffffff0000001e00000000",
            INIT_2F => X"ffffffffffffffff0000000300000000ffffffffffffffff0000000400000000",
            INIT_30 => X"00000023000000000000003700000000fffffffeffffffffffffffecffffffff",
            INIT_31 => X"ffffffd6fffffffffffffffcfffffffffffffff4ffffffffffffffdaffffffff",
            INIT_32 => X"0000000b000000000000000400000000fffffff5ffffffffffffffe9ffffffff",
            INIT_33 => X"0000001a000000000000001f0000000000000005000000000000001d00000000",
            INIT_34 => X"ffffffdafffffffffffffffcffffffff00000013000000000000000800000000",
            INIT_35 => X"ffffffedfffffffffffffffdffffffffffffffe5ffffffff0000000200000000",
            INIT_36 => X"0000001900000000fffffff0ffffffffffffffeaffffffff0000000200000000",
            INIT_37 => X"0000001500000000fffffff2ffffffff0000001100000000ffffffffffffffff",
            INIT_38 => X"ffffffefffffffff0000000b000000000000000000000000ffffffefffffffff",
            INIT_39 => X"ffffffe2fffffffffffffff1ffffffffffffffc4fffffffffffffff9ffffffff",
            INIT_3A => X"ffffffbdffffffffffffffd8ffffffffffffffc1ffffffffffffff99ffffffff",
            INIT_3B => X"0000002600000000ffffffe9ffffffffffffffb9ffffffffffffffbdffffffff",
            INIT_3C => X"ffffffeeffffffffffffffdfffffffffffffffeffffffffffffffff1ffffffff",
            INIT_3D => X"00000000000000000000001f0000000000000002000000000000001200000000",
            INIT_3E => X"ffffffb8ffffffffffffff7dffffffff00000021000000000000001000000000",
            INIT_3F => X"fffffffcffffffffffffffe4ffffffffffffffd0fffffffffffffff3ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffff68ffffffffffffffb7ffffffffffffffb9ffffffffffffff7bffffffff",
            INIT_41 => X"0000000500000000fffffff9ffffffffffffffa5ffffffffffffff8cffffffff",
            INIT_42 => X"0000000a000000000000000600000000ffffffe2fffffffffffffff5ffffffff",
            INIT_43 => X"0000001e00000000ffffffeaffffffffffffffe6ffffffffffffffd7ffffffff",
            INIT_44 => X"fffffffdfffffffffffffff0ffffffff0000000f00000000fffffffaffffffff",
            INIT_45 => X"fffffff7ffffffff00000023000000000000002a00000000fffffff7ffffffff",
            INIT_46 => X"00000013000000000000000600000000fffffffbffffffffffffffedffffffff",
            INIT_47 => X"000000260000000000000016000000000000001c000000000000003500000000",
            INIT_48 => X"ffffffe6ffffffffffffffe9ffffffff00000022000000000000001400000000",
            INIT_49 => X"0000001f00000000000000200000000000000029000000000000001500000000",
            INIT_4A => X"fffffff3fffffffffffffffcffffffff00000018000000000000002500000000",
            INIT_4B => X"000000220000000000000036000000000000004000000000fffffff8ffffffff",
            INIT_4C => X"0000000700000000000000090000000000000013000000000000002300000000",
            INIT_4D => X"0000000e00000000000000090000000000000022000000000000000c00000000",
            INIT_4E => X"fffffff4ffffffffffffffeeffffffff00000009000000000000002800000000",
            INIT_4F => X"ffffffeffffffffffffffff8ffffffff0000000700000000fffffff0ffffffff",
            INIT_50 => X"0000002c00000000fffffff0ffffffff00000033000000000000002a00000000",
            INIT_51 => X"0000001400000000ffffffe7ffffffff0000000c000000000000000000000000",
            INIT_52 => X"ffffffd2ffffffffffffffc7ffffffffffffffe2ffffffffffffffd3ffffffff",
            INIT_53 => X"ffffff9effffffffffffffbeffffffffffffffbfffffffffffffffd4ffffffff",
            INIT_54 => X"0000001c000000000000001b00000000ffffffecffffffffffffff90ffffffff",
            INIT_55 => X"0000003c000000000000004e0000000000000068000000000000003e00000000",
            INIT_56 => X"0000001b000000000000001d000000000000000a000000000000002300000000",
            INIT_57 => X"fffffff8fffffffffffffff8fffffffffffffffefffffffffffffff9ffffffff",
            INIT_58 => X"ffffffc8ffffffff0000002a000000000000002700000000fffffffbffffffff",
            INIT_59 => X"fffffff0ffffffffffffffe5ffffffffffffffeeffffffff0000000000000000",
            INIT_5A => X"ffffffb0ffffffffffffffb5ffffffffffffff99fffffffffffffffbffffffff",
            INIT_5B => X"0000000a00000000ffffffefffffffff0000000900000000ffffffd0ffffffff",
            INIT_5C => X"ffffffe4ffffffffffffffe2ffffffff0000000300000000ffffffdfffffffff",
            INIT_5D => X"0000002a000000000000000a000000000000002000000000fffffff9ffffffff",
            INIT_5E => X"fffffffcffffffff00000039000000000000004f000000000000005000000000",
            INIT_5F => X"000000170000000000000031000000000000000a00000000fffffff6ffffffff",
            INIT_60 => X"0000002f00000000000000550000000000000020000000000000003400000000",
            INIT_61 => X"0000005c00000000ffffffe7fffffffffffffffcffffffffffffffebffffffff",
            INIT_62 => X"0000009a000000000000008b0000000000000068000000000000006800000000",
            INIT_63 => X"000000730000000000000063000000000000005a000000000000006100000000",
            INIT_64 => X"0000000000000000ffffffdeffffffffffffffe8ffffffff0000002200000000",
            INIT_65 => X"0000005f000000000000001e000000000000000e00000000ffffffddffffffff",
            INIT_66 => X"000000190000000000000006000000000000001e000000000000001300000000",
            INIT_67 => X"fffffff3fffffffffffffffefffffffffffffff9fffffffffffffff6ffffffff",
            INIT_68 => X"00000023000000000000001900000000fffffff7ffffffffffffffefffffffff",
            INIT_69 => X"0000000f00000000000000350000000000000034000000000000001500000000",
            INIT_6A => X"0000000e000000000000000d000000000000001c00000000ffffffd8ffffffff",
            INIT_6B => X"00000034000000000000000b0000000000000018000000000000003300000000",
            INIT_6C => X"0000001900000000000000000000000000000014000000000000001100000000",
            INIT_6D => X"ffffffd4ffffffffffffffd6ffffffffffffffcdffffffffffffffb0ffffffff",
            INIT_6E => X"ffffffd3ffffffffffffffd6ffffffffffffffb5ffffffffffffffbfffffffff",
            INIT_6F => X"ffffffd6ffffffffffffffc0ffffffffffffffb9ffffffffffffffe4ffffffff",
            INIT_70 => X"fffffff0ffffffffffffffd0ffffffffffffffd8ffffffffffffffd9ffffffff",
            INIT_71 => X"0000002500000000fffffffafffffffffffffffcffffffff0000001900000000",
            INIT_72 => X"0000001f000000000000000e0000000000000009000000000000000000000000",
            INIT_73 => X"ffffffa8ffffffff000000260000000000000017000000000000002200000000",
            INIT_74 => X"ffffffb9ffffffffffffffd5ffffffffffffffdaffffffffffffffa2ffffffff",
            INIT_75 => X"ffffffcaffffffffffffffe2ffffffffffffffefffffffffffffffaaffffffff",
            INIT_76 => X"0000004500000000fffffff2ffffffff00000000000000000000001a00000000",
            INIT_77 => X"0000003e00000000000000420000000000000030000000000000003c00000000",
            INIT_78 => X"0000002200000000000000040000000000000006000000000000000b00000000",
            INIT_79 => X"fffffff6ffffffff000000150000000000000030000000000000003400000000",
            INIT_7A => X"fffffffbffffffffffffffe4ffffffffffffffebffffffff0000001c00000000",
            INIT_7B => X"fffffff1ffffffff0000000100000000ffffffd4ffffffff0000001100000000",
            INIT_7C => X"fffffffffffffffffffffff1ffffffffffffffe6ffffffff0000000a00000000",
            INIT_7D => X"fffffff6ffffffff0000001b0000000000000014000000000000001200000000",
            INIT_7E => X"0000000000000000fffffffbffffffff0000000a000000000000000200000000",
            INIT_7F => X"ffffffffffffffff0000000a00000000ffffffeeffffffffffffffddffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE8;


    MEM_IWGHT_LAYER1_INSTANCE9 : if BRAM_NAME = "iwght_layer1_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000ffffffe9ffffffff0000000f000000000000000500000000",
            INIT_01 => X"00000057000000000000003400000000ffffffffffffffffffffffe8ffffffff",
            INIT_02 => X"ffffffd8fffffffffffffff2ffffffffffffffbbffffffffffffffceffffffff",
            INIT_03 => X"ffffffc1ffffffffffffffcaffffffffffffffacffffffffffffffb9ffffffff",
            INIT_04 => X"ffffffdbffffffffffffffe1ffffffffffffffe8ffffffffffffffe9ffffffff",
            INIT_05 => X"ffffffcbffffffffffffffdbffffffffffffffdeffffffffffffffc4ffffffff",
            INIT_06 => X"ffffffe5ffffffffffffffefffffffff0000001200000000ffffffebffffffff",
            INIT_07 => X"fffffff1ffffffffffffffffffffffffffffffbcffffffffffffffb5ffffffff",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE9;


    MEM_IWGHT_LAYER2_INSTANCE0 : if BRAM_NAME = "iwght_layer2_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000eaf0000000000000ef700000000ffffe740ffffffffffffe193ffffffff",
            INIT_01 => X"ffffd593ffffffff000039a400000000ffffd81cffffffff0000244d00000000",
            INIT_02 => X"0000001b000000000000000700000000ffffe228ffffffff0000204700000000",
            INIT_03 => X"000000070000000000000025000000000000000d00000000ffffffefffffffff",
            INIT_04 => X"ffffffa3fffffffffffffffbffffffff00000018000000000000000800000000",
            INIT_05 => X"ffffffdeffffffff0000000600000000fffffff7ffffffff0000000400000000",
            INIT_06 => X"0000002500000000ffffffedffffffffffffffc5ffffffff0000000c00000000",
            INIT_07 => X"ffffffe9ffffffffffffffe0ffffffff0000000400000000fffffffeffffffff",
            INIT_08 => X"0000000300000000ffffffe8ffffffffffffffccffffffffffffffe1ffffffff",
            INIT_09 => X"ffffffeafffffffffffffffeffffffff0000000f00000000ffffffd5ffffffff",
            INIT_0A => X"ffffffc3fffffffffffffff3ffffffff0000000b000000000000004d00000000",
            INIT_0B => X"0000000a00000000fffffffdffffffff0000000500000000ffffffe8ffffffff",
            INIT_0C => X"ffffffedffffffffffffffe2ffffffffffffffffffffffff0000000d00000000",
            INIT_0D => X"fffffff8ffffffff0000002100000000ffffffe9fffffffffffffff7ffffffff",
            INIT_0E => X"0000003200000000000000000000000000000009000000000000001800000000",
            INIT_0F => X"ffffffbdfffffffffffffff9ffffffff0000002d000000000000000a00000000",
            INIT_10 => X"ffffffe9fffffffffffffff9ffffffffffffffc0ffffffff0000000900000000",
            INIT_11 => X"ffffffeefffffffffffffff9ffffffff0000000000000000ffffffe6ffffffff",
            INIT_12 => X"00000011000000000000002f0000000000000016000000000000000000000000",
            INIT_13 => X"00000000000000000000000b000000000000002000000000fffffff6ffffffff",
            INIT_14 => X"ffffffcbffffffff00000000000000000000000800000000ffffffedffffffff",
            INIT_15 => X"fffffff6ffffffffffffffc9ffffffff0000000000000000fffffffdffffffff",
            INIT_16 => X"0000002500000000fffffff1ffffffffffffffeeffffffff0000001600000000",
            INIT_17 => X"fffffff4ffffffff0000000600000000ffffffd4fffffffffffffffbffffffff",
            INIT_18 => X"fffffff2ffffffffffffffd6ffffffffffffffd2ffffffffffffffffffffffff",
            INIT_19 => X"0000000e00000000fffffff8ffffffff0000000500000000ffffffddffffffff",
            INIT_1A => X"000000060000000000000010000000000000000d000000000000001e00000000",
            INIT_1B => X"0000001700000000ffffffedffffffff0000000f00000000ffffffe4ffffffff",
            INIT_1C => X"ffffffebffffffffffffffffffffffff00000022000000000000000200000000",
            INIT_1D => X"0000000600000000ffffffc7ffffffff00000028000000000000001100000000",
            INIT_1E => X"00000020000000000000001f0000000000000002000000000000000d00000000",
            INIT_1F => X"ffffffcffffffffffffffffffffffffffffffff2ffffffff0000000f00000000",
            INIT_20 => X"0000001200000000ffffffdefffffffffffffffaffffffff0000000e00000000",
            INIT_21 => X"fffffffaffffffff00000006000000000000000b00000000ffffffc4ffffffff",
            INIT_22 => X"0000002d000000000000003600000000fffffffaffffffff0000000100000000",
            INIT_23 => X"fffffff8fffffffffffffff5ffffffff0000001300000000ffffffcfffffffff",
            INIT_24 => X"ffffffceffffffff00000001000000000000000600000000fffffff4ffffffff",
            INIT_25 => X"ffffffc1fffffffffffffff4ffffffff0000000b000000000000001300000000",
            INIT_26 => X"0000003200000000000000430000000000000007000000000000000b00000000",
            INIT_27 => X"ffffffebfffffffffffffffaffffffff0000000e00000000ffffffeaffffffff",
            INIT_28 => X"0000001600000000ffffffc0ffffffffffffffbfffffffff0000000000000000",
            INIT_29 => X"ffffffdeffffffff00000002000000000000000000000000fffffff2ffffffff",
            INIT_2A => X"0000000b0000000000000025000000000000000900000000ffffffedffffffff",
            INIT_2B => X"0000001400000000ffffff9fffffffff0000000800000000fffffff3ffffffff",
            INIT_2C => X"ffffffe9ffffffff0000001e00000000ffffffbbffffffff0000000200000000",
            INIT_2D => X"ffffffa4fffffffffffffff0ffffffffffffffcaffffffff0000000500000000",
            INIT_2E => X"0000001b000000000000003f00000000ffffffc9ffffffff0000000b00000000",
            INIT_2F => X"0000000b00000000ffffffeaffffffffffffffe7ffffffffffffffd6ffffffff",
            INIT_30 => X"ffffffeaffffffffffffffbcffffffffffffffd3ffffffff0000001900000000",
            INIT_31 => X"0000000500000000fffffffefffffffffffffffeffffffffffffffdbffffffff",
            INIT_32 => X"0000002b000000000000002400000000fffffffeffffffffffffffeaffffffff",
            INIT_33 => X"ffffffffffffffffffffff9effffffff0000001800000000ffffffd4ffffffff",
            INIT_34 => X"00000005000000000000000600000000ffffffecffffffffffffffffffffffff",
            INIT_35 => X"ffffffa6ffffffffffffffc8fffffffffffffffcfffffffffffffffcffffffff",
            INIT_36 => X"fffffff9ffffffff0000000a00000000ffffffe6ffffffff0000001b00000000",
            INIT_37 => X"fffffffdffffffffffffffebffffffffffffffe0fffffffffffffff7ffffffff",
            INIT_38 => X"fffffff8ffffffffffffffd0fffffffffffffff2fffffffffffffff4ffffffff",
            INIT_39 => X"00000011000000000000000a000000000000000400000000fffffffbffffffff",
            INIT_3A => X"fffffffaffffffffffffffddffffffff00000014000000000000002100000000",
            INIT_3B => X"fffffffbffffffff0000004e00000000fffffffeffffffffffffffdfffffffff",
            INIT_3C => X"0000001400000000ffffffeaffffffff0000000d000000000000001100000000",
            INIT_3D => X"ffffffefffffffff0000000000000000fffffffdffffffff0000000c00000000",
            INIT_3E => X"0000001c00000000ffffffebffffffffffffffcdffffffff0000001000000000",
            INIT_3F => X"0000001200000000ffffffeaffffffffffffffeafffffffffffffff0ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffdaffffffff0000000000000000ffffffe7fffffffffffffff0ffffffff",
            INIT_41 => X"0000001b000000000000000b00000000ffffffeeffffffffffffffe6ffffffff",
            INIT_42 => X"fffffff9ffffffffffffffd0fffffffffffffff9ffffffff0000001400000000",
            INIT_43 => X"fffffff8ffffffff00000039000000000000001100000000fffffffeffffffff",
            INIT_44 => X"ffffffcdffffffffffffffe4ffffffff0000001e000000000000000b00000000",
            INIT_45 => X"0000002f00000000fffffffeffffffff00000024000000000000000600000000",
            INIT_46 => X"0000000c00000000ffffff9efffffffffffffff9ffffffff0000001a00000000",
            INIT_47 => X"ffffffd8fffffffffffffff4ffffffff00000004000000000000000700000000",
            INIT_48 => X"0000001000000000fffffffdffffffffffffffedffffffff0000000300000000",
            INIT_49 => X"000000210000000000000007000000000000000000000000fffffff4ffffffff",
            INIT_4A => X"ffffffffffffffffffffffdeffffffffffffffefffffffff0000002300000000",
            INIT_4B => X"fffffff9ffffffff0000001e000000000000001200000000ffffffefffffffff",
            INIT_4C => X"0000000b00000000fffffff9ffffffff00000054000000000000000000000000",
            INIT_4D => X"0000004300000000ffffffeaffffffff0000000b00000000fffffff8ffffffff",
            INIT_4E => X"0000002b00000000ffffffd0ffffffffffffffd4ffffffff0000000d00000000",
            INIT_4F => X"ffffffdcfffffffffffffff9fffffffffffffff2ffffffff0000000500000000",
            INIT_50 => X"ffffffe4ffffffff0000000a00000000fffffff1fffffffffffffff1ffffffff",
            INIT_51 => X"ffffffedffffffff0000001900000000ffffffefffffffffffffffe8ffffffff",
            INIT_52 => X"0000000b00000000fffffff6ffffffff00000004000000000000000f00000000",
            INIT_53 => X"0000000a0000000000000006000000000000000f000000000000000300000000",
            INIT_54 => X"fffffffcffffffff00000008000000000000000f000000000000001400000000",
            INIT_55 => X"0000003400000000ffffffe4ffffffff00000006000000000000000e00000000",
            INIT_56 => X"0000003600000000ffffffffffffffff0000000000000000fffffff9ffffffff",
            INIT_57 => X"ffffffd5fffffffffffffff8ffffffffffffffdfffffffff0000000500000000",
            INIT_58 => X"0000000a000000000000000800000000ffffffebffffffffffffffefffffffff",
            INIT_59 => X"fffffffaffffffff0000000c000000000000000a00000000ffffffeaffffffff",
            INIT_5A => X"0000001b00000000000000000000000000000006000000000000001100000000",
            INIT_5B => X"0000000000000000fffffff2ffffffff00000003000000000000000000000000",
            INIT_5C => X"00000007000000000000000500000000ffffffe8fffffffffffffff1ffffffff",
            INIT_5D => X"ffffffd6fffffffffffffff9fffffffffffffffcfffffffffffffff5ffffffff",
            INIT_5E => X"0000002b0000000000000004000000000000001400000000ffffffeeffffffff",
            INIT_5F => X"ffffffeafffffffffffffffaffffffff0000000b00000000fffffff6ffffffff",
            INIT_60 => X"0000002c00000000fffffff4ffffffff0000000400000000ffffffffffffffff",
            INIT_61 => X"ffffffe7ffffffff0000000d000000000000000800000000fffffff3ffffffff",
            INIT_62 => X"0000002b0000000000000033000000000000001600000000fffffff4ffffffff",
            INIT_63 => X"fffffff1ffffffffffffffb1ffffffff0000000000000000ffffffefffffffff",
            INIT_64 => X"ffffffeafffffffffffffffbffffffffffffffd9ffffffffffffffefffffffff",
            INIT_65 => X"ffffff85ffffffff000000000000000000000004000000000000000000000000",
            INIT_66 => X"0000002f000000000000003700000000ffffffcdfffffffffffffffdffffffff",
            INIT_67 => X"0000001c0000000000000019000000000000000000000000fffffff3ffffffff",
            INIT_68 => X"00000015000000000000000a000000000000001000000000fffffff8ffffffff",
            INIT_69 => X"0000001a000000000000000300000000ffffffffffffffffffffffffffffffff",
            INIT_6A => X"0000001a000000000000000000000000fffffffafffffffffffffff2ffffffff",
            INIT_6B => X"fffffff8ffffffffffffffb9ffffffff0000000500000000ffffffcdffffffff",
            INIT_6C => X"00000007000000000000001a00000000ffffffdcfffffffffffffff8ffffffff",
            INIT_6D => X"ffffff82ffffffffffffffdeffffffff0000000900000000fffffff4ffffffff",
            INIT_6E => X"ffffffefffffffff0000002e000000000000002000000000fffffffbffffffff",
            INIT_6F => X"0000000200000000ffffffeafffffffffffffff0fffffffffffffffeffffffff",
            INIT_70 => X"000000060000000000000012000000000000000b00000000fffffff3ffffffff",
            INIT_71 => X"ffffffd5fffffffffffffff4ffffffffffffffe3fffffffffffffffdffffffff",
            INIT_72 => X"0000000000000000ffffffd5fffffffffffffffcffffffff0000000200000000",
            INIT_73 => X"fffffff3ffffffff0000006c000000000000000300000000ffffffedffffffff",
            INIT_74 => X"0000000e00000000ffffffd8ffffffff00000010000000000000000400000000",
            INIT_75 => X"000000030000000000000021000000000000001000000000fffffff0ffffffff",
            INIT_76 => X"0000001800000000ffffff7bffffffff0000000a00000000ffffffedffffffff",
            INIT_77 => X"0000001e00000000fffffff9ffffffff0000000400000000ffffffeeffffffff",
            INIT_78 => X"00000000000000000000000e00000000fffffff2ffffffff0000000f00000000",
            INIT_79 => X"0000000c00000000fffffff4ffffffffffffffe6fffffffffffffffeffffffff",
            INIT_7A => X"ffffffe8ffffffffffffffdbffffffff0000001500000000fffffffbffffffff",
            INIT_7B => X"000000120000000000000042000000000000000200000000ffffffffffffffff",
            INIT_7C => X"ffffffe4ffffffffffffffdaffffffff00000030000000000000000f00000000",
            INIT_7D => X"000000400000000000000045000000000000002500000000fffffff4ffffffff",
            INIT_7E => X"0000001c00000000ffffffb0ffffffff0000000000000000ffffffe2ffffffff",
            INIT_7F => X"ffffffdeffffffffffffffedffffffff00000017000000000000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE0;


    MEM_IWGHT_LAYER2_INSTANCE1 : if BRAM_NAME = "iwght_layer2_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000200000000000000017000000000000000800000000fffffff9ffffffff",
            INIT_01 => X"ffffffecffffffffffffffe9fffffffffffffffeffffffff0000001600000000",
            INIT_02 => X"0000000c00000000ffffffe3ffffffff0000000b000000000000001200000000",
            INIT_03 => X"ffffffffffffffff00000019000000000000000000000000fffffffaffffffff",
            INIT_04 => X"ffffffe3fffffffffffffffaffffffff0000001c000000000000000700000000",
            INIT_05 => X"00000014000000000000000b0000000000000017000000000000002700000000",
            INIT_06 => X"0000002f00000000ffffffe7ffffffffffffff9bffffffff0000001500000000",
            INIT_07 => X"ffffffc5ffffffff000000030000000000000002000000000000000700000000",
            INIT_08 => X"fffffffaffffffff0000000e00000000ffffffeaffffffffffffffe2ffffffff",
            INIT_09 => X"ffffffcdffffffff00000000000000000000000200000000fffffff6ffffffff",
            INIT_0A => X"fffffffdfffffffffffffff2ffffffff0000001200000000fffffffaffffffff",
            INIT_0B => X"ffffffffffffffffffffffe5fffffffffffffff4ffffffff0000002a00000000",
            INIT_0C => X"ffffffe9ffffffff0000000e0000000000000026000000000000000700000000",
            INIT_0D => X"00000025000000000000000b0000000000000005000000000000001f00000000",
            INIT_0E => X"00000043000000000000001a00000000ffffffdbffffffff0000001100000000",
            INIT_0F => X"ffffffe0ffffffffffffffe0ffffffff0000000700000000fffffffdffffffff",
            INIT_10 => X"0000000200000000ffffffd7ffffffff00000009000000000000000d00000000",
            INIT_11 => X"ffffffd3ffffffff00000015000000000000002600000000ffffffeaffffffff",
            INIT_12 => X"0000000d00000000ffffffeeffffffff0000000e00000000ffffffe5ffffffff",
            INIT_13 => X"fffffffaffffffffffffffebffffffffffffffeaffffffff0000001100000000",
            INIT_14 => X"ffffffd0ffffffff00000008000000000000000b00000000fffffffaffffffff",
            INIT_15 => X"0000001600000000000000090000000000000003000000000000000000000000",
            INIT_16 => X"0000004c000000000000000e00000000fffffff7ffffffffffffffffffffffff",
            INIT_17 => X"ffffffe2ffffffffffffffdfffffffff00000015000000000000000a00000000",
            INIT_18 => X"0000002600000000ffffffd5fffffffffffffff3ffffffffffffffffffffffff",
            INIT_19 => X"ffffffecfffffffffffffff9ffffffff0000001000000000fffffff4ffffffff",
            INIT_1A => X"0000002500000000fffffff5ffffffff0000000d00000000fffffff0ffffffff",
            INIT_1B => X"0000000b00000000ffffffb4fffffffffffffffaffffffff0000000b00000000",
            INIT_1C => X"ffffffe4ffffffff0000002400000000ffffffcffffffffffffffff2ffffffff",
            INIT_1D => X"ffffffe8ffffffff0000001e000000000000000700000000fffffff4ffffffff",
            INIT_1E => X"0000000a000000000000003a000000000000000c000000000000001200000000",
            INIT_1F => X"0000003600000000ffffffecffffffff0000000600000000fffffff6ffffffff",
            INIT_20 => X"0000002100000000fffffff8ffffffff00000023000000000000000d00000000",
            INIT_21 => X"00000000000000000000000e0000000000000010000000000000000000000000",
            INIT_22 => X"0000003c00000000000000350000000000000001000000000000001b00000000",
            INIT_23 => X"0000001200000000ffffffcafffffffffffffff9ffffffffffffffdbffffffff",
            INIT_24 => X"00000012000000000000000900000000ffffffc7ffffffff0000000700000000",
            INIT_25 => X"fffffff0ffffffff0000000a00000000fffffff3fffffffffffffff3ffffffff",
            INIT_26 => X"ffffffedffffffff0000000d00000000ffffffeeffffffffffffffefffffffff",
            INIT_27 => X"0000004400000000ffffffe8ffffffff0000000000000000ffffffeaffffffff",
            INIT_28 => X"000000480000000000000003000000000000000c00000000fffffff2ffffffff",
            INIT_29 => X"0000000b00000000ffffffeaffffffffffffffe9fffffffffffffffbffffffff",
            INIT_2A => X"ffffffe5ffffffffffffffdcffffffff00000010000000000000000e00000000",
            INIT_2B => X"fffffff8ffffffff0000004400000000ffffffe2ffffffffffffffdbffffffff",
            INIT_2C => X"0000000000000000ffffffefffffffffffffffdeffffffff0000000b00000000",
            INIT_2D => X"ffffffccffffffffffffffe1fffffffffffffffcffffffffffffffefffffffff",
            INIT_2E => X"0000001b00000000ffffffa5ffffffff0000000f00000000fffffff2ffffffff",
            INIT_2F => X"fffffffcffffffffffffffe9ffffffff00000025000000000000002b00000000",
            INIT_30 => X"ffffffe9ffffffffffffffe6ffffffffffffffffffffffffffffffeeffffffff",
            INIT_31 => X"000000040000000000000010000000000000000a000000000000001b00000000",
            INIT_32 => X"0000000400000000fffffff7fffffffffffffff0ffffffff0000000700000000",
            INIT_33 => X"fffffff8ffffffff0000003a000000000000000700000000ffffffe7ffffffff",
            INIT_34 => X"ffffffcfffffffffffffffe6ffffffff00000007000000000000000300000000",
            INIT_35 => X"ffffffc7ffffffff00000043000000000000000200000000ffffffe3ffffffff",
            INIT_36 => X"fffffffbffffffff00000002000000000000000f00000000fffffffeffffffff",
            INIT_37 => X"0000001e00000000fffffff7ffffffff0000004200000000fffffff9ffffffff",
            INIT_38 => X"0000000c00000000fffffff3ffffffff0000001f00000000fffffffaffffffff",
            INIT_39 => X"0000001100000000ffffffd7ffffffffffffffe4ffffffff0000002b00000000",
            INIT_3A => X"0000001e00000000ffffffebffffffffffffffedffffffff0000001000000000",
            INIT_3B => X"00000001000000000000001200000000fffffffaffffffffffffffeeffffffff",
            INIT_3C => X"ffffffd8fffffffffffffff2ffffffff0000000800000000fffffffcffffffff",
            INIT_3D => X"ffffffeaffffffff00000054000000000000000b000000000000000000000000",
            INIT_3E => X"ffffffeaffffffff0000000300000000ffffffdcffffffff0000000600000000",
            INIT_3F => X"0000001400000000ffffffccffffffff00000032000000000000000200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001a00000000fffffffafffffffffffffffbffffffffffffffcfffffffff",
            INIT_41 => X"ffffffb5ffffffffffffffe4ffffffff0000002f000000000000001200000000",
            INIT_42 => X"00000019000000000000001900000000fffffff5ffffffffffffffe9ffffffff",
            INIT_43 => X"fffffff4ffffffff0000001e00000000ffffffcaffffffff0000001000000000",
            INIT_44 => X"fffffff1fffffffffffffff6ffffffff00000009000000000000001500000000",
            INIT_45 => X"000000060000000000000011000000000000000f000000000000001400000000",
            INIT_46 => X"000000060000000000000003000000000000000e00000000fffffffaffffffff",
            INIT_47 => X"0000000900000000ffffffd6ffffffffffffffffffffffff0000000d00000000",
            INIT_48 => X"0000002100000000ffffffeeffffffff0000001800000000ffffffd5ffffffff",
            INIT_49 => X"ffffffdefffffffffffffff7ffffffff0000003e000000000000000000000000",
            INIT_4A => X"0000001c00000000ffffffe2ffffffff00000010000000000000000300000000",
            INIT_4B => X"00000018000000000000000100000000ffffffcffffffffffffffffeffffffff",
            INIT_4C => X"ffffffd2fffffffffffffff6ffffffff00000010000000000000000a00000000",
            INIT_4D => X"0000000a0000000000000014000000000000000800000000fffffff8ffffffff",
            INIT_4E => X"0000000f00000000000000110000000000000033000000000000000d00000000",
            INIT_4F => X"0000000100000000ffffffd2ffffffff0000001a000000000000001700000000",
            INIT_50 => X"0000002600000000ffffffcefffffffffffffff9ffffffffffffffe4ffffffff",
            INIT_51 => X"ffffffc6fffffffffffffffbffffffff00000027000000000000001d00000000",
            INIT_52 => X"00000000000000000000000500000000fffffffaffffffff0000000d00000000",
            INIT_53 => X"ffffffebffffffffffffffedffffffff0000000000000000fffffff8ffffffff",
            INIT_54 => X"ffffffd4fffffffffffffff3ffffffffffffffe2ffffffffffffffedffffffff",
            INIT_55 => X"fffffffcffffffff00000053000000000000001400000000ffffffebffffffff",
            INIT_56 => X"ffffffe5ffffffff000000230000000000000023000000000000000c00000000",
            INIT_57 => X"0000002200000000ffffffddffffffff00000015000000000000000d00000000",
            INIT_58 => X"0000003000000000ffffffdeffffffff0000000900000000ffffffdbffffffff",
            INIT_59 => X"ffffffddfffffffffffffff9ffffffff0000000c000000000000001b00000000",
            INIT_5A => X"fffffffaffffffff0000000800000000fffffffcffffffff0000001b00000000",
            INIT_5B => X"0000001300000000ffffffcaffffffff0000000d00000000ffffffd5ffffffff",
            INIT_5C => X"fffffff8ffffffff0000001700000000ffffffe2ffffffffffffffeaffffffff",
            INIT_5D => X"ffffffc1ffffffff00000029000000000000000e00000000ffffffe8ffffffff",
            INIT_5E => X"ffffffcfffffffff0000000d00000000fffffff3ffffffffffffffefffffffff",
            INIT_5F => X"0000001e00000000fffffff6ffffffff0000001a00000000ffffffe4ffffffff",
            INIT_60 => X"0000003e00000000ffffffd7fffffffffffffffcfffffffffffffff9ffffffff",
            INIT_61 => X"0000000e00000000fffffff0ffffffffffffffedffffffff0000002100000000",
            INIT_62 => X"0000000500000000ffffffeefffffffffffffff0ffffffff0000000800000000",
            INIT_63 => X"0000001600000000fffffff9ffffffff0000000c00000000ffffffeaffffffff",
            INIT_64 => X"ffffffd0ffffffff0000001500000000ffffffb6ffffffff0000001900000000",
            INIT_65 => X"ffffffceffffffff000000060000000000000000000000000000001400000000",
            INIT_66 => X"0000000600000000ffffffc9ffffffff0000003c000000000000000800000000",
            INIT_67 => X"000000020000000000000004000000000000002d000000000000002200000000",
            INIT_68 => X"0000000f00000000ffffffe8ffffffffffffffebffffffff0000001000000000",
            INIT_69 => X"00000003000000000000001500000000fffffffefffffffffffffffeffffffff",
            INIT_6A => X"0000000200000000ffffffe8ffffffff00000001000000000000000f00000000",
            INIT_6B => X"fffffff8ffffffff0000000a00000000fffffff8fffffffffffffffaffffffff",
            INIT_6C => X"fffffffdffffffff0000000300000000fffffffffffffffffffffffbffffffff",
            INIT_6D => X"ffffff73ffffffff0000003e00000000ffffffe5ffffffff0000000000000000",
            INIT_6E => X"ffffffe9ffffffffffffffe5ffffffffffffffefffffffff0000000400000000",
            INIT_6F => X"0000000c00000000ffffffe7ffffffff0000002b00000000ffffffe2ffffffff",
            INIT_70 => X"0000001700000000ffffffcdfffffffffffffff9fffffffffffffffaffffffff",
            INIT_71 => X"0000000800000000ffffffe8ffffffff00000004000000000000002300000000",
            INIT_72 => X"0000000b00000000ffffffd5ffffffffffffffe6ffffffff0000002500000000",
            INIT_73 => X"00000000000000000000000200000000ffffffeaffffffff0000001200000000",
            INIT_74 => X"ffffffd7ffffffff0000000000000000ffffffcffffffffffffffff8ffffffff",
            INIT_75 => X"ffffffd1ffffffff0000003000000000ffffffe2ffffffffffffffdbffffffff",
            INIT_76 => X"fffffff3ffffffffffffffdcffffffff0000001b000000000000000000000000",
            INIT_77 => X"0000001900000000ffffffd8ffffffff0000000400000000fffffffcffffffff",
            INIT_78 => X"0000001b00000000ffffffd5ffffffff0000000c00000000ffffffd4ffffffff",
            INIT_79 => X"ffffffe1ffffffffffffffe6ffffffff0000000b000000000000001900000000",
            INIT_7A => X"0000000d00000000ffffffecffffffffffffffeaffffffff0000000600000000",
            INIT_7B => X"00000019000000000000001e00000000ffffffdfffffffff0000002300000000",
            INIT_7C => X"fffffff8fffffffffffffffdffffffff0000000600000000fffffff6ffffffff",
            INIT_7D => X"fffffff1ffffffff0000002500000000ffffffebffffffff0000000800000000",
            INIT_7E => X"0000001900000000000000060000000000000007000000000000001a00000000",
            INIT_7F => X"ffffffe4ffffffffffffffd1ffffffff00000017000000000000001c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE1;


    MEM_IWGHT_LAYER2_INSTANCE2 : if BRAM_NAME = "iwght_layer2_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001600000000ffffffdbffffffff0000000100000000fffffff3ffffffff",
            INIT_01 => X"ffffffd0fffffffffffffff8ffffffff00000004000000000000001b00000000",
            INIT_02 => X"0000000000000000ffffffe9ffffffffffffffe9ffffffff0000000100000000",
            INIT_03 => X"0000000f000000000000000f00000000ffffffe8ffffffff0000002800000000",
            INIT_04 => X"ffffffd6fffffffffffffffeffffffff0000002a00000000fffffffeffffffff",
            INIT_05 => X"ffffffffffffffff0000000700000000ffffffe0fffffffffffffff8ffffffff",
            INIT_06 => X"fffffff5ffffffffffffffebffffffff00000023000000000000000000000000",
            INIT_07 => X"fffffff3ffffffffffffffdcfffffffffffffff2ffffffff0000002900000000",
            INIT_08 => X"0000001d00000000ffffffebffffffff0000000a000000000000000200000000",
            INIT_09 => X"ffffffd7fffffffffffffff3ffffffff0000000d000000000000001c00000000",
            INIT_0A => X"fffffffcffffffffffffffe8fffffffffffffffafffffffffffffffeffffffff",
            INIT_0B => X"0000001400000000ffffffdffffffffffffffffeffffffff0000000800000000",
            INIT_0C => X"ffffffd4ffffffff0000000900000000fffffff2fffffffffffffff4ffffffff",
            INIT_0D => X"ffffffd0ffffffff0000001e00000000fffffff7ffffffff0000000900000000",
            INIT_0E => X"0000000c00000000fffffff4ffffffffffffffdeffffffff0000001c00000000",
            INIT_0F => X"ffffffdfffffffffffffffc8ffffffff0000000b000000000000001f00000000",
            INIT_10 => X"0000002700000000fffffffbffffffffffffffdffffffffffffffff2ffffffff",
            INIT_11 => X"ffffffccffffffff000000040000000000000019000000000000001100000000",
            INIT_12 => X"ffffffe7ffffffffffffffbeffffffffffffffefffffffff0000000500000000",
            INIT_13 => X"fffffff8ffffffffffffffd6ffffffff0000001100000000ffffffe5ffffffff",
            INIT_14 => X"ffffffc5ffffffffffffffebffffffff00000000000000000000000a00000000",
            INIT_15 => X"ffffffd7ffffffff0000001000000000fffffff3ffffffff0000000000000000",
            INIT_16 => X"00000022000000000000001b0000000000000009000000000000001500000000",
            INIT_17 => X"0000001f00000000ffffffefffffffff0000004300000000fffffff1ffffffff",
            INIT_18 => X"fffffff8ffffffffffffffdbffffffffffffffd0fffffffffffffff5ffffffff",
            INIT_19 => X"0000000100000000fffffff7fffffffffffffffeffffffff0000000e00000000",
            INIT_1A => X"ffffffe8ffffffffffffffe4ffffffff00000004000000000000002300000000",
            INIT_1B => X"0000001600000000ffffffe8ffffffffffffffecffffffffffffffe0ffffffff",
            INIT_1C => X"00000005000000000000004c00000000ffffffddffffffff0000001500000000",
            INIT_1D => X"ffffffa9fffffffffffffffcffffffff0000000b000000000000001800000000",
            INIT_1E => X"ffffffeafffffffffffffff0ffffffff00000069000000000000001c00000000",
            INIT_1F => X"0000000c000000000000000c0000000000000001000000000000000200000000",
            INIT_20 => X"0000000400000000ffffffcdffffffff0000002300000000ffffffe5ffffffff",
            INIT_21 => X"0000001b000000000000001600000000ffffffdcffffffff0000002000000000",
            INIT_22 => X"0000001300000000fffffff0ffffffff00000015000000000000002700000000",
            INIT_23 => X"0000000f00000000ffffffd5fffffffffffffff7ffffffffffffffdeffffffff",
            INIT_24 => X"fffffff0ffffffff0000001700000000ffffffe1fffffffffffffff4ffffffff",
            INIT_25 => X"ffffffa0ffffffffffffffffffffffff0000001800000000fffffffdffffffff",
            INIT_26 => X"fffffff7fffffffffffffffcffffffff0000000d00000000ffffffe6ffffffff",
            INIT_27 => X"0000001f000000000000000a000000000000000e00000000fffffff6ffffffff",
            INIT_28 => X"fffffffdffffffffffffffc7fffffffffffffff3ffffffff0000000000000000",
            INIT_29 => X"fffffffbffffffff0000001600000000fffffff9ffffffff0000001b00000000",
            INIT_2A => X"0000001b00000000fffffffcffffffff0000000f000000000000000500000000",
            INIT_2B => X"0000000f000000000000000b0000000000000008000000000000002400000000",
            INIT_2C => X"fffffffdffffffff0000002c00000000ffffffccfffffffffffffff5ffffffff",
            INIT_2D => X"ffffffaeffffffffffffffe9ffffffff0000000b000000000000000700000000",
            INIT_2E => X"0000000700000000ffffffeafffffffffffffff5ffffffff0000001200000000",
            INIT_2F => X"0000002e000000000000001b000000000000000c00000000ffffffefffffffff",
            INIT_30 => X"0000001400000000fffffffbffffffff00000014000000000000000700000000",
            INIT_31 => X"ffffffefffffffff0000001800000000ffffffeeffffffff0000000a00000000",
            INIT_32 => X"0000000b00000000ffffffd9fffffffffffffff7ffffffff0000000500000000",
            INIT_33 => X"000000230000000000000000000000000000000e000000000000002a00000000",
            INIT_34 => X"fffffff8ffffffff00000022000000000000002900000000fffffff4ffffffff",
            INIT_35 => X"fffffff0ffffffff0000000a000000000000000c000000000000000f00000000",
            INIT_36 => X"00000022000000000000000200000000ffffffd2ffffffff0000001400000000",
            INIT_37 => X"fffffff3ffffffffffffffffffffffff00000017000000000000001200000000",
            INIT_38 => X"0000001800000000fffffff2ffffffff00000010000000000000000d00000000",
            INIT_39 => X"fffffffcffffffff000000130000000000000005000000000000001c00000000",
            INIT_3A => X"ffffffe7fffffffffffffff3ffffffff0000000c000000000000000200000000",
            INIT_3B => X"000000010000000000000015000000000000000b000000000000001200000000",
            INIT_3C => X"ffffffd7ffffffff0000000600000000fffffff3ffffffffffffffebffffffff",
            INIT_3D => X"ffffffd7fffffffffffffffeffffffff0000001f000000000000001000000000",
            INIT_3E => X"fffffffcffffffffffffffeeffffffffffffffa2ffffffff0000001300000000",
            INIT_3F => X"fffffffffffffffffffffffefffffffffffffff9ffffffff0000002a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001b0000000000000009000000000000000b00000000ffffffffffffffff",
            INIT_41 => X"ffffffedfffffffffffffffbffffffff00000000000000000000000700000000",
            INIT_42 => X"ffffffd3ffffffffffffffd8ffffffffffffffffffffffff0000000a00000000",
            INIT_43 => X"ffffffe0ffffffff00000052000000000000000600000000fffffff8ffffffff",
            INIT_44 => X"ffffffccffffffff0000000100000000fffffffefffffffffffffffdffffffff",
            INIT_45 => X"ffffffd6ffffffff0000000a0000000000000000000000000000001800000000",
            INIT_46 => X"0000000a000000000000000100000000ffffffbdffffffff0000000f00000000",
            INIT_47 => X"fffffff3ffffffff0000000500000000fffffff4ffffffff0000001800000000",
            INIT_48 => X"fffffff8ffffffffffffffd6ffffffffffffffe1ffffffffffffffdcffffffff",
            INIT_49 => X"fffffff1fffffffffffffff9fffffffffffffff2ffffffff0000001300000000",
            INIT_4A => X"ffffffa4ffffffffffffffe2fffffffffffffff1fffffffffffffffcffffffff",
            INIT_4B => X"0000000c000000000000001e000000000000001700000000ffffffe4ffffffff",
            INIT_4C => X"ffffffa9ffffffffffffffe0ffffffffffffffeafffffffffffffffeffffffff",
            INIT_4D => X"0000000100000000fffffffeffffffff00000029000000000000001a00000000",
            INIT_4E => X"0000001b00000000ffffffe1ffffffff00000000000000000000000b00000000",
            INIT_4F => X"fffffff8ffffffffffffffdffffffffffffffffcffffffff0000001200000000",
            INIT_50 => X"ffffffecffffffff0000000300000000ffffffe3fffffffffffffffaffffffff",
            INIT_51 => X"ffffffe7fffffffffffffffeffffffffffffffedffffffff0000000600000000",
            INIT_52 => X"fffffffbffffffffffffffecffffffff00000012000000000000000300000000",
            INIT_53 => X"0000001000000000ffffff9bffffffff0000001a00000000ffffffefffffffff",
            INIT_54 => X"00000003000000000000002100000000ffffffd3fffffffffffffff7ffffffff",
            INIT_55 => X"ffffffd5ffffffffffffffe7fffffffffffffffaffffffff0000001700000000",
            INIT_56 => X"fffffff9ffffffff0000000d000000000000002b00000000fffffff3ffffffff",
            INIT_57 => X"0000000d0000000000000012000000000000000400000000ffffffefffffffff",
            INIT_58 => X"0000000e00000000ffffff93fffffffffffffff0ffffffffffffffedffffffff",
            INIT_59 => X"00000001000000000000000600000000ffffffd8ffffffff0000000400000000",
            INIT_5A => X"0000003d00000000ffffffe1ffffffff00000004000000000000002400000000",
            INIT_5B => X"0000000a00000000ffffff9fffffffff00000014000000000000000400000000",
            INIT_5C => X"fffffffeffffffff0000002900000000ffffffe4fffffffffffffffbffffffff",
            INIT_5D => X"ffffff80fffffffffffffff4ffffffff0000000c000000000000001c00000000",
            INIT_5E => X"0000000700000000fffffff8ffffffff00000027000000000000002600000000",
            INIT_5F => X"0000000f0000000000000005000000000000000600000000fffffff7ffffffff",
            INIT_60 => X"0000000d00000000ffffffbbffffffffffffffe2fffffffffffffff2ffffffff",
            INIT_61 => X"00000005000000000000000300000000fffffff8fffffffffffffff8ffffffff",
            INIT_62 => X"0000000800000000000000040000000000000021000000000000001400000000",
            INIT_63 => X"fffffff6fffffffffffffff2fffffffffffffffaffffffff0000001d00000000",
            INIT_64 => X"00000017000000000000001e00000000ffffffe5fffffffffffffffbffffffff",
            INIT_65 => X"0000000d00000000fffffffcffffffff0000001f000000000000001e00000000",
            INIT_66 => X"0000001f000000000000000400000000fffffff5ffffffff0000002400000000",
            INIT_67 => X"00000015000000000000000e0000000000000010000000000000000000000000",
            INIT_68 => X"fffffffaffffffffffffffd6ffffffffffffffddffffffff0000000200000000",
            INIT_69 => X"00000015000000000000002200000000fffffffcfffffffffffffff3ffffffff",
            INIT_6A => X"0000001500000000000000020000000000000030000000000000000600000000",
            INIT_6B => X"0000000700000000ffffffe4ffffffff00000018000000000000000400000000",
            INIT_6C => X"0000000d000000000000000800000000fffffff3ffffffff0000002800000000",
            INIT_6D => X"fffffffcffffffffffffffe8ffffffff00000035000000000000004700000000",
            INIT_6E => X"0000002400000000ffffffefffffffffffffffcaffffffff0000001000000000",
            INIT_6F => X"ffffffe7ffffffff000000010000000000000005000000000000000200000000",
            INIT_70 => X"ffffffeaffffffffffffffb8fffffffffffffff6ffffffff0000000800000000",
            INIT_71 => X"fffffff6ffffffff00000016000000000000001300000000ffffffefffffffff",
            INIT_72 => X"0000000a00000000fffffffcffffffff00000038000000000000001100000000",
            INIT_73 => X"fffffffdffffffff0000001c0000000000000011000000000000000c00000000",
            INIT_74 => X"0000001d00000000fffffffcffffffff0000000f000000000000001200000000",
            INIT_75 => X"fffffff1ffffffff0000000c0000000000000018000000000000002200000000",
            INIT_76 => X"00000018000000000000000800000000ffffff9effffffff0000002c00000000",
            INIT_77 => X"ffffffe1ffffffff0000000c000000000000001800000000fffffff9ffffffff",
            INIT_78 => X"0000000000000000ffffffe3ffffffff0000000800000000ffffffffffffffff",
            INIT_79 => X"0000000e000000000000000f000000000000000000000000fffffff5ffffffff",
            INIT_7A => X"ffffffdaffffffffffffffd3ffffffff0000001e000000000000001200000000",
            INIT_7B => X"fffffff6ffffffff0000002f0000000000000007000000000000000200000000",
            INIT_7C => X"0000000200000000fffffff9ffffffff0000000b00000000fffffffdffffffff",
            INIT_7D => X"0000001700000000ffffffeaffffffff0000000d000000000000002b00000000",
            INIT_7E => X"fffffffeffffffffffffffc6ffffffff00000004000000000000002c00000000",
            INIT_7F => X"ffffffe4fffffffffffffffcfffffffffffffff3ffffffff0000001500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE2;


    MEM_IWGHT_LAYER2_INSTANCE3 : if BRAM_NAME = "iwght_layer2_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff1ffffffffffffffdeffffffffffffffeffffffffffffffffdffffffff",
            INIT_01 => X"fffffffcfffffffffffffff3ffffffffffffffedffffffff0000000300000000",
            INIT_02 => X"ffffffd5ffffffffffffff86ffffffff0000001b000000000000000500000000",
            INIT_03 => X"0000000c000000000000004e000000000000002d00000000fffffffcffffffff",
            INIT_04 => X"ffffffcfffffffff00000015000000000000000f000000000000000500000000",
            INIT_05 => X"ffffffeffffffffffffffffffffffffffffffffaffffffff0000000a00000000",
            INIT_06 => X"0000000b00000000ffffffc5fffffffffffffff7ffffffff0000002100000000",
            INIT_07 => X"ffffffeaffffffff0000001300000000fffffff3fffffffffffffffaffffffff",
            INIT_08 => X"ffffffc5fffffffffffffff3ffffffffffffffeafffffffffffffffcffffffff",
            INIT_09 => X"fffffffbffffffff0000000000000000ffffffdeffffffff0000001a00000000",
            INIT_0A => X"ffffffd0ffffffffffffffebffffffff00000009000000000000000700000000",
            INIT_0B => X"0000000500000000fffffffeffffffff0000000100000000ffffffebffffffff",
            INIT_0C => X"0000006600000000fffffffeffffffff00000006000000000000000300000000",
            INIT_0D => X"0000000a00000000000000320000000000000009000000000000000f00000000",
            INIT_0E => X"ffffffe0ffffffffffffffdffffffffffffffff8fffffffffffffff3ffffffff",
            INIT_0F => X"000000030000000000000005000000000000001c00000000ffffffffffffffff",
            INIT_10 => X"0000001900000000ffffffddffffffff0000001b00000000ffffffffffffffff",
            INIT_11 => X"00000010000000000000001500000000ffffffe8ffffffff0000001d00000000",
            INIT_12 => X"00000002000000000000001100000000fffffff7ffffffff0000003b00000000",
            INIT_13 => X"00000008000000000000000700000000fffffffffffffffffffffff2ffffffff",
            INIT_14 => X"0000003000000000fffffff2fffffffffffffff6ffffffff0000000500000000",
            INIT_15 => X"0000000100000000ffffffc6fffffffffffffff7ffffffff0000000600000000",
            INIT_16 => X"0000000f00000000ffffffdfffffffff0000003900000000fffffff9ffffffff",
            INIT_17 => X"fffffffcffffffff0000002500000000ffffffccffffffffffffffebffffffff",
            INIT_18 => X"0000001400000000ffffffe9ffffffff0000002f000000000000000200000000",
            INIT_19 => X"0000001400000000fffffff1ffffffffffffffe4ffffffffffffffffffffffff",
            INIT_1A => X"0000000e00000000ffffffe2ffffffffffffffffffffffff0000001500000000",
            INIT_1B => X"0000000700000000fffffff5fffffffffffffffdffffffff0000000400000000",
            INIT_1C => X"00000039000000000000001d0000000000000003000000000000000300000000",
            INIT_1D => X"ffffffe2fffffffffffffffffffffffffffffff7ffffffff0000000300000000",
            INIT_1E => X"ffffffe2ffffffff0000002100000000ffffffe6ffffffff0000000a00000000",
            INIT_1F => X"ffffffffffffffff0000001500000000fffffff2ffffffffffffffeaffffffff",
            INIT_20 => X"ffffffccffffffffffffffedffffffff00000019000000000000000000000000",
            INIT_21 => X"00000018000000000000000100000000fffffff3ffffffff0000000800000000",
            INIT_22 => X"0000002a00000000fffffff6ffffffff00000012000000000000000b00000000",
            INIT_23 => X"00000005000000000000000700000000fffffff1ffffffff0000000100000000",
            INIT_24 => X"00000002000000000000000a00000000fffffffdfffffffffffffffeffffffff",
            INIT_25 => X"ffffffd2fffffffffffffffbffffffffffffffecfffffffffffffff1ffffffff",
            INIT_26 => X"ffffffefffffffff0000000e00000000ffffffd9ffffffff0000001200000000",
            INIT_27 => X"fffffffeffffffffffffffdeffffffff0000000e00000000fffffffdffffffff",
            INIT_28 => X"0000001900000000ffffffefffffffff0000002d00000000ffffffffffffffff",
            INIT_29 => X"fffffffeffffffff0000000600000000fffffff7ffffffff0000000300000000",
            INIT_2A => X"ffffffebfffffffffffffffbffffffffffffffeaffffffff0000001200000000",
            INIT_2B => X"000000000000000000000025000000000000000d00000000fffffff8ffffffff",
            INIT_2C => X"0000000800000000fffffff3ffffffff0000000f00000000fffffff2ffffffff",
            INIT_2D => X"000000140000000000000000000000000000002600000000fffffff4ffffffff",
            INIT_2E => X"ffffffeeffffffffffffffe7ffffffffffffffdbffffffff0000000100000000",
            INIT_2F => X"ffffffdfffffffff000000000000000000000001000000000000000700000000",
            INIT_30 => X"0000000b0000000000000012000000000000002300000000fffffff0ffffffff",
            INIT_31 => X"fffffff1ffffffff0000000d00000000fffffff7fffffffffffffffaffffffff",
            INIT_32 => X"ffffffe1ffffffffffffffecffffffffffffffeaffffffffffffffedffffffff",
            INIT_33 => X"0000001e0000000000000012000000000000001200000000fffffff1ffffffff",
            INIT_34 => X"0000002000000000fffffffaffffffffffffffeefffffffffffffff5ffffffff",
            INIT_35 => X"000000210000000000000020000000000000000500000000fffffffbffffffff",
            INIT_36 => X"fffffff2ffffffffffffffe4ffffffff0000001800000000fffffff6ffffffff",
            INIT_37 => X"00000007000000000000000f00000000ffffffdbffffffff0000000f00000000",
            INIT_38 => X"0000001f000000000000001100000000fffffffcfffffffffffffff9ffffffff",
            INIT_39 => X"0000000f000000000000000300000000ffffffebfffffffffffffffcffffffff",
            INIT_3A => X"0000000900000000fffffffbfffffffffffffff5ffffffffffffffdfffffffff",
            INIT_3B => X"fffffff2ffffffff0000000b000000000000000000000000ffffffd2ffffffff",
            INIT_3C => X"0000002900000000fffffff8ffffffffffffffe2ffffffffffffffffffffffff",
            INIT_3D => X"00000011000000000000000900000000fffffff6ffffffff0000001200000000",
            INIT_3E => X"ffffffe4ffffffff0000000f000000000000001500000000fffffff7ffffffff",
            INIT_3F => X"0000002a000000000000001c00000000ffffffedfffffffffffffff1ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000d0000000000000017000000000000001c00000000fffffffeffffffff",
            INIT_41 => X"0000001a000000000000000000000000ffffffdaffffffff0000001700000000",
            INIT_42 => X"fffffff8ffffffffffffffe4ffffffffffffffe0fffffffffffffff3ffffffff",
            INIT_43 => X"0000000b00000000fffffff1ffffffff0000000a000000000000000000000000",
            INIT_44 => X"fffffffdffffffff0000000d00000000fffffff3ffffffff0000000600000000",
            INIT_45 => X"ffffffe3ffffffff0000001800000000ffffffe7fffffffffffffffbffffffff",
            INIT_46 => X"ffffffe7ffffffffffffffedffffffff0000000800000000ffffffffffffffff",
            INIT_47 => X"fffffffdffffffff00000015000000000000000300000000ffffffcbffffffff",
            INIT_48 => X"0000002600000000ffffffdaffffffffffffffe7ffffffff0000000900000000",
            INIT_49 => X"0000001c000000000000000d00000000ffffffe6ffffffff0000000300000000",
            INIT_4A => X"0000000f00000000fffffff1ffffffffffffffecffffffff0000001500000000",
            INIT_4B => X"fffffff3ffffffffffffffecffffffff00000002000000000000000800000000",
            INIT_4C => X"00000021000000000000000a0000000000000005000000000000000000000000",
            INIT_4D => X"ffffffdafffffffffffffff5ffffffff0000000a00000000fffffff6ffffffff",
            INIT_4E => X"fffffffdffffffffffffffdcffffffff0000001800000000fffffff3ffffffff",
            INIT_4F => X"00000008000000000000000600000000fffffff2ffffffffffffffddffffffff",
            INIT_50 => X"0000000a00000000fffffff1ffffffffffffffeffffffffffffffffeffffffff",
            INIT_51 => X"ffffffffffffffffffffffe9ffffffffffffffecfffffffffffffffeffffffff",
            INIT_52 => X"0000002d00000000ffffffe4fffffffffffffff8ffffffffffffffd0ffffffff",
            INIT_53 => X"ffffffe5fffffffffffffff3fffffffffffffff2ffffffff0000000300000000",
            INIT_54 => X"ffffffd7ffffffffffffffecffffffffffffffd7ffffffff0000000800000000",
            INIT_55 => X"fffffff0ffffffff0000001f00000000ffffffebffffffffffffffebffffffff",
            INIT_56 => X"fffffffaffffffff0000002400000000ffffffb5fffffffffffffffdffffffff",
            INIT_57 => X"ffffffdcfffffffffffffff2ffffffff0000002a00000000fffffff6ffffffff",
            INIT_58 => X"0000000700000000fffffff8ffffffff0000000c00000000fffffff8ffffffff",
            INIT_59 => X"0000000900000000fffffff4ffffffff0000000600000000ffffffeeffffffff",
            INIT_5A => X"0000003300000000ffffffdcffffffff0000000100000000ffffffe0ffffffff",
            INIT_5B => X"ffffffebffffffff0000000700000000ffffffeaffffffff0000000100000000",
            INIT_5C => X"ffffffd8fffffffffffffffcffffffffffffffe7fffffffffffffff0ffffffff",
            INIT_5D => X"ffffffc2ffffffff0000000a00000000fffffffefffffffffffffff8ffffffff",
            INIT_5E => X"ffffffc0ffffffff0000000600000000ffffffdfffffffff0000001400000000",
            INIT_5F => X"fffffff4ffffffffffffffe5ffffffff0000001c000000000000001900000000",
            INIT_60 => X"fffffffeffffffffffffffe7ffffffff0000000e00000000ffffffd8ffffffff",
            INIT_61 => X"ffffffceffffffffffffffd9ffffffff0000002200000000fffffff5ffffffff",
            INIT_62 => X"0000001100000000ffffffceffffffff0000001a00000000ffffffd9ffffffff",
            INIT_63 => X"ffffffffffffffff0000002900000000fffffffaffffffff0000000b00000000",
            INIT_64 => X"fffffff6ffffffffffffffebfffffffffffffff7fffffffffffffff9ffffffff",
            INIT_65 => X"fffffffaffffffff00000000000000000000001c00000000ffffffd6ffffffff",
            INIT_66 => X"0000000000000000fffffff3ffffffffffffffe5ffffffff0000000f00000000",
            INIT_67 => X"ffffffe0ffffffffffffffe1ffffffff0000002b000000000000003200000000",
            INIT_68 => X"fffffff8fffffffffffffffeffffffff0000001c00000000fffffffeffffffff",
            INIT_69 => X"fffffffbffffffffffffffddffffffff0000000a00000000ffffffecffffffff",
            INIT_6A => X"ffffffe4ffffffffffffffe7ffffffff0000001100000000ffffffcbffffffff",
            INIT_6B => X"fffffff1ffffffff000000160000000000000014000000000000000c00000000",
            INIT_6C => X"fffffff5ffffffff0000000000000000ffffffe6fffffffffffffff3ffffffff",
            INIT_6D => X"fffffffaffffffff0000000e000000000000001200000000ffffffe6ffffffff",
            INIT_6E => X"00000013000000000000000500000000fffffffffffffffffffffffcffffffff",
            INIT_6F => X"ffffffe1ffffffffffffffebfffffffffffffff3ffffffff0000001f00000000",
            INIT_70 => X"0000001a00000000fffffffbfffffffffffffff7fffffffffffffff0ffffffff",
            INIT_71 => X"0000000a00000000fffffffeffffffff0000000b000000000000000100000000",
            INIT_72 => X"fffffff8fffffffffffffff1ffffffff0000001600000000ffffffe3ffffffff",
            INIT_73 => X"000000000000000000000014000000000000001300000000ffffffefffffffff",
            INIT_74 => X"0000000600000000ffffffe6ffffffff0000000500000000fffffff2ffffffff",
            INIT_75 => X"0000000500000000fffffff9fffffffffffffff2ffffffff0000001500000000",
            INIT_76 => X"fffffff6ffffffff0000000000000000ffffffdbffffffffffffffefffffffff",
            INIT_77 => X"00000032000000000000000000000000fffffffcffffffffffffffd6ffffffff",
            INIT_78 => X"0000001200000000ffffffebffffffff0000000f000000000000000900000000",
            INIT_79 => X"0000002300000000ffffffeeffffffffffffffe1ffffffffffffffffffffffff",
            INIT_7A => X"ffffffe4fffffffffffffff8fffffffffffffff7ffffffffffffffefffffffff",
            INIT_7B => X"0000000b00000000ffffffdfffffffff0000000c000000000000002200000000",
            INIT_7C => X"fffffffeffffffff0000000a0000000000000021000000000000000900000000",
            INIT_7D => X"ffffffdeffffffff0000001900000000ffffffe5ffffffffffffffe1ffffffff",
            INIT_7E => X"fffffff9ffffffff0000000800000000ffffffa4fffffffffffffff4ffffffff",
            INIT_7F => X"0000001400000000fffffff7fffffffffffffff6ffffffffffffffe7ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE3;


    MEM_IWGHT_LAYER2_INSTANCE4 : if BRAM_NAME = "iwght_layer2_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002300000000fffffff2ffffffffffffffdcffffffff0000000200000000",
            INIT_01 => X"0000001d000000000000000100000000ffffffd5fffffffffffffffaffffffff",
            INIT_02 => X"fffffffbffffffffffffffeeffffffff0000000c000000000000000f00000000",
            INIT_03 => X"fffffffaffffffffffffffe8ffffffff00000017000000000000002800000000",
            INIT_04 => X"ffffffe4ffffffff0000000a0000000000000019000000000000000800000000",
            INIT_05 => X"0000001d000000000000001e00000000ffffffeeffffffffffffffefffffffff",
            INIT_06 => X"0000000100000000fffffff7ffffffffffffffdaffffffff0000001900000000",
            INIT_07 => X"0000000a00000000000000000000000000000033000000000000000c00000000",
            INIT_08 => X"0000001600000000ffffffdfffffffffffffffe5ffffffff0000000600000000",
            INIT_09 => X"0000002400000000fffffff1ffffffff0000000b000000000000000500000000",
            INIT_0A => X"fffffff9ffffffff00000003000000000000000900000000ffffffeeffffffff",
            INIT_0B => X"ffffffe5ffffffffffffffaefffffffffffffff2ffffffff0000002700000000",
            INIT_0C => X"ffffffd5ffffffff0000001000000000fffffff8ffffffff0000000e00000000",
            INIT_0D => X"00000025000000000000002f000000000000001500000000ffffffeeffffffff",
            INIT_0E => X"0000000900000000000000070000000000000034000000000000003a00000000",
            INIT_0F => X"fffffffeffffffffffffffecffffffff00000027000000000000001100000000",
            INIT_10 => X"0000001e00000000ffffffcaffffffffffffffd7fffffffffffffff6ffffffff",
            INIT_11 => X"0000000e00000000ffffffebffffffff00000025000000000000000300000000",
            INIT_12 => X"0000003100000000ffffffe3ffffffff0000001900000000ffffffe1ffffffff",
            INIT_13 => X"ffffffe7ffffffffffffffe2ffffffffffffffd3ffffffff0000002e00000000",
            INIT_14 => X"ffffffa6fffffffffffffff9fffffffffffffff4ffffffff0000001f00000000",
            INIT_15 => X"00000007000000000000005800000000fffffff1fffffffffffffff7ffffffff",
            INIT_16 => X"fffffffeffffffff0000002300000000ffffffe4ffffffff0000003600000000",
            INIT_17 => X"0000000800000000ffffffc7ffffffff00000043000000000000002000000000",
            INIT_18 => X"fffffffcffffffffffffffedfffffffffffffff0ffffffffffffffe3ffffffff",
            INIT_19 => X"fffffff1ffffffffffffffc0ffffffff0000004400000000fffffffaffffffff",
            INIT_1A => X"0000000200000000ffffffceffffffff0000002a00000000ffffffd6ffffffff",
            INIT_1B => X"fffffffaffffffff0000002300000000fffffffdfffffffffffffffcffffffff",
            INIT_1C => X"ffffffbffffffffffffffff6ffffffff00000002000000000000000000000000",
            INIT_1D => X"ffffffc1ffffffff00000021000000000000000500000000fffffff4ffffffff",
            INIT_1E => X"ffffffeafffffffffffffffbffffffffffffffc4ffffffff0000002100000000",
            INIT_1F => X"fffffffaffffffffffffffebffffffff0000002b000000000000002100000000",
            INIT_20 => X"0000000a00000000ffffffbfffffffffffffffd5ffffffffffffffe0ffffffff",
            INIT_21 => X"ffffffdeffffffffffffffe3ffffffff00000025000000000000000c00000000",
            INIT_22 => X"0000000100000000ffffffffffffffff0000001b00000000ffffffe5ffffffff",
            INIT_23 => X"fffffffbffffffff00000017000000000000001b000000000000000a00000000",
            INIT_24 => X"ffffffd1ffffffffffffffedffffffff0000000200000000fffffffcffffffff",
            INIT_25 => X"ffffffe5ffffffff0000002700000000ffffffe5ffffffffffffffe7ffffffff",
            INIT_26 => X"00000000000000000000001100000000ffffffa2ffffffff0000000d00000000",
            INIT_27 => X"0000000d0000000000000011000000000000002d000000000000001e00000000",
            INIT_28 => X"0000000300000000ffffffe3ffffffffffffffd8fffffffffffffff8ffffffff",
            INIT_29 => X"fffffff1fffffffffffffff0ffffffff00000016000000000000001000000000",
            INIT_2A => X"ffffffb9ffffffffffffffffffffffff0000001c00000000fffffff9ffffffff",
            INIT_2B => X"000000170000000000000025000000000000001100000000fffffff7ffffffff",
            INIT_2C => X"ffffffeeffffffff00000019000000000000003e00000000ffffffd9ffffffff",
            INIT_2D => X"fffffff1ffffffff0000001c00000000fffffffcfffffffffffffff5ffffffff",
            INIT_2E => X"fffffff5ffffffff0000000100000000ffffffa7ffffffffffffffd8ffffffff",
            INIT_2F => X"0000001400000000fffffff3fffffffffffffff6fffffffffffffffaffffffff",
            INIT_30 => X"0000001200000000ffffffffffffffffffffffe6fffffffffffffff3ffffffff",
            INIT_31 => X"0000000200000000ffffffedffffffffffffffcdffffffff0000002000000000",
            INIT_32 => X"00000013000000000000002900000000fffffff5fffffffffffffff1ffffffff",
            INIT_33 => X"00000004000000000000002500000000fffffffeffffffff0000001700000000",
            INIT_34 => X"ffffffeafffffffffffffff0ffffffff0000000e000000000000000a00000000",
            INIT_35 => X"ffffffdfffffffff0000002100000000ffffffe7ffffffff0000000000000000",
            INIT_36 => X"ffffffddffffffff0000002300000000ffffffc2ffffffffffffffefffffffff",
            INIT_37 => X"fffffff8fffffffffffffff5ffffffffffffffddffffffffffffffc0ffffffff",
            INIT_38 => X"0000002c000000000000000e00000000ffffffe9ffffffffffffffeaffffffff",
            INIT_39 => X"0000000d00000000fffffff0ffffffffffffffbafffffffffffffff1ffffffff",
            INIT_3A => X"ffffffc9fffffffffffffffeffffffffffffffffffffffffffffffd6ffffffff",
            INIT_3B => X"fffffff6ffffffffffffffd4fffffffffffffffaffffffff0000000000000000",
            INIT_3C => X"ffffffb1fffffffffffffff9ffffffff0000000f000000000000001c00000000",
            INIT_3D => X"0000003f000000000000000c00000000fffffffbffffffffffffffecffffffff",
            INIT_3E => X"ffffffcffffffffffffffff1ffffffffffffffcaffffffff0000000b00000000",
            INIT_3F => X"0000001c00000000ffffffd0fffffffffffffff6ffffffff0000001000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000b00000000ffffffc7ffffffffffffffbeffffffffffffffd0ffffffff",
            INIT_41 => X"0000000000000000ffffffe9ffffffff00000017000000000000002600000000",
            INIT_42 => X"fffffff5ffffffff000000000000000000000028000000000000002b00000000",
            INIT_43 => X"0000000200000000fffffff5fffffffffffffffeffffffff0000002000000000",
            INIT_44 => X"ffffffb6ffffffff000000230000000000000023000000000000002200000000",
            INIT_45 => X"0000000e000000000000002e000000000000001200000000fffffff5ffffffff",
            INIT_46 => X"fffffffcffffffff0000001500000000ffffffc0ffffffff0000000600000000",
            INIT_47 => X"0000000f00000000ffffffaeffffffff00000013000000000000001400000000",
            INIT_48 => X"0000001100000000ffffffa3ffffffffffffffa9ffffffffffffffe6ffffffff",
            INIT_49 => X"ffffffdfffffffffffffffe8ffffffff0000002b000000000000001700000000",
            INIT_4A => X"000000050000000000000015000000000000003600000000ffffffffffffffff",
            INIT_4B => X"0000000100000000fffffff0ffffffffffffffe3ffffffff0000001c00000000",
            INIT_4C => X"ffffffb8ffffffff0000001e0000000000000020000000000000001a00000000",
            INIT_4D => X"ffffffcdffffffff0000005300000000ffffffe9ffffffffffffffebffffffff",
            INIT_4E => X"fffffff9ffffffff0000005100000000ffffffe3ffffffff0000002400000000",
            INIT_4F => X"0000003100000000ffffffa8ffffffff0000001f000000000000001100000000",
            INIT_50 => X"00000007000000000000000300000000ffffffdaffffffffffffffeeffffffff",
            INIT_51 => X"ffffffd9ffffffffffffffbfffffffff00000047000000000000003500000000",
            INIT_52 => X"fffffff4fffffffffffffffeffffffff00000027000000000000000e00000000",
            INIT_53 => X"0000000200000000ffffffd8ffffffff00000011000000000000002c00000000",
            INIT_54 => X"ffffffbdffffffff0000002d000000000000001600000000fffffff7ffffffff",
            INIT_55 => X"ffffffa6ffffffff0000004c000000000000000200000000ffffffc8ffffffff",
            INIT_56 => X"0000001f000000000000005700000000ffffff63ffffffff0000002000000000",
            INIT_57 => X"0000001200000000ffffffc4ffffffff0000001700000000ffffffddffffffff",
            INIT_58 => X"ffffffe7ffffffffffffffc0ffffffffffffffa4ffffffff0000000100000000",
            INIT_59 => X"ffffffd8ffffffffffffffb0ffffffff0000002d000000000000000900000000",
            INIT_5A => X"fffffff6ffffffff000000030000000000000026000000000000001700000000",
            INIT_5B => X"0000001b00000000ffffffe8ffffffffffffffffffffffff0000002800000000",
            INIT_5C => X"ffffffd6ffffffff000000110000000000000005000000000000000300000000",
            INIT_5D => X"ffffffabffffffff0000000d00000000fffffffcffffffffffffffdbffffffff",
            INIT_5E => X"fffffff9ffffffff0000002200000000fffffff5ffffffff0000001300000000",
            INIT_5F => X"fffffff6ffffffffffffffd9ffffffff0000000000000000ffffffedffffffff",
            INIT_60 => X"0000000200000000ffffffc3ffffffffffffffb9ffffffffffffffdcffffffff",
            INIT_61 => X"ffffffd0ffffffffffffffcfffffffff0000002b000000000000000500000000",
            INIT_62 => X"fffffff1fffffffffffffff0ffffffff0000002a000000000000001700000000",
            INIT_63 => X"0000000f000000000000000200000000fffffffbfffffffffffffff5ffffffff",
            INIT_64 => X"00000001000000000000001d0000000000000042000000000000000600000000",
            INIT_65 => X"ffffffb5fffffffffffffffffffffffffffffff5ffffffffffffffeeffffffff",
            INIT_66 => X"ffffffe7ffffffff0000002500000000ffffff8affffffff0000000700000000",
            INIT_67 => X"fffffff4fffffffffffffff8ffffffffffffffbaffffffffffffffd7ffffffff",
            INIT_68 => X"00000032000000000000000900000000fffffffcffffffffffffffe4ffffffff",
            INIT_69 => X"fffffff9fffffffffffffff6ffffffffffffffe9ffffffff0000002500000000",
            INIT_6A => X"fffffffcfffffffffffffff9ffffffff0000000300000000fffffffaffffffff",
            INIT_6B => X"ffffffe4ffffffff0000002800000000fffffff3ffffffffffffffebffffffff",
            INIT_6C => X"0000002c00000000ffffffe9ffffffff0000003a00000000ffffffc8ffffffff",
            INIT_6D => X"ffffffd3fffffffffffffff4fffffffffffffff3ffffffff0000000700000000",
            INIT_6E => X"fffffff0ffffffffffffffe2ffffffffffffff87ffffffffffffffe3ffffffff",
            INIT_6F => X"00000002000000000000000200000000fffffff4ffffffffffffffa4ffffffff",
            INIT_70 => X"0000000500000000ffffffeeffffffffffffffe5ffffffffffffffe6ffffffff",
            INIT_71 => X"ffffffecffffffff0000000000000000ffffffd6ffffffff0000001200000000",
            INIT_72 => X"ffffffc8ffffffff0000001400000000ffffffeeffffffffffffffeaffffffff",
            INIT_73 => X"ffffffc5ffffffff0000002300000000ffffffe5fffffffffffffff7ffffffff",
            INIT_74 => X"ffffffc7ffffffffffffffdeffffffff0000006300000000fffffff8ffffffff",
            INIT_75 => X"ffffffe4ffffffff00000047000000000000003a000000000000000d00000000",
            INIT_76 => X"fffffff3ffffffffffffffebffffffffffffffdcffffffff0000001700000000",
            INIT_77 => X"0000002000000000ffffffddffffffffffffffe3ffffffff0000001500000000",
            INIT_78 => X"0000003000000000ffffffeeffffffffffffffefffffffffffffffc5ffffffff",
            INIT_79 => X"ffffffdcffffffffffffffc1ffffffff0000002a000000000000003f00000000",
            INIT_7A => X"ffffffe1ffffffff0000002a000000000000003e000000000000002400000000",
            INIT_7B => X"0000000a0000000000000011000000000000001b000000000000001d00000000",
            INIT_7C => X"ffffffddffffffff00000015000000000000002100000000fffffff6ffffffff",
            INIT_7D => X"0000000f000000000000000a000000000000002200000000fffffff2ffffffff",
            INIT_7E => X"fffffff0ffffffff000000330000000000000007000000000000000400000000",
            INIT_7F => X"fffffffcffffffffffffffe3ffffffffffffffcdffffffff0000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE4;


    MEM_IWGHT_LAYER2_INSTANCE5 : if BRAM_NAME = "iwght_layer2_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000c00000000ffffffbdfffffffffffffff7ffffffffffffffddffffffff",
            INIT_01 => X"ffffffd6ffffffffffffffdfffffffff0000002900000000fffffffcffffffff",
            INIT_02 => X"0000000800000000000000240000000000000038000000000000001200000000",
            INIT_03 => X"00000002000000000000001d000000000000000e000000000000001200000000",
            INIT_04 => X"fffffff2ffffffff00000008000000000000000900000000fffffff5ffffffff",
            INIT_05 => X"ffffffe0ffffffff00000044000000000000002200000000ffffffeaffffffff",
            INIT_06 => X"00000000000000000000001800000000fffffff3ffffffff0000001200000000",
            INIT_07 => X"0000001b00000000ffffffe5ffffffffffffffcefffffffffffffff3ffffffff",
            INIT_08 => X"0000000c00000000fffffffbffffffffffffffffffffffffffffffe7ffffffff",
            INIT_09 => X"ffffffc9ffffffffffffffd1ffffffff00000036000000000000001600000000",
            INIT_0A => X"0000001000000000000000070000000000000023000000000000003100000000",
            INIT_0B => X"00000006000000000000001300000000fffffff5ffffffff0000001700000000",
            INIT_0C => X"ffffffdfffffffff000000080000000000000028000000000000000300000000",
            INIT_0D => X"ffffffefffffffff00000022000000000000004400000000fffffffeffffffff",
            INIT_0E => X"0000003700000000fffffffcfffffffffffffff0fffffffffffffff2ffffffff",
            INIT_0F => X"0000000900000000ffffffc2ffffffffffffffb4ffffffff0000000100000000",
            INIT_10 => X"0000000e00000000ffffffffffffffff0000000500000000ffffffc7ffffffff",
            INIT_11 => X"ffffffc9ffffffffffffffcdffffffff0000003a000000000000002000000000",
            INIT_12 => X"0000000e00000000000000190000000000000016000000000000002100000000",
            INIT_13 => X"ffffffe3ffffffffffffffdbffffffff00000003000000000000001d00000000",
            INIT_14 => X"ffffffcbffffffff0000000500000000fffffff7ffffffff0000000d00000000",
            INIT_15 => X"ffffffebffffffff0000000400000000ffffffebffffffffffffffe4ffffffff",
            INIT_16 => X"ffffffebffffffff000000380000000000000022000000000000001500000000",
            INIT_17 => X"0000001c00000000ffffffd8ffffffffffffffdbffffffffffffffe9ffffffff",
            INIT_18 => X"fffffffcffffffffffffffafffffffffffffffcdffffffffffffffdbffffffff",
            INIT_19 => X"ffffffd4ffffffffffffffcaffffffff00000025000000000000000900000000",
            INIT_1A => X"0000001c000000000000001a000000000000000f000000000000003900000000",
            INIT_1B => X"ffffffd0ffffffff0000000c00000000ffffffdafffffffffffffff7ffffffff",
            INIT_1C => X"fffffff7ffffffff0000000600000000ffffffe3fffffffffffffff0ffffffff",
            INIT_1D => X"ffffffd5ffffffff0000001000000000ffffffe5ffffffffffffffdcffffffff",
            INIT_1E => X"ffffffa1ffffffff0000002f00000000ffffffd3fffffffffffffff5ffffffff",
            INIT_1F => X"0000000500000000fffffffefffffffffffffffaffffffffffffffe8ffffffff",
            INIT_20 => X"0000004400000000ffffffd3fffffffffffffffeffffffffffffffd8ffffffff",
            INIT_21 => X"fffffff5ffffffffffffffdbffffffffffffffdaffffffff0000001800000000",
            INIT_22 => X"0000002200000000fffffff6ffffffff0000002800000000ffffffe9ffffffff",
            INIT_23 => X"fffffff4ffffffff00000059000000000000001700000000ffffffe6ffffffff",
            INIT_24 => X"ffffffebffffffffffffffb4ffffffffffffffeffffffffffffffff9ffffffff",
            INIT_25 => X"0000000e00000000fffffff5ffffffff0000000000000000fffffff7ffffffff",
            INIT_26 => X"0000001300000000ffffff9dffffffffffffff52ffffffffffffffdcffffffff",
            INIT_27 => X"ffffffd2ffffffff0000000200000000ffffffd3ffffffffffffffd6ffffffff",
            INIT_28 => X"ffffffd8fffffffffffffffeffffffffffffffdeffffffff0000000300000000",
            INIT_29 => X"ffffffe0ffffffff0000000300000000ffffffddfffffffffffffffbffffffff",
            INIT_2A => X"0000000e00000000ffffffffffffffff0000001500000000ffffffc1ffffffff",
            INIT_2B => X"0000000f000000000000001100000000fffffffbfffffffffffffff7ffffffff",
            INIT_2C => X"0000002500000000ffffffd8ffffffff00000045000000000000001c00000000",
            INIT_2D => X"ffffffffffffffff0000002f000000000000000900000000ffffffffffffffff",
            INIT_2E => X"0000001e00000000fffffff9ffffffffffffffc0ffffffff0000002500000000",
            INIT_2F => X"fffffffcffffffffffffffd8ffffffff00000033000000000000003400000000",
            INIT_30 => X"0000001900000000fffffff9ffffffffffffffd7ffffffffffffffeeffffffff",
            INIT_31 => X"fffffff3ffffffffffffffd2ffffffff00000007000000000000002500000000",
            INIT_32 => X"fffffff7ffffffff000000180000000000000005000000000000002400000000",
            INIT_33 => X"fffffffeffffffff0000001300000000fffffff2ffffffff0000001100000000",
            INIT_34 => X"0000000200000000ffffffe7ffffffff0000003500000000ffffffecffffffff",
            INIT_35 => X"00000015000000000000003700000000fffffff8ffffffffffffffe6ffffffff",
            INIT_36 => X"0000000f000000000000002900000000fffffff1fffffffffffffff7ffffffff",
            INIT_37 => X"ffffffebfffffffffffffffbffffffff0000000c000000000000001e00000000",
            INIT_38 => X"0000000f000000000000000c000000000000001500000000ffffffc1ffffffff",
            INIT_39 => X"fffffff2ffffffffffffffc7ffffffff0000001e000000000000000800000000",
            INIT_3A => X"0000003e000000000000000d0000000000000009000000000000003e00000000",
            INIT_3B => X"fffffff8ffffffff0000000d00000000fffffff0ffffffff0000000d00000000",
            INIT_3C => X"0000001d00000000ffffffd6ffffffffffffffffffffffff0000001a00000000",
            INIT_3D => X"ffffffd7ffffffffffffffedffffffff0000002300000000ffffffeaffffffff",
            INIT_3E => X"0000001b000000000000000900000000fffffff6ffffffffffffffe8ffffffff",
            INIT_3F => X"fffffffbffffffff0000000700000000fffffff2ffffffff0000000b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff3ffffffffffffffa9ffffffff0000002900000000ffffffd5ffffffff",
            INIT_41 => X"ffffffdbffffffffffffffe9fffffffffffffffcffffffff0000000200000000",
            INIT_42 => X"00000024000000000000000500000000ffffffeaffffffff0000002700000000",
            INIT_43 => X"0000000300000000fffffff2fffffffffffffff0ffffffff0000001500000000",
            INIT_44 => X"0000001100000000000000050000000000000000000000000000000e00000000",
            INIT_45 => X"0000000000000000fffffffdffffffff0000001800000000fffffffcffffffff",
            INIT_46 => X"fffffffeffffffff0000000f00000000ffffffddffffffff0000000b00000000",
            INIT_47 => X"0000000400000000fffffff0ffffffff00000014000000000000000600000000",
            INIT_48 => X"0000001200000000ffffffb6ffffffff0000000c00000000ffffffe5ffffffff",
            INIT_49 => X"ffffffd1ffffffffffffffdcfffffffffffffffeffffffff0000000900000000",
            INIT_4A => X"0000004d000000000000001a00000000fffffffaffffffff0000003500000000",
            INIT_4B => X"0000000a00000000ffffffe6ffffffffffffffecffffffff0000002800000000",
            INIT_4C => X"ffffffbfffffffff000000180000000000000006000000000000002200000000",
            INIT_4D => X"ffffffd0ffffffff0000001b000000000000001b00000000fffffff4ffffffff",
            INIT_4E => X"ffffffeaffffffff0000003a00000000ffffffebffffffff0000001300000000",
            INIT_4F => X"0000000700000000ffffffe9ffffffff0000001900000000ffffffe8ffffffff",
            INIT_50 => X"0000002500000000ffffffa4fffffffffffffff3ffffffffffffffe1ffffffff",
            INIT_51 => X"ffffffe8ffffffffffffffecfffffffffffffffdffffffff0000002200000000",
            INIT_52 => X"00000052000000000000000600000000ffffffe5ffffffff0000003a00000000",
            INIT_53 => X"ffffffe9ffffffff0000000d00000000ffffffdeffffffff0000000c00000000",
            INIT_54 => X"00000028000000000000001000000000ffffffddffffffff0000000c00000000",
            INIT_55 => X"ffffffc0ffffffff0000000000000000ffffffd4ffffffffffffffeeffffffff",
            INIT_56 => X"fffffffbffffffff0000001400000000fffffff4fffffffffffffff3ffffffff",
            INIT_57 => X"0000000400000000ffffffedffffffffffffffedffffffffffffffd2ffffffff",
            INIT_58 => X"0000004c00000000ffffff90ffffffff00000003000000000000000900000000",
            INIT_59 => X"ffffffecffffffff0000001500000000ffffffccffffffff0000000600000000",
            INIT_5A => X"0000001400000000ffffffe6fffffffffffffff8ffffffffffffffffffffffff",
            INIT_5B => X"000000040000000000000080000000000000001800000000ffffffe5ffffffff",
            INIT_5C => X"ffffffe4ffffffffffffffddffffffffffffffdffffffffffffffff3ffffffff",
            INIT_5D => X"fffffff6ffffffffffffffc1ffffffff0000001c000000000000001700000000",
            INIT_5E => X"0000003300000000ffffff88ffffffffffffff94ffffffffffffffdeffffffff",
            INIT_5F => X"ffffffa6ffffffffffffffe6ffffffff0000000300000000ffffffeeffffffff",
            INIT_60 => X"ffffffbbffffffff0000002600000000ffffffadfffffffffffffff6ffffffff",
            INIT_61 => X"ffffffddffffffff0000001d00000000ffffffe8ffffffffffffffd7ffffffff",
            INIT_62 => X"fffffffbffffffffffffffddffffffffffffffefffffffffffffffbfffffffff",
            INIT_63 => X"000000170000000000000038000000000000000500000000ffffffd9ffffffff",
            INIT_64 => X"ffffffe4fffffffffffffff5ffffffff0000002a000000000000000800000000",
            INIT_65 => X"00000022000000000000002200000000ffffffd7fffffffffffffffeffffffff",
            INIT_66 => X"00000028000000000000000800000000ffffffc9fffffffffffffff3ffffffff",
            INIT_67 => X"ffffffe5fffffffffffffff5ffffffff00000039000000000000000c00000000",
            INIT_68 => X"0000000200000000fffffffdffffffffffffffe0fffffffffffffff5ffffffff",
            INIT_69 => X"ffffffe7ffffffff0000000400000000fffffffdffffffff0000000200000000",
            INIT_6A => X"0000002600000000ffffffe3ffffffffffffffd6ffffffff0000002900000000",
            INIT_6B => X"0000000a000000000000004b00000000fffffffbffffffffffffffe4ffffffff",
            INIT_6C => X"ffffffd8ffffffffffffffd4ffffffff00000004000000000000000100000000",
            INIT_6D => X"000000020000000000000013000000000000000600000000ffffffeeffffffff",
            INIT_6E => X"0000003e00000000ffffffecffffffffffffffe3ffffffffffffffffffffffff",
            INIT_6F => X"fffffff3ffffffffffffffe9ffffffff00000024000000000000003200000000",
            INIT_70 => X"fffffff8ffffffffffffffe1ffffffffffffffd6ffffffffffffffe6ffffffff",
            INIT_71 => X"ffffffdefffffffffffffff5ffffffffffffffefffffffff0000001800000000",
            INIT_72 => X"0000004400000000ffffffe4ffffffffffffffd2ffffffff0000004100000000",
            INIT_73 => X"0000002c000000000000000e00000000ffffffecfffffffffffffffdffffffff",
            INIT_74 => X"ffffffe1ffffffff0000000f0000000000000000000000000000001200000000",
            INIT_75 => X"0000000f000000000000001e00000000fffffff2ffffffff0000000100000000",
            INIT_76 => X"00000035000000000000001000000000ffffffcbfffffffffffffff3ffffffff",
            INIT_77 => X"fffffffbffffffff000000060000000000000010000000000000002700000000",
            INIT_78 => X"0000000200000000ffffffcdffffffffffffffeeffffffffffffffe3ffffffff",
            INIT_79 => X"fffffff5ffffffffffffffffffffffffffffffedffffffff0000000b00000000",
            INIT_7A => X"00000055000000000000000800000000ffffffe7ffffffff0000001500000000",
            INIT_7B => X"00000010000000000000001e000000000000000100000000ffffffeeffffffff",
            INIT_7C => X"fffffff9ffffffff00000007000000000000000000000000ffffffeaffffffff",
            INIT_7D => X"00000012000000000000000c00000000fffffffafffffffffffffff1ffffffff",
            INIT_7E => X"0000001b000000000000001f000000000000000900000000ffffffffffffffff",
            INIT_7F => X"0000000d00000000fffffff0ffffffff00000033000000000000000700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE5;


    MEM_IWGHT_LAYER2_INSTANCE6 : if BRAM_NAME = "iwght_layer2_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000500000000ffffff91fffffffffffffff1ffffffffffffffe1ffffffff",
            INIT_01 => X"fffffffdfffffffffffffff7ffffffffffffffe9ffffffff0000000800000000",
            INIT_02 => X"00000049000000000000000000000000ffffffe5ffffffff0000000900000000",
            INIT_03 => X"0000000a00000000ffffffa0ffffffff0000000d00000000fffffff2ffffffff",
            INIT_04 => X"ffffffd6ffffffff0000002800000000fffffffafffffffffffffff9ffffffff",
            INIT_05 => X"fffffff1ffffffff0000000000000000ffffffb6ffffffff0000001000000000",
            INIT_06 => X"000000510000000000000035000000000000000200000000fffffffdffffffff",
            INIT_07 => X"0000000400000000ffffffd8ffffffff0000002800000000ffffffacffffffff",
            INIT_08 => X"0000000e00000000ffffff8cffffffffffffffd9ffffffffffffffecffffffff",
            INIT_09 => X"fffffff5ffffffff0000001d00000000ffffffe5ffffffff0000001100000000",
            INIT_0A => X"0000002d000000000000002e00000000ffffffccffffffff0000001200000000",
            INIT_0B => X"00000019000000000000000e000000000000001000000000ffffffe8ffffffff",
            INIT_0C => X"00000011000000000000000d00000000ffffffc9ffffffff0000001800000000",
            INIT_0D => X"ffffffc8fffffffffffffffbffffffffffffffedffffffff0000001900000000",
            INIT_0E => X"0000004d000000000000000c00000000ffffffdcfffffffffffffff8ffffffff",
            INIT_0F => X"fffffff2ffffffffffffffeeffffffff0000002400000000ffffffadffffffff",
            INIT_10 => X"0000004200000000ffffffa9ffffffff0000000c000000000000000100000000",
            INIT_11 => X"fffffffeffffffff0000003b00000000ffffffe2ffffffffffffffd2ffffffff",
            INIT_12 => X"0000001600000000ffffffdbffffffffffffffeeffffffffffffffeaffffffff",
            INIT_13 => X"ffffffeeffffffffffffffeeffffffff00000004000000000000001600000000",
            INIT_14 => X"0000002300000000fffffff4ffffffffffffffdbfffffffffffffff7ffffffff",
            INIT_15 => X"0000001c00000000ffffffb3ffffffffffffffe8fffffffffffffff2ffffffff",
            INIT_16 => X"ffffffe1ffffffffffffffccffffffffffffffdffffffffffffffff5ffffffff",
            INIT_17 => X"00000006000000000000001400000000ffffffd6ffffffff0000000000000000",
            INIT_18 => X"ffffffc8ffffffff0000000e00000000ffffffe4fffffffffffffffeffffffff",
            INIT_19 => X"0000002200000000fffffff1ffffffff0000000000000000fffffff1ffffffff",
            INIT_1A => X"0000000f000000000000001a00000000fffffff0ffffffff0000000400000000",
            INIT_1B => X"fffffffcfffffffffffffffbfffffffffffffff6ffffffff0000000d00000000",
            INIT_1C => X"ffffffe2ffffffff00000003000000000000000e00000000ffffffcbffffffff",
            INIT_1D => X"ffffffd2ffffffffffffffebffffffff0000000000000000ffffffdaffffffff",
            INIT_1E => X"fffffffaffffffffffffffe7ffffffffffffffe1ffffffff0000000600000000",
            INIT_1F => X"00000019000000000000001d00000000ffffffe9ffffffff0000000000000000",
            INIT_20 => X"00000017000000000000000d00000000ffffffedffffffff0000000c00000000",
            INIT_21 => X"0000003600000000ffffffe3ffffffffffffffefffffffff0000000d00000000",
            INIT_22 => X"0000000600000000ffffffeafffffffffffffff1ffffffff0000000500000000",
            INIT_23 => X"0000000000000000ffffffbeffffffffffffffe7fffffffffffffff1ffffffff",
            INIT_24 => X"ffffffd1ffffffff0000001600000000fffffff8fffffffffffffff0ffffffff",
            INIT_25 => X"ffffffd3fffffffffffffff1fffffffffffffff6ffffffff0000000200000000",
            INIT_26 => X"0000000700000000000000220000000000000017000000000000000400000000",
            INIT_27 => X"0000000000000000000000020000000000000011000000000000000200000000",
            INIT_28 => X"fffffffaffffffff00000000000000000000000200000000fffffffeffffffff",
            INIT_29 => X"0000002d000000000000000200000000fffffffbfffffffffffffffdffffffff",
            INIT_2A => X"0000000d00000000fffffff2fffffffffffffffdfffffffffffffffaffffffff",
            INIT_2B => X"fffffff7ffffffffffffffe9ffffffffffffffe8ffffffffffffffe2ffffffff",
            INIT_2C => X"fffffff4ffffffffffffffebfffffffffffffffafffffffffffffff0ffffffff",
            INIT_2D => X"ffffffc6ffffffffffffffd1fffffffffffffff1ffffffff0000001100000000",
            INIT_2E => X"00000009000000000000001500000000fffffff3ffffffff0000000400000000",
            INIT_2F => X"0000000000000000000000050000000000000001000000000000001400000000",
            INIT_30 => X"ffffffeeffffffff0000000300000000ffffffe0fffffffffffffffaffffffff",
            INIT_31 => X"00000016000000000000001000000000fffffffbffffffffffffffe9ffffffff",
            INIT_32 => X"ffffffc1ffffffffffffffc8fffffffffffffffbffffffff0000000d00000000",
            INIT_33 => X"ffffffefffffffff0000001100000000ffffffebfffffffffffffffcffffffff",
            INIT_34 => X"ffffffcdfffffffffffffffbffffffff0000000100000000fffffffbffffffff",
            INIT_35 => X"ffffffeeffffffffffffffebffffffffffffffeefffffffffffffffcffffffff",
            INIT_36 => X"000000040000000000000007000000000000000400000000ffffffefffffffff",
            INIT_37 => X"ffffffeeffffffff000000070000000000000008000000000000000100000000",
            INIT_38 => X"0000000a000000000000001700000000ffffffe3ffffffff0000000600000000",
            INIT_39 => X"00000001000000000000000f00000000fffffff7fffffffffffffff3ffffffff",
            INIT_3A => X"ffffffd9ffffffffffffffc0fffffffffffffffcffffffffffffffd9ffffffff",
            INIT_3B => X"ffffffffffffffff0000002a00000000ffffffe9fffffffffffffffaffffffff",
            INIT_3C => X"ffffffdaffffffffffffffcaffffffffffffffeaffffffff0000001000000000",
            INIT_3D => X"ffffffeafffffffffffffff7ffffffff0000001000000000fffffff0ffffffff",
            INIT_3E => X"0000001200000000ffffffd9ffffffffffffffd7ffffffff0000000800000000",
            INIT_3F => X"fffffffaffffffff00000008000000000000000f000000000000002e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000008000000000000002100000000ffffffe2ffffffff0000000000000000",
            INIT_41 => X"00000016000000000000000700000000fffffffcffffffffffffffedffffffff",
            INIT_42 => X"ffffffdeffffffffffffffebfffffffffffffffdfffffffffffffff9ffffffff",
            INIT_43 => X"ffffffe6ffffffff000000270000000000000002000000000000001300000000",
            INIT_44 => X"ffffffdbfffffffffffffff6fffffffffffffff9fffffffffffffffcffffffff",
            INIT_45 => X"fffffff2ffffffffffffffe7ffffffff0000000900000000fffffffcffffffff",
            INIT_46 => X"fffffffdffffffffffffffffffffffffffffffffffffffffffffffecffffffff",
            INIT_47 => X"ffffffffffffffff0000000900000000ffffffe5ffffffff0000000000000000",
            INIT_48 => X"ffffffecffffffff000000150000000000000003000000000000000f00000000",
            INIT_49 => X"0000002a00000000fffffff8fffffffffffffffcffffffffffffffe5ffffffff",
            INIT_4A => X"0000002200000000ffffffc4ffffffffffffffffffffffff0000001100000000",
            INIT_4B => X"ffffffefffffffffffffffeefffffffffffffffafffffffffffffffaffffffff",
            INIT_4C => X"ffffffffffffffffffffffecfffffffffffffff9ffffffff0000000500000000",
            INIT_4D => X"0000002100000000ffffffdbffffffff0000001600000000ffffffe9ffffffff",
            INIT_4E => X"0000001800000000ffffffcbffffffff00000018000000000000001a00000000",
            INIT_4F => X"ffffffdbffffffff0000001400000000ffffffecffffffff0000001900000000",
            INIT_50 => X"ffffffe7ffffffff000000290000000000000016000000000000000000000000",
            INIT_51 => X"00000019000000000000000e00000000ffffffffffffffffffffffd9ffffffff",
            INIT_52 => X"0000000e000000000000000e0000000000000009000000000000000000000000",
            INIT_53 => X"fffffffffffffffffffffff9fffffffffffffffcfffffffffffffff2ffffffff",
            INIT_54 => X"ffffffffffffffffffffffe1ffffffffffffffbfffffffffffffffeaffffffff",
            INIT_55 => X"ffffffd5ffffffff00000000000000000000000400000000fffffff6ffffffff",
            INIT_56 => X"0000002500000000fffffff5ffffffff00000007000000000000001a00000000",
            INIT_57 => X"0000000a00000000fffffffaffffffff00000002000000000000001700000000",
            INIT_58 => X"00000012000000000000000000000000ffffffeffffffffffffffff1ffffffff",
            INIT_59 => X"0000001e00000000fffffff9ffffffff0000001800000000fffffff3ffffffff",
            INIT_5A => X"fffffff4ffffffff00000021000000000000000e00000000ffffffe7ffffffff",
            INIT_5B => X"0000000d00000000fffffff2ffffffff00000011000000000000000b00000000",
            INIT_5C => X"fffffff1ffffffff0000001f00000000ffffffe1fffffffffffffffaffffffff",
            INIT_5D => X"ffffffddffffffff0000000f000000000000001a00000000fffffff9ffffffff",
            INIT_5E => X"00000028000000000000001c0000000000000011000000000000000f00000000",
            INIT_5F => X"0000001e00000000fffffff5ffffffff00000001000000000000000f00000000",
            INIT_60 => X"0000001b000000000000002400000000fffffff7ffffffff0000000800000000",
            INIT_61 => X"fffffffaffffffff0000001b00000000fffffff9fffffffffffffff4ffffffff",
            INIT_62 => X"ffffffe5ffffffff0000000c00000000ffffffeeffffffff0000001200000000",
            INIT_63 => X"fffffff1ffffffff00000004000000000000000300000000fffffff9ffffffff",
            INIT_64 => X"fffffff3fffffffffffffffbfffffffffffffff0ffffffffffffffecffffffff",
            INIT_65 => X"ffffffe3fffffffffffffff8fffffffffffffff9ffffffffffffffdbffffffff",
            INIT_66 => X"0000000900000000000000150000000000000016000000000000002800000000",
            INIT_67 => X"fffffff3fffffffffffffff5fffffffffffffffefffffffffffffffdffffffff",
            INIT_68 => X"0000002e0000000000000040000000000000000200000000fffffff5ffffffff",
            INIT_69 => X"00000005000000000000000800000000ffffffd9ffffffffffffffedffffffff",
            INIT_6A => X"0000000500000000ffffffe2ffffffffffffffeeffffffffffffffdcffffffff",
            INIT_6B => X"0000001b0000000000000018000000000000000900000000fffffff0ffffffff",
            INIT_6C => X"fffffff3ffffffff0000000300000000fffffff4ffffffff0000001000000000",
            INIT_6D => X"0000002a00000000ffffffedffffffff00000002000000000000000d00000000",
            INIT_6E => X"0000000600000000fffffff1ffffffff00000011000000000000002a00000000",
            INIT_6F => X"0000000000000000ffffffe4fffffffffffffff5ffffffff0000001600000000",
            INIT_70 => X"0000000d000000000000003400000000fffffff9ffffffffffffffeaffffffff",
            INIT_71 => X"00000003000000000000000200000000fffffff5ffffffffffffffe9ffffffff",
            INIT_72 => X"0000001c00000000fffffffdffffffffffffffe2ffffffffffffffe6ffffffff",
            INIT_73 => X"00000009000000000000000f00000000ffffffeffffffffffffffff7ffffffff",
            INIT_74 => X"0000000d000000000000000100000000ffffffe9ffffffff0000000c00000000",
            INIT_75 => X"0000000200000000ffffffe3ffffffff0000000300000000fffffff8ffffffff",
            INIT_76 => X"0000000800000000fffffffaffffffffffffffd4fffffffffffffff7ffffffff",
            INIT_77 => X"0000002600000000fffffffefffffffffffffffdfffffffffffffffaffffffff",
            INIT_78 => X"ffffffebffffffff000000160000000000000026000000000000000d00000000",
            INIT_79 => X"0000000400000000fffffffcffffffff0000000300000000ffffffdaffffffff",
            INIT_7A => X"0000000b00000000ffffffe7ffffffff0000000d00000000fffffff1ffffffff",
            INIT_7B => X"fffffffefffffffffffffff0ffffffff00000013000000000000000700000000",
            INIT_7C => X"fffffff8ffffffff0000000e00000000ffffffd5ffffffff0000000500000000",
            INIT_7D => X"0000002800000000ffffffe1ffffffff00000007000000000000000900000000",
            INIT_7E => X"00000006000000000000000200000000ffffff9cffffffff0000000b00000000",
            INIT_7F => X"fffffff4ffffffff0000000b00000000ffffffcdffffffffffffffdbffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE6;


    MEM_IWGHT_LAYER2_INSTANCE7 : if BRAM_NAME = "iwght_layer2_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffedfffffffffffffffeffffffff0000000a000000000000001800000000",
            INIT_01 => X"0000001d000000000000000d000000000000000e00000000ffffffebffffffff",
            INIT_02 => X"ffffffecffffffffffffffd3ffffffff0000000d000000000000001500000000",
            INIT_03 => X"0000001500000000ffffffd7ffffffff0000001e000000000000000800000000",
            INIT_04 => X"fffffffeffffffff0000000c00000000fffffff7ffffffffffffffffffffffff",
            INIT_05 => X"0000002400000000ffffffe2ffffffff0000001f000000000000000f00000000",
            INIT_06 => X"0000001a00000000ffffffe1ffffffffffffffdfffffffff0000001100000000",
            INIT_07 => X"fffffff4ffffffff0000000700000000ffffffbcffffffff0000002a00000000",
            INIT_08 => X"ffffffefffffffff0000001b000000000000000b000000000000000900000000",
            INIT_09 => X"00000015000000000000000a000000000000000100000000ffffffc4ffffffff",
            INIT_0A => X"0000000e000000000000000a0000000000000015000000000000000700000000",
            INIT_0B => X"0000000400000000ffffffdefffffffffffffff4fffffffffffffff6ffffffff",
            INIT_0C => X"0000001b000000000000000a00000000ffffffd6ffffffff0000001800000000",
            INIT_0D => X"fffffff4fffffffffffffffaffffffff00000013000000000000000f00000000",
            INIT_0E => X"0000003500000000ffffffedffffffffffffffffffffffff0000001500000000",
            INIT_0F => X"0000001000000000fffffff9ffffffffffffffd5ffffffff0000000b00000000",
            INIT_10 => X"fffffff9ffffffff0000001b00000000fffffff7ffffffff0000000000000000",
            INIT_11 => X"fffffff8ffffffff0000001b000000000000001700000000ffffffdeffffffff",
            INIT_12 => X"0000001e00000000000000280000000000000009000000000000001b00000000",
            INIT_13 => X"0000000300000000ffffffe0ffffffff00000006000000000000001a00000000",
            INIT_14 => X"fffffff8ffffffff0000002100000000ffffffc2ffffffffffffffebffffffff",
            INIT_15 => X"ffffffeaffffffff00000015000000000000000c00000000fffffff7ffffffff",
            INIT_16 => X"00000035000000000000001200000000ffffffcfffffffff0000002d00000000",
            INIT_17 => X"fffffff0ffffffffffffffd8ffffffffffffffcdffffffff0000001100000000",
            INIT_18 => X"0000000a000000000000003a000000000000001d000000000000000b00000000",
            INIT_19 => X"fffffffdffffffff000000170000000000000004000000000000000c00000000",
            INIT_1A => X"00000016000000000000000800000000fffffff0fffffffffffffffdffffffff",
            INIT_1B => X"fffffffdffffffff0000000d000000000000002600000000ffffffdeffffffff",
            INIT_1C => X"fffffffcffffffff00000015000000000000000900000000ffffffceffffffff",
            INIT_1D => X"ffffffe4ffffffff0000001d000000000000000700000000ffffffd5ffffffff",
            INIT_1E => X"00000010000000000000000d00000000ffffffa7ffffffffffffffffffffffff",
            INIT_1F => X"fffffffaffffffffffffffe1ffffffffffffffffffffffff0000001100000000",
            INIT_20 => X"0000002d000000000000005b0000000000000026000000000000001300000000",
            INIT_21 => X"00000011000000000000000300000000ffffffbaffffffff0000000300000000",
            INIT_22 => X"ffffffe8ffffffffffffffe2ffffffff0000000300000000ffffffefffffffff",
            INIT_23 => X"000000050000000000000014000000000000000500000000fffffff0ffffffff",
            INIT_24 => X"ffffffecfffffffffffffff3fffffffffffffffcfffffffffffffff7ffffffff",
            INIT_25 => X"0000000b00000000fffffff3fffffffffffffffdffffffffffffffecffffffff",
            INIT_26 => X"0000002500000000fffffff5ffffffffffffffb7ffffffff0000001a00000000",
            INIT_27 => X"fffffff5ffffffffffffffe9ffffffffffffffdcffffffff0000002700000000",
            INIT_28 => X"0000002a000000000000004f000000000000001c000000000000000100000000",
            INIT_29 => X"0000000000000000fffffffcffffffffffffffe4fffffffffffffff3ffffffff",
            INIT_2A => X"0000001f00000000ffffffceffffffff0000000600000000ffffffeeffffffff",
            INIT_2B => X"0000001800000000fffffff1ffffffffffffffefffffffff0000000c00000000",
            INIT_2C => X"fffffff3ffffffff0000001300000000ffffffe4ffffffff0000001000000000",
            INIT_2D => X"0000001100000000fffffff7ffffffff0000000a000000000000001100000000",
            INIT_2E => X"0000001900000000fffffff5ffffffffffffffcbffffffff0000001c00000000",
            INIT_2F => X"ffffffddffffffffffffffe7ffffffffffffffd8ffffffff0000001500000000",
            INIT_30 => X"fffffffcffffffff0000000d000000000000000700000000fffffffdffffffff",
            INIT_31 => X"fffffff3ffffffffffffffffffffffff0000000e00000000ffffffedffffffff",
            INIT_32 => X"0000002b00000000ffffffe7ffffffff0000001300000000ffffffe6ffffffff",
            INIT_33 => X"0000000300000000ffffffd6ffffffff0000001d000000000000000a00000000",
            INIT_34 => X"00000000000000000000001700000000ffffffa4ffffffff0000000900000000",
            INIT_35 => X"0000001c00000000ffffffd6ffffffff0000000c000000000000000000000000",
            INIT_36 => X"0000000e000000000000000700000000ffffffedffffffffffffffebffffffff",
            INIT_37 => X"00000021000000000000001900000000fffffff0ffffffffffffffebffffffff",
            INIT_38 => X"ffffffd5ffffffff000000060000000000000005000000000000001200000000",
            INIT_39 => X"0000000d0000000000000009000000000000000000000000ffffffbaffffffff",
            INIT_3A => X"fffffff6ffffffffffffffeafffffffffffffffcfffffffffffffff4ffffffff",
            INIT_3B => X"0000000e00000000ffffffedffffffff00000012000000000000000100000000",
            INIT_3C => X"0000000500000000ffffffefffffffff0000000800000000fffffff9ffffffff",
            INIT_3D => X"0000003c00000000ffffffe0ffffffff00000021000000000000001b00000000",
            INIT_3E => X"0000002c00000000ffffffd4ffffffffffffffcbffffffff0000000c00000000",
            INIT_3F => X"ffffffefffffffff0000002300000000fffffff2fffffffffffffff9ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000ffffffecffffffffffffffd3ffffffff0000000500000000",
            INIT_41 => X"00000011000000000000000c00000000ffffffeaffffffffffffffd6ffffffff",
            INIT_42 => X"0000001000000000ffffffeffffffffffffffffefffffffffffffff4ffffffff",
            INIT_43 => X"0000000900000000ffffffd7fffffffffffffffdffffffff0000000000000000",
            INIT_44 => X"0000000300000000fffffffeffffffffffffffedffffffff0000000a00000000",
            INIT_45 => X"0000003700000000ffffffffffffffff00000009000000000000001600000000",
            INIT_46 => X"0000002300000000ffffffc3ffffffffffffffefffffffff0000000f00000000",
            INIT_47 => X"ffffffebffffffff0000000100000000ffffffe2ffffffff0000001800000000",
            INIT_48 => X"fffffffaffffffff0000000500000000fffffff9ffffffff0000000f00000000",
            INIT_49 => X"00000001000000000000002b000000000000001500000000ffffffbfffffffff",
            INIT_4A => X"0000000f00000000ffffffffffffffff0000000900000000ffffffd6ffffffff",
            INIT_4B => X"0000000000000000ffffffe3fffffffffffffffdffffffff0000000f00000000",
            INIT_4C => X"fffffff2fffffffffffffff9fffffffffffffff5ffffffffffffffe9ffffffff",
            INIT_4D => X"ffffffebffffffff0000002900000000ffffffeeffffffffffffffe0ffffffff",
            INIT_4E => X"00000023000000000000002300000000fffffff2ffffffff0000001000000000",
            INIT_4F => X"0000000000000000000000060000000000000006000000000000001800000000",
            INIT_50 => X"ffffffedffffffff00000054000000000000000800000000fffffff9ffffffff",
            INIT_51 => X"ffffffe9fffffffffffffff9ffffffffffffffe4fffffffffffffff4ffffffff",
            INIT_52 => X"00000011000000000000000000000000ffffffd8ffffffff0000000a00000000",
            INIT_53 => X"0000000800000000fffffff7ffffffff0000000d000000000000002400000000",
            INIT_54 => X"ffffffd5fffffffffffffffeffffffff0000002800000000ffffffd0ffffffff",
            INIT_55 => X"ffffffe5ffffffff0000001d00000000fffffffeffffffffffffffdaffffffff",
            INIT_56 => X"00000006000000000000003100000000fffffff3ffffffff0000001b00000000",
            INIT_57 => X"0000000000000000ffffffeaffffffff00000014000000000000001e00000000",
            INIT_58 => X"0000001a00000000000000600000000000000019000000000000001400000000",
            INIT_59 => X"fffffff8ffffffffffffffeeffffffffffffffdefffffffffffffffaffffffff",
            INIT_5A => X"ffffffefffffffffffffffe7ffffffff0000001c000000000000000000000000",
            INIT_5B => X"fffffff5ffffffff0000002a000000000000001a00000000fffffff5ffffffff",
            INIT_5C => X"ffffffedffffffff0000000d000000000000000000000000ffffffe5ffffffff",
            INIT_5D => X"fffffff9ffffffff0000000300000000fffffff9ffffffffffffffebffffffff",
            INIT_5E => X"00000000000000000000003600000000fffffffeffffffff0000002500000000",
            INIT_5F => X"ffffffbbffffffffffffffe6ffffffffffffffe8ffffffff0000001200000000",
            INIT_60 => X"0000000700000000000000410000000000000023000000000000000f00000000",
            INIT_61 => X"fffffff3ffffffff0000000800000000ffffffe3fffffffffffffff6ffffffff",
            INIT_62 => X"0000001600000000ffffffd3ffffffff0000001f00000000fffffff6ffffffff",
            INIT_63 => X"00000001000000000000000600000000fffffffeffffffff0000000100000000",
            INIT_64 => X"fffffff0ffffffff0000000d00000000fffffff1ffffffff0000001d00000000",
            INIT_65 => X"0000001600000000ffffffc4ffffffff00000013000000000000001000000000",
            INIT_66 => X"00000012000000000000002800000000ffffff7cffffffff0000003500000000",
            INIT_67 => X"ffffffddffffffffffffffecffffffffffffffefffffffff0000001200000000",
            INIT_68 => X"0000001f0000000000000036000000000000001d000000000000001100000000",
            INIT_69 => X"ffffffe3ffffffff00000016000000000000001c00000000ffffffdfffffffff",
            INIT_6A => X"fffffffdffffffffffffffe9ffffffff0000000e00000000fffffff7ffffffff",
            INIT_6B => X"00000028000000000000000a0000000000000026000000000000000a00000000",
            INIT_6C => X"ffffffe5ffffffff0000003000000000ffffffbaffffffff0000000200000000",
            INIT_6D => X"0000002600000000ffffffc7fffffffffffffff7ffffffff0000000b00000000",
            INIT_6E => X"0000001600000000000000180000000000000020000000000000002200000000",
            INIT_6F => X"00000004000000000000000100000000ffffffecffffffffffffffeaffffffff",
            INIT_70 => X"ffffffe9fffffffffffffff7ffffffffffffffffffffffff0000001d00000000",
            INIT_71 => X"00000018000000000000000f000000000000001800000000ffffffb2ffffffff",
            INIT_72 => X"0000000500000000ffffffe4ffffffff0000000500000000fffffff1ffffffff",
            INIT_73 => X"0000000700000000ffffffe9ffffffff0000000a000000000000001600000000",
            INIT_74 => X"ffffffe6ffffffff0000000600000000fffffff2fffffffffffffffbffffffff",
            INIT_75 => X"0000003100000000ffffffd0ffffffff00000037000000000000002000000000",
            INIT_76 => X"0000001300000000ffffffeaffffffffffffffc3fffffffffffffffeffffffff",
            INIT_77 => X"fffffffcffffffff000000130000000000000004000000000000001700000000",
            INIT_78 => X"fffffff0ffffffffffffffd3ffffffffffffffe0ffffffff0000001100000000",
            INIT_79 => X"000000100000000000000002000000000000000100000000ffffffc4ffffffff",
            INIT_7A => X"0000000100000000ffffffeaffffffff0000001e000000000000000f00000000",
            INIT_7B => X"fffffffcfffffffffffffff9fffffffffffffffbffffffff0000001400000000",
            INIT_7C => X"fffffff3ffffffff0000000400000000ffffffe1ffffffff0000000c00000000",
            INIT_7D => X"00000029000000000000000f0000000000000024000000000000000900000000",
            INIT_7E => X"0000003900000000ffffffebffffffffffffffe0fffffffffffffff2ffffffff",
            INIT_7F => X"ffffffedffffffff00000000000000000000002c000000000000001700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE7;


    MEM_IWGHT_LAYER2_INSTANCE8 : if BRAM_NAME = "iwght_layer2_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002b00000000fffffff2ffffffffffffffccffffffff0000001200000000",
            INIT_01 => X"fffffff6fffffffffffffff6ffffffff0000000300000000ffffffc3ffffffff",
            INIT_02 => X"ffffffdcfffffffffffffffdffffffff0000001600000000ffffffd9ffffffff",
            INIT_03 => X"fffffff2fffffffffffffff7ffffffff00000000000000000000000c00000000",
            INIT_04 => X"ffffffbfffffffffffffffecffffffff0000001700000000fffffffcffffffff",
            INIT_05 => X"0000000d000000000000004800000000ffffffebfffffffffffffff9ffffffff",
            INIT_06 => X"0000002d000000000000001a00000000ffffffe7ffffffff0000000000000000",
            INIT_07 => X"fffffff3ffffffff0000000e0000000000000031000000000000001e00000000",
            INIT_08 => X"0000002f000000000000001300000000ffffffd4ffffffff0000000000000000",
            INIT_09 => X"ffffffe9ffffffffffffffe0ffffffffffffffedffffffffffffffe8ffffffff",
            INIT_0A => X"ffffffefffffffff0000001300000000fffffff4ffffffff0000000800000000",
            INIT_0B => X"0000000c00000000ffffffe3ffffffff0000000f000000000000000900000000",
            INIT_0C => X"ffffffdafffffffffffffff5fffffffffffffff5ffffffffffffffe7ffffffff",
            INIT_0D => X"00000006000000000000001e00000000fffffff1fffffffffffffff2ffffffff",
            INIT_0E => X"0000000d000000000000002c0000000000000005000000000000003100000000",
            INIT_0F => X"fffffffbfffffffffffffffefffffffffffffff8ffffffff0000000b00000000",
            INIT_10 => X"0000000b000000000000003000000000fffffff9fffffffffffffffdffffffff",
            INIT_11 => X"0000001200000000fffffffeffffffffffffffd4fffffffffffffffbffffffff",
            INIT_12 => X"0000000500000000ffffffd4ffffffff00000012000000000000000100000000",
            INIT_13 => X"0000000000000000fffffffafffffffffffffffdfffffffffffffff1ffffffff",
            INIT_14 => X"ffffffd5fffffffffffffff1ffffffffffffffcbffffffff0000000e00000000",
            INIT_15 => X"fffffffbffffffff0000000800000000ffffffebffffffffffffffe0ffffffff",
            INIT_16 => X"00000010000000000000004700000000ffffffa6ffffffff0000001a00000000",
            INIT_17 => X"0000000500000000ffffffeaffffffff0000002d00000000ffffffe6ffffffff",
            INIT_18 => X"0000001b000000000000001a0000000000000004000000000000000700000000",
            INIT_19 => X"ffffffeffffffffffffffff8fffffffffffffff6ffffffffffffffe2ffffffff",
            INIT_1A => X"0000001c00000000ffffffd1ffffffff0000000200000000ffffffe7ffffffff",
            INIT_1B => X"00000005000000000000000c00000000fffffffeffffffff0000000b00000000",
            INIT_1C => X"ffffffeeffffffff0000000c00000000ffffffe2fffffffffffffff0ffffffff",
            INIT_1D => X"fffffffefffffffffffffffffffffffffffffff3fffffffffffffffdffffffff",
            INIT_1E => X"000000140000000000000026000000000000001d000000000000001d00000000",
            INIT_1F => X"fffffff7ffffffffffffffeeffffffff0000001100000000fffffff8ffffffff",
            INIT_20 => X"0000000b00000000fffffff6ffffffff0000000100000000fffffffaffffffff",
            INIT_21 => X"00000006000000000000000c000000000000000100000000ffffffcbffffffff",
            INIT_22 => X"0000001700000000ffffffefffffffff0000000400000000ffffffceffffffff",
            INIT_23 => X"0000001100000000ffffffdfffffffff0000000b000000000000001800000000",
            INIT_24 => X"ffffffc0ffffffff0000001300000000ffffffc0ffffffff0000001d00000000",
            INIT_25 => X"0000002400000000ffffffc4ffffffffffffffdcffffffff0000000700000000",
            INIT_26 => X"00000019000000000000001300000000ffffffd3ffffffff0000001700000000",
            INIT_27 => X"fffffffaffffffff0000000900000000ffffffebffffffffffffffdfffffffff",
            INIT_28 => X"ffffffe8ffffffffffffffeaffffffff00000002000000000000000600000000",
            INIT_29 => X"0000000d000000000000000a000000000000000600000000ffffffd0ffffffff",
            INIT_2A => X"fffffff2ffffffffffffffc3fffffffffffffff9fffffffffffffff2ffffffff",
            INIT_2B => X"0000001600000000ffffffafffffffff00000000000000000000000700000000",
            INIT_2C => X"00000011000000000000002200000000ffffffe3ffffffff0000001e00000000",
            INIT_2D => X"0000000000000000000000020000000000000014000000000000001900000000",
            INIT_2E => X"00000016000000000000001200000000ffffffcbffffffff0000000400000000",
            INIT_2F => X"fffffffeffffffff000000180000000000000024000000000000001500000000",
            INIT_30 => X"fffffff6ffffffffffffffe4fffffffffffffffdfffffffffffffff7ffffffff",
            INIT_31 => X"000000030000000000000012000000000000000600000000fffffffdffffffff",
            INIT_32 => X"fffffffaffffffffffffffd7ffffffff0000001800000000fffffff3ffffffff",
            INIT_33 => X"0000000800000000ffffffd4ffffffff00000008000000000000000800000000",
            INIT_34 => X"ffffffbeffffffffffffffffffffffffffffffd9ffffffff0000001d00000000",
            INIT_35 => X"0000000e0000000000000009000000000000000d000000000000000500000000",
            INIT_36 => X"000000180000000000000001000000000000002d00000000fffffffeffffffff",
            INIT_37 => X"fffffffdffffffff00000011000000000000000a00000000fffffff6ffffffff",
            INIT_38 => X"fffffffeffffffffffffffc3ffffffffffffffd5ffffffff0000000000000000",
            INIT_39 => X"fffffffcffffffff00000009000000000000000800000000ffffffc0ffffffff",
            INIT_3A => X"fffffffdfffffffffffffff2ffffffff0000001b00000000ffffffdfffffffff",
            INIT_3B => X"0000001400000000fffffff6fffffffffffffff9ffffffff0000001500000000",
            INIT_3C => X"ffffffcdfffffffffffffff3ffffffffffffffeeffffffff0000000d00000000",
            INIT_3D => X"000000050000000000000020000000000000000600000000fffffff1ffffffff",
            INIT_3E => X"0000002400000000ffffffe7ffffffffffffffe2ffffffff0000000e00000000",
            INIT_3F => X"0000000c0000000000000001000000000000000100000000fffffff9ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000007000000000000000800000000ffffffe2fffffffffffffff2ffffffff",
            INIT_41 => X"00000010000000000000000a000000000000001800000000ffffffd5ffffffff",
            INIT_42 => X"ffffffc5fffffffffffffffcffffffff0000002300000000ffffffe5ffffffff",
            INIT_43 => X"fffffff5ffffffffffffffd3ffffffff00000002000000000000001700000000",
            INIT_44 => X"ffffffe2ffffffffffffffe9ffffffff00000003000000000000000000000000",
            INIT_45 => X"fffffffeffffffff0000000b000000000000000a000000000000000100000000",
            INIT_46 => X"ffffffeeffffffff00000012000000000000001f00000000fffffffdffffffff",
            INIT_47 => X"0000000b00000000ffffffeaffffffff00000018000000000000000100000000",
            INIT_48 => X"ffffffdaffffffff0000002500000000ffffffd6ffffffffffffffffffffffff",
            INIT_49 => X"0000000f000000000000001a00000000ffffffefffffffff0000000500000000",
            INIT_4A => X"ffffffafffffffffffffffe1ffffffff0000000e00000000fffffff7ffffffff",
            INIT_4B => X"0000000300000000fffffff1ffffffff0000000d000000000000000900000000",
            INIT_4C => X"ffffffedffffffff00000002000000000000000000000000fffffffeffffffff",
            INIT_4D => X"000000000000000000000011000000000000001900000000ffffffecffffffff",
            INIT_4E => X"ffffffe5ffffffff0000001700000000ffffffc2ffffffff0000002a00000000",
            INIT_4F => X"ffffffeefffffffffffffffaffffffff0000000700000000fffffffcffffffff",
            INIT_50 => X"fffffffeffffffff0000001b00000000ffffffe6ffffffff0000000100000000",
            INIT_51 => X"fffffffeffffffff0000001d00000000fffffff9ffffffffffffffebffffffff",
            INIT_52 => X"ffffffc8ffffffffffffffeaffffffff0000001b00000000ffffffe1ffffffff",
            INIT_53 => X"0000000d00000000fffffff9ffffffff00000003000000000000001000000000",
            INIT_54 => X"ffffffe6ffffffff0000000e00000000ffffffc2ffffffff0000000900000000",
            INIT_55 => X"0000000100000000ffffffe8ffffffffffffffe8ffffffff0000000100000000",
            INIT_56 => X"0000001e000000000000001000000000fffffffbffffffff0000000400000000",
            INIT_57 => X"ffffffefffffffff0000000300000000fffffff7fffffffffffffffcffffffff",
            INIT_58 => X"0000000000000000fffffff1ffffffffffffffe4ffffffff0000000300000000",
            INIT_59 => X"fffffffdffffffff0000001e000000000000001d00000000fffffff0ffffffff",
            INIT_5A => X"0000000900000000ffffffc1ffffffff0000002200000000ffffffecffffffff",
            INIT_5B => X"0000002100000000fffffff4ffffffff00000000000000000000000e00000000",
            INIT_5C => X"ffffffceffffffffffffffecffffffffffffffb3ffffffff0000001900000000",
            INIT_5D => X"0000002000000000000000010000000000000027000000000000001a00000000",
            INIT_5E => X"0000001e00000000ffffffe7ffffffffffffffd2fffffffffffffffaffffffff",
            INIT_5F => X"ffffffebffffffff0000000800000000ffffffecffffffff0000000700000000",
            INIT_60 => X"ffffffd8ffffffffffffffd6ffffffffffffffd3ffffffff0000000700000000",
            INIT_61 => X"fffffff9ffffffff0000000c000000000000000900000000fffffffaffffffff",
            INIT_62 => X"0000000200000000fffffff7ffffffff0000000d00000000ffffffefffffffff",
            INIT_63 => X"0000000d00000000ffffffbefffffffffffffffeffffffff0000000f00000000",
            INIT_64 => X"00000013000000000000001a0000000000000008000000000000000500000000",
            INIT_65 => X"000000210000000000000031000000000000000100000000ffffffeeffffffff",
            INIT_66 => X"ffffffc9ffffffff00000027000000000000000300000000fffffffdffffffff",
            INIT_67 => X"00000049000000000000001f00000000fffffffdffffffffffffffdfffffffff",
            INIT_68 => X"0000003900000000ffffffdfffffffff00000041000000000000000700000000",
            INIT_69 => X"0000002000000000ffffffd4ffffffffffffffecffffffff0000001600000000",
            INIT_6A => X"0000000400000000fffffffcfffffffffffffff3fffffffffffffff1ffffffff",
            INIT_6B => X"fffffff7ffffffffffffffc9ffffffffffffffd9ffffffff0000000500000000",
            INIT_6C => X"ffffffe6ffffffff0000001500000000ffffffedffffffff0000000b00000000",
            INIT_6D => X"0000000400000000fffffff7ffffffff0000001100000000fffffffcffffffff",
            INIT_6E => X"ffffffd4ffffffff0000001f0000000000000002000000000000001000000000",
            INIT_6F => X"0000002700000000fffffff9ffffffffffffffccfffffffffffffffdffffffff",
            INIT_70 => X"0000002100000000000000260000000000000012000000000000000000000000",
            INIT_71 => X"00000001000000000000000e00000000ffffffe8ffffffffffffffd9ffffffff",
            INIT_72 => X"fffffff3ffffffff0000001700000000fffffff9fffffffffffffff8ffffffff",
            INIT_73 => X"ffffffdbffffffffffffffdcfffffffffffffffbffffffffffffffecffffffff",
            INIT_74 => X"0000004b00000000fffffff7ffffffff0000000000000000ffffffecffffffff",
            INIT_75 => X"0000001700000000ffffffd4ffffffff0000002e000000000000000000000000",
            INIT_76 => X"ffffffd0fffffffffffffff0fffffffffffffff4ffffffffffffffeeffffffff",
            INIT_77 => X"0000002400000000fffffff2ffffffffffffffbaffffffffffffffd5ffffffff",
            INIT_78 => X"ffffffe5ffffffff00000021000000000000001a000000000000001100000000",
            INIT_79 => X"fffffffcffffffffffffffecfffffffffffffff5ffffffffffffffdbffffffff",
            INIT_7A => X"ffffffddffffffff0000002b000000000000001b00000000ffffffbfffffffff",
            INIT_7B => X"ffffffddffffffffffffffedfffffffffffffff5ffffffffffffffd7ffffffff",
            INIT_7C => X"0000001000000000ffffffecfffffffffffffffafffffffffffffff0ffffffff",
            INIT_7D => X"0000002700000000ffffffc9ffffffff00000004000000000000000d00000000",
            INIT_7E => X"ffffffadffffffffffffffe4ffffffff0000001200000000fffffffaffffffff",
            INIT_7F => X"00000017000000000000000b00000000ffffffc9ffffffffffffffc2ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE8;


    MEM_IWGHT_LAYER2_INSTANCE9 : if BRAM_NAME = "iwght_layer2_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001200000000000000400000000000000025000000000000000a00000000",
            INIT_01 => X"fffffffaffffffff0000000900000000ffffffddfffffffffffffff1ffffffff",
            INIT_02 => X"ffffffd8ffffffff00000010000000000000000800000000ffffffd4ffffffff",
            INIT_03 => X"fffffff3ffffffff0000000f00000000fffffff9fffffffffffffff5ffffffff",
            INIT_04 => X"0000003e00000000ffffffd9fffffffffffffff6fffffffffffffff4ffffffff",
            INIT_05 => X"0000001f00000000ffffffe2ffffffff0000002f000000000000002000000000",
            INIT_06 => X"ffffffc0ffffffffffffffcfffffffffffffffe1ffffffff0000000d00000000",
            INIT_07 => X"00000000000000000000001400000000ffffffc0ffffffff0000000800000000",
            INIT_08 => X"00000012000000000000004a000000000000002000000000fffffffeffffffff",
            INIT_09 => X"0000000b00000000fffffff5ffffffffffffffe1ffffffff0000000500000000",
            INIT_0A => X"ffffffe1ffffffffffffffd5ffffffff0000001100000000ffffffe4ffffffff",
            INIT_0B => X"00000004000000000000002d00000000fffffffbffffffff0000000600000000",
            INIT_0C => X"0000002100000000ffffffd7ffffffff00000012000000000000000100000000",
            INIT_0D => X"00000008000000000000000a000000000000000c00000000fffffffeffffffff",
            INIT_0E => X"ffffffcbffffffffffffffdcffffffff00000002000000000000000600000000",
            INIT_0F => X"0000000a000000000000000700000000ffffffe7ffffffff0000000b00000000",
            INIT_10 => X"ffffffefffffffff00000049000000000000000a000000000000000000000000",
            INIT_11 => X"ffffffecfffffffffffffff1fffffffffffffffafffffffffffffff7ffffffff",
            INIT_12 => X"ffffffdaffffffffffffffa1ffffffff0000001800000000ffffffebffffffff",
            INIT_13 => X"fffffff3ffffffff000000120000000000000013000000000000000200000000",
            INIT_14 => X"fffffff0ffffffffffffffdcffffffff00000018000000000000000300000000",
            INIT_15 => X"0000002d000000000000001d0000000000000016000000000000000900000000",
            INIT_16 => X"ffffffecffffffffffffffdaffffffff00000008000000000000000100000000",
            INIT_17 => X"ffffffebffffffff00000017000000000000001000000000fffffff0ffffffff",
            INIT_18 => X"ffffffe7ffffffff0000000e00000000ffffffeefffffffffffffff3ffffffff",
            INIT_19 => X"fffffff9ffffffffffffffe0ffffffff00000009000000000000000000000000",
            INIT_1A => X"fffffff1ffffffff000000010000000000000003000000000000000800000000",
            INIT_1B => X"00000004000000000000000a00000000fffffffbffffffffffffffd9ffffffff",
            INIT_1C => X"0000001100000000ffffffefffffffff0000001900000000ffffffdeffffffff",
            INIT_1D => X"0000001c000000000000000000000000ffffffd9ffffffffffffffe1ffffffff",
            INIT_1E => X"0000001e00000000ffffffd8ffffffffffffffdcffffffffffffffd2ffffffff",
            INIT_1F => X"00000010000000000000000400000000fffffff3ffffffff0000000a00000000",
            INIT_20 => X"fffffffdffffffff00000008000000000000001400000000fffffffbffffffff",
            INIT_21 => X"0000000100000000fffffffdffffffff00000007000000000000001100000000",
            INIT_22 => X"ffffffd4ffffffff0000001d00000000ffffffcaffffffffffffffefffffffff",
            INIT_23 => X"fffffff8ffffffff0000000b000000000000000900000000ffffffe7ffffffff",
            INIT_24 => X"0000001e0000000000000001000000000000000300000000ffffffe8ffffffff",
            INIT_25 => X"0000002600000000ffffffdfffffffff00000009000000000000000d00000000",
            INIT_26 => X"0000001000000000ffffffe4ffffffffffffffceffffffffffffffdeffffffff",
            INIT_27 => X"00000000000000000000000a00000000fffffff3ffffffff0000002200000000",
            INIT_28 => X"fffffff0ffffffff00000049000000000000001c00000000fffffffbffffffff",
            INIT_29 => X"ffffffedfffffffffffffffdffffffffffffffe4ffffffffffffffffffffffff",
            INIT_2A => X"fffffffbffffffff0000000500000000ffffffd7fffffffffffffffcffffffff",
            INIT_2B => X"00000011000000000000001500000000fffffffaffffffff0000001500000000",
            INIT_2C => X"0000000300000000fffffffbfffffffffffffff0ffffffffffffffefffffffff",
            INIT_2D => X"0000002600000000000000030000000000000000000000000000000d00000000",
            INIT_2E => X"0000002500000000ffffffe3ffffffffffffffbbffffffffffffffebffffffff",
            INIT_2F => X"000000070000000000000005000000000000000d000000000000002b00000000",
            INIT_30 => X"fffffff8ffffffff000000050000000000000001000000000000000f00000000",
            INIT_31 => X"fffffff7ffffffff0000001100000000ffffffe7ffffffff0000001c00000000",
            INIT_32 => X"00000010000000000000002d00000000ffffffe3fffffffffffffff0ffffffff",
            INIT_33 => X"0000000300000000fffffffdffffffff00000003000000000000000000000000",
            INIT_34 => X"0000000c0000000000000005000000000000000700000000ffffffe5ffffffff",
            INIT_35 => X"00000013000000000000000000000000fffffffeffffffff0000000000000000",
            INIT_36 => X"0000000d00000000ffffffdfffffffffffffffc5ffffffff0000000600000000",
            INIT_37 => X"0000001300000000000000120000000000000000000000000000001100000000",
            INIT_38 => X"fffffff6ffffffff00000000000000000000000b000000000000001400000000",
            INIT_39 => X"fffffffbffffffff0000001300000000ffffffedffffffff0000001e00000000",
            INIT_3A => X"fffffffdffffffff0000002b00000000ffffffeeffffffffffffffffffffffff",
            INIT_3B => X"fffffff5ffffffffffffffd8ffffffffffffffe0fffffffffffffff9ffffffff",
            INIT_3C => X"00000014000000000000000000000000fffffff6ffffffff0000000e00000000",
            INIT_3D => X"0000002900000000ffffffe9ffffffffffffffcafffffffffffffff3ffffffff",
            INIT_3E => X"0000001300000000ffffffeeffffffffffffffdfffffffff0000000600000000",
            INIT_3F => X"0000000a000000000000000c00000000ffffffffffffffff0000003100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffdcffffffff0000001a0000000000000018000000000000000c00000000",
            INIT_41 => X"fffffff9ffffffff0000000d00000000fffffffcfffffffffffffffeffffffff",
            INIT_42 => X"ffffffeeffffffff0000002200000000fffffff2ffffffff0000000d00000000",
            INIT_43 => X"ffffffecffffffffffffffedfffffffffffffffbffffffffffffffffffffffff",
            INIT_44 => X"00000011000000000000000300000000fffffffefffffffffffffff4ffffffff",
            INIT_45 => X"0000000c00000000ffffffe5ffffffffffffffd6ffffffffffffffd9ffffffff",
            INIT_46 => X"fffffff1ffffffff0000000800000000ffffffbbfffffffffffffff0ffffffff",
            INIT_47 => X"00000030000000000000000100000000fffffffbfffffffffffffff8ffffffff",
            INIT_48 => X"0000001700000000ffffffe8ffffffff0000001e000000000000001400000000",
            INIT_49 => X"00000019000000000000001100000000ffffffd9fffffffffffffff7ffffffff",
            INIT_4A => X"0000003c000000000000002a00000000fffffff5fffffffffffffffdffffffff",
            INIT_4B => X"0000000900000000ffffffd7ffffffff0000000200000000ffffffebffffffff",
            INIT_4C => X"0000000f00000000ffffffedfffffffffffffffdfffffffffffffffaffffffff",
            INIT_4D => X"fffffffbffffffffffffffd4ffffffffffffffe3ffffffffffffffe8ffffffff",
            INIT_4E => X"00000000000000000000000c00000000ffffffdcffffffffffffffd7ffffffff",
            INIT_4F => X"0000000f00000000ffffffe9ffffffffffffffe9fffffffffffffff8ffffffff",
            INIT_50 => X"fffffff6ffffffff00000014000000000000002c00000000fffffff7ffffffff",
            INIT_51 => X"fffffffdffffffffffffffeffffffffffffffff7ffffffff0000000500000000",
            INIT_52 => X"fffffff5ffffffff0000001100000000ffffffe1fffffffffffffffaffffffff",
            INIT_53 => X"fffffff3ffffffff00000006000000000000000200000000ffffffcdffffffff",
            INIT_54 => X"fffffffdffffffffffffffebffffffff0000002c000000000000000000000000",
            INIT_55 => X"0000001a00000000fffffff6ffffffff0000000500000000fffffffdffffffff",
            INIT_56 => X"0000000400000000fffffffbffffffffffffffd9ffffffff0000000700000000",
            INIT_57 => X"0000001000000000fffffffbffffffff0000001d000000000000001f00000000",
            INIT_58 => X"fffffffcffffffff00000024000000000000000200000000fffffff6ffffffff",
            INIT_59 => X"0000000100000000fffffffaffffffff00000015000000000000000100000000",
            INIT_5A => X"fffffff8ffffffff0000000700000000fffffffdffffffff0000001600000000",
            INIT_5B => X"000000170000000000000024000000000000000300000000fffffff7ffffffff",
            INIT_5C => X"0000001c00000000000000070000000000000009000000000000000600000000",
            INIT_5D => X"0000001200000000ffffffdafffffffffffffff2ffffffff0000000200000000",
            INIT_5E => X"0000000b000000000000000f00000000ffffffefffffffff0000001100000000",
            INIT_5F => X"fffffff3ffffffff000000190000000000000017000000000000000200000000",
            INIT_60 => X"fffffffcffffffff0000001a000000000000001900000000fffffff7ffffffff",
            INIT_61 => X"ffffffedffffffff0000000900000000fffffff3ffffffffffffffe8ffffffff",
            INIT_62 => X"00000019000000000000001200000000ffffffccffffffff0000000700000000",
            INIT_63 => X"000000050000000000000007000000000000000000000000fffffff8ffffffff",
            INIT_64 => X"0000000200000000fffffffaffffffff0000000500000000ffffffe7ffffffff",
            INIT_65 => X"ffffffebffffffffffffffe6fffffffffffffff9fffffffffffffff7ffffffff",
            INIT_66 => X"0000000700000000ffffffebffffffffffffffbfffffffff0000001100000000",
            INIT_67 => X"ffffffe9ffffffff0000000000000000ffffffe6ffffffff0000000f00000000",
            INIT_68 => X"fffffffdffffffff000000380000000000000016000000000000000000000000",
            INIT_69 => X"00000010000000000000001400000000ffffffeaffffffff0000000000000000",
            INIT_6A => X"0000000d00000000000000040000000000000006000000000000000000000000",
            INIT_6B => X"fffffff8fffffffffffffff2fffffffffffffffcffffffffffffffd9ffffffff",
            INIT_6C => X"0000001800000000000000070000000000000010000000000000000e00000000",
            INIT_6D => X"ffffffdeffffffffffffffe8ffffffffffffffeaffffffff0000000b00000000",
            INIT_6E => X"ffffffe0ffffffffffffffedfffffffffffffff9ffffffff0000001400000000",
            INIT_6F => X"fffffff7fffffffffffffffeffffffff00000002000000000000002200000000",
            INIT_70 => X"ffffffeefffffffffffffffffffffffffffffffdffffffff0000001000000000",
            INIT_71 => X"00000018000000000000000000000000fffffffdffffffff0000000000000000",
            INIT_72 => X"00000008000000000000002200000000ffffffdffffffffffffffff6ffffffff",
            INIT_73 => X"000000210000000000000016000000000000000600000000fffffff2ffffffff",
            INIT_74 => X"ffffffffffffffff0000000f00000000fffffff5ffffffff0000000f00000000",
            INIT_75 => X"fffffff9ffffffffffffffeaffffffffffffffc3fffffffffffffff5ffffffff",
            INIT_76 => X"ffffffe4fffffffffffffffbffffffff00000011000000000000002b00000000",
            INIT_77 => X"ffffffefffffffff0000001300000000ffffffdeffffffff0000002400000000",
            INIT_78 => X"fffffffdfffffffffffffff3ffffffff00000004000000000000001900000000",
            INIT_79 => X"000000080000000000000008000000000000000700000000ffffffefffffffff",
            INIT_7A => X"0000000a000000000000001400000000ffffffdefffffffffffffff8ffffffff",
            INIT_7B => X"0000002000000000ffffffeaffffffff0000000700000000fffffff1ffffffff",
            INIT_7C => X"0000001e00000000fffffff5ffffffffffffffe0ffffffff0000000300000000",
            INIT_7D => X"ffffffe3ffffffffffffffd4fffffffffffffff8ffffffff0000001d00000000",
            INIT_7E => X"0000000900000000ffffffdeffffffffffffffb9fffffffffffffff4ffffffff",
            INIT_7F => X"0000000200000000fffffff1fffffffffffffff9ffffffff0000000d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE9;


    MEM_IWGHT_LAYER2_INSTANCE10 : if BRAM_NAME = "iwght_layer2_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff7ffffffff000000160000000000000012000000000000000b00000000",
            INIT_01 => X"ffffffffffffffff0000002700000000fffffffdffffffffffffffe5ffffffff",
            INIT_02 => X"0000001300000000000000170000000000000001000000000000000f00000000",
            INIT_03 => X"0000001200000000fffffff8fffffffffffffffaffffffffffffffe2ffffffff",
            INIT_04 => X"0000000c000000000000000e000000000000001f000000000000000d00000000",
            INIT_05 => X"fffffff6ffffffffffffffd7ffffffffffffffe6ffffffff0000000000000000",
            INIT_06 => X"fffffffeffffffffffffffe7ffffffff0000000a000000000000000200000000",
            INIT_07 => X"0000000900000000fffffffeffffffff00000007000000000000001800000000",
            INIT_08 => X"ffffffffffffffff0000001d000000000000000c00000000fffffff9ffffffff",
            INIT_09 => X"fffffffeffffffffffffffffffffffff0000000a000000000000000d00000000",
            INIT_0A => X"fffffff5ffffffff0000001700000000fffffffafffffffffffffffbffffffff",
            INIT_0B => X"000000060000000000000000000000000000000600000000ffffffe2ffffffff",
            INIT_0C => X"0000000300000000fffffffcffffffff00000000000000000000000d00000000",
            INIT_0D => X"fffffffbfffffffffffffff3ffffffffffffffe4ffffffff0000000400000000",
            INIT_0E => X"fffffff9fffffffffffffff3ffffffffffffffb9ffffffff0000000c00000000",
            INIT_0F => X"00000005000000000000001700000000ffffffdeffffffff0000001c00000000",
            INIT_10 => X"0000000c000000000000002300000000fffffff8ffffffff0000000400000000",
            INIT_11 => X"fffffff2ffffffff0000000b000000000000001d000000000000000b00000000",
            INIT_12 => X"0000001800000000ffffffe9fffffffffffffff9ffffffff0000000800000000",
            INIT_13 => X"0000000000000000fffffff1ffffffff0000000000000000fffffff2ffffffff",
            INIT_14 => X"00000005000000000000001100000000fffffff5ffffffff0000000600000000",
            INIT_15 => X"0000000d00000000ffffffc7ffffffff00000008000000000000000300000000",
            INIT_16 => X"ffffffdffffffffffffffffaffffffffffffffd3ffffffffffffffe7ffffffff",
            INIT_17 => X"fffffff1fffffffffffffff5ffffffffffffffd5ffffffffffffffe9ffffffff",
            INIT_18 => X"fffffffcffffffff00000009000000000000001500000000fffffff6ffffffff",
            INIT_19 => X"0000000a00000000fffffff4ffffffffffffffe6fffffffffffffffdffffffff",
            INIT_1A => X"0000001200000000fffffffcffffffffffffffd9ffffffff0000002200000000",
            INIT_1B => X"0000000f00000000000000090000000000000008000000000000001200000000",
            INIT_1C => X"fffffff7ffffffff0000000000000000ffffffefffffffffffffffdfffffffff",
            INIT_1D => X"ffffffebffffffffffffffb2ffffffff0000000700000000fffffff2ffffffff",
            INIT_1E => X"0000002600000000fffffff8ffffffff0000000600000000fffffff6ffffffff",
            INIT_1F => X"ffffffe3fffffffffffffff6ffffffffffffffeaffffffffffffffccffffffff",
            INIT_20 => X"0000000000000000000000290000000000000011000000000000001800000000",
            INIT_21 => X"fffffffeffffffff0000000300000000ffffffc3fffffffffffffffbffffffff",
            INIT_22 => X"ffffffffffffffffffffffefffffffffffffffcbffffffff0000000300000000",
            INIT_23 => X"fffffff8ffffffff0000000600000000ffffffe8fffffffffffffff2ffffffff",
            INIT_24 => X"0000001800000000fffffffbffffffff00000016000000000000000200000000",
            INIT_25 => X"0000000e00000000ffffffb0ffffffff00000002000000000000001800000000",
            INIT_26 => X"ffffffd7ffffffff0000000d0000000000000010000000000000004c00000000",
            INIT_27 => X"ffffffebffffffff0000001c00000000ffffffe2fffffffffffffff2ffffffff",
            INIT_28 => X"00000013000000000000001c000000000000000c000000000000002f00000000",
            INIT_29 => X"00000010000000000000002200000000ffffffc5ffffffffffffffedffffffff",
            INIT_2A => X"fffffffdfffffffffffffffbffffffffffffffd6ffffffff0000000000000000",
            INIT_2B => X"0000001b000000000000001300000000fffffffbffffffff0000001600000000",
            INIT_2C => X"fffffffdffffffff00000000000000000000000c000000000000002200000000",
            INIT_2D => X"0000002300000000ffffffd5fffffffffffffffaffffffff0000002200000000",
            INIT_2E => X"fffffff2ffffffffffffffe2ffffffff0000000b000000000000000700000000",
            INIT_2F => X"ffffffd6ffffffff0000001400000000ffffffd9ffffffff0000000f00000000",
            INIT_30 => X"00000035000000000000001600000000fffffffcffffffff0000001300000000",
            INIT_31 => X"0000000f000000000000001000000000ffffffd0ffffffffffffffcdffffffff",
            INIT_32 => X"ffffffedffffffff0000000800000000fffffffcfffffffffffffffeffffffff",
            INIT_33 => X"0000000600000000fffffffeffffffff00000001000000000000000c00000000",
            INIT_34 => X"000000000000000000000000000000000000001300000000fffffff2ffffffff",
            INIT_35 => X"0000001100000000ffffffe8ffffffff0000000300000000ffffffefffffffff",
            INIT_36 => X"fffffff5ffffffffffffffe2ffffffff0000001000000000fffffff3ffffffff",
            INIT_37 => X"fffffffcffffffff0000001800000000fffffff8ffffffff0000001800000000",
            INIT_38 => X"fffffff3ffffffff0000000b00000000ffffffecffffffff0000002300000000",
            INIT_39 => X"00000003000000000000000f00000000ffffffe8ffffffffffffffddffffffff",
            INIT_3A => X"fffffffcffffffffffffffeefffffffffffffff1fffffffffffffff2ffffffff",
            INIT_3B => X"0000001300000000fffffffbfffffffffffffffeffffffffffffffe7ffffffff",
            INIT_3C => X"0000000a0000000000000005000000000000001200000000fffffff5ffffffff",
            INIT_3D => X"0000003500000000ffffffcaffffffff0000000c000000000000001500000000",
            INIT_3E => X"0000000800000000ffffffaffffffffffffffffdffffffff0000002200000000",
            INIT_3F => X"fffffff6fffffffffffffffaffffffffffffffd7ffffffff0000002700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000900000000000000140000000000000017000000000000000300000000",
            INIT_41 => X"0000000000000000fffffff1ffffffff0000001900000000ffffffe7ffffffff",
            INIT_42 => X"ffffffffffffffff00000012000000000000001200000000ffffffe6ffffffff",
            INIT_43 => X"ffffffe8ffffffffffffffeeffffffffffffffe9ffffffff0000000500000000",
            INIT_44 => X"00000000000000000000001c000000000000001400000000ffffffebffffffff",
            INIT_45 => X"ffffffe8ffffffff00000001000000000000001600000000fffffff7ffffffff",
            INIT_46 => X"00000004000000000000002000000000ffffffedffffffff0000003a00000000",
            INIT_47 => X"fffffffdffffffff0000000500000000ffffffcdffffffff0000002600000000",
            INIT_48 => X"000000000000000000000012000000000000001c000000000000000400000000",
            INIT_49 => X"0000000700000000000000040000000000000004000000000000000400000000",
            INIT_4A => X"0000001600000000fffffff1ffffffff00000019000000000000000e00000000",
            INIT_4B => X"fffffff9ffffffffffffffdeffffffffffffffe6ffffffff0000000a00000000",
            INIT_4C => X"0000000e0000000000000002000000000000000000000000ffffffffffffffff",
            INIT_4D => X"0000000f00000000ffffffa5ffffffff0000001200000000fffffffdffffffff",
            INIT_4E => X"fffffff9ffffffffffffffdbfffffffffffffff7ffffffff0000001100000000",
            INIT_4F => X"00000009000000000000000000000000ffffffd6fffffffffffffffbffffffff",
            INIT_50 => X"00000000000000000000001b0000000000000010000000000000001300000000",
            INIT_51 => X"00000008000000000000001e00000000fffffff1ffffffffffffffe1ffffffff",
            INIT_52 => X"0000000600000000ffffffd8fffffffffffffff5fffffffffffffffcffffffff",
            INIT_53 => X"00000000000000000000000000000000fffffffbfffffffffffffff9ffffffff",
            INIT_54 => X"00000000000000000000000e00000000fffffff4fffffffffffffff2ffffffff",
            INIT_55 => X"0000000400000000ffffffb4ffffffff0000001c000000000000000300000000",
            INIT_56 => X"ffffffdeffffffff00000009000000000000000e000000000000000700000000",
            INIT_57 => X"ffffffe2ffffffffffffffffffffffff0000000200000000ffffffc5ffffffff",
            INIT_58 => X"ffffffeeffffffff000000270000000000000015000000000000000300000000",
            INIT_59 => X"00000001000000000000001000000000ffffffd0ffffffffffffffd2ffffffff",
            INIT_5A => X"ffffffe3ffffffffffffffdefffffffffffffff9ffffffffffffffe3ffffffff",
            INIT_5B => X"fffffff2ffffffff0000001200000000fffffffeffffffff0000000200000000",
            INIT_5C => X"00000006000000000000001400000000ffffffedffffffff0000000500000000",
            INIT_5D => X"0000000c00000000ffffffe1ffffffff00000025000000000000000f00000000",
            INIT_5E => X"ffffffd8ffffffffffffffd9ffffffff0000002c000000000000001b00000000",
            INIT_5F => X"ffffffd9ffffffff0000000f00000000ffffffe0ffffffffffffffecffffffff",
            INIT_60 => X"0000000f000000000000000b0000000000000011000000000000000c00000000",
            INIT_61 => X"0000000f000000000000000e00000000ffffffbdffffffffffffffc7ffffffff",
            INIT_62 => X"ffffffeeffffffffffffffd1ffffffffffffffe4ffffffffffffffdbffffffff",
            INIT_63 => X"fffffff9ffffffff0000000c00000000fffffffaffffffff0000001000000000",
            INIT_64 => X"0000000c00000000ffffffe0ffffffff00000007000000000000002400000000",
            INIT_65 => X"0000002400000000ffffffdbffffffff0000001a000000000000001d00000000",
            INIT_66 => X"ffffffdaffffffffffffffc4ffffffff00000017000000000000000900000000",
            INIT_67 => X"00000005000000000000001900000000ffffffb4ffffffff0000000c00000000",
            INIT_68 => X"0000000000000000000000220000000000000016000000000000000500000000",
            INIT_69 => X"0000000e000000000000001a00000000ffffffdbffffffffffffffdbffffffff",
            INIT_6A => X"0000001900000000fffffff5fffffffffffffff3ffffffffffffffd2ffffffff",
            INIT_6B => X"000000150000000000000006000000000000000000000000fffffffbffffffff",
            INIT_6C => X"000000080000000000000000000000000000000e00000000fffffff8ffffffff",
            INIT_6D => X"0000001d00000000ffffffbeffffffff0000000900000000fffffffcffffffff",
            INIT_6E => X"0000001300000000ffffffc7ffffffff0000003f000000000000001e00000000",
            INIT_6F => X"0000000400000000fffffffafffffffffffffff1fffffffffffffffeffffffff",
            INIT_70 => X"ffffffdfffffffff000000160000000000000002000000000000002a00000000",
            INIT_71 => X"00000010000000000000001b00000000ffffffe9ffffffffffffffdfffffffff",
            INIT_72 => X"ffffffffffffffffffffffefffffffffffffffeffffffffffffffff1ffffffff",
            INIT_73 => X"ffffffe5ffffffff0000002200000000fffffffcffffffff0000000000000000",
            INIT_74 => X"0000000100000000fffffff2fffffffffffffffcfffffffffffffffbffffffff",
            INIT_75 => X"0000001200000000ffffffd6ffffffffffffffffffffffff0000002e00000000",
            INIT_76 => X"ffffffe9ffffffffffffffd8ffffffffffffffc7ffffffff0000000400000000",
            INIT_77 => X"ffffffebffffffff0000000f00000000ffffffd5ffffffff0000001500000000",
            INIT_78 => X"ffffffddffffffff00000016000000000000001f000000000000000c00000000",
            INIT_79 => X"0000000f000000000000000d00000000fffffffdffffffff0000000500000000",
            INIT_7A => X"ffffffecffffffff000000040000000000000014000000000000000c00000000",
            INIT_7B => X"fffffff7ffffffffffffffdafffffffffffffff5fffffffffffffff7ffffffff",
            INIT_7C => X"ffffffddffffffff0000000000000000ffffffd1ffffffff0000000c00000000",
            INIT_7D => X"0000001900000000ffffffe8fffffffffffffff8fffffffffffffffcffffffff",
            INIT_7E => X"ffffffe1ffffffff0000001000000000ffffffeeffffffff0000000000000000",
            INIT_7F => X"0000000000000000fffffff2ffffffffffffffedfffffffffffffff2ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE10;


    MEM_IWGHT_LAYER2_INSTANCE11 : if BRAM_NAME = "iwght_layer2_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000e0000000000000026000000000000000e00000000ffffffeaffffffff",
            INIT_01 => X"0000000d0000000000000019000000000000001000000000fffffffeffffffff",
            INIT_02 => X"ffffffdcffffffffffffffddfffffffffffffff7ffffffff0000000100000000",
            INIT_03 => X"fffffff9fffffffffffffff2ffffffff0000000000000000fffffff1ffffffff",
            INIT_04 => X"ffffffe2fffffffffffffffcfffffffffffffff0ffffffff0000000d00000000",
            INIT_05 => X"0000001100000000ffffffdbffffffff0000002200000000ffffffeaffffffff",
            INIT_06 => X"fffffffcffffffffffffffe7ffffffff0000000800000000fffffffeffffffff",
            INIT_07 => X"ffffffd4fffffffffffffff8ffffffffffffffe0ffffffffffffffebffffffff",
            INIT_08 => X"00000000000000000000001d0000000000000005000000000000000200000000",
            INIT_09 => X"0000001400000000fffffffefffffffffffffff3ffffffffffffffc6ffffffff",
            INIT_0A => X"ffffffdeffffffffffffffe4ffffffff0000000900000000fffffff4ffffffff",
            INIT_0B => X"fffffff1fffffffffffffff2fffffffffffffffdffffffffffffffeeffffffff",
            INIT_0C => X"00000006000000000000002000000000fffffff4ffffffff0000000f00000000",
            INIT_0D => X"0000001700000000ffffffaeffffffff0000001c000000000000000300000000",
            INIT_0E => X"ffffffdeffffffff00000011000000000000002600000000ffffffccffffffff",
            INIT_0F => X"fffffff2ffffffff0000000100000000ffffffe1ffffffffffffffe4ffffffff",
            INIT_10 => X"ffffffe7ffffffff0000003a000000000000000a000000000000000c00000000",
            INIT_11 => X"00000008000000000000000b00000000ffffffe4ffffffffffffffecffffffff",
            INIT_12 => X"ffffffcfffffffffffffffe9fffffffffffffff5ffffffffffffffd6ffffffff",
            INIT_13 => X"ffffffeefffffffffffffffaffffffff0000000500000000ffffffdaffffffff",
            INIT_14 => X"0000000b00000000fffffff4ffffffff0000000c000000000000000d00000000",
            INIT_15 => X"0000002f00000000ffffffd8ffffffff0000004a000000000000000d00000000",
            INIT_16 => X"ffffffcdffffffff0000001100000000ffffffafffffffffffffffd7ffffffff",
            INIT_17 => X"fffffff2ffffffffffffffecffffffffffffffe3ffffffffffffffd2ffffffff",
            INIT_18 => X"ffffffe6ffffffff0000002b00000000fffffff5ffffffff0000000000000000",
            INIT_19 => X"00000004000000000000000500000000ffffffebffffffffffffffe9ffffffff",
            INIT_1A => X"fffffff4ffffffffffffffefffffffff0000000200000000fffffffcffffffff",
            INIT_1B => X"fffffff7ffffffffffffffebfffffffffffffffcffffffffffffffecffffffff",
            INIT_1C => X"fffffff5fffffffffffffff3ffffffff00000004000000000000000200000000",
            INIT_1D => X"0000000f00000000fffffff8ffffffff0000001b000000000000000c00000000",
            INIT_1E => X"0000000500000000ffffffdeffffffffffffffeffffffffffffffff0ffffffff",
            INIT_1F => X"0000000d0000000000000005000000000000000800000000ffffffe2ffffffff",
            INIT_20 => X"fffffff7ffffffff0000002e0000000000000009000000000000000200000000",
            INIT_21 => X"00000014000000000000001000000000ffffffffffffffffffffffc8ffffffff",
            INIT_22 => X"fffffff7ffffffffffffffe9fffffffffffffffdffffffffffffffeaffffffff",
            INIT_23 => X"0000000e00000000fffffff8fffffffffffffffcfffffffffffffffaffffffff",
            INIT_24 => X"fffffff7ffffffff000000010000000000000007000000000000000000000000",
            INIT_25 => X"fffffff8ffffffffffffffc8ffffffff0000001300000000fffffff1ffffffff",
            INIT_26 => X"fffffff1ffffffffffffffebffffffff0000000e00000000ffffffe4ffffffff",
            INIT_27 => X"ffffffe3ffffffff0000001300000000ffffffeffffffffffffffffdffffffff",
            INIT_28 => X"ffffffd8ffffffff0000001e000000000000000b000000000000000800000000",
            INIT_29 => X"0000001100000000fffffff6ffffffffffffffe6ffffffffffffffd7ffffffff",
            INIT_2A => X"0000000000000000ffffffeeffffffffffffffe4ffffffffffffffe0ffffffff",
            INIT_2B => X"0000001900000000ffffffdbffffffff0000001e00000000ffffffeeffffffff",
            INIT_2C => X"fffffffdffffffff00000011000000000000000e000000000000000300000000",
            INIT_2D => X"fffffffeffffffffffffffebffffffff0000000b000000000000002500000000",
            INIT_2E => X"fffffffbffffffffffffffe6ffffffffffffffcbfffffffffffffff2ffffffff",
            INIT_2F => X"00000011000000000000000000000000ffffffeafffffffffffffff8ffffffff",
            INIT_30 => X"fffffff0ffffffff0000002800000000fffffff2ffffffff0000001300000000",
            INIT_31 => X"0000000b000000000000001700000000fffffff7ffffffffffffffffffffffff",
            INIT_32 => X"fffffff6ffffffffffffffffffffffff0000001000000000fffffff6ffffffff",
            INIT_33 => X"0000000300000000ffffffefffffffff00000000000000000000000f00000000",
            INIT_34 => X"fffffff5ffffffff0000001f0000000000000012000000000000000f00000000",
            INIT_35 => X"0000002400000000fffffffdffffffff00000009000000000000000100000000",
            INIT_36 => X"fffffffcffffffff000000300000000000000016000000000000002600000000",
            INIT_37 => X"fffffff9ffffffffffffffe4ffffffffffffffe4ffffffff0000002000000000",
            INIT_38 => X"0000000a000000000000001b0000000000000000000000000000000000000000",
            INIT_39 => X"0000000d00000000fffffffbffffffff0000002600000000fffffffaffffffff",
            INIT_3A => X"ffffffc9fffffffffffffff3ffffffff00000024000000000000002b00000000",
            INIT_3B => X"0000000000000000fffffff6ffffffff0000000a00000000ffffffffffffffff",
            INIT_3C => X"00000002000000000000000d000000000000000f00000000fffffff7ffffffff",
            INIT_3D => X"0000001900000000ffffffd8ffffffff0000001100000000ffffffeeffffffff",
            INIT_3E => X"000000090000000000000002000000000000003b00000000ffffffe5ffffffff",
            INIT_3F => X"fffffff6ffffffff00000005000000000000000000000000ffffffe2ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffffcffffffff0000003e000000000000001000000000fffffff9ffffffff",
            INIT_41 => X"ffffffffffffffff0000000200000000ffffffffffffffffffffffd3ffffffff",
            INIT_42 => X"ffffffb8fffffffffffffffefffffffffffffff3fffffffffffffff2ffffffff",
            INIT_43 => X"fffffff7fffffffffffffffdffffffff0000001300000000fffffff8ffffffff",
            INIT_44 => X"0000000500000000ffffffefffffffff00000011000000000000001300000000",
            INIT_45 => X"fffffff9fffffffffffffff9ffffffff0000002c000000000000000c00000000",
            INIT_46 => X"0000000100000000fffffff7ffffffffffffffd9ffffffff0000000e00000000",
            INIT_47 => X"fffffff4ffffffff000000090000000000000004000000000000001000000000",
            INIT_48 => X"fffffffbffffffff0000002c00000000fffffffcffffffff0000000300000000",
            INIT_49 => X"0000001100000000fffffff5ffffffffffffffe2fffffffffffffff1ffffffff",
            INIT_4A => X"ffffffe8fffffffffffffff6ffffffff0000000c000000000000000300000000",
            INIT_4B => X"fffffff8ffffffffffffffefffffffff0000000000000000ffffffd4ffffffff",
            INIT_4C => X"ffffffeaffffffff0000001c00000000fffffff4ffffffff0000000b00000000",
            INIT_4D => X"fffffffdfffffffffffffffbffffffff00000003000000000000001100000000",
            INIT_4E => X"ffffffefffffffff0000000b000000000000001a000000000000001a00000000",
            INIT_4F => X"0000000b000000000000000a00000000fffffff6ffffffff0000001100000000",
            INIT_50 => X"fffffff8ffffffff000000340000000000000008000000000000000100000000",
            INIT_51 => X"0000001000000000fffffff3ffffffff0000001400000000fffffff8ffffffff",
            INIT_52 => X"fffffffbfffffffffffffffcffffffff0000000400000000ffffffefffffffff",
            INIT_53 => X"fffffffcffffffffffffffeffffffffffffffff4fffffffffffffff6ffffffff",
            INIT_54 => X"fffffff0ffffffff0000000a0000000000000006000000000000000f00000000",
            INIT_55 => X"0000001200000000000000040000000000000001000000000000000f00000000",
            INIT_56 => X"0000001e000000000000001300000000fffffff8ffffffff0000000600000000",
            INIT_57 => X"0000000900000000fffffff9ffffffffffffffe9ffffffffffffffcfffffffff",
            INIT_58 => X"fffffff2ffffffff0000002100000000fffffff0ffffffff0000000400000000",
            INIT_59 => X"00000002000000000000000200000000fffffff5ffffffffffffffe5ffffffff",
            INIT_5A => X"ffffffe4ffffffffffffffe6ffffffff0000000a00000000ffffffeaffffffff",
            INIT_5B => X"0000000300000000ffffffbcffffffff0000001000000000fffffff8ffffffff",
            INIT_5C => X"0000000600000000fffffffaffffffffffffffd1ffffffff0000000c00000000",
            INIT_5D => X"0000000100000000fffffffcffffffff0000002800000000fffffff9ffffffff",
            INIT_5E => X"0000001200000000ffffffdeffffffff0000002200000000ffffffd5ffffffff",
            INIT_5F => X"fffffff1ffffffff0000000100000000fffffff4ffffffffffffffefffffffff",
            INIT_60 => X"ffffffffffffffff00000034000000000000000a000000000000001900000000",
            INIT_61 => X"00000004000000000000001700000000ffffffe6ffffffffffffffcaffffffff",
            INIT_62 => X"00000006000000000000000900000000fffffff9fffffffffffffff2ffffffff",
            INIT_63 => X"0000000500000000ffffffeaffffffff0000000c00000000fffffff6ffffffff",
            INIT_64 => X"fffffff8ffffffff00000001000000000000000c000000000000000300000000",
            INIT_65 => X"fffffff9ffffffffffffffe1ffffffff00000000000000000000001f00000000",
            INIT_66 => X"000000080000000000000000000000000000002e00000000fffffffaffffffff",
            INIT_67 => X"fffffffaffffffffffffffeaffffffff00000000000000000000000800000000",
            INIT_68 => X"fffffffcffffffff00000017000000000000000e000000000000000700000000",
            INIT_69 => X"0000000f00000000fffffff2ffffffffffffffffffffffffffffffd7ffffffff",
            INIT_6A => X"fffffff5ffffffff00000000000000000000001a000000000000001000000000",
            INIT_6B => X"ffffffe8ffffffffffffffddfffffffffffffff6ffffffff0000000000000000",
            INIT_6C => X"fffffffaffffffff00000015000000000000002400000000fffffff8ffffffff",
            INIT_6D => X"0000002c000000000000001700000000fffffffdffffffff0000001700000000",
            INIT_6E => X"fffffffbffffffff0000000f0000000000000025000000000000001b00000000",
            INIT_6F => X"0000002e00000000ffffffeaffffffffffffffefffffffff0000002000000000",
            INIT_70 => X"0000002a0000000000000012000000000000003700000000fffffffcffffffff",
            INIT_71 => X"0000000800000000ffffffeeffffffff00000023000000000000001b00000000",
            INIT_72 => X"ffffffd9ffffffff000000140000000000000019000000000000002c00000000",
            INIT_73 => X"fffffffdffffffff0000001700000000fffffff0ffffffffffffffebffffffff",
            INIT_74 => X"fffffff3fffffffffffffffcffffffff0000001300000000ffffffffffffffff",
            INIT_75 => X"0000001b00000000ffffffeffffffffffffffffafffffffffffffffdffffffff",
            INIT_76 => X"0000000b0000000000000001000000000000000200000000ffffffe8ffffffff",
            INIT_77 => X"0000000800000000fffffff7fffffffffffffff0fffffffffffffffeffffffff",
            INIT_78 => X"0000001c00000000000000290000000000000012000000000000000200000000",
            INIT_79 => X"fffffffcffffffffffffffeefffffffffffffffffffffffffffffff9ffffffff",
            INIT_7A => X"ffffffbdffffffff00000005000000000000000a00000000fffffffbffffffff",
            INIT_7B => X"000000150000000000000004000000000000002700000000ffffffe9ffffffff",
            INIT_7C => X"ffffffe6ffffffff000000060000000000000007000000000000002100000000",
            INIT_7D => X"fffffff9ffffffffffffffdfffffffffffffffd9ffffffff0000000b00000000",
            INIT_7E => X"fffffff3ffffffff0000000e00000000ffffffeefffffffffffffff8ffffffff",
            INIT_7F => X"ffffffeaffffffff0000000a0000000000000000000000000000000d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE11;


    MEM_IWGHT_LAYER2_INSTANCE12 : if BRAM_NAME = "iwght_layer2_instance12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff7ffffffff0000002f000000000000000a000000000000001500000000",
            INIT_01 => X"fffffff6fffffffffffffffafffffffffffffffbffffffffffffffedffffffff",
            INIT_02 => X"ffffffe3fffffffffffffff5ffffffffffffffd0ffffffffffffffbdffffffff",
            INIT_03 => X"0000000e00000000ffffffeaffffffff0000000100000000fffffff2ffffffff",
            INIT_04 => X"fffffff4fffffffffffffff9ffffffff00000016000000000000000d00000000",
            INIT_05 => X"ffffffe6fffffffffffffffbffffffff0000000300000000fffffff0ffffffff",
            INIT_06 => X"00000000000000000000000600000000fffffffbffffffff0000001e00000000",
            INIT_07 => X"fffffffcffffffffffffffeefffffffffffffff0ffffffff0000002200000000",
            INIT_08 => X"0000000c00000000fffffff2ffffffffffffffe2ffffffff0000001200000000",
            INIT_09 => X"0000000e00000000fffffff0ffffffff0000000500000000ffffffedffffffff",
            INIT_0A => X"00000011000000000000000100000000fffffffbfffffffffffffff5ffffffff",
            INIT_0B => X"0000000e00000000ffffffdaffffffffffffffeefffffffffffffff4ffffffff",
            INIT_0C => X"00000004000000000000002e000000000000001800000000fffffffdffffffff",
            INIT_0D => X"ffffffeefffffffffffffffcffffffff0000001900000000fffffffaffffffff",
            INIT_0E => X"fffffff9ffffffff00000008000000000000003d000000000000001b00000000",
            INIT_0F => X"0000001300000000000000000000000000000008000000000000000300000000",
            INIT_10 => X"fffffffdffffffff0000001100000000ffffffd6ffffffff0000001d00000000",
            INIT_11 => X"fffffff5ffffffffffffffe8ffffffff0000000800000000fffffff1ffffffff",
            INIT_12 => X"00000021000000000000000600000000fffffff0ffffffffffffffe7ffffffff",
            INIT_13 => X"0000001200000000ffffffd8fffffffffffffff8fffffffffffffff9ffffffff",
            INIT_14 => X"fffffff2ffffffff0000001700000000ffffffddffffffff0000001900000000",
            INIT_15 => X"0000000600000000000000030000000000000016000000000000000000000000",
            INIT_16 => X"fffffffdffffffff0000000e00000000fffffff2fffffffffffffff8ffffffff",
            INIT_17 => X"0000001800000000ffffffebffffffffffffffe4fffffffffffffff3ffffffff",
            INIT_18 => X"ffffffe8ffffffff00000017000000000000000b00000000fffffffbffffffff",
            INIT_19 => X"0000000400000000fffffffdfffffffffffffffdffffffff0000000400000000",
            INIT_1A => X"fffffffdffffffff0000000700000000fffffff9ffffffff0000000f00000000",
            INIT_1B => X"0000000100000000ffffffe7fffffffffffffff2ffffffffffffffdfffffffff",
            INIT_1C => X"fffffff4ffffffff0000000f0000000000000023000000000000000c00000000",
            INIT_1D => X"0000001100000000000000030000000000000000000000000000000400000000",
            INIT_1E => X"00000013000000000000000e00000000fffffffbffffffffffffffe8ffffffff",
            INIT_1F => X"0000001700000000fffffff0ffffffffffffffebffffffff0000003000000000",
            INIT_20 => X"ffffffe4ffffffff00000046000000000000003000000000fffffff9ffffffff",
            INIT_21 => X"ffffffe8fffffffffffffff1ffffffff00000025000000000000002200000000",
            INIT_22 => X"0000000a00000000ffffffcaffffffff00000017000000000000000900000000",
            INIT_23 => X"0000000c000000000000001800000000fffffffaffffffff0000000900000000",
            INIT_24 => X"0000000b00000000fffffff6ffffffff0000001e00000000fffffffaffffffff",
            INIT_25 => X"0000001e000000000000002600000000ffffffeaffffffffffffffdeffffffff",
            INIT_26 => X"ffffffc6fffffffffffffff0ffffffff0000001f00000000fffffff5ffffffff",
            INIT_27 => X"0000000b00000000ffffffe8ffffffff0000001700000000ffffffe7ffffffff",
            INIT_28 => X"ffffffd0ffffffffffffffc6ffffffff0000001d000000000000000000000000",
            INIT_29 => X"0000000300000000ffffffe4ffffffffffffffe4ffffffff0000001e00000000",
            INIT_2A => X"0000000a00000000fffffff0fffffffffffffff9ffffffffffffffefffffffff",
            INIT_2B => X"fffffffeffffffff0000000c00000000ffffffeeffffffff0000000000000000",
            INIT_2C => X"0000000400000000fffffff7fffffffffffffff7ffffffff0000000300000000",
            INIT_2D => X"00000019000000000000000f00000000fffffff1ffffffffffffffe7ffffffff",
            INIT_2E => X"ffffffecffffffffffffffd0ffffffffffffffedffffffff0000001200000000",
            INIT_2F => X"fffffffbffffffff000000070000000000000028000000000000000500000000",
            INIT_30 => X"ffffffd7ffffffffffffffdeffffffff00000015000000000000000a00000000",
            INIT_31 => X"fffffff8ffffffff0000000500000000fffffffcfffffffffffffffcffffffff",
            INIT_32 => X"fffffff4ffffffffffffffefffffffff0000000600000000ffffffdaffffffff",
            INIT_33 => X"ffffffe4fffffffffffffffdffffffffffffffddffffffff0000000000000000",
            INIT_34 => X"0000003b00000000ffffffcfffffffffffffffefffffffff0000000100000000",
            INIT_35 => X"0000001a00000000fffffff1ffffffffffffffeefffffffffffffff7ffffffff",
            INIT_36 => X"fffffff2ffffffffffffffd4ffffffffffffffecffffffffffffffefffffffff",
            INIT_37 => X"fffffff1ffffffff0000001400000000fffffff4ffffffffffffffd1ffffffff",
            INIT_38 => X"ffffffdaffffffffffffffdcffffffff0000000100000000ffffffffffffffff",
            INIT_39 => X"0000000a0000000000000002000000000000000d00000000ffffffd8ffffffff",
            INIT_3A => X"ffffffe3ffffffff00000006000000000000000d00000000ffffffccffffffff",
            INIT_3B => X"fffffff3ffffffff0000001500000000fffffff7ffffffff0000001700000000",
            INIT_3C => X"00000027000000000000000000000000ffffffdcfffffffffffffff3ffffffff",
            INIT_3D => X"fffffffeffffffffffffffe1ffffffff0000001600000000ffffffe8ffffffff",
            INIT_3E => X"ffffffeaffffffffffffffd1ffffffff0000001a000000000000000300000000",
            INIT_3F => X"fffffffaffffffff0000000200000000ffffffe5fffffffffffffff0ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffd4ffffffffffffffc6ffffffff0000001d000000000000000300000000",
            INIT_41 => X"fffffffcffffffff00000007000000000000001300000000fffffff3ffffffff",
            INIT_42 => X"0000003d0000000000000003000000000000001800000000ffffffd1ffffffff",
            INIT_43 => X"0000000b00000000ffffffd1ffffffffffffffe7ffffffff0000001700000000",
            INIT_44 => X"0000002200000000ffffffebffffffffffffffeffffffffffffffff6ffffffff",
            INIT_45 => X"000000170000000000000001000000000000001900000000ffffffe7ffffffff",
            INIT_46 => X"ffffffeeffffffffffffffeffffffffffffffffaffffffff0000000c00000000",
            INIT_47 => X"0000000d0000000000000000000000000000000900000000fffffff6ffffffff",
            INIT_48 => X"ffffffb2ffffffffffffffb8ffffffff00000010000000000000000e00000000",
            INIT_49 => X"0000000b0000000000000003000000000000001100000000fffffff8ffffffff",
            INIT_4A => X"000000400000000000000011000000000000000000000000ffffffd2ffffffff",
            INIT_4B => X"ffffffedffffffffffffffd4ffffffffffffffe2ffffffff0000001600000000",
            INIT_4C => X"0000001f00000000fffffff2ffffffffffffffcefffffffffffffff6ffffffff",
            INIT_4D => X"ffffffe9ffffffff00000009000000000000000100000000ffffffebffffffff",
            INIT_4E => X"ffffffebffffffff00000014000000000000002500000000ffffffddffffffff",
            INIT_4F => X"0000000e000000000000000d000000000000000400000000ffffffd4ffffffff",
            INIT_50 => X"ffffffcfffffffffffffffe5ffffffffffffffd4ffffffffffffffffffffffff",
            INIT_51 => X"0000000100000000fffffff6ffffffff0000000f00000000fffffff0ffffffff",
            INIT_52 => X"00000028000000000000000400000000fffffffbffffffffffffffc6ffffffff",
            INIT_53 => X"ffffffeaffffffff0000000500000000ffffffd3ffffffff0000000600000000",
            INIT_54 => X"0000004600000000ffffffd6ffffffff0000001200000000ffffffdcffffffff",
            INIT_55 => X"ffffffecffffffff0000003400000000fffffff3ffffffff0000000b00000000",
            INIT_56 => X"fffffff4ffffffff0000000000000000ffffffbeffffffffffffffe0ffffffff",
            INIT_57 => X"000000210000000000000015000000000000002f00000000ffffffd6ffffffff",
            INIT_58 => X"ffffffe5ffffffff0000000a00000000ffffffdeffffffff0000000a00000000",
            INIT_59 => X"0000000200000000ffffffe2ffffffffffffffebffffffff0000000600000000",
            INIT_5A => X"ffffffffffffffff0000000800000000fffffffbfffffffffffffff7ffffffff",
            INIT_5B => X"00000014000000000000002a00000000ffffffe1fffffffffffffffcffffffff",
            INIT_5C => X"fffffff6ffffffff00000015000000000000001400000000fffffffaffffffff",
            INIT_5D => X"00000045000000000000000e0000000000000001000000000000000100000000",
            INIT_5E => X"ffffffd5fffffffffffffffbffffffffffffffc1ffffffffffffffe4ffffffff",
            INIT_5F => X"ffffffe9ffffffff00000003000000000000001d000000000000002f00000000",
            INIT_60 => X"ffffffcfffffffffffffffebffffffff0000001000000000ffffffffffffffff",
            INIT_61 => X"fffffff2fffffffffffffffefffffffffffffff6ffffffff0000000f00000000",
            INIT_62 => X"ffffffefffffffffffffffe6fffffffffffffff7fffffffffffffff4ffffffff",
            INIT_63 => X"00000012000000000000001d00000000fffffffafffffffffffffff1ffffffff",
            INIT_64 => X"fffffffdfffffffffffffff6ffffffff0000000d000000000000001000000000",
            INIT_65 => X"0000001500000000fffffffeffffffff00000022000000000000000000000000",
            INIT_66 => X"ffffffdfffffffffffffffdeffffffffffffffcbffffffffffffffefffffffff",
            INIT_67 => X"fffffff5ffffffffffffffffffffffffffffffe9fffffffffffffff7ffffffff",
            INIT_68 => X"ffffffbfffffffffffffffdcffffffff00000005000000000000000500000000",
            INIT_69 => X"fffffffcffffffff0000001200000000fffffffdfffffffffffffffaffffffff",
            INIT_6A => X"ffffffdefffffffffffffffeffffffff0000000900000000fffffffbffffffff",
            INIT_6B => X"ffffffdfffffffff0000001d0000000000000009000000000000000200000000",
            INIT_6C => X"0000000c00000000fffffff1ffffffffffffffddfffffffffffffffbffffffff",
            INIT_6D => X"fffffffcffffffffffffffefffffffff0000002b000000000000003000000000",
            INIT_6E => X"ffffffdeffffffffffffffddffffffffffffffd2ffffffff0000000a00000000",
            INIT_6F => X"000000060000000000000017000000000000000400000000ffffffd5ffffffff",
            INIT_70 => X"ffffffc4ffffffffffffffbbfffffffffffffff0ffffffff0000000d00000000",
            INIT_71 => X"00000000000000000000001e0000000000000014000000000000000000000000",
            INIT_72 => X"0000000700000000fffffff6ffffffff0000001200000000fffffff0ffffffff",
            INIT_73 => X"fffffff2fffffffffffffff6ffffffff00000003000000000000001900000000",
            INIT_74 => X"00000023000000000000000500000000ffffffbcffffffffffffffeeffffffff",
            INIT_75 => X"ffffffdfffffffffffffffd9ffffffff00000003000000000000003000000000",
            INIT_76 => X"0000000900000000ffffffeeffffffffffffffcefffffffffffffffeffffffff",
            INIT_77 => X"fffffffcffffffff0000000900000000ffffffd9fffffffffffffff1ffffffff",
            INIT_78 => X"ffffffd9ffffffffffffffaaffffffff0000000d000000000000001200000000",
            INIT_79 => X"fffffffbffffffff00000025000000000000000a00000000fffffff7ffffffff",
            INIT_7A => X"fffffffbffffffff000000110000000000000016000000000000000800000000",
            INIT_7B => X"ffffffe2ffffffffffffffe9ffffffffffffffecffffffff0000001d00000000",
            INIT_7C => X"0000002800000000fffffff0ffffffffffffff98ffffffffffffffe6ffffffff",
            INIT_7D => X"ffffffcdffffffffffffffedffffffff00000029000000000000002b00000000",
            INIT_7E => X"0000001300000000ffffffe9ffffffffffffffeaffffffffffffffc3ffffffff",
            INIT_7F => X"00000001000000000000000a00000000ffffffe2ffffffffffffffcaffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE12;


    MEM_IWGHT_LAYER2_INSTANCE13 : if BRAM_NAME = "iwght_layer2_instance13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffb7ffffffffffffffc6fffffffffffffff5ffffffff0000001100000000",
            INIT_01 => X"fffffff7ffffffff00000014000000000000000d00000000ffffffddffffffff",
            INIT_02 => X"0000002400000000000000100000000000000011000000000000000c00000000",
            INIT_03 => X"0000000100000000ffffffaafffffffffffffff2ffffffff0000000900000000",
            INIT_04 => X"00000010000000000000000a00000000ffffffeaffffffffffffffe1ffffffff",
            INIT_05 => X"ffffffe5ffffffffffffffefffffffff0000001b000000000000001700000000",
            INIT_06 => X"fffffff9ffffffff000000180000000000000015000000000000001300000000",
            INIT_07 => X"00000033000000000000001200000000ffffffebffffffffffffffffffffffff",
            INIT_08 => X"ffffffdfffffffffffffffbaffffffffffffffe9ffffffff0000000f00000000",
            INIT_09 => X"fffffff0ffffffff00000004000000000000000a00000000ffffffefffffffff",
            INIT_0A => X"000000220000000000000039000000000000001a00000000fffffffaffffffff",
            INIT_0B => X"fffffff4ffffffffffffffaefffffffffffffffbfffffffffffffff2ffffffff",
            INIT_0C => X"0000001f00000000fffffff3fffffffffffffff1fffffffffffffff6ffffffff",
            INIT_0D => X"fffffff4ffffffff0000000a0000000000000009000000000000000400000000",
            INIT_0E => X"ffffffe8ffffffff0000001d000000000000001c000000000000000a00000000",
            INIT_0F => X"0000001800000000fffffffaffffffff00000029000000000000000900000000",
            INIT_10 => X"ffffffd3fffffffffffffffefffffffffffffffdfffffffffffffff2ffffffff",
            INIT_11 => X"0000000200000000ffffffe3fffffffffffffff4ffffffffffffffedffffffff",
            INIT_12 => X"0000000d00000000ffffffe2fffffffffffffffaffffffffffffffddffffffff",
            INIT_13 => X"0000001e0000000000000014000000000000000a000000000000001100000000",
            INIT_14 => X"fffffff7ffffffff000000100000000000000000000000000000001a00000000",
            INIT_15 => X"0000001d00000000fffffff1ffffffff0000000000000000fffffff8ffffffff",
            INIT_16 => X"fffffffbffffffffffffffd3ffffffff00000044000000000000000700000000",
            INIT_17 => X"ffffffedfffffffffffffff3ffffffff00000020000000000000003800000000",
            INIT_18 => X"ffffffc6fffffffffffffffdfffffffffffffff3ffffffff0000000800000000",
            INIT_19 => X"fffffffaffffffff00000009000000000000001900000000fffffff3ffffffff",
            INIT_1A => X"ffffffefffffffffffffffecfffffffffffffff4ffffffffffffffdfffffffff",
            INIT_1B => X"0000000100000000000000380000000000000031000000000000000200000000",
            INIT_1C => X"ffffffe8fffffffffffffffeffffffff0000000f000000000000000d00000000",
            INIT_1D => X"ffffffdefffffffffffffff2ffffffff0000000c00000000fffffff2ffffffff",
            INIT_1E => X"fffffff2fffffffffffffff7ffffffff00000016000000000000000200000000",
            INIT_1F => X"fffffffdffffffff0000000a000000000000001b000000000000001100000000",
            INIT_20 => X"ffffffe8ffffffffffffffe3ffffffffffffffe9ffffffff0000000600000000",
            INIT_21 => X"0000000d00000000fffffff2ffffffff0000001500000000fffffffeffffffff",
            INIT_22 => X"fffffff5ffffffffffffffe0ffffffff0000000800000000fffffff4ffffffff",
            INIT_23 => X"00000005000000000000002b0000000000000011000000000000001b00000000",
            INIT_24 => X"00000009000000000000000200000000fffffff2ffffffff0000000600000000",
            INIT_25 => X"ffffffe4ffffffffffffffe0ffffffff0000001a000000000000001300000000",
            INIT_26 => X"0000001500000000ffffffd4ffffffffffffffb5fffffffffffffff6ffffffff",
            INIT_27 => X"fffffff0fffffffffffffff7ffffffffffffffeaffffffff0000000e00000000",
            INIT_28 => X"fffffff2ffffffffffffffdeffffffffffffffd8ffffffff0000000000000000",
            INIT_29 => X"fffffffefffffffffffffff9ffffffff00000001000000000000000c00000000",
            INIT_2A => X"fffffff2ffffffffffffffd6fffffffffffffff8ffffffff0000001200000000",
            INIT_2B => X"ffffffeefffffffffffffff2ffffffff00000008000000000000002e00000000",
            INIT_2C => X"ffffffe6ffffffff0000000000000000ffffffcaffffffff0000000900000000",
            INIT_2D => X"fffffff3fffffffffffffffefffffffffffffff8ffffffff0000001500000000",
            INIT_2E => X"0000002900000000ffffffecffffffff0000001300000000ffffffe9ffffffff",
            INIT_2F => X"fffffffeffffffff000000150000000000000005000000000000001000000000",
            INIT_30 => X"fffffffdfffffffffffffff6ffffffffffffffe5ffffffff0000000600000000",
            INIT_31 => X"0000001c000000000000000000000000ffffffe9fffffffffffffffdffffffff",
            INIT_32 => X"0000000c00000000ffffffffffffffff00000010000000000000001c00000000",
            INIT_33 => X"ffffffe1ffffffffffffffcaffffffff00000002000000000000002300000000",
            INIT_34 => X"fffffff8ffffffff0000002300000000ffffffbfffffffff0000000000000000",
            INIT_35 => X"fffffff5ffffffff0000001a00000000ffffffeaffffffff0000002700000000",
            INIT_36 => X"0000000a000000000000000500000000fffffff3fffffffffffffff2ffffffff",
            INIT_37 => X"0000000700000000fffffffeffffffff0000001900000000ffffffe4ffffffff",
            INIT_38 => X"ffffffe3ffffffffffffffafffffffffffffffe5ffffffff0000001400000000",
            INIT_39 => X"000000220000000000000002000000000000000f000000000000000b00000000",
            INIT_3A => X"00000020000000000000001a0000000000000000000000000000000900000000",
            INIT_3B => X"fffffff2ffffffffffffffe1ffffffff00000005000000000000001a00000000",
            INIT_3C => X"ffffffecffffffff000000150000000000000007000000000000001200000000",
            INIT_3D => X"fffffff2fffffffffffffff3ffffffffffffffecffffffff0000001300000000",
            INIT_3E => X"000000000000000000000003000000000000001400000000fffffff9ffffffff",
            INIT_3F => X"0000002b00000000fffffffaffffffff0000003800000000ffffffd3ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff4ffffffffffffffddffffffffffffffe4ffffffff0000000300000000",
            INIT_41 => X"000000080000000000000007000000000000000100000000ffffffeaffffffff",
            INIT_42 => X"0000000b000000000000000500000000fffffff8fffffffffffffffaffffffff",
            INIT_43 => X"ffffffffffffffffffffffb6ffffffffffffffecffffffff0000001e00000000",
            INIT_44 => X"ffffffeffffffffffffffff2ffffffffffffffebffffffff0000000300000000",
            INIT_45 => X"0000001a000000000000000c00000000fffffff0ffffffff0000000400000000",
            INIT_46 => X"00000008000000000000002f00000000fffffff1ffffffff0000000300000000",
            INIT_47 => X"0000000000000000fffffff7ffffffff00000015000000000000000300000000",
            INIT_48 => X"ffffffeaffffffffffffffceffffffffffffffeeffffffff0000000200000000",
            INIT_49 => X"ffffffe9ffffffff00000004000000000000001800000000ffffffceffffffff",
            INIT_4A => X"ffffffe7ffffffffffffffd7ffffffffffffffe4fffffffffffffff5ffffffff",
            INIT_4B => X"fffffff5ffffffffffffffffffffffffffffffe2ffffffff0000000f00000000",
            INIT_4C => X"ffffffe7ffffffff0000001400000000ffffffdaffffffff0000002b00000000",
            INIT_4D => X"0000001500000000fffffff1ffffffff00000004000000000000001f00000000",
            INIT_4E => X"ffffffe5ffffffff0000001e00000000fffffff4ffffffff0000001900000000",
            INIT_4F => X"fffffff0fffffffffffffff9ffffffff00000003000000000000003a00000000",
            INIT_50 => X"ffffffbffffffffffffffffdfffffffffffffff8fffffffffffffffeffffffff",
            INIT_51 => X"fffffff1ffffffff00000011000000000000003a00000000ffffffe1ffffffff",
            INIT_52 => X"fffffffbffffffff00000016000000000000000500000000ffffffffffffffff",
            INIT_53 => X"000000270000000000000022000000000000001500000000fffffff4ffffffff",
            INIT_54 => X"0000000c00000000000000230000000000000027000000000000001a00000000",
            INIT_55 => X"0000000300000000ffffffe9fffffffffffffff5fffffffffffffff6ffffffff",
            INIT_56 => X"00000010000000000000000800000000ffffffe8ffffffff0000001100000000",
            INIT_57 => X"ffffffe8fffffffffffffffeffffffffffffffe9ffffffff0000001f00000000",
            INIT_58 => X"ffffffe7ffffffff0000001100000000ffffffccffffffff0000001500000000",
            INIT_59 => X"0000000800000000ffffffe7ffffffff00000007000000000000000a00000000",
            INIT_5A => X"ffffffe8fffffffffffffffbfffffffffffffff6ffffffff0000000000000000",
            INIT_5B => X"fffffff9ffffffff0000001e000000000000001b00000000fffffff9ffffffff",
            INIT_5C => X"0000001900000000000000210000000000000035000000000000000900000000",
            INIT_5D => X"fffffffefffffffffffffff2ffffffffffffffd4ffffffff0000001f00000000",
            INIT_5E => X"0000002700000000fffffff8ffffffffffffffcdffffffff0000000400000000",
            INIT_5F => X"0000000f000000000000001d00000000ffffffffffffffff0000000a00000000",
            INIT_60 => X"fffffffaffffffff0000000e00000000ffffffe7ffffffff0000000900000000",
            INIT_61 => X"0000001900000000fffffff1ffffffffffffffd5ffffffff0000001c00000000",
            INIT_62 => X"00000015000000000000001700000000fffffff6fffffffffffffff4ffffffff",
            INIT_63 => X"fffffff0ffffffff00000002000000000000001000000000ffffffe5ffffffff",
            INIT_64 => X"fffffffbfffffffffffffff9ffffffff0000003c00000000fffffff8ffffffff",
            INIT_65 => X"fffffffbfffffffffffffff0ffffffffffffffd3ffffffffffffffd8ffffffff",
            INIT_66 => X"00000006000000000000000200000000ffffff9dfffffffffffffff0ffffffff",
            INIT_67 => X"ffffffe3ffffffff0000000d00000000ffffffebffffffffffffffadffffffff",
            INIT_68 => X"0000001b000000000000000f00000000ffffffddffffffffffffffffffffffff",
            INIT_69 => X"0000002200000000ffffffefffffffffffffff6dffffffff0000001100000000",
            INIT_6A => X"00000004000000000000001800000000ffffffe7ffffffffffffffe9ffffffff",
            INIT_6B => X"fffffff9fffffffffffffffeffffffff0000001000000000fffffffaffffffff",
            INIT_6C => X"ffffffffffffffff00000000000000000000000500000000ffffffedffffffff",
            INIT_6D => X"fffffff5ffffffff0000000f00000000ffffffcbfffffffffffffffaffffffff",
            INIT_6E => X"0000000b00000000ffffffefffffffffffffffc6ffffffff0000000500000000",
            INIT_6F => X"fffffffcffffffff0000000000000000fffffff4ffffffffffffffebffffffff",
            INIT_70 => X"fffffff9fffffffffffffffbffffffffffffffe3ffffffff0000000500000000",
            INIT_71 => X"00000021000000000000000a00000000ffffffceffffffff0000001900000000",
            INIT_72 => X"fffffffcfffffffffffffffcffffffff0000001000000000ffffffffffffffff",
            INIT_73 => X"0000000000000000ffffffebffffffff0000000200000000fffffff4ffffffff",
            INIT_74 => X"fffffffaffffffff0000002a0000000000000025000000000000002f00000000",
            INIT_75 => X"00000021000000000000000d00000000ffffffeaffffffffffffffffffffffff",
            INIT_76 => X"0000001600000000000000250000000000000011000000000000001700000000",
            INIT_77 => X"0000000000000000000000150000000000000011000000000000000e00000000",
            INIT_78 => X"fffffff7fffffffffffffff9fffffffffffffff7fffffffffffffffbffffffff",
            INIT_79 => X"0000002600000000fffffff7ffffffff0000000000000000ffffffffffffffff",
            INIT_7A => X"fffffff1ffffffff0000000300000000fffffff8ffffffffffffffebffffffff",
            INIT_7B => X"0000000700000000ffffffa7fffffffffffffff5ffffffff0000001a00000000",
            INIT_7C => X"ffffffefffffffff0000002600000000ffffffddffffffff0000001700000000",
            INIT_7D => X"0000004c000000000000001400000000fffffff0fffffffffffffffcffffffff",
            INIT_7E => X"0000001d000000000000003100000000ffffffedffffffff0000001900000000",
            INIT_7F => X"ffffffe4fffffffffffffffcffffffff0000000c000000000000002b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE13;


    MEM_IWGHT_LAYER2_INSTANCE14 : if BRAM_NAME = "iwght_layer2_instance14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffaefffffffffffffffbfffffffffffffffcffffffff0000001700000000",
            INIT_01 => X"fffffff5ffffffff00000001000000000000002b00000000ffffffecffffffff",
            INIT_02 => X"0000002500000000ffffffd5ffffffff0000000c00000000ffffffe9ffffffff",
            INIT_03 => X"0000000d00000000ffffffe7fffffffffffffffafffffffffffffffcffffffff",
            INIT_04 => X"0000000100000000fffffff8ffffffff0000001c000000000000000c00000000",
            INIT_05 => X"fffffff7ffffffff0000001500000000fffffff4ffffffff0000000f00000000",
            INIT_06 => X"fffffffeffffffff0000001b00000000fffffff3ffffffff0000000200000000",
            INIT_07 => X"ffffffeffffffffffffffffafffffffffffffff4ffffffff0000002400000000",
            INIT_08 => X"ffffffc8fffffffffffffff6ffffffffffffffeeffffffff0000001000000000",
            INIT_09 => X"fffffffaffffffff00000008000000000000001600000000ffffffdeffffffff",
            INIT_0A => X"000000110000000000000012000000000000000c00000000fffffffbffffffff",
            INIT_0B => X"0000000e00000000fffffff1ffffffff00000012000000000000000200000000",
            INIT_0C => X"00000000000000000000001200000000ffffffedffffffff0000001300000000",
            INIT_0D => X"0000000800000000ffffffeaffffffffffffffd0ffffffff0000002f00000000",
            INIT_0E => X"00000001000000000000002000000000ffffffd8ffffffff0000000000000000",
            INIT_0F => X"fffffffaffffffff0000000400000000ffffffdfffffffff0000000b00000000",
            INIT_10 => X"ffffffc2fffffffffffffffcffffffffffffffe6ffffffff0000002200000000",
            INIT_11 => X"000000220000000000000014000000000000000c00000000fffffffdffffffff",
            INIT_12 => X"fffffff6ffffffff0000001600000000fffffffbfffffffffffffff3ffffffff",
            INIT_13 => X"fffffff2fffffffffffffff9ffffffff0000000c00000000ffffffe4ffffffff",
            INIT_14 => X"000000120000000000000009000000000000003200000000fffffff9ffffffff",
            INIT_15 => X"0000000300000000fffffff2ffffffffffffffddffffffff0000002200000000",
            INIT_16 => X"0000001600000000fffffff5ffffffffffffffd2ffffffff0000002000000000",
            INIT_17 => X"ffffffe9ffffffff0000001900000000fffffffaffffffffffffffe7ffffffff",
            INIT_18 => X"ffffffc8ffffffff0000001b00000000fffffffffffffffffffffffeffffffff",
            INIT_19 => X"0000001c000000000000001e00000000fffffff2ffffffff0000001a00000000",
            INIT_1A => X"fffffff8ffffffff0000001e00000000ffffffceffffffff0000000300000000",
            INIT_1B => X"fffffff4ffffffff0000001500000000fffffff7ffffffffffffffdfffffffff",
            INIT_1C => X"0000002f000000000000000c000000000000001d00000000ffffffdcffffffff",
            INIT_1D => X"0000000a00000000ffffffd0ffffffffffffffdcffffffff0000001300000000",
            INIT_1E => X"0000002600000000ffffffebfffffffffffffffefffffffffffffff4ffffffff",
            INIT_1F => X"ffffffe7ffffffff0000001c00000000ffffffc5ffffffffffffffa6ffffffff",
            INIT_20 => X"fffffff6ffffffff000000500000000000000012000000000000000700000000",
            INIT_21 => X"00000016000000000000000e00000000ffffffb8ffffffff0000001300000000",
            INIT_22 => X"00000001000000000000001300000000ffffffa9ffffffffffffffc4ffffffff",
            INIT_23 => X"ffffffe6fffffffffffffff9ffffffff0000000700000000ffffffd8ffffffff",
            INIT_24 => X"000000330000000000000014000000000000001500000000ffffffe5ffffffff",
            INIT_25 => X"0000000300000000ffffffecffffffffffffffdbffffffff0000001400000000",
            INIT_26 => X"00000016000000000000000300000000ffffffebffffffff0000001a00000000",
            INIT_27 => X"fffffff5ffffffff0000001a00000000ffffffb7ffffffffffffffd2ffffffff",
            INIT_28 => X"ffffffebffffffff0000002a0000000000000010000000000000000600000000",
            INIT_29 => X"00000006000000000000001300000000ffffffc1ffffffff0000001400000000",
            INIT_2A => X"fffffff2fffffffffffffffcfffffffffffffff0ffffffffffffffcdffffffff",
            INIT_2B => X"0000000300000000ffffffd7ffffffff0000000800000000ffffffe8ffffffff",
            INIT_2C => X"0000000c0000000000000018000000000000001b00000000fffffff8ffffffff",
            INIT_2D => X"ffffffdbfffffffffffffff6fffffffffffffff6ffffffff0000001900000000",
            INIT_2E => X"00000010000000000000000700000000ffffffcfffffffff0000002500000000",
            INIT_2F => X"fffffffcffffffff0000000e00000000ffffffe4ffffffffffffffe7ffffffff",
            INIT_30 => X"ffffffefffffffffffffffd1ffffffffffffffe7ffffffff0000000400000000",
            INIT_31 => X"00000004000000000000001e00000000ffffffecfffffffffffffffeffffffff",
            INIT_32 => X"ffffffd1ffffffff000000010000000000000006000000000000000900000000",
            INIT_33 => X"0000000600000000ffffffedffffffff00000002000000000000000600000000",
            INIT_34 => X"0000002600000000ffffffe6fffffffffffffff3fffffffffffffffdffffffff",
            INIT_35 => X"0000000300000000fffffff8ffffffff00000031000000000000001000000000",
            INIT_36 => X"0000002900000000ffffffd2ffffffff0000000800000000fffffff6ffffffff",
            INIT_37 => X"fffffff0ffffffff0000000600000000ffffffe1ffffffff0000001a00000000",
            INIT_38 => X"fffffff1fffffffffffffff7fffffffffffffffaffffffff0000000100000000",
            INIT_39 => X"0000000700000000fffffff6ffffffff0000002200000000ffffffe8ffffffff",
            INIT_3A => X"fffffff6ffffffff00000020000000000000001000000000ffffffeaffffffff",
            INIT_3B => X"0000000600000000ffffffc7fffffffffffffff0ffffffff0000000d00000000",
            INIT_3C => X"0000000000000000fffffffcffffffff00000025000000000000000d00000000",
            INIT_3D => X"ffffffe5ffffffff0000002c00000000fffffff4ffffffff0000002100000000",
            INIT_3E => X"ffffffdfffffffff0000002300000000fffffff0ffffffffffffffe2ffffffff",
            INIT_3F => X"fffffffeffffffff000000180000000000000006000000000000001000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffd5ffffffffffffffebffffffffffffffe5ffffffff0000000300000000",
            INIT_41 => X"0000001200000000fffffff8ffffffff0000001e00000000fffffff0ffffffff",
            INIT_42 => X"0000001b000000000000004000000000fffffff7ffffffff0000001100000000",
            INIT_43 => X"ffffffffffffffffffffffc5ffffffff00000007000000000000000800000000",
            INIT_44 => X"00000021000000000000000a0000000000000011000000000000000000000000",
            INIT_45 => X"0000000500000000fffffff2ffffffffffffffe6ffffffff0000001400000000",
            INIT_46 => X"fffffff9ffffffff00000025000000000000001100000000ffffffe5ffffffff",
            INIT_47 => X"0000000b000000000000002800000000ffffffe1ffffffff0000000200000000",
            INIT_48 => X"ffffffbeffffffffffffffd5fffffffffffffff9ffffffff0000001700000000",
            INIT_49 => X"0000001700000000fffffffbffffffff0000001d00000000ffffffecffffffff",
            INIT_4A => X"00000005000000000000001900000000fffffff9ffffffff0000001400000000",
            INIT_4B => X"0000002200000000ffffffd6ffffffff0000000400000000ffffffeeffffffff",
            INIT_4C => X"0000003a0000000000000007000000000000001c000000000000001c00000000",
            INIT_4D => X"0000000600000000fffffff8fffffffffffffffeffffffff0000003d00000000",
            INIT_4E => X"fffffffeffffffff00000010000000000000001800000000fffffff8ffffffff",
            INIT_4F => X"0000000100000000ffffffffffffffffffffffd2fffffffffffffff2ffffffff",
            INIT_50 => X"ffffffb8ffffffff0000000600000000fffffffdffffffff0000000000000000",
            INIT_51 => X"000000080000000000000018000000000000004100000000ffffffeaffffffff",
            INIT_52 => X"fffffff1ffffffff00000046000000000000000000000000fffffff3ffffffff",
            INIT_53 => X"0000001400000000fffffff7fffffffffffffff4ffffffffffffffedffffffff",
            INIT_54 => X"0000004500000000fffffff2ffffffff0000000e000000000000000100000000",
            INIT_55 => X"0000001100000000ffffffe4ffffffffffffffdbffffffff0000002b00000000",
            INIT_56 => X"fffffffeffffffffffffffd7ffffffffffffffe2ffffffff0000000400000000",
            INIT_57 => X"ffffffecffffffff0000000e00000000ffffff98ffffffffffffffe2ffffffff",
            INIT_58 => X"ffffffcfffffffff000000050000000000000009000000000000001c00000000",
            INIT_59 => X"fffffffbffffffff00000023000000000000000600000000fffffff4ffffffff",
            INIT_5A => X"fffffff1ffffffff0000001a00000000fffffff9ffffffffffffffe1ffffffff",
            INIT_5B => X"0000000900000000ffffffeeffffffffffffffe9ffffffffffffffe9ffffffff",
            INIT_5C => X"00000047000000000000001500000000fffffff2fffffffffffffff4ffffffff",
            INIT_5D => X"0000002000000000ffffffcefffffffffffffffbffffffff0000002c00000000",
            INIT_5E => X"00000012000000000000000600000000ffffffb2ffffffff0000000d00000000",
            INIT_5F => X"fffffffbffffffff0000000400000000ffffffc4ffffffffffffffeeffffffff",
            INIT_60 => X"ffffffe8ffffffff00000008000000000000001f000000000000000000000000",
            INIT_61 => X"00000000000000000000000d000000000000002200000000ffffffe6ffffffff",
            INIT_62 => X"ffffffc4ffffffff00000017000000000000000b00000000ffffffdaffffffff",
            INIT_63 => X"0000000400000000fffffffbffffffff0000000d00000000ffffffedffffffff",
            INIT_64 => X"0000002800000000ffffffebffffffff0000003c000000000000000a00000000",
            INIT_65 => X"0000001b00000000000000000000000000000027000000000000002100000000",
            INIT_66 => X"fffffff6fffffffffffffff5ffffffffffffffdcfffffffffffffff9ffffffff",
            INIT_67 => X"00000023000000000000001300000000ffffffe7ffffffffffffffd8ffffffff",
            INIT_68 => X"ffffffcdfffffffffffffff0fffffffffffffff7ffffffff0000000000000000",
            INIT_69 => X"fffffff8ffffffff00000002000000000000001100000000fffffff5ffffffff",
            INIT_6A => X"ffffffbfffffffffffffffe8ffffffff0000000800000000fffffff1ffffffff",
            INIT_6B => X"000000040000000000000031000000000000000c000000000000000b00000000",
            INIT_6C => X"000000360000000000000000000000000000000800000000fffffff5ffffffff",
            INIT_6D => X"0000000000000000ffffffffffffffff0000001400000000fffffff8ffffffff",
            INIT_6E => X"fffffffcffffffffffffffceffffffffffffffb5fffffffffffffff5ffffffff",
            INIT_6F => X"fffffff9ffffffff0000000d00000000ffffffe7fffffffffffffff9ffffffff",
            INIT_70 => X"ffffff94ffffffff0000000800000000ffffffe3ffffffff0000000100000000",
            INIT_71 => X"0000000000000000fffffffaffffffff0000000d000000000000000500000000",
            INIT_72 => X"00000033000000000000000b00000000fffffff0ffffffff0000001600000000",
            INIT_73 => X"fffffff9ffffffffffffffd9ffffffff00000009000000000000002600000000",
            INIT_74 => X"ffffffffffffffffffffffedffffffff0000000a00000000ffffffffffffffff",
            INIT_75 => X"ffffffe9ffffffff0000001f00000000ffffffc8fffffffffffffffcffffffff",
            INIT_76 => X"ffffffd0ffffffff0000004f00000000ffffffbdffffffff0000000900000000",
            INIT_77 => X"00000005000000000000001d000000000000001d000000000000000400000000",
            INIT_78 => X"ffffffbcfffffffffffffffafffffffffffffff3ffffffff0000000a00000000",
            INIT_79 => X"0000002200000000fffffffcffffffffffffffffffffffff0000001c00000000",
            INIT_7A => X"00000014000000000000000300000000ffffffffffffffff0000000d00000000",
            INIT_7B => X"fffffffbffffffffffffffbdffffffff00000023000000000000002d00000000",
            INIT_7C => X"0000001e00000000fffffff0ffffffff0000001600000000ffffffe2ffffffff",
            INIT_7D => X"ffffffdffffffffffffffff7fffffffffffffff1ffffffffffffffffffffffff",
            INIT_7E => X"ffffffe1ffffffffffffffeafffffffffffffff9ffffffffffffffebffffffff",
            INIT_7F => X"0000000b000000000000001000000000fffffffbffffffff0000000c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE14;


    MEM_IWGHT_LAYER2_INSTANCE15 : if BRAM_NAME = "iwght_layer2_instance15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffc3fffffffffffffffefffffffffffffff4ffffffff0000002500000000",
            INIT_01 => X"0000001e00000000ffffffecffffffff0000001900000000ffffffcfffffffff",
            INIT_02 => X"ffffffe3ffffffff0000001400000000ffffffd2fffffffffffffffeffffffff",
            INIT_03 => X"fffffff8ffffffffffffffacffffffff00000002000000000000001f00000000",
            INIT_04 => X"0000003700000000ffffffd5fffffffffffffff5ffffffffffffffe7ffffffff",
            INIT_05 => X"0000000f000000000000000200000000ffffffe2ffffffff0000000a00000000",
            INIT_06 => X"ffffffeafffffffffffffffdfffffffffffffff7ffffffff0000000000000000",
            INIT_07 => X"fffffffbffffffff0000002400000000ffffffe9ffffffff0000000b00000000",
            INIT_08 => X"ffffffcbffffffff00000008000000000000000e000000000000001a00000000",
            INIT_09 => X"0000002a000000000000000a000000000000001600000000ffffffe0ffffffff",
            INIT_0A => X"ffffffffffffffff0000001a000000000000000a00000000fffffff0ffffffff",
            INIT_0B => X"0000001800000000ffffffeaffffffff00000004000000000000000d00000000",
            INIT_0C => X"0000005000000000ffffffcbffffffffffffffe5ffffffffffffffd6ffffffff",
            INIT_0D => X"0000001100000000fffffff3fffffffffffffffefffffffffffffffeffffffff",
            INIT_0E => X"ffffffffffffffffffffffe1fffffffffffffffbffffffffffffffecffffffff",
            INIT_0F => X"fffffff3ffffffff0000002900000000ffffffddffffffffffffffe2ffffffff",
            INIT_10 => X"ffffffcaffffffffffffffe2fffffffffffffff7ffffffff0000000c00000000",
            INIT_11 => X"000000040000000000000024000000000000000700000000ffffffebffffffff",
            INIT_12 => X"ffffffd0ffffffff0000001000000000ffffffe8ffffffff0000001400000000",
            INIT_13 => X"ffffffedfffffffffffffff5ffffffff00000015000000000000001500000000",
            INIT_14 => X"0000002800000000ffffffe2ffffffffffffffe0ffffffffffffffe9ffffffff",
            INIT_15 => X"fffffff8ffffffffffffffe7fffffffffffffffaffffffff0000001100000000",
            INIT_16 => X"0000000400000000ffffffefffffffff0000001400000000fffffff5ffffffff",
            INIT_17 => X"fffffffaffffffff0000001100000000ffffffebffffffffffffffe1ffffffff",
            INIT_18 => X"ffffffb8ffffffffffffffe2ffffffff0000003b000000000000001b00000000",
            INIT_19 => X"0000000100000000fffffffcffffffff0000001f00000000ffffffd1ffffffff",
            INIT_1A => X"ffffffd0ffffffff0000000700000000fffffff1fffffffffffffff6ffffffff",
            INIT_1B => X"fffffffffffffffffffffffbffffffff0000000d000000000000001f00000000",
            INIT_1C => X"0000001b00000000ffffffd7ffffffff0000000e00000000fffffffdffffffff",
            INIT_1D => X"ffffffe5ffffffffffffffedfffffffffffffffcffffffff0000000500000000",
            INIT_1E => X"fffffff9ffffffffffffffe8ffffffffffffff8cffffffff0000000e00000000",
            INIT_1F => X"ffffffeeffffffff0000002200000000ffffffe1fffffffffffffffeffffffff",
            INIT_20 => X"ffffffeaffffffffffffffc2fffffffffffffffaffffffff0000000c00000000",
            INIT_21 => X"0000001200000000000000000000000000000000000000000000000f00000000",
            INIT_22 => X"ffffffdfffffffff0000001700000000ffffffd9fffffffffffffffbffffffff",
            INIT_23 => X"fffffff4ffffffff000000080000000000000020000000000000001a00000000",
            INIT_24 => X"0000002000000000ffffffd9fffffffffffffff0ffffffffffffffb5ffffffff",
            INIT_25 => X"0000002f00000000fffffff6ffffffff00000033000000000000000000000000",
            INIT_26 => X"ffffffefffffffff0000000400000000ffffffe2ffffffff0000001f00000000",
            INIT_27 => X"0000000d000000000000001f00000000fffffff9ffffffff0000000e00000000",
            INIT_28 => X"ffffffd6ffffffffffffffcaffffffffffffffc5ffffffff0000000f00000000",
            INIT_29 => X"0000000800000000ffffffe3ffffffffffffffefffffffff0000002b00000000",
            INIT_2A => X"0000001e000000000000004a00000000ffffffe9ffffffff0000002400000000",
            INIT_2B => X"ffffffb9ffffffffffffffc3ffffffffffffffceffffffff0000001000000000",
            INIT_2C => X"0000000f00000000ffffffceffffffff0000000400000000ffffffbeffffffff",
            INIT_2D => X"ffffffd2ffffffffffffffdbffffffff0000000b000000000000000000000000",
            INIT_2E => X"00000039000000000000001300000000fffffff0ffffffffffffffe4ffffffff",
            INIT_2F => X"00000017000000000000000a00000000ffffffccffffffff0000002300000000",
            INIT_30 => X"ffffffdfffffffff00000027000000000000000a000000000000001f00000000",
            INIT_31 => X"00000007000000000000001800000000ffffffedffffffffffffffebffffffff",
            INIT_32 => X"0000001a000000000000001e00000000fffffff4ffffffffffffffe5ffffffff",
            INIT_33 => X"ffffffeaffffffffffffffb9ffffffffffffffeeffffffff0000000800000000",
            INIT_34 => X"ffffffcefffffffffffffffbffffffff0000001c00000000ffffffdfffffffff",
            INIT_35 => X"ffffffd5ffffffff00000000000000000000001300000000fffffff2ffffffff",
            INIT_36 => X"00000001000000000000002e00000000fffffff4ffffffffffffffd6ffffffff",
            INIT_37 => X"0000002200000000ffffffeeffffffff00000000000000000000000400000000",
            INIT_38 => X"0000001e00000000000000090000000000000000000000000000000600000000",
            INIT_39 => X"fffffff6ffffffffffffffffffffffffffffffddffffffff0000002800000000",
            INIT_3A => X"00000016000000000000002700000000fffffff5ffffffff0000000b00000000",
            INIT_3B => X"0000000600000000ffffffd8ffffffff0000000e00000000fffffffeffffffff",
            INIT_3C => X"00000000000000000000002000000000fffffff1fffffffffffffffeffffffff",
            INIT_3D => X"0000000100000000fffffff7ffffffffffffffe3ffffffffffffffeeffffffff",
            INIT_3E => X"fffffffdffffffff0000002700000000ffffffa0ffffffffffffffc6ffffffff",
            INIT_3F => X"000000250000000000000005000000000000000600000000ffffffe9ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000031000000000000001a0000000000000005000000000000000200000000",
            INIT_41 => X"fffffffafffffffffffffff1fffffffffffffffcffffffff0000000200000000",
            INIT_42 => X"0000000900000000fffffff2fffffffffffffffaffffffff0000000a00000000",
            INIT_43 => X"0000002a00000000fffffff2ffffffff0000002e000000000000000b00000000",
            INIT_44 => X"ffffffc7ffffffff000000060000000000000021000000000000001e00000000",
            INIT_45 => X"ffffffd9ffffffff0000003900000000ffffffdafffffffffffffffeffffffff",
            INIT_46 => X"00000022000000000000001700000000ffffffacffffffffffffffe5ffffffff",
            INIT_47 => X"0000000f00000000000000080000000000000008000000000000000e00000000",
            INIT_48 => X"00000029000000000000002800000000ffffffffffffffff0000001200000000",
            INIT_49 => X"fffffff3ffffffff0000000700000000ffffffffffffffff0000000400000000",
            INIT_4A => X"fffffff7ffffffffffffffe0ffffffff0000000f00000000ffffffebffffffff",
            INIT_4B => X"0000003300000000fffffff5ffffffff0000003c00000000fffffffcffffffff",
            INIT_4C => X"ffffffe9ffffffffffffffebffffffff00000028000000000000000700000000",
            INIT_4D => X"ffffffeeffffffffffffffeafffffffffffffff8ffffffff0000000900000000",
            INIT_4E => X"0000000700000000ffffffdcfffffffffffffffbffffffff0000000100000000",
            INIT_4F => X"ffffffffffffffff0000000d00000000ffffffdeffffffff0000000400000000",
            INIT_50 => X"fffffffaffffffff0000003900000000fffffff9fffffffffffffff7ffffffff",
            INIT_51 => X"0000000000000000fffffff8ffffffffffffffedffffffff0000000600000000",
            INIT_52 => X"0000000c000000000000000a00000000ffffffeeffffffff0000000e00000000",
            INIT_53 => X"000000210000000000000034000000000000000600000000fffffffaffffffff",
            INIT_54 => X"fffffff0ffffffffffffffedffffffff0000003b000000000000001000000000",
            INIT_55 => X"ffffffedffffffff0000000a0000000000000000000000000000000400000000",
            INIT_56 => X"0000001d00000000fffffff2fffffffffffffff8ffffffff0000000a00000000",
            INIT_57 => X"ffffffe8ffffffff0000000300000000fffffff5ffffffff0000003800000000",
            INIT_58 => X"0000000b000000000000003f000000000000000300000000fffffff6ffffffff",
            INIT_59 => X"ffffffdbffffffffffffffe1fffffffffffffff4ffffffff0000002900000000",
            INIT_5A => X"ffffffd0ffffffff0000002800000000ffffffcfffffffff0000000d00000000",
            INIT_5B => X"fffffffeffffffff0000000c00000000fffffffaffffffff0000001e00000000",
            INIT_5C => X"ffffffe7ffffffffffffffdbffffffff0000003200000000fffffff9ffffffff",
            INIT_5D => X"00000026000000000000000d00000000ffffffd3ffffffff0000000000000000",
            INIT_5E => X"0000003700000000ffffffffffffffffffffffd2ffffffff0000001300000000",
            INIT_5F => X"fffffff0ffffffff0000001100000000ffffffeeffffffff0000002f00000000",
            INIT_60 => X"fffffff5ffffffff0000003200000000fffffff8ffffffff0000000400000000",
            INIT_61 => X"ffffffeefffffffffffffffcffffffff00000003000000000000000500000000",
            INIT_62 => X"0000001f000000000000003500000000ffffffdbffffffff0000001100000000",
            INIT_63 => X"ffffffe8ffffffffffffffcbffffffff00000002000000000000000000000000",
            INIT_64 => X"fffffff3ffffffffffffffe2ffffffffffffffceffffffffffffffe6ffffffff",
            INIT_65 => X"ffffffddffffffffffffffccffffffff0000000000000000ffffffebffffffff",
            INIT_66 => X"00000016000000000000000100000000fffffff4fffffffffffffffeffffffff",
            INIT_67 => X"0000000400000000ffffffdbffffffffffffffd5ffffffff0000001700000000",
            INIT_68 => X"000000070000000000000012000000000000001200000000fffffff2ffffffff",
            INIT_69 => X"ffffffdaffffffff0000000000000000fffffff5ffffffff0000001900000000",
            INIT_6A => X"00000022000000000000000f00000000fffffffbffffffffffffffdfffffffff",
            INIT_6B => X"ffffffddffffffffffffffdaffffffffffffffedffffffffffffffebffffffff",
            INIT_6C => X"0000000100000000fffffff5ffffffffffffffe8ffffffffffffffe8ffffffff",
            INIT_6D => X"00000014000000000000000d00000000ffffffe3fffffffffffffffbffffffff",
            INIT_6E => X"ffffffdbffffffff0000002000000000ffffffa8ffffffffffffffdcffffffff",
            INIT_6F => X"0000001400000000ffffffecffffffffffffffdeffffffffffffffedffffffff",
            INIT_70 => X"000000140000000000000023000000000000001c00000000fffffffdffffffff",
            INIT_71 => X"0000001200000000ffffffedffffffffffffffe8ffffffff0000000000000000",
            INIT_72 => X"0000001700000000fffffffaffffffff0000000500000000ffffffedffffffff",
            INIT_73 => X"0000001e00000000ffffffe1ffffffff0000000e00000000fffffff4ffffffff",
            INIT_74 => X"00000007000000000000000d000000000000001f00000000fffffffeffffffff",
            INIT_75 => X"0000001b000000000000001300000000fffffff3ffffffff0000000500000000",
            INIT_76 => X"00000002000000000000002c00000000ffffff95ffffffffffffffabffffffff",
            INIT_77 => X"0000000200000000fffffff9ffffffffffffffe6fffffffffffffffdffffffff",
            INIT_78 => X"000000290000000000000008000000000000001e000000000000000500000000",
            INIT_79 => X"0000003400000000ffffffd6ffffffffffffffe4ffffffff0000000300000000",
            INIT_7A => X"0000001900000000fffffffafffffffffffffffdfffffffffffffffcffffffff",
            INIT_7B => X"0000001e00000000fffffff0fffffffffffffffdffffffff0000000400000000",
            INIT_7C => X"fffffff9ffffffff000000200000000000000012000000000000001400000000",
            INIT_7D => X"00000035000000000000001200000000fffffff0ffffffff0000001000000000",
            INIT_7E => X"fffffff7ffffffff00000025000000000000000800000000ffffffa5ffffffff",
            INIT_7F => X"00000012000000000000000300000000fffffff3ffffffffffffffdfffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE15;


    MEM_IWGHT_LAYER2_INSTANCE16 : if BRAM_NAME = "iwght_layer2_instance16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000d0000000000000015000000000000001200000000fffffff4ffffffff",
            INIT_01 => X"0000001000000000ffffffd6ffffffffffffffeeffffffff0000001300000000",
            INIT_02 => X"fffffff0ffffffffffffffe3ffffffff0000000c00000000fffffffbffffffff",
            INIT_03 => X"00000019000000000000001f000000000000001a000000000000001500000000",
            INIT_04 => X"0000000000000000000000130000000000000007000000000000001b00000000",
            INIT_05 => X"0000000400000000000000180000000000000016000000000000001b00000000",
            INIT_06 => X"fffffff2ffffffff0000001a000000000000001300000000ffffffd4ffffffff",
            INIT_07 => X"00000010000000000000000900000000fffffffbffffffff0000000700000000",
            INIT_08 => X"fffffffdffffffff0000002d000000000000000300000000fffffff0ffffffff",
            INIT_09 => X"0000001b00000000fffffff5ffffffff0000000d000000000000001700000000",
            INIT_0A => X"ffffffeefffffffffffffff6ffffffffffffffebffffffff0000002400000000",
            INIT_0B => X"0000001f00000000000000230000000000000004000000000000000100000000",
            INIT_0C => X"fffffffaffffffff000000120000000000000031000000000000002100000000",
            INIT_0D => X"00000037000000000000000d00000000fffffffdffffffff0000000000000000",
            INIT_0E => X"0000000300000000ffffffd9ffffffffffffffdbfffffffffffffff0ffffffff",
            INIT_0F => X"0000000600000000fffffff0ffffffffffffffdcffffffff0000000000000000",
            INIT_10 => X"000000090000000000000019000000000000000d00000000fffffffeffffffff",
            INIT_11 => X"ffffffefffffffffffffffeeffffffffffffffebffffffff0000000b00000000",
            INIT_12 => X"ffffffeaffffffff0000000600000000ffffffc4fffffffffffffffeffffffff",
            INIT_13 => X"fffffff5ffffffff0000000e00000000fffffff8ffffffff0000000100000000",
            INIT_14 => X"000000000000000000000004000000000000000b00000000fffffffaffffffff",
            INIT_15 => X"fffffffafffffffffffffffcffffffff0000001c000000000000000400000000",
            INIT_16 => X"0000000900000000ffffffc8ffffffffffffffd3fffffffffffffff6ffffffff",
            INIT_17 => X"ffffffeffffffffffffffff7ffffffffffffffccffffffff0000003000000000",
            INIT_18 => X"ffffffffffffffff0000002c0000000000000012000000000000000000000000",
            INIT_19 => X"fffffff6ffffffff0000001a0000000000000008000000000000000700000000",
            INIT_1A => X"00000000000000000000001800000000fffffff5ffffffffffffffdeffffffff",
            INIT_1B => X"ffffffd4ffffffffffffffccfffffffffffffff0ffffffff0000001d00000000",
            INIT_1C => X"0000000100000000fffffff1ffffffffffffffd3fffffffffffffffaffffffff",
            INIT_1D => X"0000000300000000ffffffc2ffffffff00000004000000000000000100000000",
            INIT_1E => X"0000003400000000fffffff6ffffffffffffffd0ffffffff0000002c00000000",
            INIT_1F => X"ffffffeaffffffffffffffe4ffffffffffffffb7fffffffffffffff8ffffffff",
            INIT_20 => X"00000012000000000000002300000000fffffff7ffffffff0000000900000000",
            INIT_21 => X"00000004000000000000000800000000fffffff9ffffffff0000000100000000",
            INIT_22 => X"0000001300000000000000090000000000000018000000000000002300000000",
            INIT_23 => X"ffffffe8ffffffffffffffd3ffffffffffffffddffffffff0000000a00000000",
            INIT_24 => X"0000000f00000000fffffffbffffffffffffffebffffffff0000000000000000",
            INIT_25 => X"fffffffcffffffffffffffe3ffffffffffffffd6ffffffff0000000800000000",
            INIT_26 => X"0000000d00000000ffffffe6ffffffffffffffd7ffffffffffffffd8ffffffff",
            INIT_27 => X"fffffffdffffffff0000000d00000000ffffffc2ffffffffffffffcfffffffff",
            INIT_28 => X"ffffffe7ffffffff000000100000000000000025000000000000000700000000",
            INIT_29 => X"0000000100000000fffffffafffffffffffffff0ffffffffffffffe5ffffffff",
            INIT_2A => X"00000015000000000000001300000000fffffffdfffffffffffffff5ffffffff",
            INIT_2B => X"ffffffffffffffff0000001100000000ffffffceffffffffffffffcfffffffff",
            INIT_2C => X"0000001e00000000fffffffaffffffffffffffeefffffffffffffffaffffffff",
            INIT_2D => X"00000010000000000000000700000000ffffffc2ffffffff0000000200000000",
            INIT_2E => X"ffffffd8ffffffff00000006000000000000000e00000000ffffffc3ffffffff",
            INIT_2F => X"000000110000000000000009000000000000000500000000ffffffebffffffff",
            INIT_30 => X"000000110000000000000002000000000000002600000000fffffff8ffffffff",
            INIT_31 => X"0000001c00000000ffffffedffffffffffffffedffffffffffffffeaffffffff",
            INIT_32 => X"0000002a00000000fffffffdffffffff0000001400000000ffffffe2ffffffff",
            INIT_33 => X"00000000000000000000002900000000ffffffdbffffffffffffffc2ffffffff",
            INIT_34 => X"0000002800000000ffffffd6ffffffffffffffe6fffffffffffffffaffffffff",
            INIT_35 => X"0000000e000000000000001700000000ffffffdcffffffffffffffedffffffff",
            INIT_36 => X"ffffffd3ffffffffffffffeaffffffff0000001d00000000ffffffa1ffffffff",
            INIT_37 => X"0000000e000000000000000e000000000000001000000000ffffffcfffffffff",
            INIT_38 => X"ffffffdbffffffff00000008000000000000002700000000ffffffefffffffff",
            INIT_39 => X"fffffffdfffffffffffffffaffffffffffffffd1ffffffff0000000500000000",
            INIT_3A => X"fffffffeffffffff0000001400000000ffffffd4fffffffffffffff5ffffffff",
            INIT_3B => X"00000019000000000000000c00000000ffffffe9ffffffffffffffe5ffffffff",
            INIT_3C => X"00000013000000000000000e000000000000000b00000000fffffffaffffffff",
            INIT_3D => X"0000003d00000000fffffff8fffffffffffffff9fffffffffffffff2ffffffff",
            INIT_3E => X"ffffffb6fffffffffffffff7ffffffff0000000800000000ffffffbdffffffff",
            INIT_3F => X"fffffffcfffffffffffffff5fffffffffffffff2ffffffffffffffd3ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001e00000000fffffff4ffffffff0000001e000000000000000300000000",
            INIT_41 => X"0000000000000000ffffffd0fffffffffffffff1fffffffffffffff2ffffffff",
            INIT_42 => X"ffffffe9ffffffff0000001a00000000ffffffd0ffffffff0000001100000000",
            INIT_43 => X"00000001000000000000002d000000000000000600000000ffffffe8ffffffff",
            INIT_44 => X"0000001d00000000fffffffdffffffffffffffd6ffffffff0000000b00000000",
            INIT_45 => X"0000001100000000ffffffe8ffffffff0000000a000000000000000000000000",
            INIT_46 => X"fffffffeffffffffffffffaeffffffffffffffdbffffffffffffffedffffffff",
            INIT_47 => X"ffffffdeffffffff0000001200000000fffffff5ffffffffffffffefffffffff",
            INIT_48 => X"ffffffffffffffff00000020000000000000001f000000000000000000000000",
            INIT_49 => X"0000001f00000000fffffffdffffffffffffffd8fffffffffffffff4ffffffff",
            INIT_4A => X"ffffffd4ffffffff0000003900000000ffffffe8ffffffffffffffecffffffff",
            INIT_4B => X"000000000000000000000018000000000000000e00000000fffffffdffffffff",
            INIT_4C => X"fffffffdffffffff0000000500000000ffffffe2fffffffffffffffbffffffff",
            INIT_4D => X"fffffff2fffffffffffffff0fffffffffffffff4ffffffffffffffeaffffffff",
            INIT_4E => X"00000028000000000000001b00000000ffffffb4ffffffff0000001c00000000",
            INIT_4F => X"ffffffe8ffffffff0000000800000000fffffff1ffffffff0000000700000000",
            INIT_50 => X"0000000f00000000000000210000000000000014000000000000000500000000",
            INIT_51 => X"0000001c000000000000001a000000000000000200000000fffffffdffffffff",
            INIT_52 => X"ffffffe8ffffffff00000025000000000000000100000000ffffffefffffffff",
            INIT_53 => X"ffffffdcffffffffffffffeeffffffff00000005000000000000000b00000000",
            INIT_54 => X"0000000600000000fffffffbffffffff00000002000000000000000800000000",
            INIT_55 => X"fffffff8ffffffffffffffadfffffffffffffffcfffffffffffffffbffffffff",
            INIT_56 => X"0000003500000000ffffffe6fffffffffffffff9fffffffffffffff9ffffffff",
            INIT_57 => X"fffffff7ffffffffffffffedffffffffffffffd7ffffffff0000000000000000",
            INIT_58 => X"0000001c000000000000002300000000fffffff4fffffffffffffff1ffffffff",
            INIT_59 => X"fffffff1ffffffff0000001600000000fffffff8ffffffffffffffdcffffffff",
            INIT_5A => X"fffffffaffffffff0000001d00000000fffffffaffffffff0000002500000000",
            INIT_5B => X"0000000600000000ffffffe9ffffffff0000000a00000000ffffffeeffffffff",
            INIT_5C => X"00000010000000000000000d000000000000000200000000ffffffe1ffffffff",
            INIT_5D => X"0000002500000000fffffff5fffffffffffffffcfffffffffffffffaffffffff",
            INIT_5E => X"0000000000000000ffffffeaffffffffffffffb8ffffffff0000000000000000",
            INIT_5F => X"0000000100000000ffffffe0ffffffffffffffddffffffffffffffceffffffff",
            INIT_60 => X"0000000c000000000000002f000000000000000400000000fffffffdffffffff",
            INIT_61 => X"fffffff2ffffffff0000000600000000ffffffe6ffffffffffffffe0ffffffff",
            INIT_62 => X"0000000e000000000000000400000000fffffff0ffffffffffffffd8ffffffff",
            INIT_63 => X"00000023000000000000000500000000fffffff0ffffffffffffffdfffffffff",
            INIT_64 => X"0000002a000000000000000800000000ffffffe3ffffffffffffffecffffffff",
            INIT_65 => X"0000002200000000ffffffe5ffffffffffffffd4ffffffff0000000900000000",
            INIT_66 => X"0000001100000000ffffffd8ffffffffffffffdcffffffffffffffc7ffffffff",
            INIT_67 => X"fffffff9ffffffff0000000400000000fffffff5ffffffffffffffbaffffffff",
            INIT_68 => X"0000000d00000000000000090000000000000017000000000000000600000000",
            INIT_69 => X"0000001e000000000000000c00000000ffffffc4ffffffffffffffd1ffffffff",
            INIT_6A => X"0000000d000000000000000000000000ffffffecffffffffffffffdcffffffff",
            INIT_6B => X"0000000a000000000000002700000000ffffffd7ffffffffffffffd7ffffffff",
            INIT_6C => X"00000025000000000000001c00000000ffffffd9ffffffff0000000100000000",
            INIT_6D => X"000000200000000000000020000000000000000500000000fffffffdffffffff",
            INIT_6E => X"ffffffffffffffffffffffdfffffffff0000001b00000000ffffffafffffffff",
            INIT_6F => X"fffffff9ffffffff0000000b000000000000000a00000000ffffffddffffffff",
            INIT_70 => X"0000000c0000000000000017000000000000003900000000ffffffedffffffff",
            INIT_71 => X"fffffff4ffffffff0000001400000000ffffffcafffffffffffffff8ffffffff",
            INIT_72 => X"00000006000000000000001100000000ffffffe7ffffffffffffffcfffffffff",
            INIT_73 => X"00000018000000000000004600000000ffffffe7ffffffffffffffdeffffffff",
            INIT_74 => X"0000001200000000000000030000000000000009000000000000000d00000000",
            INIT_75 => X"00000010000000000000001100000000ffffffe6ffffffff0000000100000000",
            INIT_76 => X"fffffff9ffffffffffffffdbffffffff0000000100000000ffffffd7ffffffff",
            INIT_77 => X"0000000900000000000000000000000000000022000000000000000000000000",
            INIT_78 => X"fffffff6ffffffff0000001f000000000000000900000000fffffffdffffffff",
            INIT_79 => X"0000000d000000000000000e00000000ffffffeffffffffffffffff5ffffffff",
            INIT_7A => X"ffffffdcffffffff0000002600000000fffffffcffffffffffffffd0ffffffff",
            INIT_7B => X"00000012000000000000001d000000000000000600000000fffffff3ffffffff",
            INIT_7C => X"000000270000000000000008000000000000000e000000000000000e00000000",
            INIT_7D => X"0000002500000000ffffffbefffffffffffffff0ffffffff0000002c00000000",
            INIT_7E => X"ffffffd0ffffffffffffffd7ffffffffffffffe1ffffffffffffffd4ffffffff",
            INIT_7F => X"ffffffe8ffffffff0000000200000000ffffffb9ffffffffffffffeaffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE16;


    MEM_IWGHT_LAYER2_INSTANCE17 : if BRAM_NAME = "iwght_layer2_instance17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff1ffffffff0000000e0000000000000014000000000000000400000000",
            INIT_01 => X"00000013000000000000000100000000ffffffecffffffffffffffceffffffff",
            INIT_02 => X"00000000000000000000000c00000000fffffff0ffffffffffffffcfffffffff",
            INIT_03 => X"fffffffcffffffff0000000700000000fffffff4ffffffff0000000700000000",
            INIT_04 => X"0000001e00000000fffffff8ffffffff00000029000000000000001000000000",
            INIT_05 => X"fffffff6ffffffffffffffaeffffffff0000000b000000000000000400000000",
            INIT_06 => X"0000001f00000000ffffffeafffffffffffffffdffffffff0000002600000000",
            INIT_07 => X"ffffffe3ffffffff0000000b00000000ffffffd6ffffffff0000004300000000",
            INIT_08 => X"ffffffeaffffffff00000021000000000000000a000000000000000800000000",
            INIT_09 => X"00000018000000000000001a000000000000000c00000000fffffff1ffffffff",
            INIT_0A => X"ffffffebfffffffffffffff3ffffffff0000001200000000ffffffe1ffffffff",
            INIT_0B => X"ffffffe5ffffffffffffffdaffffffff00000018000000000000001100000000",
            INIT_0C => X"ffffffecffffffff00000006000000000000001300000000fffffffaffffffff",
            INIT_0D => X"ffffffe8ffffffffffffffdfffffffff0000000d000000000000000000000000",
            INIT_0E => X"00000025000000000000000a000000000000000600000000fffffffdffffffff",
            INIT_0F => X"ffffffd3fffffffffffffff2ffffffffffffffb8ffffffff0000001f00000000",
            INIT_10 => X"000000030000000000000018000000000000000f00000000fffffff7ffffffff",
            INIT_11 => X"0000000e0000000000000006000000000000000c00000000ffffffd6ffffffff",
            INIT_12 => X"0000000600000000fffffff9ffffffff0000000f000000000000000800000000",
            INIT_13 => X"0000000600000000fffffff5ffffffff0000000500000000fffffffaffffffff",
            INIT_14 => X"0000000e000000000000000c0000000000000012000000000000000b00000000",
            INIT_15 => X"0000001c00000000ffffffb5fffffffffffffffeffffffff0000000a00000000",
            INIT_16 => X"0000000000000000fffffffdfffffffffffffffbffffffffffffffdeffffffff",
            INIT_17 => X"ffffffeffffffffffffffffeffffffffffffffcafffffffffffffff6ffffffff",
            INIT_18 => X"ffffffebffffffff00000027000000000000002800000000fffffffbffffffff",
            INIT_19 => X"fffffff3ffffffff0000001100000000ffffffe6ffffffffffffffe1ffffffff",
            INIT_1A => X"0000001200000000ffffffe7fffffffffffffff7ffffffffffffffd5ffffffff",
            INIT_1B => X"0000002100000000ffffffd5fffffffffffffffdffffffffffffffd1ffffffff",
            INIT_1C => X"00000029000000000000000a000000000000001300000000ffffffedffffffff",
            INIT_1D => X"0000000200000000ffffffe0fffffffffffffff6ffffffff0000001000000000",
            INIT_1E => X"0000000200000000ffffffcbfffffffffffffff9ffffffffffffffd6ffffffff",
            INIT_1F => X"ffffffe4ffffffff0000000d00000000fffffff8ffffffffffffffebffffffff",
            INIT_20 => X"ffffffd5ffffffff00000015000000000000000c000000000000000f00000000",
            INIT_21 => X"00000008000000000000001d00000000fffffff6ffffffffffffffe2ffffffff",
            INIT_22 => X"fffffff4fffffffffffffff2fffffffffffffff9ffffffffffffffd0ffffffff",
            INIT_23 => X"00000016000000000000000d00000000fffffffbffffffffffffffd2ffffffff",
            INIT_24 => X"00000004000000000000002400000000ffffffe2ffffffff0000001100000000",
            INIT_25 => X"0000001f000000000000000a00000000fffffffcffffffff0000001700000000",
            INIT_26 => X"ffffffebfffffffffffffffbffffffff00000001000000000000000300000000",
            INIT_27 => X"ffffffe1fffffffffffffffaffffffff0000001800000000ffffffd6ffffffff",
            INIT_28 => X"ffffffedfffffffffffffffbffffffffffffffd7ffffffff0000000500000000",
            INIT_29 => X"00000001000000000000001e00000000fffffff0ffffffffffffffdcffffffff",
            INIT_2A => X"fffffffeffffffff0000000900000000ffffffe1ffffffffffffffc2ffffffff",
            INIT_2B => X"0000001b000000000000000900000000fffffff3ffffffffffffffdbffffffff",
            INIT_2C => X"0000001200000000000000320000000000000003000000000000000f00000000",
            INIT_2D => X"0000001f00000000fffffffaffffffff00000003000000000000001000000000",
            INIT_2E => X"ffffffd5ffffffff0000000e00000000fffffffeffffffffffffffeeffffffff",
            INIT_2F => X"ffffffeefffffffffffffffdffffffffffffffdcffffffffffffffe7ffffffff",
            INIT_30 => X"fffffff2ffffffff0000000d0000000000000013000000000000001500000000",
            INIT_31 => X"00000013000000000000000700000000ffffffdcffffffffffffffd5ffffffff",
            INIT_32 => X"ffffffeaffffffff0000000600000000fffffff3ffffffffffffffceffffffff",
            INIT_33 => X"00000029000000000000000d000000000000001300000000fffffff4ffffffff",
            INIT_34 => X"000000180000000000000005000000000000001b000000000000002100000000",
            INIT_35 => X"0000002c00000000fffffff1fffffffffffffffcffffffffffffffffffffffff",
            INIT_36 => X"0000000900000000ffffffdeffffffffffffffbfffffffffffffffdaffffffff",
            INIT_37 => X"ffffffd8ffffffff0000001d00000000ffffffdaffffffff0000000200000000",
            INIT_38 => X"ffffffecffffffff00000046000000000000000500000000fffffffeffffffff",
            INIT_39 => X"00000010000000000000001900000000ffffffdeffffffffffffffc9ffffffff",
            INIT_3A => X"000000010000000000000014000000000000000800000000fffffff0ffffffff",
            INIT_3B => X"0000000100000000000000180000000000000001000000000000000500000000",
            INIT_3C => X"000000070000000000000003000000000000000e000000000000000000000000",
            INIT_3D => X"fffffff7ffffffffffffffdffffffffffffffffaffffffff0000000000000000",
            INIT_3E => X"0000002800000000ffffffedffffffffffffff81ffffffff0000001a00000000",
            INIT_3F => X"ffffffddffffffffffffffefffffffffffffffe5ffffffff0000004300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffefffffffff0000002e000000000000001600000000fffffff7ffffffff",
            INIT_41 => X"ffffffe4ffffffff0000000d000000000000003000000000ffffffe3ffffffff",
            INIT_42 => X"00000015000000000000001a000000000000001300000000fffffff0ffffffff",
            INIT_43 => X"ffffffecfffffffffffffff4fffffffffffffffdffffffff0000001200000000",
            INIT_44 => X"fffffffbffffffffffffffe9fffffffffffffff7fffffffffffffff5ffffffff",
            INIT_45 => X"fffffff1ffffffffffffffd6ffffffff0000000700000000ffffffe9ffffffff",
            INIT_46 => X"0000001b000000000000004a00000000ffffffc9ffffffff0000000e00000000",
            INIT_47 => X"0000000200000000ffffffe3ffffffffffffffa4ffffffff0000000900000000",
            INIT_48 => X"0000001e000000000000001f0000000000000010000000000000000000000000",
            INIT_49 => X"fffffff1fffffffffffffffdffffffff0000000800000000ffffffd8ffffffff",
            INIT_4A => X"ffffffe5ffffffff0000000500000000fffffffbffffffff0000000d00000000",
            INIT_4B => X"0000000300000000ffffffe7fffffffffffffff9fffffffffffffff3ffffffff",
            INIT_4C => X"0000000100000000fffffffcffffffff0000002900000000ffffffefffffffff",
            INIT_4D => X"0000000000000000ffffffccffffffff00000016000000000000000400000000",
            INIT_4E => X"ffffffd5fffffffffffffff2ffffffffffffffbefffffffffffffff0ffffffff",
            INIT_4F => X"fffffff2ffffffffffffffe3ffffffffffffffe3ffffffff0000000000000000",
            INIT_50 => X"000000260000000000000020000000000000001e000000000000001800000000",
            INIT_51 => X"fffffff3ffffffff0000000400000000ffffffe2ffffffffffffffdcffffffff",
            INIT_52 => X"ffffffe7ffffffff00000001000000000000000800000000ffffffdcffffffff",
            INIT_53 => X"00000008000000000000000300000000fffffff8ffffffffffffffddffffffff",
            INIT_54 => X"0000000f00000000fffffffdffffffff0000000800000000fffffffaffffffff",
            INIT_55 => X"0000002600000000ffffffd6ffffffff0000002500000000ffffffe3ffffffff",
            INIT_56 => X"ffffffd4ffffffffffffffddffffffff0000004200000000ffffffd1ffffffff",
            INIT_57 => X"ffffffe1ffffffff0000001400000000ffffffdcffffffffffffffd2ffffffff",
            INIT_58 => X"000000030000000000000017000000000000002700000000ffffffefffffffff",
            INIT_59 => X"0000000000000000fffffff3fffffffffffffff0ffffffffffffffd3ffffffff",
            INIT_5A => X"fffffff2ffffffff00000006000000000000001a00000000fffffff0ffffffff",
            INIT_5B => X"00000016000000000000001a000000000000000400000000ffffffebffffffff",
            INIT_5C => X"00000002000000000000000c000000000000000c00000000ffffffffffffffff",
            INIT_5D => X"fffffff7ffffffff00000017000000000000000c00000000ffffffe1ffffffff",
            INIT_5E => X"ffffffc9fffffffffffffffcffffffff0000001e00000000ffffffeaffffffff",
            INIT_5F => X"ffffffe8fffffffffffffffefffffffffffffffbffffffffffffffe7ffffffff",
            INIT_60 => X"00000003000000000000000e000000000000000800000000ffffffeeffffffff",
            INIT_61 => X"fffffff0ffffffff0000000a00000000fffffff7ffffffffffffffd7ffffffff",
            INIT_62 => X"fffffff2ffffffff0000000500000000fffffff4fffffffffffffff4ffffffff",
            INIT_63 => X"fffffffdffffffffffffffe9fffffffffffffff2ffffffffffffffe1ffffffff",
            INIT_64 => X"fffffffaffffffff00000000000000000000000a00000000fffffff9ffffffff",
            INIT_65 => X"ffffffe1fffffffffffffffcfffffffffffffff7ffffffffffffffffffffffff",
            INIT_66 => X"fffffff3fffffffffffffff1ffffffff0000000f00000000ffffffb7ffffffff",
            INIT_67 => X"fffffff0fffffffffffffffeffffffff0000000100000000ffffffe0ffffffff",
            INIT_68 => X"fffffff5ffffffff00000029000000000000000000000000fffffff3ffffffff",
            INIT_69 => X"ffffffecffffffff0000000a00000000ffffffe9fffffffffffffff7ffffffff",
            INIT_6A => X"ffffffbeffffffff0000001800000000ffffffe4ffffffffffffffe6ffffffff",
            INIT_6B => X"0000000400000000fffffffaffffffff0000000400000000ffffffedffffffff",
            INIT_6C => X"0000000d0000000000000011000000000000002700000000fffffff7ffffffff",
            INIT_6D => X"0000000900000000ffffffccffffffff0000000a00000000ffffffdaffffffff",
            INIT_6E => X"fffffff3ffffffff0000000000000000ffffffe8fffffffffffffff2ffffffff",
            INIT_6F => X"fffffff3ffffffff0000000700000000ffffffb9ffffffff0000000300000000",
            INIT_70 => X"000000100000000000000034000000000000000f000000000000000600000000",
            INIT_71 => X"0000002800000000ffffffecffffffffffffffd3ffffffffffffffe1ffffffff",
            INIT_72 => X"ffffffd0fffffffffffffff2ffffffffffffffe1ffffffffffffffe0ffffffff",
            INIT_73 => X"00000009000000000000000e0000000000000000000000000000001200000000",
            INIT_74 => X"ffffffe2fffffffffffffff4ffffffff0000001c000000000000002200000000",
            INIT_75 => X"fffffff9ffffffffffffffceffffffff00000000000000000000000400000000",
            INIT_76 => X"fffffff9ffffffffffffffe8ffffffffffffffceffffffff0000002200000000",
            INIT_77 => X"fffffffefffffffffffffffbffffffffffffffe2ffffffff0000002700000000",
            INIT_78 => X"fffffff8ffffffff0000003900000000ffffffffffffffff0000000400000000",
            INIT_79 => X"ffffffe0fffffffffffffff8ffffffff0000001200000000fffffff3ffffffff",
            INIT_7A => X"ffffffd9ffffffff0000003000000000ffffffeeffffffff0000000d00000000",
            INIT_7B => X"ffffffc9ffffffffffffffc9ffffffff00000005000000000000001500000000",
            INIT_7C => X"fffffff0ffffffffffffffe4fffffffffffffff3fffffffffffffffdffffffff",
            INIT_7D => X"ffffffdffffffffffffffff6ffffffff0000001a000000000000000400000000",
            INIT_7E => X"00000029000000000000001500000000ffffffc6ffffffff0000004700000000",
            INIT_7F => X"0000000300000000ffffffd3ffffffffffffffe7ffffffff0000001400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE17;


    MEM_IWGHT_LAYER2_INSTANCE18 : if BRAM_NAME = "iwght_layer2_instance18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff9ffffffff00000017000000000000000000000000fffffff8ffffffff",
            INIT_01 => X"0000000a000000000000001f000000000000000f00000000fffffff9ffffffff",
            INIT_02 => X"ffffffc8ffffffff0000002a000000000000001b000000000000003600000000",
            INIT_03 => X"0000000b00000000ffffffe1ffffffff00000011000000000000001300000000",
            INIT_04 => X"fffffff7ffffffff0000000c000000000000001a00000000fffffff8ffffffff",
            INIT_05 => X"0000002b00000000ffffffdcffffffff00000006000000000000000000000000",
            INIT_06 => X"00000006000000000000000000000000fffffff8fffffffffffffff9ffffffff",
            INIT_07 => X"0000000c000000000000000600000000ffffffc5ffffffff0000000400000000",
            INIT_08 => X"00000006000000000000000b000000000000000f00000000ffffffe3ffffffff",
            INIT_09 => X"0000001100000000ffffffffffffffff0000002000000000ffffffe8ffffffff",
            INIT_0A => X"ffffffc5ffffffff0000001e00000000fffffff9fffffffffffffff1ffffffff",
            INIT_0B => X"0000000700000000fffffff2ffffffff0000001400000000fffffff4ffffffff",
            INIT_0C => X"00000024000000000000001e000000000000001d000000000000000800000000",
            INIT_0D => X"ffffffe2fffffffffffffff7ffffffff00000006000000000000000000000000",
            INIT_0E => X"0000002200000000ffffffe5ffffffffffffffdeffffffff0000002200000000",
            INIT_0F => X"0000000f000000000000000000000000ffffffcefffffffffffffff9ffffffff",
            INIT_10 => X"ffffffe8ffffffff000000040000000000000000000000000000000900000000",
            INIT_11 => X"00000001000000000000000400000000fffffff7fffffffffffffff5ffffffff",
            INIT_12 => X"ffffffe1ffffffff000000120000000000000000000000000000000a00000000",
            INIT_13 => X"fffffff2ffffffff00000005000000000000001c000000000000001600000000",
            INIT_14 => X"fffffffcffffffff00000024000000000000001e00000000fffffff9ffffffff",
            INIT_15 => X"fffffffaffffffffffffffe5ffffffff0000000d00000000fffffffdffffffff",
            INIT_16 => X"ffffffecffffffff0000001500000000ffffffdbffffffff0000001700000000",
            INIT_17 => X"fffffff9ffffffff0000000200000000ffffffebffffffff0000001b00000000",
            INIT_18 => X"000000000000000000000033000000000000001800000000fffffff7ffffffff",
            INIT_19 => X"fffffffafffffffffffffff5ffffffffffffffefffffffff0000000600000000",
            INIT_1A => X"ffffffdfffffffff0000000900000000fffffffbffffffffffffffe6ffffffff",
            INIT_1B => X"fffffffeffffffffffffffefffffffff0000001e000000000000000500000000",
            INIT_1C => X"000000110000000000000014000000000000001e00000000ffffffe9ffffffff",
            INIT_1D => X"fffffffdfffffffffffffffbfffffffffffffffeffffffffffffffe9ffffffff",
            INIT_1E => X"ffffffebffffffff0000000900000000ffffffefffffffffffffffffffffffff",
            INIT_1F => X"00000006000000000000000200000000ffffffdbffffffff0000003400000000",
            INIT_20 => X"fffffff0ffffffff0000001a000000000000000500000000fffffff5ffffffff",
            INIT_21 => X"fffffff1fffffffffffffffeffffffff0000001200000000ffffffe6ffffffff",
            INIT_22 => X"ffffffb1ffffffff0000002800000000ffffffffffffffffffffffd9ffffffff",
            INIT_23 => X"ffffffecffffffff0000002600000000ffffffffffffffff0000001100000000",
            INIT_24 => X"0000003000000000fffffff7ffffffff0000002300000000ffffffe6ffffffff",
            INIT_25 => X"ffffffffffffffffffffffbdffffffff0000000a00000000fffffff6ffffffff",
            INIT_26 => X"00000003000000000000001100000000ffffffe9ffffffff0000001800000000",
            INIT_27 => X"ffffffe9ffffffff0000000300000000ffffffc6ffffffff0000002200000000",
            INIT_28 => X"fffffffdffffffff00000038000000000000001e000000000000001100000000",
            INIT_29 => X"fffffffbfffffffffffffff3ffffffff0000001a00000000ffffffdbffffffff",
            INIT_2A => X"ffffffc6ffffffff00000005000000000000000300000000ffffffc8ffffffff",
            INIT_2B => X"fffffff7fffffffffffffff9ffffffff00000017000000000000000a00000000",
            INIT_2C => X"ffffffe5ffffffff00000000000000000000002b000000000000001600000000",
            INIT_2D => X"ffffffedffffffffffffffdcfffffffffffffff2ffffffff0000000000000000",
            INIT_2E => X"ffffffefffffffffffffffe7ffffffffffffffe6ffffffff0000002800000000",
            INIT_2F => X"ffffffe8fffffffffffffff1ffffffffffffffdaffffffff0000003e00000000",
            INIT_30 => X"000000050000000000000037000000000000000300000000fffffffeffffffff",
            INIT_31 => X"00000008000000000000000f000000000000001800000000ffffffedffffffff",
            INIT_32 => X"fffffff0ffffffff0000000e000000000000002e000000000000000c00000000",
            INIT_33 => X"fffffffcffffffffffffffc2ffffffff00000006000000000000001900000000",
            INIT_34 => X"ffffffe5ffffffff0000001000000000ffffffc2ffffffffffffffc4ffffffff",
            INIT_35 => X"fffffffbffffffffffffffdfffffffffffffffd3ffffffffffffffd8ffffffff",
            INIT_36 => X"ffffffedfffffffffffffff2ffffffffffffffdfffffffffffffffcbffffffff",
            INIT_37 => X"00000017000000000000002300000000ffffffe6fffffffffffffff0ffffffff",
            INIT_38 => X"ffffffefffffffffffffffe5ffffffffffffffeeffffffff0000001d00000000",
            INIT_39 => X"fffffffbffffffff0000001300000000ffffffe4ffffffffffffffeeffffffff",
            INIT_3A => X"00000036000000000000000700000000ffffffb2ffffffff0000000800000000",
            INIT_3B => X"ffffffefffffffff0000001800000000fffffff5ffffffff0000001400000000",
            INIT_3C => X"0000002900000000fffffffeffffffffffffffe9ffffffffffffffe4ffffffff",
            INIT_3D => X"fffffff2fffffffffffffff6ffffffffffffffd8fffffffffffffff7ffffffff",
            INIT_3E => X"fffffffeffffffffffffffdaffffffffffffffebfffffffffffffff6ffffffff",
            INIT_3F => X"0000003a000000000000001c000000000000000c00000000fffffffeffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffe7ffffffffffffffb1ffffffff0000000b000000000000001c00000000",
            INIT_41 => X"ffffffffffffffff0000000c00000000fffffff3ffffffff0000000300000000",
            INIT_42 => X"00000006000000000000000400000000ffffffb6ffffffff0000001200000000",
            INIT_43 => X"fffffffeffffffff0000000600000000fffffffcffffffff0000000200000000",
            INIT_44 => X"fffffffdffffffff00000012000000000000000000000000ffffffe5ffffffff",
            INIT_45 => X"ffffffffffffffffffffffe7ffffffffffffffebfffffffffffffff2ffffffff",
            INIT_46 => X"0000000900000000ffffffebffffffff00000042000000000000001100000000",
            INIT_47 => X"fffffffefffffffffffffff4ffffffff00000004000000000000001500000000",
            INIT_48 => X"fffffff9ffffffffffffffd9ffffffffffffffffffffffff0000000d00000000",
            INIT_49 => X"fffffff9ffffffff00000014000000000000000b000000000000000800000000",
            INIT_4A => X"ffffffcbffffffff0000001100000000ffffffc6fffffffffffffffdffffffff",
            INIT_4B => X"fffffff6ffffffffffffffceffffffff00000005000000000000000e00000000",
            INIT_4C => X"fffffff9fffffffffffffff7ffffffff0000000200000000ffffffefffffffff",
            INIT_4D => X"00000045000000000000000800000000ffffffeaffffffffffffffe0ffffffff",
            INIT_4E => X"ffffffffffffffffffffffd2ffffffff0000003600000000fffffffaffffffff",
            INIT_4F => X"fffffffaffffffff00000003000000000000000a000000000000001e00000000",
            INIT_50 => X"ffffffecffffffffffffffebffffffff0000000f000000000000000c00000000",
            INIT_51 => X"00000010000000000000001c000000000000000c000000000000001900000000",
            INIT_52 => X"ffffffe4ffffffff0000002000000000ffffffddffffffff0000000700000000",
            INIT_53 => X"fffffffbfffffffffffffff1ffffffff00000004000000000000000600000000",
            INIT_54 => X"fffffff0ffffffff0000001e00000000fffffffbffffffff0000000000000000",
            INIT_55 => X"0000001e000000000000001200000000ffffffd1ffffffff0000000100000000",
            INIT_56 => X"ffffffdbffffffff000000050000000000000004000000000000001700000000",
            INIT_57 => X"00000041000000000000001e00000000fffffffefffffffffffffffcffffffff",
            INIT_58 => X"0000001100000000ffffffddffffffff0000001d000000000000000400000000",
            INIT_59 => X"0000001b000000000000000600000000fffffffcffffffff0000000800000000",
            INIT_5A => X"ffffffbcffffffff0000000300000000ffffffd8ffffffff0000001800000000",
            INIT_5B => X"ffffffdbffffffff000000150000000000000001000000000000001200000000",
            INIT_5C => X"000000090000000000000000000000000000000700000000fffffff7ffffffff",
            INIT_5D => X"00000021000000000000000800000000ffffffe6ffffffff0000000e00000000",
            INIT_5E => X"ffffffebffffffffffffffb7ffffffff0000000800000000ffffffd6ffffffff",
            INIT_5F => X"fffffff6ffffffff000000110000000000000013000000000000000a00000000",
            INIT_60 => X"0000000700000000ffffffe6ffffffffffffffe6fffffffffffffffbffffffff",
            INIT_61 => X"0000001e00000000000000110000000000000013000000000000000500000000",
            INIT_62 => X"ffffff9fffffffffffffffe0ffffffffffffffe8ffffffff0000001400000000",
            INIT_63 => X"ffffffffffffffff0000003a00000000fffffff7ffffffff0000001200000000",
            INIT_64 => X"0000001500000000fffffffaffffffffffffffd7ffffffffffffffd3ffffffff",
            INIT_65 => X"ffffffeefffffffffffffff8ffffffffffffffc2ffffffffffffffe9ffffffff",
            INIT_66 => X"0000001500000000ffffffc6ffffffff0000005300000000ffffffd4ffffffff",
            INIT_67 => X"fffffff6ffffffff0000001500000000ffffffe8ffffffff0000000900000000",
            INIT_68 => X"00000003000000000000000600000000ffffffe9ffffffff0000000c00000000",
            INIT_69 => X"fffffffaffffffff0000001b0000000000000009000000000000001b00000000",
            INIT_6A => X"0000000a000000000000001f00000000ffffffd0ffffffff0000001300000000",
            INIT_6B => X"0000000f00000000ffffffe6ffffffff00000016000000000000000500000000",
            INIT_6C => X"00000009000000000000002100000000ffffffceffffffffffffffefffffffff",
            INIT_6D => X"fffffff3fffffffffffffff9fffffffffffffff4ffffffff0000000e00000000",
            INIT_6E => X"0000000900000000fffffff1ffffffff00000008000000000000001300000000",
            INIT_6F => X"0000001a000000000000000c00000000fffffff4fffffffffffffff7ffffffff",
            INIT_70 => X"00000012000000000000000300000000ffffffffffffffff0000001200000000",
            INIT_71 => X"fffffffdffffffff000000140000000000000009000000000000000400000000",
            INIT_72 => X"0000000e000000000000001200000000ffffffe8ffffffffffffffefffffffff",
            INIT_73 => X"ffffffeaffffffffffffffebffffffffffffffdcffffffff0000000700000000",
            INIT_74 => X"fffffffefffffffffffffff9fffffffffffffff3ffffffff0000000900000000",
            INIT_75 => X"fffffff4fffffffffffffff6ffffffff0000000c000000000000000800000000",
            INIT_76 => X"ffffffe8ffffffffffffffecffffffffffffffefffffffff0000001200000000",
            INIT_77 => X"0000000b000000000000000d000000000000000500000000fffffff1ffffffff",
            INIT_78 => X"0000001400000000ffffffeeffffffff00000007000000000000000000000000",
            INIT_79 => X"0000000800000000fffffff9ffffffff0000000a000000000000001500000000",
            INIT_7A => X"000000000000000000000008000000000000000b00000000ffffffe7ffffffff",
            INIT_7B => X"fffffff7ffffffffffffffe0ffffffff00000004000000000000000600000000",
            INIT_7C => X"ffffffe0ffffffffffffffeeffffffffffffffe2fffffffffffffff9ffffffff",
            INIT_7D => X"fffffff8ffffffff0000000c000000000000000500000000ffffffb9ffffffff",
            INIT_7E => X"ffffffb5ffffffffffffffedffffffffffffffecfffffffffffffffbffffffff",
            INIT_7F => X"0000001e000000000000001b00000000ffffffe5ffffffffffffffe4ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE18;


    MEM_IWGHT_LAYER2_INSTANCE19 : if BRAM_NAME = "iwght_layer2_instance19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff6ffffffffffffff98ffffffffffffffd6ffffffff0000000f00000000",
            INIT_01 => X"0000000200000000000000010000000000000017000000000000001600000000",
            INIT_02 => X"ffffffc5ffffffffffffffffffffffffffffffe9ffffffffffffffe9ffffffff",
            INIT_03 => X"fffffff0ffffffffffffffdeffffffff00000040000000000000000f00000000",
            INIT_04 => X"ffffffa3ffffffffffffffeafffffffffffffff7ffffffff0000000100000000",
            INIT_05 => X"0000000000000000fffffff0ffffffffffffffe3ffffffffffffffb6ffffffff",
            INIT_06 => X"fffffff5fffffffffffffff0ffffffffffffffa3ffffffff0000002500000000",
            INIT_07 => X"0000002b00000000fffffffdffffffff00000002000000000000001700000000",
            INIT_08 => X"0000000e00000000ffffffe2ffffffffffffffcdffffffff0000001a00000000",
            INIT_09 => X"0000001f000000000000000a00000000fffffff1ffffffff0000000d00000000",
            INIT_0A => X"ffffffa3ffffffff0000000700000000fffffff1ffffffff0000002800000000",
            INIT_0B => X"ffffffccffffffff00000000000000000000001c000000000000001900000000",
            INIT_0C => X"ffffffc6ffffffffffffffc5ffffffff0000004800000000ffffffddffffffff",
            INIT_0D => X"ffffffe2ffffffff0000000d00000000ffffffceffffffffffffffceffffffff",
            INIT_0E => X"ffffffd4ffffffffffffffbeffffffffffffffe8ffffffff0000002200000000",
            INIT_0F => X"fffffffeffffffff0000001f000000000000001400000000fffffff0ffffffff",
            INIT_10 => X"fffffff8ffffffffffffffcdffffffffffffff9effffffff0000000e00000000",
            INIT_11 => X"0000002900000000fffffffcffffffffffffffdfffffffff0000001300000000",
            INIT_12 => X"ffffffa7ffffffffffffffdefffffffffffffffbfffffffffffffff8ffffffff",
            INIT_13 => X"ffffffe4ffffffff000000260000000000000014000000000000000e00000000",
            INIT_14 => X"fffffff7ffffffffffffffcdffffffffffffffdffffffffffffffffeffffffff",
            INIT_15 => X"fffffffbffffffff0000000f00000000ffffffc7fffffffffffffff9ffffffff",
            INIT_16 => X"ffffffddffffffffffffffddfffffffffffffffcffffffffffffffebffffffff",
            INIT_17 => X"fffffff4ffffffff0000001a000000000000000000000000fffffff8ffffffff",
            INIT_18 => X"0000001a000000000000000e00000000ffffffdaffffffff0000000500000000",
            INIT_19 => X"0000000a000000000000001b00000000fffffffdffffffff0000000f00000000",
            INIT_1A => X"ffffffdeffffffffffffffe2ffffffff0000000a000000000000000200000000",
            INIT_1B => X"ffffffedffffffff0000003e00000000fffffff6ffffffff0000000300000000",
            INIT_1C => X"ffffffeafffffffffffffffcffffffff0000001000000000fffffff9ffffffff",
            INIT_1D => X"00000010000000000000001e0000000000000003000000000000001800000000",
            INIT_1E => X"0000000a00000000ffffffa7fffffffffffffff8ffffffffffffffb6ffffffff",
            INIT_1F => X"00000002000000000000000200000000ffffffe1ffffffff0000000300000000",
            INIT_20 => X"0000001a00000000fffffff3ffffffffffffffecffffffff0000000000000000",
            INIT_21 => X"ffffffe7ffffffff00000012000000000000003100000000fffffff7ffffffff",
            INIT_22 => X"ffffffe0ffffffff00000009000000000000000700000000fffffff6ffffffff",
            INIT_23 => X"0000002000000000fffffffafffffffffffffff2fffffffffffffff1ffffffff",
            INIT_24 => X"ffffffccffffffff0000002100000000ffffffc6ffffffff0000000d00000000",
            INIT_25 => X"ffffffeeffffffffffffffd3ffffffffffffffe5ffffffff0000001200000000",
            INIT_26 => X"0000000300000000ffffffdeffffffffffffffd0fffffffffffffff2ffffffff",
            INIT_27 => X"00000015000000000000000a00000000ffffffd8fffffffffffffff1ffffffff",
            INIT_28 => X"0000000800000000fffffff8fffffffffffffffffffffffffffffff8ffffffff",
            INIT_29 => X"fffffff7ffffffff0000002e000000000000000e000000000000002400000000",
            INIT_2A => X"ffffffdfffffffffffffffe9ffffffffffffffd4ffffffffffffffcaffffffff",
            INIT_2B => X"fffffffdffffffff0000000300000000fffffff3ffffffff0000001200000000",
            INIT_2C => X"fffffff4ffffffff0000001800000000ffffffe1fffffffffffffff5ffffffff",
            INIT_2D => X"ffffffe7ffffffff0000000b00000000fffffff0ffffffffffffffebffffffff",
            INIT_2E => X"ffffffc6ffffffffffffffe6ffffffff00000002000000000000003000000000",
            INIT_2F => X"0000000300000000ffffffeaffffffffffffffeffffffffffffffff1ffffffff",
            INIT_30 => X"0000000f0000000000000012000000000000000400000000fffffffaffffffff",
            INIT_31 => X"0000000600000000000000110000000000000001000000000000000900000000",
            INIT_32 => X"ffffffe6ffffffff00000008000000000000003a00000000ffffffd3ffffffff",
            INIT_33 => X"fffffff3fffffffffffffff9ffffffff0000000e000000000000001300000000",
            INIT_34 => X"ffffffecffffffffffffffc9ffffffff0000001e000000000000001100000000",
            INIT_35 => X"ffffffadffffffffffffffecffffffff0000000600000000ffffffb0ffffffff",
            INIT_36 => X"ffffffbaffffffffffffffcfffffffffffffffe2ffffffff0000002100000000",
            INIT_37 => X"0000000d000000000000001c0000000000000000000000000000000000000000",
            INIT_38 => X"0000001c00000000ffffffc9ffffffffffffffeeffffffff0000001e00000000",
            INIT_39 => X"0000001b00000000fffffff4ffffffffffffffe9ffffffff0000000200000000",
            INIT_3A => X"ffffffd5ffffffffffffffffffffffff0000003f000000000000000500000000",
            INIT_3B => X"ffffffefffffffffffffffc3ffffffff00000013000000000000004800000000",
            INIT_3C => X"ffffffa6ffffffffffffffd3ffffffff0000002200000000fffffffeffffffff",
            INIT_3D => X"ffffff8cffffffffffffffdaffffffff0000000200000000ffffffa8ffffffff",
            INIT_3E => X"0000000c00000000ffffffb1ffffffffffffff50fffffffffffffffcffffffff",
            INIT_3F => X"ffffffffffffffff0000001000000000fffffff1ffffffff0000002b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff8ffffffffffffffd4ffffffffffffffceffffffff0000001f00000000",
            INIT_41 => X"0000002000000000000000080000000000000003000000000000000200000000",
            INIT_42 => X"ffffffd8ffffffffffffffedffffffffffffffd0ffffffff0000001400000000",
            INIT_43 => X"0000001700000000ffffffdcffffffff00000025000000000000001e00000000",
            INIT_44 => X"fffffff3ffffffffffffffc9ffffffff0000003b00000000ffffffedffffffff",
            INIT_45 => X"ffffffc0ffffffffffffffedfffffffffffffff7ffffffffffffffbeffffffff",
            INIT_46 => X"0000000e00000000ffffffa4fffffffffffffffdffffffff0000000800000000",
            INIT_47 => X"fffffff8ffffffff0000001b000000000000000300000000fffffff2ffffffff",
            INIT_48 => X"00000005000000000000000b00000000ffffffd1ffffffff0000001a00000000",
            INIT_49 => X"0000002b000000000000000700000000ffffffeeffffffff0000000e00000000",
            INIT_4A => X"0000000e00000000ffffffdbffffffffffffffffffffffff0000001100000000",
            INIT_4B => X"ffffffe2ffffffff0000000700000000ffffffeefffffffffffffffdffffffff",
            INIT_4C => X"0000000a00000000ffffffd6ffffffff0000001800000000ffffffe2ffffffff",
            INIT_4D => X"fffffff2ffffffff0000000600000000fffffff8fffffffffffffffbffffffff",
            INIT_4E => X"fffffff2ffffffffffffffb4fffffffffffffff6ffffffffffffffb7ffffffff",
            INIT_4F => X"00000003000000000000001700000000fffffff1ffffffff0000000000000000",
            INIT_50 => X"00000034000000000000001b000000000000001200000000fffffffcffffffff",
            INIT_51 => X"0000001300000000fffffffbffffffffffffffebffffffff0000002300000000",
            INIT_52 => X"000000110000000000000001000000000000001c00000000ffffffdaffffffff",
            INIT_53 => X"fffffff3ffffffff0000002200000000ffffffebffffffffffffffe2ffffffff",
            INIT_54 => X"fffffff5ffffffff0000001100000000ffffffdcffffffff0000002e00000000",
            INIT_55 => X"fffffff4ffffffff0000000400000000fffffff8ffffffff0000001e00000000",
            INIT_56 => X"ffffffd4fffffffffffffff3ffffffffffffffcfffffffffffffffcfffffffff",
            INIT_57 => X"fffffffafffffffffffffff1fffffffffffffffaffffffff0000002700000000",
            INIT_58 => X"0000001c00000000ffffffe6ffffffff0000001c00000000fffffff8ffffffff",
            INIT_59 => X"000000000000000000000017000000000000002a000000000000000b00000000",
            INIT_5A => X"0000000a000000000000001a000000000000000700000000ffffffe3ffffffff",
            INIT_5B => X"0000000f000000000000000000000000fffffffbffffffffffffffe3ffffffff",
            INIT_5C => X"ffffffebffffffff0000002100000000ffffffb3ffffffff0000002900000000",
            INIT_5D => X"ffffffffffffffffffffffe0ffffffffffffffe1ffffffff0000001200000000",
            INIT_5E => X"ffffffedffffffffffffffd0ffffffffffffffcfffffffff0000001c00000000",
            INIT_5F => X"0000001400000000ffffffecffffffffffffffdaffffffff0000000700000000",
            INIT_60 => X"0000001b000000000000000c00000000fffffff0fffffffffffffff2ffffffff",
            INIT_61 => X"ffffffd8ffffffff000000070000000000000018000000000000000d00000000",
            INIT_62 => X"ffffffc3ffffffffffffffd2fffffffffffffff8ffffffffffffffeaffffffff",
            INIT_63 => X"00000005000000000000005100000000fffffff1ffffffff0000000800000000",
            INIT_64 => X"0000000000000000fffffff1ffffffffffffffcbffffffff0000000300000000",
            INIT_65 => X"ffffffe0ffffffffffffffccffffffffffffffe8fffffffffffffff8ffffffff",
            INIT_66 => X"ffffffdeffffffffffffffc5ffffffffffffff9cffffffffffffffd9ffffffff",
            INIT_67 => X"fffffffaffffffff0000000d000000000000002f00000000fffffff8ffffffff",
            INIT_68 => X"0000002500000000000000190000000000000019000000000000000900000000",
            INIT_69 => X"000000080000000000000005000000000000000f000000000000000800000000",
            INIT_6A => X"ffffffd9ffffffffffffffc2ffffffff0000003000000000ffffffc6ffffffff",
            INIT_6B => X"ffffffd5ffffffff0000001f00000000ffffffecffffffff0000004600000000",
            INIT_6C => X"ffffffd1ffffffffffffffc9ffffffffffffffeeffffffffffffffebffffffff",
            INIT_6D => X"ffffffd2ffffffffffffffc8ffffffff0000000600000000ffffffc8ffffffff",
            INIT_6E => X"fffffff4ffffffffffffffb4ffffffffffffffc0ffffffffffffffe5ffffffff",
            INIT_6F => X"fffffffbffffffff0000000700000000ffffffdbffffffff0000001200000000",
            INIT_70 => X"0000001200000000000000030000000000000000000000000000002000000000",
            INIT_71 => X"000000110000000000000014000000000000000100000000ffffffe3ffffffff",
            INIT_72 => X"ffffffbdffffffffffffff94ffffffff0000001800000000ffffffdeffffffff",
            INIT_73 => X"fffffff0ffffffffffffffc0ffffffff00000022000000000000006200000000",
            INIT_74 => X"ffffffd2ffffffffffffffe9ffffffffffffffe0ffffffffffffffe8ffffffff",
            INIT_75 => X"ffffffa4ffffffffffffffa1fffffffffffffff2ffffffffffffffd6ffffffff",
            INIT_76 => X"0000003700000000ffffffb3ffffffffffffff26ffffffff0000002c00000000",
            INIT_77 => X"ffffffefffffffff0000001200000000ffffffc2ffffffff0000001200000000",
            INIT_78 => X"ffffffe0ffffffffffffffd7ffffffffffffffb3ffffffff0000004000000000",
            INIT_79 => X"0000001e000000000000002a00000000fffffffaffffffffffffffe2ffffffff",
            INIT_7A => X"0000001900000000ffffffd9fffffffffffffff7ffffffffffffffecffffffff",
            INIT_7B => X"0000000500000000ffffffd9ffffffff00000017000000000000005300000000",
            INIT_7C => X"ffffffe0ffffffffffffffeafffffffffffffff5ffffffffffffffe5ffffffff",
            INIT_7D => X"ffffffa7ffffffffffffffddffffffff0000000e00000000ffffffe3ffffffff",
            INIT_7E => X"0000003400000000ffffff9dffffffffffffffd6ffffffffffffffc6ffffffff",
            INIT_7F => X"fffffff6ffffffff0000002800000000ffffffebffffffffffffffcaffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE19;


    MEM_IWGHT_LAYER2_INSTANCE20 : if BRAM_NAME = "iwght_layer2_instance20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffffefffffffffffffffaffffffff0000000d000000000000002300000000",
            INIT_01 => X"00000017000000000000000500000000ffffffe2ffffffff0000000c00000000",
            INIT_02 => X"0000001800000000fffffff9ffffffffffffffe9fffffffffffffff1ffffffff",
            INIT_03 => X"ffffffe2fffffffffffffff7ffffffffffffffdeffffffff0000001100000000",
            INIT_04 => X"0000000000000000ffffffe6ffffffffffffffa8ffffffff0000000b00000000",
            INIT_05 => X"ffffffcfffffffff0000002600000000fffffff4ffffffffffffffd7ffffffff",
            INIT_06 => X"fffffff5ffffffffffffffbeffffffffffffffecffffffffffffffd9ffffffff",
            INIT_07 => X"00000006000000000000001e00000000fffffffaffffffffffffffd3ffffffff",
            INIT_08 => X"00000000000000000000002b000000000000002300000000fffffffbffffffff",
            INIT_09 => X"ffffffffffffffff0000000200000000fffffff2ffffffff0000000700000000",
            INIT_0A => X"000000070000000000000009000000000000001e00000000ffffffdbffffffff",
            INIT_0B => X"fffffffcffffffff0000000700000000fffffff6ffffffffffffffdeffffffff",
            INIT_0C => X"ffffffd6ffffffff0000000b00000000fffffffaffffffff0000002800000000",
            INIT_0D => X"ffffffe3ffffffff0000000300000000ffffffe7fffffffffffffffeffffffff",
            INIT_0E => X"ffffffd9ffffffffffffffdaffffffffffffffceffffffffffffffc0ffffffff",
            INIT_0F => X"0000000c00000000ffffffecffffffff0000000700000000fffffff7ffffffff",
            INIT_10 => X"0000003b000000000000000a000000000000000900000000ffffffefffffffff",
            INIT_11 => X"fffffff6fffffffffffffff5ffffffff00000012000000000000000d00000000",
            INIT_12 => X"ffffffdeffffffff0000001000000000fffffffbffffffffffffffddffffffff",
            INIT_13 => X"000000230000000000000010000000000000001100000000ffffffeeffffffff",
            INIT_14 => X"00000000000000000000002200000000ffffffc2ffffffff0000001300000000",
            INIT_15 => X"0000000900000000ffffffdfffffffffffffffebffffffffffffffe5ffffffff",
            INIT_16 => X"fffffff4ffffffffffffff86ffffffffffffffeaffffffffffffffdcffffffff",
            INIT_17 => X"0000000e00000000fffffff9ffffffffffffffc3ffffffff0000000800000000",
            INIT_18 => X"ffffffebffffffffffffffffffffffff0000001e000000000000001200000000",
            INIT_19 => X"fffffff9ffffffff00000010000000000000002000000000fffffff7ffffffff",
            INIT_1A => X"fffffff0fffffffffffffffeffffffff0000000900000000ffffffeaffffffff",
            INIT_1B => X"000000060000000000000045000000000000000700000000fffffffcffffffff",
            INIT_1C => X"00000001000000000000000400000000ffffffceffffffff0000000700000000",
            INIT_1D => X"0000003b00000000ffffffe1ffffffffffffffddffffffffffffffd1ffffffff",
            INIT_1E => X"ffffffc2ffffffffffffffd1ffffffff0000000400000000fffffff9ffffffff",
            INIT_1F => X"00000014000000000000000a000000000000002700000000ffffffbaffffffff",
            INIT_20 => X"0000000900000000000000000000000000000006000000000000001100000000",
            INIT_21 => X"0000001800000000000000070000000000000002000000000000000a00000000",
            INIT_22 => X"ffffffe4fffffffffffffff0ffffffff0000001300000000ffffffd5ffffffff",
            INIT_23 => X"ffffffeeffffffff0000002e00000000fffffff5ffffffff0000000f00000000",
            INIT_24 => X"0000000e00000000fffffffaffffffffffffffddffffffff0000000800000000",
            INIT_25 => X"ffffffe4ffffffffffffffeefffffffffffffffdffffffffffffffdaffffffff",
            INIT_26 => X"ffffffe6ffffffffffffffb8ffffffffffffffcfffffffff0000001e00000000",
            INIT_27 => X"00000010000000000000001a000000000000000e00000000fffffff8ffffffff",
            INIT_28 => X"00000023000000000000001d000000000000000a000000000000000700000000",
            INIT_29 => X"0000001e000000000000000000000000ffffffe0ffffffff0000002000000000",
            INIT_2A => X"fffffff5ffffffffffffffb9ffffffff0000003500000000ffffffe8ffffffff",
            INIT_2B => X"ffffffe9ffffffff0000002000000000fffffffdffffffff0000003100000000",
            INIT_2C => X"fffffff4ffffffffffffffd5ffffffffffffffb7ffffffffffffffd4ffffffff",
            INIT_2D => X"ffffffffffffffffffffffc4fffffffffffffffcfffffffffffffff0ffffffff",
            INIT_2E => X"0000000800000000ffffff89ffffffff0000001100000000ffffffb2ffffffff",
            INIT_2F => X"0000000c000000000000001500000000ffffffebffffffffffffffc0ffffffff",
            INIT_30 => X"fffffffeffffffffffffffe6fffffffffffffff3ffffffff0000001100000000",
            INIT_31 => X"000000130000000000000004000000000000001700000000fffffff9ffffffff",
            INIT_32 => X"fffffffefffffffffffffff0ffffffff0000004300000000ffffffe4ffffffff",
            INIT_33 => X"0000002a00000000000000050000000000000008000000000000001f00000000",
            INIT_34 => X"0000000e000000000000000b00000000ffffffbaffffffff0000001700000000",
            INIT_35 => X"ffffffacffffffff0000000800000000ffffffe2ffffffffffffffcbffffffff",
            INIT_36 => X"0000000a00000000ffffffd5ffffffffffffff81ffffffffffffffd9ffffffff",
            INIT_37 => X"0000001d0000000000000024000000000000003600000000ffffffdaffffffff",
            INIT_38 => X"0000002d00000000000000030000000000000019000000000000001900000000",
            INIT_39 => X"0000001e00000000ffffffe9fffffffffffffffdfffffffffffffffdffffffff",
            INIT_3A => X"ffffffefffffffff0000001c00000000fffffffdffffffffffffffe6ffffffff",
            INIT_3B => X"fffffff2ffffffff0000000b00000000fffffff5ffffffff0000001500000000",
            INIT_3C => X"fffffff9fffffffffffffff2ffffffffffffffb6fffffffffffffffdffffffff",
            INIT_3D => X"fffffffcffffffff0000002900000000ffffffeaffffffffffffffdaffffffff",
            INIT_3E => X"ffffffedffffffffffffffe5ffffffffffffff92ffffffffffffffdeffffffff",
            INIT_3F => X"000000240000000000000012000000000000002700000000fffffff0ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002a00000000fffffff4ffffffff00000005000000000000000400000000",
            INIT_41 => X"0000001c00000000ffffffeffffffffffffffff0ffffffffffffffe8ffffffff",
            INIT_42 => X"ffffffd8ffffffff00000005000000000000001600000000ffffffdaffffffff",
            INIT_43 => X"ffffffe2fffffffffffffff7fffffffffffffffdffffffff0000000500000000",
            INIT_44 => X"00000001000000000000002200000000fffffff3ffffffff0000003800000000",
            INIT_45 => X"00000025000000000000000200000000fffffff3fffffffffffffffaffffffff",
            INIT_46 => X"ffffffb8ffffffffffffffb8ffffffff0000001d00000000ffffffd3ffffffff",
            INIT_47 => X"0000000e000000000000001900000000ffffffc4ffffffffffffffefffffffff",
            INIT_48 => X"00000016000000000000001a000000000000000e000000000000000b00000000",
            INIT_49 => X"0000000700000000fffffffcffffffff0000001300000000ffffffdcffffffff",
            INIT_4A => X"ffffffdaffffffffffffffe9ffffffff0000000f00000000ffffffe9ffffffff",
            INIT_4B => X"00000025000000000000004c00000000ffffffecffffffff0000000600000000",
            INIT_4C => X"0000000c000000000000000600000000ffffffd3ffffffff0000001200000000",
            INIT_4D => X"0000003700000000ffffffe6ffffffffffffffe8ffffffff0000000000000000",
            INIT_4E => X"ffffffe3ffffffffffffff5cffffffffffffffd8fffffffffffffff4ffffffff",
            INIT_4F => X"0000000d000000000000000000000000ffffffbdffffffff0000000800000000",
            INIT_50 => X"0000000b0000000000000015000000000000001a00000000ffffffffffffffff",
            INIT_51 => X"0000000100000000fffffff7ffffffff0000001000000000ffffffcdffffffff",
            INIT_52 => X"ffffffb2ffffffffffffffe2ffffffff0000000100000000ffffffcdffffffff",
            INIT_53 => X"000000000000000000000052000000000000000000000000fffffff7ffffffff",
            INIT_54 => X"ffffffeeffffffffffffffddffffffffffffffe9ffffffff0000001300000000",
            INIT_55 => X"0000000c00000000ffffffcfffffffffffffffd9ffffffff0000000000000000",
            INIT_56 => X"ffffffe9ffffffffffffffa9ffffffffffffffc9ffffffffffffffeeffffffff",
            INIT_57 => X"fffffffbffffffff0000001c00000000fffffff7ffffffff0000001900000000",
            INIT_58 => X"ffffffdbffffffff0000000900000000fffffff8ffffffff0000000200000000",
            INIT_59 => X"0000001000000000fffffff6ffffffff0000001b000000000000000000000000",
            INIT_5A => X"ffffffc9ffffffffffffffeeffffffff0000002b00000000ffffffbaffffffff",
            INIT_5B => X"0000000300000000000000320000000000000008000000000000000c00000000",
            INIT_5C => X"0000000000000000fffffff8ffffffffffffffe3ffffffffffffffeeffffffff",
            INIT_5D => X"00000010000000000000001600000000ffffffb8fffffffffffffff7ffffffff",
            INIT_5E => X"ffffffc0ffffffffffffffd2ffffffffffffffb6ffffffffffffffb5ffffffff",
            INIT_5F => X"00000006000000000000000e000000000000001e00000000ffffffcbffffffff",
            INIT_60 => X"000000150000000000000002000000000000000c00000000fffffffaffffffff",
            INIT_61 => X"0000000300000000fffffffeffffffffffffffefffffffff0000000e00000000",
            INIT_62 => X"0000000400000000fffffff4fffffffffffffff5ffffffffffffffecffffffff",
            INIT_63 => X"ffffffffffffffff00000039000000000000000200000000ffffffe9ffffffff",
            INIT_64 => X"0000001d000000000000002a00000000ffffffe3fffffffffffffff3ffffffff",
            INIT_65 => X"0000002a00000000ffffffe9ffffffff0000000100000000ffffffd6ffffffff",
            INIT_66 => X"ffffffcbffffffffffffffefffffffffffffffe3ffffffffffffffc3ffffffff",
            INIT_67 => X"0000002c000000000000000900000000fffffff5ffffffffffffffd5ffffffff",
            INIT_68 => X"000000310000000000000026000000000000002400000000ffffffebffffffff",
            INIT_69 => X"0000000900000000ffffffe1ffffffffffffffe1ffffffff0000000f00000000",
            INIT_6A => X"0000000100000000fffffffefffffffffffffffdffffffffffffffe1ffffffff",
            INIT_6B => X"00000000000000000000001e00000000fffffffaffffffff0000000c00000000",
            INIT_6C => X"0000000e00000000ffffffe8ffffffff00000006000000000000003200000000",
            INIT_6D => X"00000020000000000000002000000000ffffffedfffffffffffffff4ffffffff",
            INIT_6E => X"ffffffcdffffffffffffffe9ffffffff0000002500000000ffffffdcffffffff",
            INIT_6F => X"00000032000000000000001a000000000000000b00000000ffffffd0ffffffff",
            INIT_70 => X"0000003b0000000000000019000000000000001200000000fffffff1ffffffff",
            INIT_71 => X"0000002200000000fffffff8fffffffffffffff3ffffffff0000000000000000",
            INIT_72 => X"ffffffe6ffffffff0000000c000000000000002900000000fffffff7ffffffff",
            INIT_73 => X"ffffffedfffffffffffffffcfffffffffffffff6ffffffff0000000800000000",
            INIT_74 => X"00000005000000000000002500000000ffffffefffffffff0000001a00000000",
            INIT_75 => X"fffffff3fffffffffffffff6ffffffffffffffc9ffffffff0000000100000000",
            INIT_76 => X"ffffffe5ffffffff00000009000000000000000f00000000ffffffc5ffffffff",
            INIT_77 => X"00000007000000000000001400000000fffffffcfffffffffffffff0ffffffff",
            INIT_78 => X"0000001800000000fffffffafffffffffffffff5ffffffff0000000c00000000",
            INIT_79 => X"0000000e00000000fffffffbfffffffffffffffeffffffff0000000b00000000",
            INIT_7A => X"0000001a0000000000000012000000000000001500000000ffffffdbffffffff",
            INIT_7B => X"ffffffe8ffffffffffffffb9ffffffffffffffe1ffffffff0000000300000000",
            INIT_7C => X"00000002000000000000001700000000ffffffd9ffffffff0000001d00000000",
            INIT_7D => X"0000000f00000000ffffffeaffffffffffffffcaffffffff0000001800000000",
            INIT_7E => X"ffffffceffffffff0000001300000000ffffffdcffffffffffffffd2ffffffff",
            INIT_7F => X"00000012000000000000001200000000ffffffe5fffffffffffffff4ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE20;


    MEM_IWGHT_LAYER2_INSTANCE21 : if BRAM_NAME = "iwght_layer2_instance21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000008000000000000000600000000fffffff6ffffffff0000000f00000000",
            INIT_01 => X"0000002400000000fffffffcffffffff0000001200000000ffffffe8ffffffff",
            INIT_02 => X"ffffffacffffffff00000017000000000000001100000000ffffffe8ffffffff",
            INIT_03 => X"00000005000000000000001700000000fffffff8ffffffff0000002100000000",
            INIT_04 => X"00000029000000000000001b00000000ffffffffffffffff0000001e00000000",
            INIT_05 => X"0000001300000000fffffffaffffffffffffffe8ffffffff0000004900000000",
            INIT_06 => X"ffffffd9ffffffffffffffb9ffffffffffffffb8ffffffffffffffd4ffffffff",
            INIT_07 => X"00000021000000000000000400000000ffffffdfffffffff0000003500000000",
            INIT_08 => X"0000000c00000000fffffff5ffffffff00000029000000000000000e00000000",
            INIT_09 => X"fffffff3ffffffff0000000c000000000000001300000000fffffff3ffffffff",
            INIT_0A => X"ffffffc6fffffffffffffff1ffffffffffffffedfffffffffffffff2ffffffff",
            INIT_0B => X"0000000b000000000000002a000000000000000000000000fffffff9ffffffff",
            INIT_0C => X"fffffff9fffffffffffffffcffffffffffffffe1ffffffff0000002700000000",
            INIT_0D => X"0000001300000000fffffffeffffffffffffffddffffffff0000003f00000000",
            INIT_0E => X"ffffffe0ffffffffffffffa8fffffffffffffffbffffffffffffffdcffffffff",
            INIT_0F => X"ffffffebfffffffffffffff8ffffffffffffffcbffffffff0000001b00000000",
            INIT_10 => X"ffffffedffffffff00000004000000000000000900000000fffffffaffffffff",
            INIT_11 => X"fffffff1fffffffffffffffdffffffff00000019000000000000000600000000",
            INIT_12 => X"0000000200000000fffffff2ffffffffffffffffffffffffffffffe5ffffffff",
            INIT_13 => X"0000000b000000000000001700000000ffffffe5ffffffffffffffecffffffff",
            INIT_14 => X"fffffff5ffffffff0000003500000000fffffff6ffffffffffffffffffffffff",
            INIT_15 => X"ffffffdfffffffff0000001700000000ffffffdcffffffff0000001e00000000",
            INIT_16 => X"fffffffbfffffffffffffff6fffffffffffffff4ffffffffffffffc6ffffffff",
            INIT_17 => X"00000016000000000000000000000000ffffffe5fffffffffffffff7ffffffff",
            INIT_18 => X"00000021000000000000000b00000000fffffff1fffffffffffffff4ffffffff",
            INIT_19 => X"fffffff1ffffffffffffffebffffffff0000001d000000000000000000000000",
            INIT_1A => X"ffffffc2ffffffff00000021000000000000001f00000000ffffffe9ffffffff",
            INIT_1B => X"00000000000000000000000e00000000ffffffeefffffffffffffffdffffffff",
            INIT_1C => X"ffffffdbffffffff0000001000000000ffffffdeffffffff0000002200000000",
            INIT_1D => X"fffffff9ffffffff0000000600000000ffffffb1fffffffffffffffeffffffff",
            INIT_1E => X"ffffffd2fffffffffffffff6ffffffffffffffb9ffffffffffffffddffffffff",
            INIT_1F => X"0000001f00000000fffffff3ffffffff00000008000000000000000300000000",
            INIT_20 => X"0000001600000000fffffff8fffffffffffffff8fffffffffffffffaffffffff",
            INIT_21 => X"0000000400000000fffffff1ffffffff0000001300000000fffffffaffffffff",
            INIT_22 => X"ffffffe5ffffffff00000000000000000000000600000000fffffff0ffffffff",
            INIT_23 => X"0000000400000000fffffff9ffffffffffffffe6fffffffffffffff7ffffffff",
            INIT_24 => X"ffffffc6ffffffff0000000c0000000000000007000000000000001f00000000",
            INIT_25 => X"ffffffe1fffffffffffffff5ffffffffffffffa4ffffffff0000001500000000",
            INIT_26 => X"ffffffd1ffffffffffffffeaffffffffffffffd8fffffffffffffff6ffffffff",
            INIT_27 => X"0000001e000000000000000b00000000ffffffdfffffffffffffffddffffffff",
            INIT_28 => X"0000001800000000fffffff0fffffffffffffff6ffffffff0000000600000000",
            INIT_29 => X"0000000800000000fffffffcffffffff0000000f000000000000000200000000",
            INIT_2A => X"00000006000000000000001c00000000fffffffcfffffffffffffff6ffffffff",
            INIT_2B => X"0000000000000000ffffffedfffffffffffffff1ffffffff0000000e00000000",
            INIT_2C => X"ffffffd8ffffffff0000001b00000000ffffffbbffffffff0000001c00000000",
            INIT_2D => X"ffffffe6fffffffffffffff3ffffffffffffffc9ffffffff0000002600000000",
            INIT_2E => X"ffffffccffffffff0000000200000000fffffff0ffffffffffffffbfffffffff",
            INIT_2F => X"0000000b000000000000000100000000fffffffaffffffff0000000400000000",
            INIT_30 => X"0000002800000000000000070000000000000019000000000000001100000000",
            INIT_31 => X"00000002000000000000000a000000000000001900000000ffffffdbffffffff",
            INIT_32 => X"00000009000000000000001b000000000000000600000000ffffffddffffffff",
            INIT_33 => X"fffffffeffffffffffffffd9ffffffffffffffe0ffffffff0000002700000000",
            INIT_34 => X"0000001a000000000000002300000000ffffffd0ffffffff0000002800000000",
            INIT_35 => X"ffffffe3ffffffff0000000a00000000ffffff9bffffffff0000001400000000",
            INIT_36 => X"ffffffdffffffffffffffff6ffffffffffffffc6ffffffffffffffd9ffffffff",
            INIT_37 => X"00000016000000000000001900000000ffffffdfffffffff0000000000000000",
            INIT_38 => X"0000000c00000000ffffffe7ffffffff00000012000000000000001600000000",
            INIT_39 => X"0000000c000000000000000b000000000000002b00000000ffffffdbffffffff",
            INIT_3A => X"ffffffeffffffffffffffff4ffffffff0000000900000000ffffffdbffffffff",
            INIT_3B => X"0000000a00000000fffffff4fffffffffffffffafffffffffffffffeffffffff",
            INIT_3C => X"0000000b00000000000000150000000000000002000000000000000600000000",
            INIT_3D => X"ffffffdcffffffff000000160000000000000014000000000000001d00000000",
            INIT_3E => X"0000000f000000000000003600000000fffffff5fffffffffffffffeffffffff",
            INIT_3F => X"ffffffdeffffffffffffffddffffffff00000010000000000000000100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffffafffffffffffffffafffffffffffffffcffffffffffffffd3ffffffff",
            INIT_41 => X"ffffffe4ffffffffffffffebffffffff0000001500000000fffffff2ffffffff",
            INIT_42 => X"ffffffeeffffffffffffffcdffffffff0000001d00000000ffffffb4ffffffff",
            INIT_43 => X"0000000400000000000000220000000000000009000000000000000d00000000",
            INIT_44 => X"ffffffdcfffffffffffffff9ffffffff00000027000000000000002200000000",
            INIT_45 => X"ffffffe2ffffffff0000001300000000fffffffaffffffff0000000700000000",
            INIT_46 => X"fffffffcffffffff0000002e0000000000000004000000000000001a00000000",
            INIT_47 => X"ffffffeaffffffffffffffdafffffffffffffffeffffffff0000001e00000000",
            INIT_48 => X"00000019000000000000000000000000ffffffd6ffffffffffffffd2ffffffff",
            INIT_49 => X"ffffffdfffffffffffffffeafffffffffffffffaffffffff0000000800000000",
            INIT_4A => X"ffffffd1ffffffffffffffe9ffffffff0000000700000000ffffffddffffffff",
            INIT_4B => X"00000000000000000000003f00000000fffffff3ffffffff0000002000000000",
            INIT_4C => X"0000000d00000000fffffff3ffffffff00000037000000000000000f00000000",
            INIT_4D => X"00000000000000000000001400000000fffffff3ffffffff0000001700000000",
            INIT_4E => X"fffffffcfffffffffffffff5ffffffff0000003a00000000fffffffdffffffff",
            INIT_4F => X"ffffffdfffffffffffffffeffffffffffffffff4ffffffff0000001d00000000",
            INIT_50 => X"00000012000000000000003e00000000ffffffffffffffffffffffe7ffffffff",
            INIT_51 => X"ffffffc7ffffffff00000000000000000000000400000000ffffffecffffffff",
            INIT_52 => X"000000020000000000000000000000000000000800000000fffffff1ffffffff",
            INIT_53 => X"ffffffceffffffff0000001b00000000ffffffd3ffffffff0000002300000000",
            INIT_54 => X"0000004900000000ffffffe8ffffffff0000000e000000000000000300000000",
            INIT_55 => X"ffffffb0ffffffff0000000a0000000000000019000000000000002400000000",
            INIT_56 => X"ffffffe5ffffffff00000007000000000000000a000000000000000400000000",
            INIT_57 => X"ffffffebffffffff0000000700000000ffffffddffffffffffffffebffffffff",
            INIT_58 => X"000000120000000000000003000000000000002400000000ffffffe3ffffffff",
            INIT_59 => X"fffffff0fffffffffffffff4ffffffff0000000c00000000fffffff9ffffffff",
            INIT_5A => X"0000001e000000000000000e000000000000001500000000ffffffe0ffffffff",
            INIT_5B => X"ffffffecffffffffffffffd7ffffffffffffffd5ffffffff0000002900000000",
            INIT_5C => X"0000000b0000000000000000000000000000002600000000ffffffeaffffffff",
            INIT_5D => X"ffffffb9ffffffff000000030000000000000021000000000000001900000000",
            INIT_5E => X"fffffff3ffffffff0000002200000000ffffffd5ffffffffffffffe2ffffffff",
            INIT_5F => X"fffffffdfffffffffffffffcfffffffffffffff9ffffffffffffffe8ffffffff",
            INIT_60 => X"000000090000000000000000000000000000001e00000000ffffffdaffffffff",
            INIT_61 => X"ffffffe1ffffffffffffffefffffffff0000001900000000fffffff1ffffffff",
            INIT_62 => X"0000002600000000ffffffe9ffffffff0000001b00000000fffffff4ffffffff",
            INIT_63 => X"fffffff8ffffffff0000000000000000fffffff8ffffffff0000001800000000",
            INIT_64 => X"ffffffbeffffffff000000210000000000000005000000000000000200000000",
            INIT_65 => X"ffffffd4ffffffff000000190000000000000010000000000000000200000000",
            INIT_66 => X"fffffff1ffffffff0000001b0000000000000011000000000000000b00000000",
            INIT_67 => X"0000000800000000ffffffddffffffff0000001900000000ffffffeaffffffff",
            INIT_68 => X"0000001600000000ffffffd4ffffffff0000000600000000ffffffcfffffffff",
            INIT_69 => X"ffffffe7ffffffff00000008000000000000001600000000fffffff5ffffffff",
            INIT_6A => X"0000000800000000ffffffe9ffffffff00000013000000000000001700000000",
            INIT_6B => X"ffffffefffffffff000000200000000000000021000000000000001000000000",
            INIT_6C => X"ffffffd1ffffffff0000000200000000ffffffeaffffffff0000000c00000000",
            INIT_6D => X"ffffffc6ffffffff00000032000000000000002500000000ffffffe7ffffffff",
            INIT_6E => X"fffffff6ffffffffffffffd5ffffffff00000029000000000000003600000000",
            INIT_6F => X"ffffffe5ffffffffffffffe3ffffffff0000001f00000000fffffff4ffffffff",
            INIT_70 => X"0000002a00000000ffffffbfffffffffffffffe0ffffffffffffffe5ffffffff",
            INIT_71 => X"fffffff3ffffffffffffffecffffffff0000001300000000ffffffbfffffffff",
            INIT_72 => X"000000080000000000000020000000000000000b00000000ffffffc9ffffffff",
            INIT_73 => X"fffffff6ffffffffffffffdfffffffffffffffdbffffffff0000001300000000",
            INIT_74 => X"fffffff6ffffffff0000000000000000ffffffd2fffffffffffffff0ffffffff",
            INIT_75 => X"ffffff8fffffffff00000028000000000000000d000000000000000700000000",
            INIT_76 => X"00000008000000000000002d00000000ffffffc9ffffffffffffffd9ffffffff",
            INIT_77 => X"000000100000000000000001000000000000000000000000fffffff8ffffffff",
            INIT_78 => X"ffffffecffffffff0000000000000000ffffffeeffffffff0000000800000000",
            INIT_79 => X"fffffffafffffffffffffff8ffffffff0000000d00000000fffffffdffffffff",
            INIT_7A => X"ffffffd6ffffffff00000013000000000000000b00000000ffffffefffffffff",
            INIT_7B => X"fffffff2ffffffff000000100000000000000001000000000000001300000000",
            INIT_7C => X"fffffffeffffffff00000000000000000000001300000000fffffffdffffffff",
            INIT_7D => X"0000000000000000000000110000000000000003000000000000000700000000",
            INIT_7E => X"000000170000000000000026000000000000001200000000ffffffefffffffff",
            INIT_7F => X"0000001800000000fffffff5ffffffff00000024000000000000001500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE21;


    MEM_IWGHT_LAYER2_INSTANCE22 : if BRAM_NAME = "iwght_layer2_instance22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffeefffffffffffffffffffffffffffffffefffffffffffffff7ffffffff",
            INIT_01 => X"0000000000000000ffffffd3ffffffffffffffe3ffffffff0000002100000000",
            INIT_02 => X"ffffffccfffffffffffffff7fffffffffffffff1ffffffff0000002000000000",
            INIT_03 => X"ffffffecffffffff000000390000000000000019000000000000000800000000",
            INIT_04 => X"ffffffe5ffffffffffffffebffffffff00000049000000000000002400000000",
            INIT_05 => X"ffffffe3ffffffffffffffffffffffffffffffeafffffffffffffff4ffffffff",
            INIT_06 => X"0000001d00000000ffffffd3ffffffff0000004e000000000000000400000000",
            INIT_07 => X"ffffffd4ffffffff000000040000000000000009000000000000001a00000000",
            INIT_08 => X"00000009000000000000004000000000ffffffe9ffffffffffffffedffffffff",
            INIT_09 => X"fffffff9ffffffffffffffd3fffffffffffffff2ffffffffffffffe0ffffffff",
            INIT_0A => X"ffffffeeffffffff0000002b000000000000000000000000ffffffedffffffff",
            INIT_0B => X"ffffffe8ffffffff0000000100000000fffffffffffffffffffffffeffffffff",
            INIT_0C => X"0000001600000000000000040000000000000026000000000000000600000000",
            INIT_0D => X"0000002200000000ffffffeefffffffffffffffcffffffff0000000400000000",
            INIT_0E => X"0000000a00000000ffffffceffffffffffffffd3ffffffffffffffe6ffffffff",
            INIT_0F => X"fffffff0fffffffffffffffaffffffffffffffe7ffffffff0000000200000000",
            INIT_10 => X"ffffffdeffffffff0000004b000000000000001f00000000fffffff0ffffffff",
            INIT_11 => X"fffffffafffffffffffffffcfffffffffffffffeffffffff0000001700000000",
            INIT_12 => X"0000001f000000000000003f000000000000000700000000ffffffe6ffffffff",
            INIT_13 => X"0000000400000000ffffffcdfffffffffffffff2ffffffff0000000400000000",
            INIT_14 => X"fffffffeffffffff00000028000000000000000d00000000ffffffe3ffffffff",
            INIT_15 => X"0000001c00000000fffffff8ffffffffffffffecffffffff0000000800000000",
            INIT_16 => X"ffffffd9ffffffff0000003100000000ffffffb4fffffffffffffffdffffffff",
            INIT_17 => X"0000000d00000000ffffffe1ffffffffffffffe6ffffffffffffffc0ffffffff",
            INIT_18 => X"0000001200000000000000320000000000000012000000000000000000000000",
            INIT_19 => X"fffffff3ffffffffffffffebffffffffffffffd5ffffffff0000000d00000000",
            INIT_1A => X"fffffff1ffffffff0000001000000000ffffffeaffffffffffffffcdffffffff",
            INIT_1B => X"000000000000000000000008000000000000001b000000000000000d00000000",
            INIT_1C => X"ffffffe7ffffffff000000210000000000000041000000000000002b00000000",
            INIT_1D => X"ffffffe0fffffffffffffffbffffffffffffffefffffffff0000001400000000",
            INIT_1E => X"00000016000000000000002d000000000000001900000000fffffff6ffffffff",
            INIT_1F => X"fffffff7ffffffffffffffebffffffff00000009000000000000000500000000",
            INIT_20 => X"00000000000000000000000a00000000ffffffeafffffffffffffff8ffffffff",
            INIT_21 => X"0000001000000000ffffffdffffffffffffffffeffffffffffffffdbffffffff",
            INIT_22 => X"ffffffefffffffffffffffe7ffffffff00000008000000000000000200000000",
            INIT_23 => X"ffffffd6ffffffff0000002c00000000ffffffe6ffffffff0000000000000000",
            INIT_24 => X"0000000600000000ffffffe1ffffffff0000000c000000000000000f00000000",
            INIT_25 => X"ffffffeaffffffff0000001800000000fffffffbffffffffffffffeeffffffff",
            INIT_26 => X"fffffff7fffffffffffffff5ffffffff00000015000000000000001200000000",
            INIT_27 => X"ffffffcbffffffff0000000d0000000000000013000000000000002700000000",
            INIT_28 => X"000000120000000000000000000000000000000000000000fffffffaffffffff",
            INIT_29 => X"0000000a00000000ffffffdfffffffffffffffe7ffffffff0000002a00000000",
            INIT_2A => X"0000001a000000000000003800000000ffffffffffffffff0000000d00000000",
            INIT_2B => X"fffffff6ffffffffffffffdeffffffffffffffe0ffffffff0000000e00000000",
            INIT_2C => X"0000000900000000fffffffbfffffffffffffff5ffffffffffffffceffffffff",
            INIT_2D => X"ffffffbaffffffff00000044000000000000001100000000fffffff1ffffffff",
            INIT_2E => X"ffffffd2ffffffff00000059000000000000000a00000000ffffffd1ffffffff",
            INIT_2F => X"0000001a000000000000001e0000000000000053000000000000000900000000",
            INIT_30 => X"fffffff0ffffffffffffffeafffffffffffffffcffffffff0000000c00000000",
            INIT_31 => X"ffffffe4fffffffffffffff1fffffffffffffff0ffffffff0000001400000000",
            INIT_32 => X"0000001c000000000000002c000000000000000f00000000ffffffccffffffff",
            INIT_33 => X"0000000700000000fffffffcfffffffffffffff2ffffffff0000000700000000",
            INIT_34 => X"0000001b00000000fffffff9ffffffff0000004000000000ffffffe0ffffffff",
            INIT_35 => X"000000000000000000000009000000000000000a00000000fffffffbffffffff",
            INIT_36 => X"ffffffe4ffffffff00000028000000000000001e00000000ffffffecffffffff",
            INIT_37 => X"0000002200000000fffffff9ffffffff0000002000000000fffffff8ffffffff",
            INIT_38 => X"ffffffebffffffff0000000d0000000000000014000000000000001000000000",
            INIT_39 => X"0000000b00000000ffffffedffffffffffffffddffffffff0000000b00000000",
            INIT_3A => X"ffffffe5fffffffffffffff9ffffffffffffffffffffffffffffffefffffffff",
            INIT_3B => X"0000000b0000000000000019000000000000001300000000ffffff85ffffffff",
            INIT_3C => X"0000000c0000000000000006000000000000004d000000000000002a00000000",
            INIT_3D => X"0000003600000000ffffffc8ffffffffffffffe0ffffffff0000000f00000000",
            INIT_3E => X"ffffffaffffffffffffffffbffffffffffffffe1ffffffffffffffc3ffffffff",
            INIT_3F => X"0000000000000000fffffffeffffffffffffffe1ffffffffffffffc7ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffddffffffff0000001e00000000fffffffaffffffffffffffe6ffffffff",
            INIT_41 => X"0000001300000000ffffffd5fffffffffffffffbffffffff0000000600000000",
            INIT_42 => X"fffffff0ffffffff0000002d00000000fffffffdffffffffffffffe8ffffffff",
            INIT_43 => X"000000120000000000000011000000000000001e00000000ffffff7affffffff",
            INIT_44 => X"00000014000000000000001e0000000000000035000000000000002800000000",
            INIT_45 => X"0000000600000000ffffffc8ffffffff00000016000000000000004f00000000",
            INIT_46 => X"ffffffe0ffffffffffffffd5ffffffffffffffabffffffffffffffd6ffffffff",
            INIT_47 => X"ffffffeafffffffffffffff2ffffffffffffffc9ffffffffffffffc8ffffffff",
            INIT_48 => X"fffffff6ffffffff00000033000000000000001600000000ffffffbbffffffff",
            INIT_49 => X"0000000400000000fffffffaffffffff00000008000000000000001700000000",
            INIT_4A => X"00000000000000000000002b000000000000002100000000fffffff4ffffffff",
            INIT_4B => X"0000002300000000ffffffdafffffffffffffffcffffffffffffff8fffffffff",
            INIT_4C => X"fffffffbffffffff000000450000000000000013000000000000001800000000",
            INIT_4D => X"ffffffbfffffffffffffffb3fffffffffffffff8ffffffff0000003f00000000",
            INIT_4E => X"ffffffcbffffffff0000004700000000ffffffb6ffffffffffffffbcffffffff",
            INIT_4F => X"fffffff4fffffffffffffff0ffffffffffffffc5ffffffffffffffbbffffffff",
            INIT_50 => X"ffffffe8ffffffff0000003a00000000fffffff9ffffffffffffffe6ffffffff",
            INIT_51 => X"00000005000000000000000c00000000ffffffe6ffffffffffffffffffffffff",
            INIT_52 => X"fffffff3ffffffff0000001900000000fffffffcffffffffffffffe0ffffffff",
            INIT_53 => X"0000000a00000000fffffff8fffffffffffffffeffffffffffffffd1ffffffff",
            INIT_54 => X"0000001a00000000000000100000000000000026000000000000002f00000000",
            INIT_55 => X"0000000300000000ffffffb9ffffffffffffffefffffffff0000000b00000000",
            INIT_56 => X"ffffffe4ffffffff0000003400000000ffffffc8ffffffff0000000400000000",
            INIT_57 => X"ffffffe1ffffffff0000000500000000ffffffb4fffffffffffffff3ffffffff",
            INIT_58 => X"ffffffe1ffffffff0000001b000000000000000c00000000ffffffeaffffffff",
            INIT_59 => X"0000000800000000fffffff2fffffffffffffff3ffffffffffffffffffffffff",
            INIT_5A => X"fffffffcffffffffffffffc8ffffffff0000001a00000000ffffffffffffffff",
            INIT_5B => X"ffffffe0ffffffff0000003d00000000fffffffdffffffff0000000600000000",
            INIT_5C => X"0000002700000000ffffffccffffffff0000002e000000000000001c00000000",
            INIT_5D => X"ffffffd6ffffffff0000002900000000ffffffdeffffffff0000000200000000",
            INIT_5E => X"ffffffdcffffffffffffffe6ffffffff00000032000000000000000e00000000",
            INIT_5F => X"ffffffe8ffffffff000000010000000000000035000000000000002c00000000",
            INIT_60 => X"fffffff6ffffffff00000018000000000000000100000000fffffff6ffffffff",
            INIT_61 => X"0000000f00000000ffffffdbffffffff00000007000000000000001400000000",
            INIT_62 => X"000000470000000000000012000000000000000d00000000ffffffe8ffffffff",
            INIT_63 => X"fffffffdffffffffffffffc7ffffffff0000000d000000000000001700000000",
            INIT_64 => X"0000000b00000000ffffffebffffffff0000001e00000000ffffffd0ffffffff",
            INIT_65 => X"ffffffc7ffffffff00000039000000000000000c00000000ffffffe9ffffffff",
            INIT_66 => X"0000002d000000000000000d00000000ffffffefffffffffffffffe5ffffffff",
            INIT_67 => X"fffffffdffffffff000000150000000000000026000000000000000c00000000",
            INIT_68 => X"ffffffd5ffffffffffffffffffffffffffffffe2ffffffff0000000d00000000",
            INIT_69 => X"00000000000000000000001700000000fffffff9fffffffffffffffdffffffff",
            INIT_6A => X"000000280000000000000037000000000000000700000000ffffffdfffffffff",
            INIT_6B => X"0000000200000000ffffffd8fffffffffffffff1fffffffffffffff3ffffffff",
            INIT_6C => X"0000003a0000000000000000000000000000000400000000fffffff3ffffffff",
            INIT_6D => X"ffffffc7fffffffffffffffcffffffffffffffe2fffffffffffffff2ffffffff",
            INIT_6E => X"00000005000000000000004a000000000000004500000000ffffffbaffffffff",
            INIT_6F => X"fffffff3ffffffff0000001b00000000ffffffd2ffffffffffffffc9ffffffff",
            INIT_70 => X"00000021000000000000001d0000000000000023000000000000000b00000000",
            INIT_71 => X"00000001000000000000000000000000ffffffe6ffffffffffffffe1ffffffff",
            INIT_72 => X"fffffff0ffffffff0000002500000000ffffffe5ffffffffffffffcbffffffff",
            INIT_73 => X"00000017000000000000002000000000fffffffcffffffffffffffa1ffffffff",
            INIT_74 => X"0000001d0000000000000003000000000000003f000000000000000c00000000",
            INIT_75 => X"0000004b00000000ffffffc5ffffffff00000019000000000000001600000000",
            INIT_76 => X"ffffffd7ffffffff0000001700000000ffffffe9ffffffffffffffbcffffffff",
            INIT_77 => X"ffffffe7ffffffff0000000e00000000ffffffe3ffffffffffffffecffffffff",
            INIT_78 => X"ffffffd7ffffffff00000021000000000000001a00000000fffffff5ffffffff",
            INIT_79 => X"fffffff6ffffffffffffffc4ffffffffffffffdeffffffff0000000300000000",
            INIT_7A => X"ffffffebffffffff00000021000000000000001100000000ffffffffffffffff",
            INIT_7B => X"0000002400000000fffffff7ffffffff0000001600000000ffffff84ffffffff",
            INIT_7C => X"000000230000000000000016000000000000001b000000000000003f00000000",
            INIT_7D => X"0000004700000000ffffffecffffffff0000001a000000000000002100000000",
            INIT_7E => X"ffffffc3fffffffffffffffcffffffffffffffc2ffffffffffffffc5ffffffff",
            INIT_7F => X"ffffffe7ffffffffffffffffffffffffffffffecffffffffffffffcaffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE22;


    MEM_IWGHT_LAYER2_INSTANCE23 : if BRAM_NAME = "iwght_layer2_instance23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffe7ffffffffffffffe2ffffffffffffffe7ffffffffffffffc3ffffffff",
            INIT_01 => X"ffffffe3ffffffffffffffd3ffffffffffffffcffffffffffffffffdffffffff",
            INIT_02 => X"0000000b0000000000000030000000000000000c000000000000001e00000000",
            INIT_03 => X"0000002200000000ffffffc7ffffffff0000000b00000000ffffffa6ffffffff",
            INIT_04 => X"0000001b000000000000002d0000000000000023000000000000003800000000",
            INIT_05 => X"0000003000000000ffffffb6ffffffffffffffffffffffff0000000000000000",
            INIT_06 => X"ffffff8bffffffff0000003f00000000ffffffbcfffffffffffffff9ffffffff",
            INIT_07 => X"ffffffeeffffffff0000000500000000ffffffb5ffffffffffffffcbffffffff",
            INIT_08 => X"ffffffe0ffffffffffffffe4ffffffffffffffebffffffffffffffdaffffffff",
            INIT_09 => X"0000001700000000ffffffd5ffffffffffffffd8ffffffffffffffdfffffffff",
            INIT_0A => X"0000000900000000000000020000000000000017000000000000000700000000",
            INIT_0B => X"fffffffcffffffff0000001400000000ffffffffffffffffffffffceffffffff",
            INIT_0C => X"0000000d00000000ffffffd6ffffffff00000059000000000000001000000000",
            INIT_0D => X"fffffffeffffffffffffffd4ffffffff0000000c00000000ffffffecffffffff",
            INIT_0E => X"0000000700000000fffffff0ffffffffffffffcbffffffffffffffecffffffff",
            INIT_0F => X"fffffff1fffffffffffffffdffffffffffffffc3ffffffff0000000200000000",
            INIT_10 => X"fffffffeffffffff00000018000000000000000500000000ffffffe9ffffffff",
            INIT_11 => X"0000000700000000ffffffe4ffffffff00000000000000000000000800000000",
            INIT_12 => X"ffffffe5ffffffff0000000100000000fffffff3ffffffffffffffe3ffffffff",
            INIT_13 => X"ffffffe4ffffffff000000350000000000000002000000000000001400000000",
            INIT_14 => X"0000000400000000ffffffc5fffffffffffffffdffffffff0000001000000000",
            INIT_15 => X"000000190000000000000011000000000000000400000000fffffffbffffffff",
            INIT_16 => X"0000001100000000ffffffaefffffffffffffff4fffffffffffffff0ffffffff",
            INIT_17 => X"ffffffedffffffff000000130000000000000000000000000000002300000000",
            INIT_18 => X"ffffffd9ffffffff0000000e0000000000000001000000000000000c00000000",
            INIT_19 => X"00000014000000000000000400000000fffffff3ffffffffffffffe9ffffffff",
            INIT_1A => X"00000029000000000000001f00000000ffffffe5fffffffffffffff3ffffffff",
            INIT_1B => X"0000001a00000000ffffffd0ffffffff0000000e000000000000001500000000",
            INIT_1C => X"00000016000000000000001d000000000000000200000000ffffffd3ffffffff",
            INIT_1D => X"ffffffecffffffff0000001b00000000fffffffeffffffffffffffe8ffffffff",
            INIT_1E => X"00000026000000000000003d000000000000001b000000000000001000000000",
            INIT_1F => X"ffffffecffffffff0000001c000000000000001f000000000000000000000000",
            INIT_20 => X"ffffffedfffffffffffffff1ffffffffffffffedffffffff0000001e00000000",
            INIT_21 => X"ffffffebffffffff00000001000000000000001200000000fffffffcffffffff",
            INIT_22 => X"0000003b000000000000003600000000fffffffdfffffffffffffff3ffffffff",
            INIT_23 => X"fffffff4ffffffffffffffb6fffffffffffffffeffffffff0000002200000000",
            INIT_24 => X"00000029000000000000002b00000000ffffffe0fffffffffffffff8ffffffff",
            INIT_25 => X"0000000100000000ffffffc4fffffffffffffff4ffffffff0000001300000000",
            INIT_26 => X"000000090000000000000037000000000000000a00000000ffffffeaffffffff",
            INIT_27 => X"fffffffcffffffff0000000d00000000ffffffa8ffffffffffffffd1ffffffff",
            INIT_28 => X"ffffffd3ffffffff000000080000000000000031000000000000001c00000000",
            INIT_29 => X"00000009000000000000002d00000000ffffffffffffffffffffffb9ffffffff",
            INIT_2A => X"0000002f000000000000002600000000ffffffe4ffffffffffffffc5ffffffff",
            INIT_2B => X"ffffffe4fffffffffffffff5ffffffff00000009000000000000001d00000000",
            INIT_2C => X"0000002700000000ffffffdeffffffff00000009000000000000000700000000",
            INIT_2D => X"ffffffe6ffffffffffffffc6ffffffffffffffefffffffff0000001300000000",
            INIT_2E => X"00000009000000000000003900000000ffffffb1ffffffffffffffeaffffffff",
            INIT_2F => X"ffffffefffffffff0000000200000000ffffffb8ffffffff0000000600000000",
            INIT_30 => X"ffffffdbffffffffffffffc1ffffffff0000001a000000000000001400000000",
            INIT_31 => X"0000000800000000fffffff1fffffffffffffff6ffffffffffffffd4ffffffff",
            INIT_32 => X"0000003a000000000000000c00000000fffffff6ffffffffffffffd9ffffffff",
            INIT_33 => X"ffffffeaffffffff0000001300000000fffffffeffffffff0000001800000000",
            INIT_34 => X"0000002a00000000ffffffd2ffffffff0000004800000000fffffffdffffffff",
            INIT_35 => X"fffffffaffffffff0000000500000000ffffffe9ffffffff0000000a00000000",
            INIT_36 => X"fffffff8ffffffff0000002e00000000ffffffddffffffff0000001c00000000",
            INIT_37 => X"fffffff5ffffffff00000021000000000000001d000000000000002600000000",
            INIT_38 => X"fffffff3ffffffffffffffd8ffffffff0000001400000000ffffffffffffffff",
            INIT_39 => X"0000001800000000ffffffc4ffffffffffffffdafffffffffffffff1ffffffff",
            INIT_3A => X"000000140000000000000025000000000000000000000000fffffffdffffffff",
            INIT_3B => X"fffffff3fffffffffffffffdffffffff00000004000000000000000400000000",
            INIT_3C => X"0000003e00000000ffffffd2ffffffff0000002b00000000fffffff0ffffffff",
            INIT_3D => X"0000001f00000000fffffff6ffffffff00000015000000000000001800000000",
            INIT_3E => X"0000000f000000000000000f00000000ffffffe9ffffffffffffffd6ffffffff",
            INIT_3F => X"000000070000000000000003000000000000000500000000ffffffd7ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffebffffffffffffffc0fffffffffffffff7ffffffff0000000000000000",
            INIT_41 => X"0000001300000000fffffffeffffffffffffffe4fffffffffffffff8ffffffff",
            INIT_42 => X"fffffff9ffffffff0000000200000000fffffff9ffffffff0000001a00000000",
            INIT_43 => X"ffffffdbffffffff0000003100000000fffffff2ffffffff0000001600000000",
            INIT_44 => X"0000002200000000ffffffd3ffffffff00000034000000000000001c00000000",
            INIT_45 => X"0000002900000000ffffffc2ffffffff0000001b000000000000000e00000000",
            INIT_46 => X"0000001600000000ffffffadfffffffffffffffaffffffffffffffcaffffffff",
            INIT_47 => X"fffffff7fffffffffffffff8ffffffffffffffc4fffffffffffffffaffffffff",
            INIT_48 => X"ffffffeeffffffff00000004000000000000002800000000fffffffbffffffff",
            INIT_49 => X"fffffffefffffffffffffffaffffffff0000000800000000ffffffdcffffffff",
            INIT_4A => X"ffffffddffffffffffffffebffffffffffffffffffffffff0000000600000000",
            INIT_4B => X"000000090000000000000031000000000000000e00000000fffffffeffffffff",
            INIT_4C => X"0000000700000000ffffffe1fffffffffffffff9ffffffff0000001200000000",
            INIT_4D => X"0000003500000000ffffffe0ffffffff0000002f000000000000001200000000",
            INIT_4E => X"0000000c00000000ffffffa4fffffffffffffff1fffffffffffffff1ffffffff",
            INIT_4F => X"fffffffeffffffff0000001000000000ffffffdfffffffff0000000600000000",
            INIT_50 => X"ffffffbaffffffffffffffe0fffffffffffffffcffffffff0000001600000000",
            INIT_51 => X"0000000b00000000ffffffffffffffff0000000c00000000ffffffddffffffff",
            INIT_52 => X"0000002a0000000000000033000000000000002400000000fffffff8ffffffff",
            INIT_53 => X"0000002100000000ffffffb9ffffffff0000001a00000000fffffffeffffffff",
            INIT_54 => X"000000150000000000000013000000000000002100000000ffffffe4ffffffff",
            INIT_55 => X"ffffffd6ffffffff0000001b00000000fffffff8ffffffff0000000b00000000",
            INIT_56 => X"0000001a000000000000002200000000ffffffd4ffffffff0000002200000000",
            INIT_57 => X"00000025000000000000001f000000000000003f00000000ffffffefffffffff",
            INIT_58 => X"fffffffcffffffffffffffe1fffffffffffffffdffffffff0000000800000000",
            INIT_59 => X"00000000000000000000000300000000ffffffeeffffffff0000000e00000000",
            INIT_5A => X"0000002e000000000000002400000000ffffffe8ffffffff0000000c00000000",
            INIT_5B => X"ffffffffffffffffffffffb4ffffffffffffffe7ffffffff0000000700000000",
            INIT_5C => X"0000003a000000000000002300000000ffffffe2fffffffffffffffdffffffff",
            INIT_5D => X"ffffffb9ffffffffffffffe1ffffffffffffffdfffffffff0000002000000000",
            INIT_5E => X"fffffff2ffffffff0000001d00000000ffffffb4ffffffff0000001000000000",
            INIT_5F => X"fffffff9fffffffffffffffcffffffffffffffedffffffffffffffd9ffffffff",
            INIT_60 => X"ffffffedffffffffffffffd1ffffffff00000003000000000000000e00000000",
            INIT_61 => X"00000001000000000000001e000000000000001c00000000fffffff0ffffffff",
            INIT_62 => X"00000035000000000000001900000000ffffffe9ffffffffffffffddffffffff",
            INIT_63 => X"ffffffeaffffffffffffffe8ffffffffffffffebffffffff0000002c00000000",
            INIT_64 => X"00000031000000000000000500000000ffffffdffffffffffffffff5ffffffff",
            INIT_65 => X"ffffffbfffffffffffffffd5ffffffffffffffecffffffff0000001c00000000",
            INIT_66 => X"0000000a000000000000001700000000ffffffa5ffffffff0000000f00000000",
            INIT_67 => X"0000000600000000ffffffffffffffffffffffe2ffffffffffffffefffffffff",
            INIT_68 => X"ffffffddffffffffffffffbcffffffff0000000b000000000000002200000000",
            INIT_69 => X"00000007000000000000001c000000000000001e00000000ffffffcfffffffff",
            INIT_6A => X"0000002300000000ffffffeeffffffff0000001000000000ffffffc2ffffffff",
            INIT_6B => X"fffffff3ffffffff000000000000000000000004000000000000004e00000000",
            INIT_6C => X"0000001100000000ffffffcfffffffff0000000200000000ffffffe1ffffffff",
            INIT_6D => X"ffffffdfffffffffffffffe8ffffffff00000011000000000000001100000000",
            INIT_6E => X"0000001200000000fffffff0ffffffffffffffa1ffffffff0000003500000000",
            INIT_6F => X"fffffff0ffffffff0000000c00000000ffffffe9ffffffff0000001800000000",
            INIT_70 => X"ffffffc6ffffffffffffffc4ffffffff00000021000000000000002900000000",
            INIT_71 => X"000000270000000000000000000000000000000d00000000ffffffe1ffffffff",
            INIT_72 => X"00000001000000000000000000000000fffffffaffffffffffffffdfffffffff",
            INIT_73 => X"ffffffe0ffffffff0000002c000000000000000e000000000000002000000000",
            INIT_74 => X"0000002900000000ffffffbbffffffff0000000100000000fffffffbffffffff",
            INIT_75 => X"ffffffeffffffffffffffff5ffffffff0000000b000000000000002800000000",
            INIT_76 => X"0000001a00000000ffffff9affffffffffffffe9ffffffffffffffffffffffff",
            INIT_77 => X"fffffff9ffffffff0000001500000000fffffffdffffffff0000003e00000000",
            INIT_78 => X"ffffffd5ffffffffffffffc3ffffffff00000000000000000000001000000000",
            INIT_79 => X"00000006000000000000002a000000000000001300000000ffffffcfffffffff",
            INIT_7A => X"0000001900000000ffffffe7ffffffffffffffdffffffffffffffff4ffffffff",
            INIT_7B => X"00000007000000000000002400000000fffffff3ffffffff0000000500000000",
            INIT_7C => X"0000003b00000000ffffffdaffffffff0000001000000000ffffffe3ffffffff",
            INIT_7D => X"0000004300000000ffffffe4ffffffff0000000a000000000000001400000000",
            INIT_7E => X"fffffffbffffffffffffffbeffffffffffffffbffffffffffffffff4ffffffff",
            INIT_7F => X"fffffffdfffffffffffffff8ffffffffffffffd5fffffffffffffffdffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE23;


    MEM_IWGHT_LAYER2_INSTANCE24 : if BRAM_NAME = "iwght_layer2_instance24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffff9cffffffffffffffc9ffffffff00000021000000000000001300000000",
            INIT_01 => X"ffffffe9ffffffff00000005000000000000001600000000ffffffd0ffffffff",
            INIT_02 => X"fffffff9ffffffff0000000e00000000ffffffedffffffffffffffd6ffffffff",
            INIT_03 => X"0000001f0000000000000028000000000000002500000000ffffffeaffffffff",
            INIT_04 => X"0000002c00000000fffffff9ffffffff00000014000000000000001200000000",
            INIT_05 => X"0000003100000000fffffff9ffffffff0000000f000000000000001900000000",
            INIT_06 => X"ffffffeeffffffffffffffdeffffffffffffff91ffffffff0000000b00000000",
            INIT_07 => X"000000210000000000000013000000000000000200000000fffffffaffffffff",
            INIT_08 => X"ffffffeaffffffffffffffb1ffffffff00000006000000000000001000000000",
            INIT_09 => X"00000009000000000000001000000000ffffffe4ffffffff0000000100000000",
            INIT_0A => X"ffffffeaffffffff0000002b00000000ffffffeeffffffff0000001900000000",
            INIT_0B => X"000000340000000000000000000000000000002300000000fffffff3ffffffff",
            INIT_0C => X"0000000e000000000000002b000000000000001d00000000fffffff3ffffffff",
            INIT_0D => X"fffffff1ffffffff00000008000000000000000900000000ffffffdaffffffff",
            INIT_0E => X"000000110000000000000008000000000000002900000000fffffff6ffffffff",
            INIT_0F => X"fffffff8ffffffff00000032000000000000001c00000000ffffffdeffffffff",
            INIT_10 => X"fffffffbffffffffffffffc9ffffffffffffffd3fffffffffffffffeffffffff",
            INIT_11 => X"0000000d00000000fffffff4ffffffffffffffc1ffffffff0000001c00000000",
            INIT_12 => X"00000011000000000000002f00000000fffffff5ffffffff0000001000000000",
            INIT_13 => X"0000000c00000000ffffffc9ffffffff0000001c00000000fffffffaffffffff",
            INIT_14 => X"00000025000000000000001200000000ffffffd8ffffffff0000000e00000000",
            INIT_15 => X"ffffffbdfffffffffffffff0ffffffff0000003300000000ffffffefffffffff",
            INIT_16 => X"ffffffd8ffffffff000000070000000000000033000000000000001100000000",
            INIT_17 => X"00000019000000000000000f00000000fffffff3ffffffffffffffbeffffffff",
            INIT_18 => X"ffffffe4ffffffffffffffbaffffffffffffffe5ffffffff0000001400000000",
            INIT_19 => X"0000000d000000000000001600000000ffffffd3fffffffffffffff3ffffffff",
            INIT_1A => X"0000001400000000fffffffafffffffffffffffeffffffffffffffe3ffffffff",
            INIT_1B => X"fffffff9fffffffffffffffbffffffff00000010000000000000000700000000",
            INIT_1C => X"0000000b00000000ffffffecffffffffffffffddfffffffffffffff0ffffffff",
            INIT_1D => X"ffffffbdffffffffffffffedffffffff00000005000000000000000200000000",
            INIT_1E => X"fffffff9fffffffffffffffaffffffffffffffb9ffffffffffffffebffffffff",
            INIT_1F => X"00000010000000000000001f00000000fffffffaffffffffffffffd1ffffffff",
            INIT_20 => X"ffffffe5ffffffffffffffe6ffffffff00000002000000000000000200000000",
            INIT_21 => X"fffffffdffffffff0000000d00000000ffffffddffffffffffffffbdffffffff",
            INIT_22 => X"00000000000000000000000500000000ffffffe2ffffffff0000001800000000",
            INIT_23 => X"ffffffeeffffffff0000000900000000fffffffcffffffff0000000c00000000",
            INIT_24 => X"0000003100000000ffffffe0ffffffffffffffe9ffffffff0000000a00000000",
            INIT_25 => X"ffffffcffffffffffffffff3ffffffff0000003300000000ffffffeeffffffff",
            INIT_26 => X"ffffffdfffffffffffffffddffffffff0000002800000000ffffffedffffffff",
            INIT_27 => X"00000023000000000000000c00000000fffffff4fffffffffffffff0ffffffff",
            INIT_28 => X"ffffffd9fffffffffffffffcffffffff00000016000000000000000800000000",
            INIT_29 => X"00000000000000000000000400000000fffffff8ffffffffffffffd9ffffffff",
            INIT_2A => X"ffffffdbffffffff0000001800000000fffffffcffffffffffffffffffffffff",
            INIT_2B => X"ffffffd9ffffffff000000280000000000000020000000000000001000000000",
            INIT_2C => X"0000003900000000ffffffc0fffffffffffffff9ffffffff0000000d00000000",
            INIT_2D => X"ffffffd7fffffffffffffff6ffffffff0000001200000000ffffffdeffffffff",
            INIT_2E => X"fffffff5ffffffffffffffabffffffffffffffeafffffffffffffff2ffffffff",
            INIT_2F => X"0000000a000000000000001d000000000000001300000000fffffff2ffffffff",
            INIT_30 => X"ffffffc3ffffffffffffffd6ffffffff00000012000000000000000f00000000",
            INIT_31 => X"0000001a000000000000000b00000000fffffff5ffffffffffffffd9ffffffff",
            INIT_32 => X"ffffffe4ffffffffffffffefffffffffffffffebffffffff0000002100000000",
            INIT_33 => X"ffffffe9ffffffff000000330000000000000023000000000000000a00000000",
            INIT_34 => X"0000001700000000ffffffbefffffffffffffffffffffffffffffff6ffffffff",
            INIT_35 => X"0000000700000000000000010000000000000050000000000000000700000000",
            INIT_36 => X"0000000e00000000ffffff8dffffffff0000001400000000ffffffdeffffffff",
            INIT_37 => X"fffffff3ffffffff0000000c00000000fffffffaffffffff0000001400000000",
            INIT_38 => X"ffffffc2ffffffffffffffbeffffffff00000000000000000000000900000000",
            INIT_39 => X"ffffffefffffffff00000007000000000000000200000000fffffff3ffffffff",
            INIT_3A => X"fffffffaffffffff0000001f00000000ffffffdbfffffffffffffff3ffffffff",
            INIT_3B => X"000000180000000000000016000000000000003200000000fffffff5ffffffff",
            INIT_3C => X"0000002d00000000fffffff9ffffffff00000011000000000000000d00000000",
            INIT_3D => X"fffffffdffffffff00000009000000000000000600000000ffffffe7ffffffff",
            INIT_3E => X"ffffffeaffffffffffffffc0ffffffffffffffb3ffffffff0000000100000000",
            INIT_3F => X"000000290000000000000018000000000000000400000000fffffffdffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffe8ffffffffffffffc0fffffffffffffffaffffffff0000001d00000000",
            INIT_41 => X"0000000b00000000ffffffeeffffffffffffffb1ffffffff0000000f00000000",
            INIT_42 => X"0000001f00000000ffffffdbffffffffffffffd3ffffffff0000002a00000000",
            INIT_43 => X"000000150000000000000018000000000000000500000000ffffffe7ffffffff",
            INIT_44 => X"ffffff88ffffffff0000000a0000000000000035000000000000001400000000",
            INIT_45 => X"0000000f000000000000000c0000000000000007000000000000000900000000",
            INIT_46 => X"fffffff2ffffffff0000004300000000ffffffafffffffff0000001300000000",
            INIT_47 => X"ffffffe4ffffffffffffffeeffffffff00000037000000000000000700000000",
            INIT_48 => X"0000001b00000000ffffff96ffffffffffffffc8ffffffffffffffe0ffffffff",
            INIT_49 => X"fffffffffffffffffffffff0ffffffff00000015000000000000001b00000000",
            INIT_4A => X"0000001f00000000ffffffcaffffffff0000001700000000ffffffe6ffffffff",
            INIT_4B => X"0000001300000000ffffffecffffffff0000001200000000ffffffd9ffffffff",
            INIT_4C => X"ffffffecffffffff0000001f0000000000000026000000000000002500000000",
            INIT_4D => X"0000001900000000fffffff6ffffffff00000002000000000000001700000000",
            INIT_4E => X"00000004000000000000000600000000ffffffacffffffff0000000800000000",
            INIT_4F => X"ffffffe4ffffffff00000009000000000000000700000000ffffffe7ffffffff",
            INIT_50 => X"0000001600000000ffffffe6fffffffffffffff2fffffffffffffff1ffffffff",
            INIT_51 => X"fffffff5ffffffff0000000c000000000000000f000000000000000000000000",
            INIT_52 => X"0000000000000000ffffffebffffffff0000001f00000000fffffff9ffffffff",
            INIT_53 => X"0000001700000000fffffff1ffffffff00000002000000000000000700000000",
            INIT_54 => X"ffffffe4ffffffff0000001700000000ffffffb3ffffffff0000001500000000",
            INIT_55 => X"fffffff7ffffffffffffffe4ffffffff0000001c000000000000001000000000",
            INIT_56 => X"0000000a00000000fffffff5ffffffffffffffbeffffffff0000000600000000",
            INIT_57 => X"ffffffbcfffffffffffffff3fffffffffffffffefffffffffffffff5ffffffff",
            INIT_58 => X"fffffff6ffffffffffffffcaffffffffffffffccfffffffffffffff1ffffffff",
            INIT_59 => X"fffffff6ffffffff0000000a000000000000001a00000000ffffffeaffffffff",
            INIT_5A => X"fffffffeffffffffffffffc9ffffffff0000000f00000000ffffffdeffffffff",
            INIT_5B => X"0000000b00000000fffffffbfffffffffffffffaffffffff0000000100000000",
            INIT_5C => X"00000026000000000000000d00000000ffffffbaffffffff0000000900000000",
            INIT_5D => X"fffffff4ffffffffffffffd0ffffffff0000001a000000000000000100000000",
            INIT_5E => X"fffffffaffffffffffffffedffffffffffffffe9ffffffffffffffebffffffff",
            INIT_5F => X"ffffffecfffffffffffffffbfffffffffffffff1ffffffffffffffe7ffffffff",
            INIT_60 => X"ffffffe3ffffffffffffffdaffffffffffffffe0ffffffff0000000100000000",
            INIT_61 => X"fffffff2ffffffff0000001000000000ffffffffffffffffffffffe2ffffffff",
            INIT_62 => X"0000002500000000ffffffdaffffffff00000012000000000000000e00000000",
            INIT_63 => X"0000001b0000000000000025000000000000000200000000ffffffeaffffffff",
            INIT_64 => X"0000000a000000000000001d00000000ffffffc7fffffffffffffff1ffffffff",
            INIT_65 => X"ffffffffffffffffffffffc9ffffffff00000004000000000000001500000000",
            INIT_66 => X"fffffffbffffffff0000002000000000fffffff4fffffffffffffff6ffffffff",
            INIT_67 => X"fffffff0ffffffffffffffe8fffffffffffffff0ffffffffffffffddffffffff",
            INIT_68 => X"ffffffd1ffffffffffffffc7ffffffffffffffd7fffffffffffffffbffffffff",
            INIT_69 => X"ffffffefffffffff00000011000000000000000400000000fffffff6ffffffff",
            INIT_6A => X"0000002900000000000000050000000000000001000000000000001900000000",
            INIT_6B => X"000000270000000000000005000000000000000b00000000ffffffedffffffff",
            INIT_6C => X"00000006000000000000001200000000fffffff4ffffffff0000000e00000000",
            INIT_6D => X"ffffffecffffffffffffffb8ffffffff00000018000000000000001200000000",
            INIT_6E => X"ffffffffffffffff0000004600000000ffffffa8fffffffffffffff7ffffffff",
            INIT_6F => X"ffffffe4fffffffffffffff8ffffffff0000000800000000ffffffe3ffffffff",
            INIT_70 => X"0000000000000000ffffffc9ffffffffffffffc7ffffffff0000000700000000",
            INIT_71 => X"00000017000000000000001c00000000fffffff3ffffffff0000000300000000",
            INIT_72 => X"0000002000000000fffffff8ffffffff00000008000000000000000d00000000",
            INIT_73 => X"0000002c00000000fffffffeffffffff0000000900000000ffffffe5ffffffff",
            INIT_74 => X"ffffffd0ffffffff0000001f000000000000001e000000000000000a00000000",
            INIT_75 => X"ffffffffffffffffffffffc6fffffffffffffff7ffffffff0000001200000000",
            INIT_76 => X"fffffffaffffffff0000002800000000ffffff98ffffffff0000001700000000",
            INIT_77 => X"ffffffdaffffffff00000001000000000000000000000000fffffff4ffffffff",
            INIT_78 => X"0000000000000000ffffffbeffffffffffffffd3fffffffffffffffbffffffff",
            INIT_79 => X"000000040000000000000006000000000000000b000000000000001e00000000",
            INIT_7A => X"fffffff4ffffffffffffffa9ffffffff00000019000000000000002000000000",
            INIT_7B => X"0000002a00000000ffffffd9ffffffff0000000500000000fffffff6ffffffff",
            INIT_7C => X"ffffffe3ffffffff0000000a0000000000000025000000000000000a00000000",
            INIT_7D => X"fffffffbfffffffffffffff8fffffffffffffff0ffffffff0000000400000000",
            INIT_7E => X"00000019000000000000001700000000ffffffd1ffffffff0000001500000000",
            INIT_7F => X"ffffffccffffffffffffffe2fffffffffffffffbffffffff0000000f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE24;


    MEM_IWGHT_LAYER2_INSTANCE25 : if BRAM_NAME = "iwght_layer2_instance25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001b00000000ffffffdbfffffffffffffffcffffffff0000000a00000000",
            INIT_01 => X"fffffff3ffffffff0000000200000000ffffffffffffffff0000001300000000",
            INIT_02 => X"0000001100000000fffffff1ffffffff0000000700000000fffffffaffffffff",
            INIT_03 => X"0000000c00000000ffffffebffffffff00000003000000000000001200000000",
            INIT_04 => X"fffffff6ffffffff00000001000000000000000200000000fffffffeffffffff",
            INIT_05 => X"fffffffcfffffffffffffffdffffffff00000010000000000000001000000000",
            INIT_06 => X"0000000e000000000000001700000000ffffffc6ffffffff0000000200000000",
            INIT_07 => X"ffffffeeffffffff0000001a0000000000000000000000000000000100000000",
            INIT_08 => X"fffffffaffffffffffffffd0fffffffffffffff6ffffffff0000000f00000000",
            INIT_09 => X"0000000d000000000000001300000000fffffffafffffffffffffff5ffffffff",
            INIT_0A => X"0000000c00000000ffffffe5ffffffff00000023000000000000002300000000",
            INIT_0B => X"fffffffdffffffffffffffe7ffffffffffffffe0ffffffff0000001800000000",
            INIT_0C => X"0000000800000000fffffffaffffffffffffffe7ffffffff0000000900000000",
            INIT_0D => X"ffffffe4fffffffffffffff7ffffffff00000005000000000000001200000000",
            INIT_0E => X"0000001c000000000000000900000000fffffff8ffffffffffffffebffffffff",
            INIT_0F => X"fffffffaffffffff000000180000000000000004000000000000000600000000",
            INIT_10 => X"ffffffd3fffffffffffffff3ffffffff00000001000000000000000000000000",
            INIT_11 => X"ffffffd6ffffffff0000000c000000000000000c00000000fffffff8ffffffff",
            INIT_12 => X"ffffffe6fffffffffffffff5ffffffff0000000600000000fffffff5ffffffff",
            INIT_13 => X"ffffffeaffffffff0000002e00000000fffffff2fffffffffffffffdffffffff",
            INIT_14 => X"0000000e00000000ffffffeeffffffffffffffe5fffffffffffffffaffffffff",
            INIT_15 => X"fffffff7ffffffff0000001d0000000000000005000000000000000d00000000",
            INIT_16 => X"00000005000000000000000e000000000000001a00000000ffffffebffffffff",
            INIT_17 => X"0000000600000000000000080000000000000030000000000000001000000000",
            INIT_18 => X"ffffffdbffffffffffffffdbfffffffffffffff2ffffffff0000000000000000",
            INIT_19 => X"ffffffd9ffffffff0000000d00000000fffffffdfffffffffffffff3ffffffff",
            INIT_1A => X"ffffffd8ffffffffffffffe0fffffffffffffff4ffffffffffffffe1ffffffff",
            INIT_1B => X"fffffff5ffffffffffffffe6ffffffffffffffecfffffffffffffff7ffffffff",
            INIT_1C => X"0000000a00000000fffffff0ffffffffffffffe6fffffffffffffff4ffffffff",
            INIT_1D => X"0000000800000000fffffffdffffffff00000018000000000000002300000000",
            INIT_1E => X"0000002000000000fffffffcffffffff0000000000000000ffffffdbffffffff",
            INIT_1F => X"fffffff2ffffffff00000017000000000000002200000000fffffffcffffffff",
            INIT_20 => X"ffffffeaffffffffffffffe2ffffffffffffffdcffffffff0000000c00000000",
            INIT_21 => X"ffffffe7ffffffff00000013000000000000000900000000fffffffbffffffff",
            INIT_22 => X"0000000f000000000000000d00000000fffffff8ffffffff0000000b00000000",
            INIT_23 => X"0000000b00000000fffffff5fffffffffffffff0ffffffff0000000e00000000",
            INIT_24 => X"0000000b000000000000000000000000ffffffe0ffffffff0000000800000000",
            INIT_25 => X"fffffffdffffffff0000001700000000fffffff4ffffffff0000000700000000",
            INIT_26 => X"ffffffeeffffffff000000120000000000000005000000000000000200000000",
            INIT_27 => X"000000260000000000000002000000000000000300000000ffffffdfffffffff",
            INIT_28 => X"ffffffc8ffffffffffffff97ffffffffffffffd6fffffffffffffffaffffffff",
            INIT_29 => X"ffffffdbffffffff0000000200000000fffffff7ffffffff0000001400000000",
            INIT_2A => X"0000003000000000ffffffc8ffffffff0000000b000000000000001400000000",
            INIT_2B => X"0000001400000000fffffff4fffffffffffffff8fffffffffffffffbffffffff",
            INIT_2C => X"ffffffcaffffffff000000030000000000000008000000000000000000000000",
            INIT_2D => X"0000001500000000fffffff9ffffffffffffffe5ffffffff0000002000000000",
            INIT_2E => X"0000001e000000000000004600000000ffffffffffffffff0000000600000000",
            INIT_2F => X"ffffffecffffffffffffffe8ffffffff0000001800000000ffffffeaffffffff",
            INIT_30 => X"ffffffe6ffffffffffffffb5ffffffffffffffd5ffffffff0000000c00000000",
            INIT_31 => X"ffffffeeffffffff000000150000000000000015000000000000000400000000",
            INIT_32 => X"ffffffe7ffffffffffffffcdffffffff00000010000000000000001d00000000",
            INIT_33 => X"0000000300000000ffffffdffffffffffffffffbffffffffffffffe8ffffffff",
            INIT_34 => X"ffffffdffffffffffffffffdffffffff0000004500000000fffffff1ffffffff",
            INIT_35 => X"0000002100000000fffffffdffffffffffffffffffffffff0000002c00000000",
            INIT_36 => X"00000000000000000000005200000000ffffffe1fffffffffffffff8ffffffff",
            INIT_37 => X"ffffffdfffffffffffffffe9ffffffff0000000f000000000000000600000000",
            INIT_38 => X"0000000200000000ffffffbdffffffffffffffd6fffffffffffffffcffffffff",
            INIT_39 => X"ffffffe1ffffffff0000000f000000000000000700000000fffffff6ffffffff",
            INIT_3A => X"ffffffebfffffffffffffff8ffffffff00000018000000000000000e00000000",
            INIT_3B => X"ffffffffffffffff0000000000000000fffffff6ffffffff0000000000000000",
            INIT_3C => X"ffffffe9ffffffffffffffe5ffffffffffffffebffffffffffffffebffffffff",
            INIT_3D => X"ffffffacffffffffffffffd7ffffffffffffffe2ffffffff0000001300000000",
            INIT_3E => X"00000005000000000000000b00000000ffffffe3ffffffff0000000000000000",
            INIT_3F => X"fffffffdffffffff0000001b000000000000000b00000000fffffff1ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffffffffffffffffff95ffffffffffffffd9ffffffff0000001100000000",
            INIT_41 => X"ffffffe7ffffffff0000000e00000000fffffffcffffffff0000001000000000",
            INIT_42 => X"ffffffe9fffffffffffffffefffffffffffffffdffffffff0000001300000000",
            INIT_43 => X"fffffff9fffffffffffffffaffffffff0000000600000000ffffffe3ffffffff",
            INIT_44 => X"ffffffeefffffffffffffff9ffffffffffffffc8fffffffffffffff6ffffffff",
            INIT_45 => X"ffffffe6ffffffff000000060000000000000017000000000000001600000000",
            INIT_46 => X"ffffffe6ffffffff0000001e00000000ffffffd1fffffffffffffff7ffffffff",
            INIT_47 => X"0000002500000000000000120000000000000007000000000000001200000000",
            INIT_48 => X"ffffffe2fffffffffffffff8fffffffffffffffeffffffff0000000d00000000",
            INIT_49 => X"ffffffd5ffffffff0000000700000000fffffffbffffffff0000000200000000",
            INIT_4A => X"fffffffcfffffffffffffffdffffffffffffffe6fffffffffffffffdffffffff",
            INIT_4B => X"fffffff3ffffffff0000000d00000000fffffff5ffffffffffffffc9ffffffff",
            INIT_4C => X"0000002300000000ffffffe3ffffffffffffffedffffffffffffffe5ffffffff",
            INIT_4D => X"ffffffc9ffffffffffffffebffffffff0000002e000000000000000e00000000",
            INIT_4E => X"ffffffe8ffffffff00000000000000000000005a00000000fffffff8ffffffff",
            INIT_4F => X"0000001e000000000000001c0000000000000025000000000000000900000000",
            INIT_50 => X"ffffffedffffffffffffffcafffffffffffffffdffffffffffffffefffffffff",
            INIT_51 => X"ffffffd1fffffffffffffffaffffffff00000003000000000000000500000000",
            INIT_52 => X"0000000800000000fffffffeffffffffffffffedffffffff0000000e00000000",
            INIT_53 => X"ffffffdbffffffff00000015000000000000000000000000ffffffedffffffff",
            INIT_54 => X"0000003b00000000fffffff1fffffffffffffff0ffffffffffffffe8ffffffff",
            INIT_55 => X"ffffffc2ffffffff000000160000000000000018000000000000001b00000000",
            INIT_56 => X"0000001100000000000000020000000000000004000000000000000900000000",
            INIT_57 => X"000000170000000000000008000000000000002400000000ffffffffffffffff",
            INIT_58 => X"ffffffc6ffffffffffffffeaffffffff00000018000000000000000a00000000",
            INIT_59 => X"ffffffdeffffffff0000001700000000fffffffbffffffff0000001100000000",
            INIT_5A => X"fffffff3ffffffffffffffe8fffffffffffffffbffffffff0000000d00000000",
            INIT_5B => X"fffffffbffffffffffffffe3ffffffff00000000000000000000000d00000000",
            INIT_5C => X"0000000b00000000fffffff0ffffffff00000024000000000000000400000000",
            INIT_5D => X"ffffffbeffffffff0000000400000000fffffffbffffffff0000000b00000000",
            INIT_5E => X"0000003300000000ffffffedfffffffffffffff0ffffffff0000000000000000",
            INIT_5F => X"0000001300000000000000180000000000000008000000000000000000000000",
            INIT_60 => X"ffffffe8ffffffffffffffceffffffffffffffe9ffffffff0000001000000000",
            INIT_61 => X"ffffffddffffffff000000140000000000000006000000000000000100000000",
            INIT_62 => X"0000002b00000000ffffffc3fffffffffffffff0ffffffff0000000900000000",
            INIT_63 => X"0000000700000000ffffffc6ffffffff0000000d000000000000000800000000",
            INIT_64 => X"ffffffceffffffff000000250000000000000018000000000000001000000000",
            INIT_65 => X"ffffffacfffffffffffffff4ffffffff00000011000000000000002500000000",
            INIT_66 => X"0000001e000000000000003100000000fffffff3ffffffff0000001100000000",
            INIT_67 => X"fffffffaffffffff0000001d000000000000001900000000ffffffeaffffffff",
            INIT_68 => X"fffffff0ffffffffffffffb3ffffffffffffffcfffffffff0000002200000000",
            INIT_69 => X"ffffffeeffffffff00000021000000000000000e000000000000001400000000",
            INIT_6A => X"ffffffeeffffffffffffffe8ffffffff00000007000000000000000600000000",
            INIT_6B => X"0000000c00000000fffffffcffffffffffffffecffffffffffffffe3ffffffff",
            INIT_6C => X"ffffffedffffffff00000010000000000000000f000000000000001800000000",
            INIT_6D => X"fffffffdfffffffffffffffeffffffff0000001600000000fffffffdffffffff",
            INIT_6E => X"fffffffaffffffff0000003d00000000ffffffb1ffffffff0000002400000000",
            INIT_6F => X"fffffff1fffffffffffffffcffffffff0000001b00000000fffffffbffffffff",
            INIT_70 => X"fffffffbfffffffffffffffffffffffffffffff5fffffffffffffff3ffffffff",
            INIT_71 => X"ffffffc8fffffffffffffff8fffffffffffffffdffffffff0000000500000000",
            INIT_72 => X"fffffff3ffffffffffffffeaffffffff0000001100000000fffffff8ffffffff",
            INIT_73 => X"00000019000000000000000d000000000000000400000000fffffffdffffffff",
            INIT_74 => X"fffffff7fffffffffffffffeffffffff00000016000000000000000000000000",
            INIT_75 => X"0000002400000000000000020000000000000012000000000000000800000000",
            INIT_76 => X"ffffffedffffffff0000001e000000000000000b000000000000001300000000",
            INIT_77 => X"ffffffffffffffff0000001b00000000fffffffafffffffffffffff8ffffffff",
            INIT_78 => X"ffffffeaffffffffffffffe1ffffffffffffffefffffffff0000000700000000",
            INIT_79 => X"fffffff8ffffffff0000001200000000ffffffe6ffffffff0000000800000000",
            INIT_7A => X"ffffffe0ffffffffffffffd9fffffffffffffff5fffffffffffffffdffffffff",
            INIT_7B => X"fffffffafffffffffffffffbfffffffffffffff7ffffffffffffffefffffffff",
            INIT_7C => X"0000000300000000ffffffeffffffffffffffff3fffffffffffffff4ffffffff",
            INIT_7D => X"ffffffe8fffffffffffffffafffffffffffffffdffffffff0000000700000000",
            INIT_7E => X"ffffffe7ffffffff0000000a0000000000000018000000000000000d00000000",
            INIT_7F => X"0000000b00000000000000040000000000000000000000000000001d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE25;


    MEM_IWGHT_LAYER2_INSTANCE26 : if BRAM_NAME = "iwght_layer2_instance26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000ffffffd1ffffffffffffffebffffffff0000000000000000",
            INIT_01 => X"ffffffe4ffffffff0000000300000000fffffff7ffffffff0000001900000000",
            INIT_02 => X"fffffffbfffffffffffffff1fffffffffffffff0ffffffff0000001300000000",
            INIT_03 => X"ffffffe7ffffffff0000000500000000ffffffebffffffffffffffe1ffffffff",
            INIT_04 => X"0000001200000000ffffffe0ffffffffffffffebffffffffffffffcdffffffff",
            INIT_05 => X"ffffffc5ffffffff00000009000000000000000000000000fffffff0ffffffff",
            INIT_06 => X"ffffffe3ffffffffffffffdcfffffffffffffffeffffffff0000002800000000",
            INIT_07 => X"0000000000000000000000030000000000000026000000000000001a00000000",
            INIT_08 => X"ffffffe7ffffffffffffffc9fffffffffffffff2fffffffffffffff6ffffffff",
            INIT_09 => X"ffffffdcfffffffffffffffcffffffff00000002000000000000001a00000000",
            INIT_0A => X"fffffff7ffffffffffffffe8fffffffffffffffbffffffff0000001a00000000",
            INIT_0B => X"ffffffddfffffffffffffffeffffffff0000000200000000ffffffd8ffffffff",
            INIT_0C => X"0000000f00000000ffffffc5fffffffffffffffcffffffff0000000200000000",
            INIT_0D => X"ffffffadffffffff000000220000000000000005000000000000000600000000",
            INIT_0E => X"0000000d00000000ffffffdbffffffff00000020000000000000000200000000",
            INIT_0F => X"0000000d0000000000000013000000000000003e000000000000000700000000",
            INIT_10 => X"fffffffaffffffffffffffd5fffffffffffffff9ffffffffffffffffffffffff",
            INIT_11 => X"ffffffe4fffffffffffffffafffffffffffffff2ffffffff0000000700000000",
            INIT_12 => X"fffffff8fffffffffffffff0ffffffffffffffe6ffffffff0000001f00000000",
            INIT_13 => X"fffffffaffffffffffffffd5ffffffff0000000400000000fffffff8ffffffff",
            INIT_14 => X"0000000e00000000ffffffe0ffffffff00000005000000000000000600000000",
            INIT_15 => X"ffffffbfffffffff0000002c00000000ffffffedffffffff0000000b00000000",
            INIT_16 => X"0000000400000000ffffffe6ffffffffffffffc0fffffffffffffffeffffffff",
            INIT_17 => X"0000000a000000000000001d000000000000004100000000ffffffe7ffffffff",
            INIT_18 => X"fffffff2ffffffffffffffd7ffffffffffffffe0ffffffff0000001a00000000",
            INIT_19 => X"ffffffe4ffffffffffffffedffffffffffffffeeffffffff0000000d00000000",
            INIT_1A => X"0000001800000000ffffffddffffffffffffffd7ffffffff0000002500000000",
            INIT_1B => X"0000000900000000ffffffb9ffffffffffffffdbfffffffffffffff4ffffffff",
            INIT_1C => X"0000000f0000000000000006000000000000002c000000000000000800000000",
            INIT_1D => X"ffffffc6ffffffff000000200000000000000013000000000000002000000000",
            INIT_1E => X"0000000d000000000000000f0000000000000010000000000000000600000000",
            INIT_1F => X"0000000600000000ffffffdfffffffff0000005400000000fffffff6ffffffff",
            INIT_20 => X"ffffffe8ffffffff0000000700000000ffffffedffffffff0000001500000000",
            INIT_21 => X"ffffffe4ffffffff0000000f0000000000000008000000000000000800000000",
            INIT_22 => X"0000000d00000000fffffffffffffffffffffff0fffffffffffffffaffffffff",
            INIT_23 => X"ffffffeeffffffff0000002100000000ffffffecffffffffffffffc9ffffffff",
            INIT_24 => X"ffffffcdffffffffffffffd9ffffffff0000000d00000000fffffffaffffffff",
            INIT_25 => X"00000000000000000000001b00000000fffffff6fffffffffffffff2ffffffff",
            INIT_26 => X"ffffffddffffffff0000005c00000000ffffffd4ffffffff0000002700000000",
            INIT_27 => X"0000000b00000000ffffffcdffffffff00000019000000000000002200000000",
            INIT_28 => X"00000024000000000000002e000000000000001500000000fffffff8ffffffff",
            INIT_29 => X"ffffffc8ffffffff00000005000000000000000e000000000000000000000000",
            INIT_2A => X"ffffffd7ffffffffffffffd8fffffffffffffff1ffffffffffffffefffffffff",
            INIT_2B => X"00000011000000000000000b000000000000002a00000000ffffffe9ffffffff",
            INIT_2C => X"ffffffeafffffffffffffff0fffffffffffffffdffffffffffffffeaffffffff",
            INIT_2D => X"0000002000000000fffffffcffffffff0000001c00000000ffffffd6ffffffff",
            INIT_2E => X"00000024000000000000001700000000ffffff9dffffffff0000001500000000",
            INIT_2F => X"fffffff5fffffffffffffff2ffffffff0000003b000000000000002000000000",
            INIT_30 => X"fffffff8ffffffff0000001b00000000fffffffbffffffff0000001500000000",
            INIT_31 => X"fffffffdffffffff0000000000000000ffffffe3ffffffff0000001f00000000",
            INIT_32 => X"ffffffeeffffffffffffffc0fffffffffffffff0ffffffff0000001200000000",
            INIT_33 => X"fffffff7ffffffffffffffebffffffff0000001000000000ffffffe8ffffffff",
            INIT_34 => X"ffffffd1ffffffffffffffe8ffffffffffffffd0ffffffff0000001200000000",
            INIT_35 => X"00000003000000000000001a000000000000000b00000000fffffff7ffffffff",
            INIT_36 => X"ffffffd8ffffffff0000000400000000ffffffe0ffffffff0000001b00000000",
            INIT_37 => X"00000000000000000000000b0000000000000044000000000000002700000000",
            INIT_38 => X"fffffff8ffffffff0000001000000000ffffffddffffffff0000000d00000000",
            INIT_39 => X"fffffffcfffffffffffffff5ffffffff00000009000000000000001900000000",
            INIT_3A => X"ffffffe8ffffffffffffffe4ffffffffffffffe7ffffffff0000002d00000000",
            INIT_3B => X"0000000800000000ffffffd5ffffffff0000001d00000000fffffff5ffffffff",
            INIT_3C => X"ffffffa0fffffffffffffff7ffffffffffffffdfffffffff0000002500000000",
            INIT_3D => X"ffffffddffffffff00000026000000000000000400000000fffffff9ffffffff",
            INIT_3E => X"fffffff6ffffffffffffffd9ffffffff0000001c000000000000001e00000000",
            INIT_3F => X"0000002000000000fffffff0ffffffff0000001f000000000000002300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000900000000ffffffaeffffffffffffffe0ffffffffffffffedffffffff",
            INIT_41 => X"fffffff2ffffffff000000170000000000000020000000000000001d00000000",
            INIT_42 => X"fffffff5ffffffffffffffdeffffffffffffffecffffffff0000002900000000",
            INIT_43 => X"ffffffe7ffffffffffffffc0ffffffff0000000e00000000ffffffeaffffffff",
            INIT_44 => X"ffffffd2ffffffff0000000400000000fffffff5ffffffff0000002300000000",
            INIT_45 => X"ffffffb8ffffffff00000018000000000000000200000000fffffffdffffffff",
            INIT_46 => X"0000001600000000fffffff4ffffffff0000004e000000000000001e00000000",
            INIT_47 => X"0000002200000000fffffffdffffffff0000003d000000000000000900000000",
            INIT_48 => X"ffffffd6ffffffffffffffcdffffffffffffffcbffffffff0000001100000000",
            INIT_49 => X"fffffffaffffffff0000000d000000000000000c000000000000002100000000",
            INIT_4A => X"fffffffeffffffffffffffedffffffffffffffecffffffff0000002900000000",
            INIT_4B => X"fffffff5ffffffffffffffe2ffffffff0000000600000000fffffff8ffffffff",
            INIT_4C => X"ffffffe0ffffffffffffffe9ffffffff00000029000000000000000500000000",
            INIT_4D => X"fffffff9ffffffff0000003400000000fffffff8ffffffffffffffe6ffffffff",
            INIT_4E => X"fffffffffffffffffffffffdffffffff00000043000000000000000600000000",
            INIT_4F => X"000000190000000000000024000000000000003d000000000000000600000000",
            INIT_50 => X"fffffffcffffffff000000170000000000000003000000000000001d00000000",
            INIT_51 => X"0000000900000000ffffffe8fffffffffffffff3ffffffff0000002400000000",
            INIT_52 => X"0000000c000000000000000500000000ffffffe8ffffffff0000001400000000",
            INIT_53 => X"0000001000000000ffffffdeffffffffffffffeeffffffffffffffc4ffffffff",
            INIT_54 => X"fffffff6ffffffff000000060000000000000059000000000000000700000000",
            INIT_55 => X"0000000900000000000000410000000000000011000000000000000500000000",
            INIT_56 => X"ffffffeaffffffff00000009000000000000006300000000fffffff5ffffffff",
            INIT_57 => X"ffffffecffffffffffffffdfffffffff0000002700000000fffffff6ffffffff",
            INIT_58 => X"ffffffe7ffffffff00000015000000000000002000000000fffffffdffffffff",
            INIT_59 => X"ffffffd6ffffffff000000170000000000000000000000000000001e00000000",
            INIT_5A => X"fffffff7fffffffffffffff5ffffffffffffffe2fffffffffffffff4ffffffff",
            INIT_5B => X"ffffffdeffffffff0000001d00000000ffffffcfffffffffffffffc4ffffffff",
            INIT_5C => X"ffffffdeffffffffffffffdeffffffffffffffdffffffffffffffff8ffffffff",
            INIT_5D => X"0000000f000000000000001400000000ffffffdffffffffffffffff7ffffffff",
            INIT_5E => X"00000007000000000000001e000000000000000e000000000000000300000000",
            INIT_5F => X"0000001a00000000ffffff92ffffffff00000005000000000000002100000000",
            INIT_60 => X"000000170000000000000038000000000000002e00000000ffffffdaffffffff",
            INIT_61 => X"ffffffc5ffffffffffffffe5ffffffff00000024000000000000000200000000",
            INIT_62 => X"fffffff4ffffffffffffffc6fffffffffffffff9fffffffffffffff2ffffffff",
            INIT_63 => X"fffffff4ffffffff00000021000000000000001200000000fffffffaffffffff",
            INIT_64 => X"ffffffb8ffffffff00000013000000000000000400000000ffffffe7ffffffff",
            INIT_65 => X"00000030000000000000003c000000000000001c00000000ffffffd2ffffffff",
            INIT_66 => X"0000002400000000fffffff8fffffffffffffffdffffffff0000000600000000",
            INIT_67 => X"ffffffecffffffffffffffe8ffffffffffffffffffffffff0000000800000000",
            INIT_68 => X"0000001900000000000000570000000000000002000000000000000600000000",
            INIT_69 => X"ffffffebffffffffffffffebffffffff00000000000000000000001000000000",
            INIT_6A => X"ffffffe4ffffffffffffffd0ffffffffffffffdbffffffff0000002000000000",
            INIT_6B => X"0000001100000000ffffffeaffffffff0000001b00000000fffffffcffffffff",
            INIT_6C => X"ffffff7dffffffff0000001c000000000000000800000000fffffff6ffffffff",
            INIT_6D => X"00000036000000000000001500000000fffffffcffffffffffffffe2ffffffff",
            INIT_6E => X"0000004800000000000000260000000000000029000000000000001500000000",
            INIT_6F => X"fffffffdffffffffffffffe3ffffffff0000001c000000000000000f00000000",
            INIT_70 => X"00000018000000000000003400000000ffffffbafffffffffffffffaffffffff",
            INIT_71 => X"fffffff8ffffffffffffffd4fffffffffffffff9ffffffff0000003500000000",
            INIT_72 => X"ffffffd0ffffffffffffffcaffffffffffffffe7ffffffff0000004500000000",
            INIT_73 => X"0000000800000000ffffffb3ffffffff0000003a000000000000002000000000",
            INIT_74 => X"ffffff4cffffffff0000002100000000fffffff6ffffffff0000001900000000",
            INIT_75 => X"00000031000000000000002700000000ffffffefffffffffffffffdeffffffff",
            INIT_76 => X"0000002500000000000000180000000000000011000000000000003100000000",
            INIT_77 => X"fffffff3ffffffffffffffdfffffffff00000027000000000000002800000000",
            INIT_78 => X"fffffff4ffffffffffffffedffffffffffffff8dffffffffffffffe9ffffffff",
            INIT_79 => X"fffffffaffffffffffffffd8ffffffff00000015000000000000002000000000",
            INIT_7A => X"ffffffdeffffffffffffffebfffffffffffffff6ffffffff0000003900000000",
            INIT_7B => X"fffffff5ffffffffffffffd6ffffffff0000003400000000fffffff1ffffffff",
            INIT_7C => X"ffffff7bffffffff0000001e00000000ffffffd8ffffffff0000000f00000000",
            INIT_7D => X"ffffffe3ffffffff0000002e00000000ffffffd8ffffffffffffffd8ffffffff",
            INIT_7E => X"0000000400000000000000220000000000000049000000000000003a00000000",
            INIT_7F => X"0000001100000000ffffffe8ffffffff0000001c000000000000000900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE26;


    MEM_IWGHT_LAYER2_INSTANCE27 : if BRAM_NAME = "iwght_layer2_instance27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffefffffffff0000001c00000000ffffffceffffffff0000000000000000",
            INIT_01 => X"ffffffffffffffff00000000000000000000001c000000000000002b00000000",
            INIT_02 => X"0000000300000000ffffffdeffffffffffffffd9fffffffffffffffdffffffff",
            INIT_03 => X"0000001e00000000ffffffa9ffffffff0000004700000000ffffffe5ffffffff",
            INIT_04 => X"ffffffc2ffffffff0000001b0000000000000010000000000000000800000000",
            INIT_05 => X"00000008000000000000003000000000ffffffe5ffffffffffffffddffffffff",
            INIT_06 => X"00000001000000000000000a00000000ffffffffffffffff0000000200000000",
            INIT_07 => X"0000001200000000ffffffecffffffff00000034000000000000000200000000",
            INIT_08 => X"00000012000000000000003f00000000ffffffeaffffffffffffffffffffffff",
            INIT_09 => X"fffffff8ffffffffffffffefffffffff00000000000000000000003300000000",
            INIT_0A => X"0000000900000000ffffffe8fffffffffffffff3ffffffff0000001e00000000",
            INIT_0B => X"fffffff7ffffffffffffffc7ffffffffffffffd3ffffffffffffffb9ffffffff",
            INIT_0C => X"000000080000000000000033000000000000002600000000ffffffe5ffffffff",
            INIT_0D => X"00000004000000000000001500000000ffffffefffffffffffffffdeffffffff",
            INIT_0E => X"ffffffeaffffffff0000000d000000000000002800000000fffffffcffffffff",
            INIT_0F => X"fffffff9ffffffffffffffe0ffffffff0000001d000000000000000e00000000",
            INIT_10 => X"ffffffe8ffffffff0000005b000000000000002b00000000ffffffe4ffffffff",
            INIT_11 => X"ffffffeaffffffff0000000a000000000000001b000000000000001a00000000",
            INIT_12 => X"ffffffe2ffffffff00000009000000000000000000000000ffffffeaffffffff",
            INIT_13 => X"ffffffdbffffffff0000002400000000ffffff9effffffffffffffb9ffffffff",
            INIT_14 => X"0000001600000000ffffffeaffffffffffffffc7fffffffffffffff1ffffffff",
            INIT_15 => X"ffffffddffffffffffffffd0ffffffff0000002500000000ffffffd7ffffffff",
            INIT_16 => X"00000028000000000000003d00000000ffffffd9ffffffff0000000600000000",
            INIT_17 => X"fffffff0ffffffffffffffafffffffffffffffd7ffffffff0000003400000000",
            INIT_18 => X"000000250000000000000045000000000000003900000000ffffffd3ffffffff",
            INIT_19 => X"ffffffc5fffffffffffffffeffffffff0000005f00000000fffffff3ffffffff",
            INIT_1A => X"fffffff2fffffffffffffffaffffffff0000001d00000000ffffff88ffffffff",
            INIT_1B => X"ffffffeaffffffffffffffffffffffff0000000000000000ffffffeeffffffff",
            INIT_1C => X"ffffffc9fffffffffffffff1ffffffff0000000100000000ffffffe7ffffffff",
            INIT_1D => X"0000003c00000000fffffff0ffffffff0000002800000000ffffffd1ffffffff",
            INIT_1E => X"00000036000000000000001b00000000ffffffd2ffffffff0000000400000000",
            INIT_1F => X"ffffffe6ffffffffffffffe1ffffffffffffffe4ffffffff0000000d00000000",
            INIT_20 => X"000000140000000000000036000000000000001900000000fffffff3ffffffff",
            INIT_21 => X"0000001800000000ffffffddffffffff0000000c000000000000002d00000000",
            INIT_22 => X"ffffffecffffffffffffffccffffffff00000015000000000000000300000000",
            INIT_23 => X"ffffffe6ffffffffffffffdcffffffff0000000d000000000000000800000000",
            INIT_24 => X"ffffff85ffffffff000000080000000000000009000000000000000000000000",
            INIT_25 => X"0000002b0000000000000003000000000000002e00000000ffffffc6ffffffff",
            INIT_26 => X"0000003e000000000000001100000000fffffff3fffffffffffffff8ffffffff",
            INIT_27 => X"ffffffccfffffffffffffffafffffffffffffff2ffffffff0000002f00000000",
            INIT_28 => X"0000002b000000000000004f00000000fffffff1fffffffffffffff5ffffffff",
            INIT_29 => X"0000001600000000ffffffe1ffffffff0000001a000000000000004300000000",
            INIT_2A => X"fffffff3ffffffffffffffcbffffffff00000000000000000000000400000000",
            INIT_2B => X"ffffffecffffffffffffffccffffffff00000015000000000000002600000000",
            INIT_2C => X"ffffff62ffffffff00000029000000000000001600000000fffffff9ffffffff",
            INIT_2D => X"fffffffcffffffff0000001400000000ffffffd8ffffffffffffffcfffffffff",
            INIT_2E => X"0000002a000000000000004700000000ffffffeaffffffff0000001100000000",
            INIT_2F => X"fffffff2ffffffffffffffcbffffffff00000002000000000000001100000000",
            INIT_30 => X"0000002d000000000000004200000000ffffffdcfffffffffffffff0ffffffff",
            INIT_31 => X"0000000c00000000ffffffefffffffff0000000c000000000000003200000000",
            INIT_32 => X"ffffffd3ffffffffffffffdbfffffffffffffff5ffffffff0000002400000000",
            INIT_33 => X"0000000900000000ffffffdeffffffff00000005000000000000001500000000",
            INIT_34 => X"ffffff58ffffffff0000002e000000000000001400000000fffffffdffffffff",
            INIT_35 => X"000000050000000000000011000000000000000400000000ffffffc8ffffffff",
            INIT_36 => X"00000010000000000000001d00000000fffffff2ffffffff0000001c00000000",
            INIT_37 => X"ffffffd7ffffffffffffffedfffffffffffffffbffffffff0000001100000000",
            INIT_38 => X"fffffffaffffffff0000004900000000ffffffe6fffffffffffffffdffffffff",
            INIT_39 => X"0000000400000000000000060000000000000015000000000000002600000000",
            INIT_3A => X"0000000000000000fffffff9ffffffff00000007000000000000002800000000",
            INIT_3B => X"0000000100000000ffffffd2fffffffffffffff3fffffffffffffff4ffffffff",
            INIT_3C => X"ffffffbcffffffff00000031000000000000001f00000000ffffffeaffffffff",
            INIT_3D => X"ffffffe2ffffffff0000000000000000fffffff8ffffffffffffffcfffffffff",
            INIT_3E => X"0000003d000000000000003a00000000fffffff5ffffffff0000002100000000",
            INIT_3F => X"ffffffe3ffffffffffffffecffffffffffffffebfffffffffffffffcffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000000000000000000006200000000ffffffefffffffff0000000600000000",
            INIT_41 => X"ffffffeaffffffff000000090000000000000015000000000000003800000000",
            INIT_42 => X"0000002700000000fffffff2ffffffff0000000a000000000000002100000000",
            INIT_43 => X"ffffffebffffffffffffffa6ffffffffffffff8dffffffffffffff92ffffffff",
            INIT_44 => X"ffffffe7ffffffff000000000000000000000029000000000000000200000000",
            INIT_45 => X"fffffff1ffffffffffffffd6ffffffff0000001c00000000fffffff5ffffffff",
            INIT_46 => X"ffffffebffffffff0000002a00000000ffffffeaffffffff0000000600000000",
            INIT_47 => X"ffffffa2ffffffffffffffc0ffffffffffffffd6ffffffff0000001e00000000",
            INIT_48 => X"ffffffe9ffffffff0000005a000000000000001d00000000ffffffc8ffffffff",
            INIT_49 => X"ffffffbaffffffff00000008000000000000005200000000ffffffffffffffff",
            INIT_4A => X"ffffffe9ffffffff00000001000000000000001e00000000ffffffb1ffffffff",
            INIT_4B => X"000000070000000000000003000000000000002b000000000000000300000000",
            INIT_4C => X"ffffffe8ffffffff0000002100000000ffffffbcffffffff0000003400000000",
            INIT_4D => X"ffffffcfffffffffffffffeaffffffff00000007000000000000001900000000",
            INIT_4E => X"0000000400000000ffffffe8ffffffff00000017000000000000003400000000",
            INIT_4F => X"fffffff2ffffffffffffffceffffffff0000000000000000fffffff9ffffffff",
            INIT_50 => X"0000002a000000000000002e00000000fffffffdfffffffffffffff1ffffffff",
            INIT_51 => X"ffffffd9ffffffff0000000d000000000000000d00000000fffffff3ffffffff",
            INIT_52 => X"0000000500000000ffffffeaffffffff0000001200000000ffffffbaffffffff",
            INIT_53 => X"0000000900000000ffffffddffffffff00000023000000000000001400000000",
            INIT_54 => X"fffffffaffffffff0000000b00000000ffffffbdffffffff0000001200000000",
            INIT_55 => X"ffffffd8ffffffff000000100000000000000019000000000000001d00000000",
            INIT_56 => X"00000012000000000000000a00000000ffffffdcffffffff0000001200000000",
            INIT_57 => X"fffffffaffffffffffffffe9ffffffffffffffc5ffffffffffffffe2ffffffff",
            INIT_58 => X"ffffffe6ffffffff00000050000000000000002000000000fffffffcffffffff",
            INIT_59 => X"ffffffffffffffff00000000000000000000000600000000fffffffeffffffff",
            INIT_5A => X"ffffffefffffffffffffffecffffffff0000000400000000ffffffd9ffffffff",
            INIT_5B => X"0000000100000000fffffffcfffffffffffffff8ffffffff0000000300000000",
            INIT_5C => X"ffffffe2fffffffffffffffdffffffff00000009000000000000002300000000",
            INIT_5D => X"ffffffc9ffffffff00000040000000000000001000000000ffffffecffffffff",
            INIT_5E => X"ffffffecfffffffffffffff7ffffffffffffffdbffffffff0000000100000000",
            INIT_5F => X"0000000300000000fffffff0fffffffffffffff4ffffffff0000000200000000",
            INIT_60 => X"000000260000000000000015000000000000000400000000ffffffecffffffff",
            INIT_61 => X"ffffffe9ffffffffffffffebfffffffffffffff9ffffffff0000001700000000",
            INIT_62 => X"ffffffefffffffffffffffe2fffffffffffffffeffffffffffffffdaffffffff",
            INIT_63 => X"0000000b00000000000000070000000000000025000000000000000400000000",
            INIT_64 => X"ffffffdbffffffff0000000a0000000000000003000000000000000b00000000",
            INIT_65 => X"00000006000000000000004400000000fffffff7ffffffffffffffefffffffff",
            INIT_66 => X"ffffffd0ffffffff0000002100000000fffffffaffffffff0000000300000000",
            INIT_67 => X"0000002b00000000fffffff6ffffffff00000001000000000000000400000000",
            INIT_68 => X"ffffffffffffffff0000001100000000fffffff8ffffffff0000000400000000",
            INIT_69 => X"0000000b00000000ffffffd5fffffffffffffffdffffffff0000002d00000000",
            INIT_6A => X"fffffff4ffffffffffffffd1ffffffff00000004000000000000000d00000000",
            INIT_6B => X"fffffffbffffffff000000160000000000000029000000000000001f00000000",
            INIT_6C => X"00000009000000000000000200000000ffffffd4ffffffff0000002500000000",
            INIT_6D => X"ffffffdfffffffff00000026000000000000000600000000ffffffedffffffff",
            INIT_6E => X"0000001200000000ffffffe4ffffffffffffffd1ffffffff0000001000000000",
            INIT_6F => X"fffffff3fffffffffffffff8ffffffff00000008000000000000000a00000000",
            INIT_70 => X"000000350000000000000027000000000000000b00000000fffffff6ffffffff",
            INIT_71 => X"0000000900000000ffffffdfffffffffffffffeeffffffff0000001b00000000",
            INIT_72 => X"fffffff1ffffffffffffffbdfffffffffffffff7ffffffffffffffeeffffffff",
            INIT_73 => X"0000000300000000000000130000000000000013000000000000001400000000",
            INIT_74 => X"fffffffbffffffff00000000000000000000001a000000000000001500000000",
            INIT_75 => X"fffffff1ffffffff00000030000000000000000d00000000fffffffcffffffff",
            INIT_76 => X"fffffffeffffffffffffffdcffffffffffffffc0ffffffff0000002000000000",
            INIT_77 => X"ffffffcdfffffffffffffffaffffffffffffffe2ffffffff0000000300000000",
            INIT_78 => X"0000000600000000000000460000000000000036000000000000000900000000",
            INIT_79 => X"fffffff7fffffffffffffff6ffffffff0000000b00000000fffffff3ffffffff",
            INIT_7A => X"ffffffe2ffffffffffffffc7ffffffff0000001900000000ffffffd0ffffffff",
            INIT_7B => X"0000000500000000000000110000000000000008000000000000000e00000000",
            INIT_7C => X"00000010000000000000002600000000fffffff3ffffffff0000002c00000000",
            INIT_7D => X"fffffffaffffffff000000000000000000000047000000000000000c00000000",
            INIT_7E => X"ffffffddffffffffffffffe8ffffffffffffff8bffffffff0000001600000000",
            INIT_7F => X"ffffffe5ffffffffffffffe6fffffffffffffff3ffffffff0000000300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE27;


    MEM_IWGHT_LAYER2_INSTANCE28 : if BRAM_NAME = "iwght_layer2_instance28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffffffffffff00000018000000000000002500000000ffffffeaffffffff",
            INIT_01 => X"fffffffeffffffff00000012000000000000000b00000000fffffff4ffffffff",
            INIT_02 => X"fffffffaffffffffffffffd4ffffffff0000001b00000000ffffffcfffffffff",
            INIT_03 => X"fffffffbffffffff0000000100000000fffffffbffffffff0000001a00000000",
            INIT_04 => X"0000000400000000fffffffeffffffff0000003500000000fffffff9ffffffff",
            INIT_05 => X"0000000000000000000000070000000000000001000000000000002200000000",
            INIT_06 => X"ffffffe8ffffffffffffffd6ffffffff0000004800000000fffffff1ffffffff",
            INIT_07 => X"fffffffafffffffffffffffbffffffffffffffecfffffffffffffffbffffffff",
            INIT_08 => X"0000001e0000000000000001000000000000000a000000000000000300000000",
            INIT_09 => X"0000000600000000fffffff8fffffffffffffffbffffffff0000000c00000000",
            INIT_0A => X"0000000700000000ffffffebfffffffffffffffefffffffffffffffaffffffff",
            INIT_0B => X"0000000100000000fffffffffffffffffffffff6ffffffff0000002b00000000",
            INIT_0C => X"000000120000000000000000000000000000000c000000000000001700000000",
            INIT_0D => X"ffffffd6ffffffff00000005000000000000000500000000ffffffffffffffff",
            INIT_0E => X"0000001f00000000fffffff1ffffffff0000000b000000000000000400000000",
            INIT_0F => X"fffffff7ffffffffffffffe4ffffffff0000000700000000fffffffbffffffff",
            INIT_10 => X"ffffffe7fffffffffffffffeffffffff0000001e00000000ffffffebffffffff",
            INIT_11 => X"fffffffcffffffff000000020000000000000002000000000000000600000000",
            INIT_12 => X"0000000e0000000000000000000000000000000a00000000fffffff7ffffffff",
            INIT_13 => X"0000000000000000ffffffd6ffffffff00000002000000000000000100000000",
            INIT_14 => X"0000001e00000000000000000000000000000008000000000000001100000000",
            INIT_15 => X"ffffffeffffffffffffffff9ffffffff0000000700000000fffffff8ffffffff",
            INIT_16 => X"ffffffe5ffffffff000000100000000000000006000000000000000900000000",
            INIT_17 => X"0000001200000000ffffffe4ffffffff00000004000000000000000e00000000",
            INIT_18 => X"ffffffe8ffffffffffffffeeffffffff0000000a00000000fffffffdffffffff",
            INIT_19 => X"ffffffdffffffffffffffff1fffffffffffffff1ffffffff0000001f00000000",
            INIT_1A => X"fffffff3fffffffffffffffffffffffffffffff8ffffffff0000001100000000",
            INIT_1B => X"0000000500000000ffffffedffffffffffffffe0ffffffff0000001000000000",
            INIT_1C => X"0000001300000000000000080000000000000000000000000000001200000000",
            INIT_1D => X"ffffffd7ffffffff00000005000000000000001e00000000fffffffcffffffff",
            INIT_1E => X"0000001200000000000000070000000000000027000000000000000c00000000",
            INIT_1F => X"fffffff7ffffffff0000000100000000fffffff2fffffffffffffffbffffffff",
            INIT_20 => X"ffffffe5ffffffffffffffe7ffffffff00000000000000000000000600000000",
            INIT_21 => X"ffffffe6ffffffffffffffeeffffffff0000000a000000000000002800000000",
            INIT_22 => X"0000001900000000fffffff4ffffffff0000000c00000000fffffff0ffffffff",
            INIT_23 => X"fffffff3ffffffffffffffefffffffffffffffeaffffffffffffffecffffffff",
            INIT_24 => X"fffffff4fffffffffffffff4ffffffff0000002500000000ffffffffffffffff",
            INIT_25 => X"ffffffceffffffff00000020000000000000000e00000000fffffffbffffffff",
            INIT_26 => X"00000005000000000000000200000000ffffff82ffffffff0000001c00000000",
            INIT_27 => X"fffffff0fffffffffffffff3ffffffff0000000a000000000000000300000000",
            INIT_28 => X"fffffff1ffffffff00000000000000000000000100000000ffffffe9ffffffff",
            INIT_29 => X"ffffffdbffffffffffffffedfffffffffffffff7ffffffff0000001d00000000",
            INIT_2A => X"fffffff7ffffffffffffffd5ffffffff0000000c000000000000000000000000",
            INIT_2B => X"0000000e000000000000000100000000fffffff4ffffffff0000000e00000000",
            INIT_2C => X"fffffffeffffffff00000001000000000000001300000000fffffff3ffffffff",
            INIT_2D => X"00000001000000000000001d000000000000001100000000fffffffbffffffff",
            INIT_2E => X"0000000900000000ffffffd9ffffffff0000001c000000000000000100000000",
            INIT_2F => X"fffffff1fffffffffffffff3fffffffffffffffcffffffff0000000e00000000",
            INIT_30 => X"ffffffffffffffff00000027000000000000000600000000ffffffefffffffff",
            INIT_31 => X"ffffffdafffffffffffffffcfffffffffffffffdffffffff0000000000000000",
            INIT_32 => X"fffffffcfffffffffffffff4ffffffff0000001900000000ffffffe8ffffffff",
            INIT_33 => X"fffffffafffffffffffffffdffffffff0000001e000000000000004300000000",
            INIT_34 => X"fffffffeffffffff0000001b00000000fffffff5ffffffff0000000000000000",
            INIT_35 => X"fffffff4ffffffff00000018000000000000001500000000fffffffdffffffff",
            INIT_36 => X"00000008000000000000000900000000ffffffc6ffffffff0000001900000000",
            INIT_37 => X"ffffffe5ffffffff0000000c00000000ffffffe2ffffffff0000001e00000000",
            INIT_38 => X"ffffffe1ffffffff0000000600000000fffffffefffffffffffffff8ffffffff",
            INIT_39 => X"0000000f000000000000000c00000000fffffffdffffffff0000001c00000000",
            INIT_3A => X"0000001100000000ffffffddffffffff00000022000000000000001300000000",
            INIT_3B => X"0000000e000000000000000800000000ffffffedffffffff0000000600000000",
            INIT_3C => X"0000001400000000fffffff7fffffffffffffff6ffffffff0000000000000000",
            INIT_3D => X"0000000b000000000000000100000000ffffffeefffffffffffffff2ffffffff",
            INIT_3E => X"ffffffbdffffffffffffffe3ffffffff0000001a00000000fffffff6ffffffff",
            INIT_3F => X"0000000700000000fffffff8ffffffff0000001700000000ffffffe0ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001100000000000000060000000000000048000000000000000500000000",
            INIT_41 => X"0000000500000000ffffffd0ffffffffffffffebffffffff0000001700000000",
            INIT_42 => X"fffffffefffffffffffffff1ffffffffffffffeefffffffffffffffeffffffff",
            INIT_43 => X"00000019000000000000000b00000000ffffffe9ffffffffffffffebffffffff",
            INIT_44 => X"0000000500000000fffffffeffffffffffffffcdffffffff0000000b00000000",
            INIT_45 => X"ffffffd0fffffffffffffffeffffffff00000005000000000000000400000000",
            INIT_46 => X"ffffffeeffffffff0000001000000000ffffffe1ffffffff0000000e00000000",
            INIT_47 => X"ffffffffffffffffffffffeefffffffffffffff9ffffffff0000000600000000",
            INIT_48 => X"0000000000000000fffffffbffffffff0000000700000000fffffffdffffffff",
            INIT_49 => X"fffffff3ffffffff0000000a0000000000000002000000000000000a00000000",
            INIT_4A => X"0000000d000000000000000000000000fffffff8ffffffffffffffe4ffffffff",
            INIT_4B => X"0000000900000000fffffffbffffffffffffffe8ffffffff0000000a00000000",
            INIT_4C => X"0000001400000000fffffff1ffffffff0000000b00000000fffffff9ffffffff",
            INIT_4D => X"ffffffdfffffffff0000001700000000fffffffdffffffffffffffefffffffff",
            INIT_4E => X"0000000d000000000000001000000000ffffffbaffffffffffffffe9ffffffff",
            INIT_4F => X"fffffff5fffffffffffffff3ffffffffffffffd5ffffffff0000002200000000",
            INIT_50 => X"0000000000000000ffffffe5ffffffff0000000e00000000ffffffefffffffff",
            INIT_51 => X"ffffffecffffffff000000000000000000000020000000000000001000000000",
            INIT_52 => X"ffffffeaffffffff0000001800000000fffffff3ffffffff0000001200000000",
            INIT_53 => X"00000024000000000000000800000000fffffffcfffffffffffffffcffffffff",
            INIT_54 => X"0000004400000000fffffffeffffffffffffffd8ffffffffffffffe3ffffffff",
            INIT_55 => X"0000000100000000fffffff4ffffffff0000001000000000fffffffbffffffff",
            INIT_56 => X"fffffffdfffffffffffffff0ffffffffffffffc1ffffffff0000000700000000",
            INIT_57 => X"00000009000000000000001100000000ffffffbefffffffffffffffdffffffff",
            INIT_58 => X"0000000000000000ffffffebffffffff0000000400000000fffffff6ffffffff",
            INIT_59 => X"ffffffe2ffffffff00000012000000000000002500000000fffffff8ffffffff",
            INIT_5A => X"0000000b000000000000003f00000000fffffff4fffffffffffffff1ffffffff",
            INIT_5B => X"0000000800000000fffffffefffffffffffffff5ffffffff0000001700000000",
            INIT_5C => X"0000002d000000000000000c00000000ffffffbbfffffffffffffff2ffffffff",
            INIT_5D => X"0000000d00000000fffffffffffffffffffffffbffffffff0000001e00000000",
            INIT_5E => X"0000002500000000ffffffe2ffffffffffffff85ffffffff0000000d00000000",
            INIT_5F => X"0000000a000000000000000000000000ffffffcdffffffff0000000d00000000",
            INIT_60 => X"ffffffe6ffffffffffffffe9ffffffff0000001300000000fffffff9ffffffff",
            INIT_61 => X"ffffffd6ffffffff0000001d000000000000001b000000000000000000000000",
            INIT_62 => X"0000000800000000fffffff3ffffffff00000005000000000000000200000000",
            INIT_63 => X"0000000000000000fffffffcffffffff0000000100000000fffffff1ffffffff",
            INIT_64 => X"0000000f00000000fffffff7fffffffffffffff4fffffffffffffff0ffffffff",
            INIT_65 => X"ffffffe0fffffffffffffff6ffffffff0000001e000000000000000c00000000",
            INIT_66 => X"ffffffeeffffffffffffffc7fffffffffffffffdffffffff0000000e00000000",
            INIT_67 => X"fffffff8ffffffffffffffd0ffffffffffffffe4ffffffff0000001c00000000",
            INIT_68 => X"ffffffdbffffffff0000000600000000fffffffcffffffffffffffe8ffffffff",
            INIT_69 => X"ffffffcfffffffff00000003000000000000001a000000000000000c00000000",
            INIT_6A => X"ffffffc9ffffffff00000002000000000000000a000000000000001600000000",
            INIT_6B => X"ffffffe7fffffffffffffff5ffffffff0000000d00000000ffffffdcffffffff",
            INIT_6C => X"0000001600000000fffffff4ffffffff0000001400000000ffffffdeffffffff",
            INIT_6D => X"ffffffeafffffffffffffff7ffffffff0000002600000000fffffffaffffffff",
            INIT_6E => X"ffffffe2ffffffff000000070000000000000027000000000000000800000000",
            INIT_6F => X"ffffffdaffffffff0000000000000000fffffff0ffffffff0000001100000000",
            INIT_70 => X"ffffffdaffffffff0000000200000000fffffff0ffffffffffffffe9ffffffff",
            INIT_71 => X"ffffffeaffffffffffffffdffffffffffffffff6ffffffff0000001300000000",
            INIT_72 => X"ffffffe3ffffffffffffffe3fffffffffffffffcffffffff0000001600000000",
            INIT_73 => X"ffffffecfffffffffffffff2fffffffffffffff0ffffffffffffffdeffffffff",
            INIT_74 => X"0000001900000000fffffff7ffffffff0000001300000000ffffffb8ffffffff",
            INIT_75 => X"00000013000000000000001c00000000ffffffe4ffffffffffffffe2ffffffff",
            INIT_76 => X"ffffff9afffffffffffffff8ffffffff0000003400000000ffffffe3ffffffff",
            INIT_77 => X"0000000a00000000fffffff6ffffffff0000003500000000ffffffe2ffffffff",
            INIT_78 => X"fffffff4fffffffffffffff1ffffffff0000002e00000000ffffffebffffffff",
            INIT_79 => X"0000001400000000ffffffbdfffffffffffffff8ffffffff0000001b00000000",
            INIT_7A => X"0000001a0000000000000015000000000000000900000000fffffff1ffffffff",
            INIT_7B => X"0000000000000000ffffffe7fffffffffffffff8ffffffffffffffffffffffff",
            INIT_7C => X"0000001300000000ffffffe4ffffffffffffffb7ffffffff0000000300000000",
            INIT_7D => X"ffffffb9ffffffff00000006000000000000000b000000000000002d00000000",
            INIT_7E => X"0000001200000000ffffffebffffffffffffffb6fffffffffffffff8ffffffff",
            INIT_7F => X"0000001200000000fffffff3ffffffff00000014000000000000001400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE28;


    MEM_IWGHT_LAYER2_INSTANCE29 : if BRAM_NAME = "iwght_layer2_instance29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffc2ffffffffffffffc4ffffffff0000000700000000ffffffe1ffffffff",
            INIT_01 => X"ffffffeeffffffff000000210000000000000027000000000000000e00000000",
            INIT_02 => X"00000025000000000000002d000000000000001f000000000000000b00000000",
            INIT_03 => X"0000000900000000ffffffccffffffff00000029000000000000001d00000000",
            INIT_04 => X"0000002100000000fffffffaffffffffffffffe3ffffffff0000000800000000",
            INIT_05 => X"ffffffc8ffffffffffffffcdffffffffffffffebffffffff0000001000000000",
            INIT_06 => X"0000002900000000ffffffe4ffffffffffffffaefffffffffffffff0ffffffff",
            INIT_07 => X"00000002000000000000001400000000ffffffdeffffffff0000002200000000",
            INIT_08 => X"fffffff8ffffffffffffffafffffffff0000002100000000fffffff2ffffffff",
            INIT_09 => X"0000000f0000000000000014000000000000001d00000000fffffff0ffffffff",
            INIT_0A => X"0000000d000000000000002f0000000000000002000000000000003900000000",
            INIT_0B => X"fffffffaffffffffffffffeaffffffff00000014000000000000002600000000",
            INIT_0C => X"0000003800000000ffffffdcffffffffffffffbeffffffff0000000200000000",
            INIT_0D => X"ffffffe4ffffffffffffffddffffffff0000001d000000000000002300000000",
            INIT_0E => X"0000003c00000000ffffffd0ffffffffffffff8bffffffff0000000000000000",
            INIT_0F => X"00000022000000000000003200000000ffffffe8ffffffff0000003c00000000",
            INIT_10 => X"ffffffeeffffffffffffffc5ffffffff0000001400000000ffffffebffffffff",
            INIT_11 => X"fffffffdffffffff0000001f000000000000002e000000000000000000000000",
            INIT_12 => X"00000022000000000000002800000000fffffff4ffffffff0000002c00000000",
            INIT_13 => X"ffffffe4ffffffff00000006000000000000001f000000000000001300000000",
            INIT_14 => X"0000003100000000fffffff7ffffffffffffffd2ffffffffffffffedffffffff",
            INIT_15 => X"0000002900000000ffffffccfffffffffffffff8ffffffff0000004c00000000",
            INIT_16 => X"0000001c00000000ffffffd9ffffffffffffffabffffffff0000000b00000000",
            INIT_17 => X"0000000a00000000fffffffbffffffffffffffd6ffffffff0000002500000000",
            INIT_18 => X"ffffffe7fffffffffffffffffffffffffffffff8ffffffffffffffedffffffff",
            INIT_19 => X"ffffffeaffffffff0000003d0000000000000019000000000000000900000000",
            INIT_1A => X"00000000000000000000001f00000000fffffff9ffffffff0000002e00000000",
            INIT_1B => X"fffffffaffffffff000000030000000000000011000000000000001d00000000",
            INIT_1C => X"0000000c00000000ffffffefffffffffffffffc3ffffffff0000001300000000",
            INIT_1D => X"ffffffe7ffffffff0000000c0000000000000005000000000000002b00000000",
            INIT_1E => X"0000002100000000ffffffe5ffffffffffffffbbffffffff0000000d00000000",
            INIT_1F => X"0000000c00000000000000050000000000000007000000000000003800000000",
            INIT_20 => X"ffffffcbffffffffffffffe2ffffffffffffffdfffffffffffffffdcffffffff",
            INIT_21 => X"ffffffd7ffffffff000000140000000000000012000000000000000400000000",
            INIT_22 => X"fffffff1ffffffff000000190000000000000007000000000000001e00000000",
            INIT_23 => X"ffffffe1ffffffff0000000a000000000000001b00000000ffffffeeffffffff",
            INIT_24 => X"0000001a00000000ffffffe7fffffffffffffffbffffffffffffffe1ffffffff",
            INIT_25 => X"ffffffddffffffff0000000f00000000ffffffefffffffff0000000000000000",
            INIT_26 => X"ffffffd4ffffffff00000006000000000000001f00000000fffffffcffffffff",
            INIT_27 => X"000000160000000000000016000000000000000a000000000000000400000000",
            INIT_28 => X"00000000000000000000000900000000ffffffe1fffffffffffffffbffffffff",
            INIT_29 => X"ffffffe8ffffffffffffffebffffffffffffffe6ffffffff0000001300000000",
            INIT_2A => X"ffffffecffffffffffffffffffffffffffffffc4ffffffff0000000f00000000",
            INIT_2B => X"fffffff4ffffffff0000001300000000ffffffedffffffffffffffceffffffff",
            INIT_2C => X"0000001200000000fffffff0ffffffff0000002e00000000ffffffc4ffffffff",
            INIT_2D => X"000000230000000000000014000000000000000300000000ffffffd2ffffffff",
            INIT_2E => X"ffffffcffffffffffffffff8ffffffffffffffa3ffffffffffffffefffffffff",
            INIT_2F => X"0000000a000000000000000c000000000000003c00000000ffffffdfffffffff",
            INIT_30 => X"0000001a0000000000000016000000000000001700000000ffffffdaffffffff",
            INIT_31 => X"0000000400000000ffffffa8ffffffffffffffb9ffffffff0000002a00000000",
            INIT_32 => X"00000024000000000000001000000000ffffffe6fffffffffffffff6ffffffff",
            INIT_33 => X"ffffffeeffffffff0000001000000000fffffff9fffffffffffffff4ffffffff",
            INIT_34 => X"0000001200000000ffffffeafffffffffffffff3ffffffff0000001200000000",
            INIT_35 => X"ffffffd2ffffffff0000000f000000000000000e00000000fffffffcffffffff",
            INIT_36 => X"ffffffd6ffffffff0000000900000000ffffffc0fffffffffffffff2ffffffff",
            INIT_37 => X"0000000e00000000ffffffdeffffffff0000000e000000000000000e00000000",
            INIT_38 => X"0000000900000000ffffffdfffffffff0000000e00000000ffffffd6ffffffff",
            INIT_39 => X"ffffffecffffffff000000030000000000000002000000000000000a00000000",
            INIT_3A => X"00000041000000000000001c00000000ffffffedffffffff0000002000000000",
            INIT_3B => X"fffffffbfffffffffffffffdffffffffffffffefffffffff0000001000000000",
            INIT_3C => X"00000000000000000000000500000000ffffffceffffffff0000001300000000",
            INIT_3D => X"ffffffd5ffffffffffffffdcffffffff00000017000000000000001f00000000",
            INIT_3E => X"00000023000000000000000200000000ffffffc1fffffffffffffff9ffffffff",
            INIT_3F => X"0000001600000000ffffffffffffffff00000010000000000000000600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002000000000ffffffb2fffffffffffffff4ffffffffffffffe1ffffffff",
            INIT_41 => X"00000025000000000000001600000000fffffffdffffffff0000000800000000",
            INIT_42 => X"0000001700000000000000190000000000000000000000000000001300000000",
            INIT_43 => X"00000009000000000000000d0000000000000012000000000000001300000000",
            INIT_44 => X"00000011000000000000000000000000ffffffdaffffffffffffffeaffffffff",
            INIT_45 => X"ffffffb9ffffffffffffffb3ffffffff0000001b00000000fffffff1ffffffff",
            INIT_46 => X"0000002500000000ffffffceffffffffffffff52fffffffffffffffeffffffff",
            INIT_47 => X"0000002500000000fffffffaffffffffffffffdcffffffff0000003100000000",
            INIT_48 => X"ffffffefffffffffffffffceffffffffffffffffffffffffffffffd8ffffffff",
            INIT_49 => X"00000007000000000000000e0000000000000027000000000000000c00000000",
            INIT_4A => X"00000003000000000000001d0000000000000007000000000000001300000000",
            INIT_4B => X"fffffff4ffffffff0000000b0000000000000006000000000000000b00000000",
            INIT_4C => X"0000000a00000000ffffffecffffffffffffffd1fffffffffffffffaffffffff",
            INIT_4D => X"ffffffebffffffffffffffc4fffffffffffffffeffffffff0000001800000000",
            INIT_4E => X"fffffffcffffffffffffffbeffffffffffffff97fffffffffffffffdffffffff",
            INIT_4F => X"fffffff4ffffffff00000015000000000000000a000000000000001f00000000",
            INIT_50 => X"0000000000000000ffffffd1ffffffffffffffe5ffffffffffffffd7ffffffff",
            INIT_51 => X"ffffffe5fffffffffffffff7ffffffff0000000d000000000000000e00000000",
            INIT_52 => X"00000000000000000000000d0000000000000010000000000000001200000000",
            INIT_53 => X"ffffffddffffffff0000001800000000ffffffeeffffffff0000000500000000",
            INIT_54 => X"0000001500000000fffffff1ffffffffffffffe3ffffffffffffffeeffffffff",
            INIT_55 => X"ffffffd2ffffffffffffffdeffffffffffffffe5ffffffff0000002800000000",
            INIT_56 => X"ffffffe3ffffffff0000000100000000ffffff6bfffffffffffffff9ffffffff",
            INIT_57 => X"ffffffeffffffffffffffff7ffffffff0000002c000000000000001e00000000",
            INIT_58 => X"0000000c00000000ffffffdfffffffffffffffe6ffffffffffffffe2ffffffff",
            INIT_59 => X"ffffffe3ffffffff0000000e00000000fffffff8ffffffff0000001b00000000",
            INIT_5A => X"0000001c0000000000000027000000000000001b000000000000000400000000",
            INIT_5B => X"fffffff1ffffffff0000002e000000000000000b00000000fffffff3ffffffff",
            INIT_5C => X"0000001a0000000000000006000000000000000600000000ffffffbfffffffff",
            INIT_5D => X"ffffffabffffffffffffffe8ffffffffffffffdaffffffffffffffbfffffffff",
            INIT_5E => X"ffffff8cffffffff0000003a000000000000000a00000000fffffff8ffffffff",
            INIT_5F => X"0000000f000000000000000d00000000fffffff8ffffffff0000002100000000",
            INIT_60 => X"0000001400000000ffffffdeffffffff0000000100000000fffffff4ffffffff",
            INIT_61 => X"0000000d000000000000000a00000000ffffffbfffffffff0000002200000000",
            INIT_62 => X"0000000800000000fffffff8ffffffffffffffb1ffffffff0000000f00000000",
            INIT_63 => X"ffffffedffffffff0000002e000000000000000300000000ffffffefffffffff",
            INIT_64 => X"0000000f00000000ffffffe3ffffffff0000003300000000ffffffd3ffffffff",
            INIT_65 => X"ffffffceffffffff00000019000000000000000100000000ffffffd1ffffffff",
            INIT_66 => X"fffffff2ffffffffffffffd5ffffffffffffffc5ffffffffffffffc2ffffffff",
            INIT_67 => X"ffffffc9ffffffff00000013000000000000003400000000ffffffcfffffffff",
            INIT_68 => X"fffffffdffffffff0000000500000000ffffffe9fffffffffffffff9ffffffff",
            INIT_69 => X"0000000200000000fffffffbffffffffffffffabffffffff0000002000000000",
            INIT_6A => X"0000002b000000000000000200000000ffffffd9ffffffffffffffd5ffffffff",
            INIT_6B => X"ffffffd9ffffffff0000002100000000ffffffddffffffffffffffe6ffffffff",
            INIT_6C => X"0000001900000000ffffffe2ffffffff0000000d00000000ffffffeeffffffff",
            INIT_6D => X"fffffffeffffffff0000001500000000ffffffdaffffffff0000001700000000",
            INIT_6E => X"ffffffe5fffffffffffffff1ffffffffffffffb7ffffffff0000000800000000",
            INIT_6F => X"ffffffd8ffffffffffffffd0ffffffff0000001600000000fffffff8ffffffff",
            INIT_70 => X"0000000d00000000ffffffe4fffffffffffffff1ffffffffffffffd8ffffffff",
            INIT_71 => X"ffffffefffffffff0000000000000000ffffffe7ffffffff0000002200000000",
            INIT_72 => X"0000005d0000000000000010000000000000000600000000ffffffe6ffffffff",
            INIT_73 => X"fffffff1ffffffff0000001300000000ffffffc5ffffffffffffffd6ffffffff",
            INIT_74 => X"000000010000000000000008000000000000001e00000000fffffff6ffffffff",
            INIT_75 => X"ffffffe7fffffffffffffff2ffffffffffffffb5ffffffff0000001400000000",
            INIT_76 => X"fffffffffffffffffffffff5ffffffffffffff90ffffffffffffffedffffffff",
            INIT_77 => X"fffffffcffffffffffffffe8ffffffff0000001100000000fffffffdffffffff",
            INIT_78 => X"0000001800000000ffffffcaffffffff0000000000000000fffffff7ffffffff",
            INIT_79 => X"00000005000000000000000400000000ffffffedffffffff0000002c00000000",
            INIT_7A => X"0000001d000000000000001800000000fffffff0ffffffffffffffd9ffffffff",
            INIT_7B => X"fffffff1ffffffff0000002a00000000ffffffe4fffffffffffffff1ffffffff",
            INIT_7C => X"ffffffe9ffffffffffffffecfffffffffffffffcffffffff0000000f00000000",
            INIT_7D => X"ffffffc4ffffffffffffffdafffffffffffffff1ffffffff0000000c00000000",
            INIT_7E => X"0000004700000000ffffffd1ffffffffffffff84fffffffffffffff4ffffffff",
            INIT_7F => X"0000000f00000000ffffffe6ffffffff0000000b00000000fffffffeffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE29;


    MEM_IWGHT_LAYER2_INSTANCE30 : if BRAM_NAME = "iwght_layer2_instance30" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003400000000fffffff1fffffffffffffff9ffffffffffffffe8ffffffff",
            INIT_01 => X"0000001400000000fffffff0ffffffffffffffdfffffffff0000000200000000",
            INIT_02 => X"0000003100000000fffffff3ffffffffffffffe7ffffffffffffffd3ffffffff",
            INIT_03 => X"000000050000000000000026000000000000001000000000fffffff0ffffffff",
            INIT_04 => X"ffffffdafffffffffffffff4ffffffff0000000800000000ffffffdcffffffff",
            INIT_05 => X"00000016000000000000000100000000fffffff0ffffffff0000000800000000",
            INIT_06 => X"0000004900000000ffffffeeffffffffffffffabffffffffffffffecffffffff",
            INIT_07 => X"0000000200000000ffffffecffffffff0000000d00000000fffffff5ffffffff",
            INIT_08 => X"0000001e00000000ffffffb4fffffffffffffff3ffffffffffffffe1ffffffff",
            INIT_09 => X"ffffffecfffffffffffffffffffffffffffffffeffffffff0000001200000000",
            INIT_0A => X"000000450000000000000006000000000000000000000000ffffffecffffffff",
            INIT_0B => X"00000005000000000000002600000000ffffffdeffffffffffffffe8ffffffff",
            INIT_0C => X"0000000100000000ffffffe2ffffffff0000000500000000ffffffebffffffff",
            INIT_0D => X"ffffffe1ffffffff0000000600000000ffffffe2ffffffff0000001000000000",
            INIT_0E => X"00000019000000000000000200000000ffffffcaffffffff0000001000000000",
            INIT_0F => X"ffffffe9fffffffffffffff0ffffffff0000001b00000000fffffff7ffffffff",
            INIT_10 => X"0000001000000000ffffffb1ffffffffffffffdeffffffffffffffe6ffffffff",
            INIT_11 => X"ffffffeafffffffffffffff8ffffffff00000002000000000000001f00000000",
            INIT_12 => X"000000210000000000000029000000000000002400000000fffffff0ffffffff",
            INIT_13 => X"000000030000000000000016000000000000000b00000000fffffff8ffffffff",
            INIT_14 => X"0000000d00000000fffffff5ffffffff0000001200000000ffffffebffffffff",
            INIT_15 => X"ffffffdcffffffff0000000000000000ffffffddffffffffffffffe5ffffffff",
            INIT_16 => X"fffffff6ffffffff0000002900000000fffffff7ffffffffffffffe5ffffffff",
            INIT_17 => X"0000000f000000000000001e000000000000003400000000fffffff0ffffffff",
            INIT_18 => X"0000001600000000ffffffeafffffffffffffff2ffffffff0000000400000000",
            INIT_19 => X"00000016000000000000000d00000000ffffffaaffffffff0000001600000000",
            INIT_1A => X"0000003f00000000ffffffc3ffffffffffffffecffffffffffffffecffffffff",
            INIT_1B => X"00000011000000000000003c000000000000000500000000fffffff7ffffffff",
            INIT_1C => X"ffffffbcffffffffffffffe3ffffffff0000000a00000000fffffffdffffffff",
            INIT_1D => X"fffffffaffffffff00000000000000000000001a00000000ffffffe6ffffffff",
            INIT_1E => X"0000004200000000ffffffcbffffffffffffffebffffffffffffffe0ffffffff",
            INIT_1F => X"ffffff95ffffffff00000026000000000000002700000000ffffff88ffffffff",
            INIT_20 => X"fffffffdffffffff0000001000000000ffffff8dffffffff0000000400000000",
            INIT_21 => X"fffffff9ffffffff0000000200000000ffffffbffffffffffffffff9ffffffff",
            INIT_22 => X"00000044000000000000000000000000ffffffd3ffffffffffffffd8ffffffff",
            INIT_23 => X"0000000b000000000000004700000000ffffffcbffffffffffffffe7ffffffff",
            INIT_24 => X"0000001b00000000ffffffd1ffffffff0000000400000000ffffffedffffffff",
            INIT_25 => X"ffffffdcffffffff0000001a00000000ffffffc8fffffffffffffff9ffffffff",
            INIT_26 => X"00000033000000000000000000000000ffffff41ffffffff0000000000000000",
            INIT_27 => X"ffffffccffffffffffffffebffffffff0000002900000000fffffff7ffffffff",
            INIT_28 => X"fffffffaffffffffffffffe4ffffffffffffffcaffffffffffffffedffffffff",
            INIT_29 => X"fffffff3ffffffff0000000a00000000ffffffd3ffffffff0000003100000000",
            INIT_2A => X"0000003a00000000fffffffeffffffff0000000d00000000ffffffefffffffff",
            INIT_2B => X"00000010000000000000003400000000ffffffd2ffffffffffffffd3ffffffff",
            INIT_2C => X"fffffff9ffffffff00000017000000000000001700000000fffffff6ffffffff",
            INIT_2D => X"ffffffe1ffffffff0000001000000000ffffffc3ffffffff0000000300000000",
            INIT_2E => X"0000002400000000fffffff8fffffffffffffffaffffffff0000000f00000000",
            INIT_2F => X"0000000000000000ffffffe4ffffffff0000002500000000ffffffe4ffffffff",
            INIT_30 => X"0000003300000000ffffffbdffffffffffffffd9ffffffffffffffeeffffffff",
            INIT_31 => X"00000005000000000000000800000000fffffff9ffffffff0000000d00000000",
            INIT_32 => X"0000005700000000ffffffcefffffffffffffffffffffffffffffff8ffffffff",
            INIT_33 => X"00000022000000000000001300000000ffffffdbffffffffffffffe5ffffffff",
            INIT_34 => X"ffffffd2ffffffffffffffffffffffff00000009000000000000001400000000",
            INIT_35 => X"fffffffbffffffff0000002300000000ffffffecffffffff0000000100000000",
            INIT_36 => X"0000003e000000000000001700000000ffffffe3ffffffffffffffe5ffffffff",
            INIT_37 => X"fffffffdffffffffffffffcdffffffff0000001a00000000ffffffe9ffffffff",
            INIT_38 => X"0000001300000000fffffffaffffffff0000000000000000ffffffeeffffffff",
            INIT_39 => X"fffffff9ffffffff0000000a00000000ffffffffffffffff0000000000000000",
            INIT_3A => X"0000003e00000000fffffff9ffffffffffffffe3ffffffffffffffd6ffffffff",
            INIT_3B => X"00000022000000000000001300000000ffffffe5ffffffffffffffd7ffffffff",
            INIT_3C => X"fffffff2ffffffff0000000c00000000ffffffe0fffffffffffffffaffffffff",
            INIT_3D => X"00000016000000000000000900000000ffffffe8ffffffff0000001d00000000",
            INIT_3E => X"0000004a000000000000000000000000ffffffa9ffffffffffffffccffffffff",
            INIT_3F => X"0000000300000000ffffffdfffffffff0000001c00000000ffffffe1ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001500000000fffffffbffffffffffffffe5ffffffffffffffe6ffffffff",
            INIT_41 => X"ffffffe6ffffffff0000002100000000ffffffdaffffffff0000000d00000000",
            INIT_42 => X"0000005f00000000ffffffeaffffffffffffffedfffffffffffffffbffffffff",
            INIT_43 => X"0000002e000000000000000a00000000ffffffdfffffffffffffffd6ffffffff",
            INIT_44 => X"fffffff2ffffffff000000140000000000000008000000000000000f00000000",
            INIT_45 => X"ffffffd9ffffffff0000000f00000000fffffffeffffffff0000000a00000000",
            INIT_46 => X"00000033000000000000000b00000000ffffffb9ffffffffffffffd7ffffffff",
            INIT_47 => X"fffffff1fffffffffffffff0ffffffff00000016000000000000000300000000",
            INIT_48 => X"0000003000000000ffffffb7ffffffffffffffdeffffffffffffffe8ffffffff",
            INIT_49 => X"0000000000000000ffffffffffffffffffffffe6ffffffff0000001100000000",
            INIT_4A => X"00000038000000000000000200000000ffffffecffffffff0000000400000000",
            INIT_4B => X"0000000000000000ffffffebffffffff0000000800000000fffffffcffffffff",
            INIT_4C => X"ffffffccfffffffffffffffffffffffffffffffaffffffffffffffd6ffffffff",
            INIT_4D => X"ffffffcdffffffff00000016000000000000000000000000ffffffd8ffffffff",
            INIT_4E => X"0000003d0000000000000021000000000000000200000000ffffffaeffffffff",
            INIT_4F => X"0000000f00000000fffffff9ffffffff0000002a00000000ffffffb3ffffffff",
            INIT_50 => X"0000003e00000000ffffffa1ffffffff0000000600000000fffffff8ffffffff",
            INIT_51 => X"00000019000000000000000500000000ffffffadfffffffffffffff8ffffffff",
            INIT_52 => X"ffffffc4ffffffffffffffdcffffffff",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE30;


    MEM_IFMAP_LAYER0_INSTANCE0 : if BRAM_NAME = "ifmap_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a600000000000000a5000000000000009f000000000000009e00000000",
            INIT_01 => X"0000009f00000000000000a2000000000000009c00000000000000a000000000",
            INIT_02 => X"000000a000000000000000a1000000000000009f000000000000009e00000000",
            INIT_03 => X"000000aa00000000000000a900000000000000a600000000000000a100000000",
            INIT_04 => X"000000a000000000000000a000000000000000a200000000000000a700000000",
            INIT_05 => X"0000009400000000000000960000000000000095000000000000009c00000000",
            INIT_06 => X"0000008d000000000000008c000000000000008f000000000000009500000000",
            INIT_07 => X"00000074000000000000007e0000000000000089000000000000008f00000000",
            INIT_08 => X"000000a6000000000000009f0000000000000097000000000000009800000000",
            INIT_09 => X"000000a200000000000000a400000000000000a000000000000000a200000000",
            INIT_0A => X"0000009f000000000000009b000000000000009c00000000000000a300000000",
            INIT_0B => X"000000ab00000000000000ab00000000000000aa00000000000000a300000000",
            INIT_0C => X"00000097000000000000009a00000000000000a000000000000000a900000000",
            INIT_0D => X"0000008d000000000000008c000000000000008b000000000000009100000000",
            INIT_0E => X"0000008e00000000000000910000000000000093000000000000009500000000",
            INIT_0F => X"00000077000000000000007d0000000000000088000000000000008f00000000",
            INIT_10 => X"000000a7000000000000009e0000000000000097000000000000009700000000",
            INIT_11 => X"000000a500000000000000a500000000000000a300000000000000a000000000",
            INIT_12 => X"0000009d000000000000009e00000000000000a200000000000000a300000000",
            INIT_13 => X"000000a900000000000000a700000000000000a600000000000000a100000000",
            INIT_14 => X"000000790000000000000091000000000000009f00000000000000aa00000000",
            INIT_15 => X"0000007200000000000000650000000000000062000000000000006e00000000",
            INIT_16 => X"0000008c000000000000008f0000000000000086000000000000007800000000",
            INIT_17 => X"000000780000000000000082000000000000008b000000000000008e00000000",
            INIT_18 => X"000000ae00000000000000a0000000000000009b000000000000009b00000000",
            INIT_19 => X"000000a900000000000000a900000000000000a700000000000000a700000000",
            INIT_1A => X"000000bf00000000000000a700000000000000a500000000000000a500000000",
            INIT_1B => X"000000a400000000000000a2000000000000009d00000000000000b100000000",
            INIT_1C => X"0000006700000000000000680000000000000095000000000000009e00000000",
            INIT_1D => X"0000004a0000000000000050000000000000005c000000000000006200000000",
            INIT_1E => X"0000008400000000000000710000000000000053000000000000005600000000",
            INIT_1F => X"0000007f0000000000000088000000000000008c000000000000008c00000000",
            INIT_20 => X"000000aa00000000000000a1000000000000009c000000000000009b00000000",
            INIT_21 => X"000000a600000000000000a900000000000000a300000000000000a900000000",
            INIT_22 => X"000000f600000000000000ad00000000000000a400000000000000a400000000",
            INIT_23 => X"0000008e0000000000000092000000000000009700000000000000c300000000",
            INIT_24 => X"000000710000000000000055000000000000004e000000000000006f00000000",
            INIT_25 => X"0000005d0000000000000061000000000000006a000000000000007000000000",
            INIT_26 => X"0000006900000000000000550000000000000054000000000000004a00000000",
            INIT_27 => X"000000810000000000000085000000000000008a000000000000008000000000",
            INIT_28 => X"0000009300000000000000820000000000000085000000000000009400000000",
            INIT_29 => X"000000a700000000000000a700000000000000a500000000000000a100000000",
            INIT_2A => X"000000b400000000000000a300000000000000a500000000000000a300000000",
            INIT_2B => X"0000004200000000000000610000000000000080000000000000009d00000000",
            INIT_2C => X"0000007600000000000000590000000000000042000000000000004500000000",
            INIT_2D => X"0000005e00000000000000720000000000000077000000000000007a00000000",
            INIT_2E => X"00000043000000000000003a000000000000005b000000000000006300000000",
            INIT_2F => X"00000086000000000000008a000000000000008c000000000000006c00000000",
            INIT_30 => X"00000058000000000000002f000000000000006d000000000000007f00000000",
            INIT_31 => X"000000aa00000000000000a800000000000000aa000000000000009900000000",
            INIT_32 => X"0000009300000000000000a400000000000000a600000000000000a900000000",
            INIT_33 => X"000000440000000000000064000000000000007f000000000000008100000000",
            INIT_34 => X"0000008400000000000000530000000000000048000000000000004e00000000",
            INIT_35 => X"0000006b0000000000000069000000000000007c000000000000009200000000",
            INIT_36 => X"0000002e000000000000003f0000000000000055000000000000007300000000",
            INIT_37 => X"00000086000000000000008d0000000000000084000000000000004f00000000",
            INIT_38 => X"00000046000000000000002a0000000000000063000000000000008300000000",
            INIT_39 => X"000000a800000000000000a500000000000000a7000000000000008f00000000",
            INIT_3A => X"00000078000000000000008c00000000000000a100000000000000ab00000000",
            INIT_3B => X"0000005800000000000000740000000000000090000000000000008200000000",
            INIT_3C => X"0000007c000000000000004d0000000000000055000000000000005b00000000",
            INIT_3D => X"0000006a0000000000000066000000000000008800000000000000a300000000",
            INIT_3E => X"0000003100000000000000360000000000000055000000000000006400000000",
            INIT_3F => X"00000088000000000000008a000000000000006b000000000000003900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007c0000000000000036000000000000006700000000000000aa00000000",
            INIT_41 => X"000000a600000000000000a300000000000000a1000000000000009900000000",
            INIT_42 => X"0000007d000000000000007100000000000000ae00000000000000a500000000",
            INIT_43 => X"000000560000000000000079000000000000009c000000000000009d00000000",
            INIT_44 => X"0000005100000000000000500000000000000054000000000000005200000000",
            INIT_45 => X"0000005700000000000000710000000000000092000000000000008a00000000",
            INIT_46 => X"0000003800000000000000470000000000000056000000000000005300000000",
            INIT_47 => X"000000890000000000000085000000000000004a000000000000002800000000",
            INIT_48 => X"0000009a000000000000005e000000000000008600000000000000b400000000",
            INIT_49 => X"00000099000000000000009c000000000000009e00000000000000ae00000000",
            INIT_4A => X"0000009c00000000000000cf00000000000000ed00000000000000cf00000000",
            INIT_4B => X"0000005d000000000000007d000000000000009400000000000000ae00000000",
            INIT_4C => X"0000004c000000000000003b000000000000004a000000000000005600000000",
            INIT_4D => X"0000006a0000000000000085000000000000008f000000000000008900000000",
            INIT_4E => X"0000004b00000000000000540000000000000057000000000000005600000000",
            INIT_4F => X"00000084000000000000005f0000000000000028000000000000003200000000",
            INIT_50 => X"000000a5000000000000008e000000000000006c00000000000000b700000000",
            INIT_51 => X"0000007a000000000000009f000000000000009b00000000000000b100000000",
            INIT_52 => X"000000a400000000000000dc00000000000000ed00000000000000d500000000",
            INIT_53 => X"00000078000000000000007d000000000000009c00000000000000b700000000",
            INIT_54 => X"0000005b000000000000002d0000000000000050000000000000004e00000000",
            INIT_55 => X"0000006b000000000000009b000000000000009d00000000000000af00000000",
            INIT_56 => X"0000004e00000000000000580000000000000067000000000000005700000000",
            INIT_57 => X"00000068000000000000003b0000000000000029000000000000003b00000000",
            INIT_58 => X"000000aa0000000000000087000000000000006400000000000000bc00000000",
            INIT_59 => X"0000008600000000000000ad00000000000000a600000000000000bb00000000",
            INIT_5A => X"000000aa00000000000000c700000000000000c2000000000000007500000000",
            INIT_5B => X"00000075000000000000008600000000000000bd00000000000000b900000000",
            INIT_5C => X"0000007d00000000000000260000000000000054000000000000006600000000",
            INIT_5D => X"0000005d000000000000009200000000000000a000000000000000d200000000",
            INIT_5E => X"000000550000000000000068000000000000005e000000000000005300000000",
            INIT_5F => X"0000004c000000000000003e0000000000000037000000000000004900000000",
            INIT_60 => X"000000af000000000000007f000000000000005a00000000000000bd00000000",
            INIT_61 => X"0000009f00000000000000b200000000000000a600000000000000ae00000000",
            INIT_62 => X"0000008900000000000000a800000000000000a8000000000000006100000000",
            INIT_63 => X"0000007b00000000000000a000000000000000d800000000000000ba00000000",
            INIT_64 => X"0000009600000000000000320000000000000073000000000000007800000000",
            INIT_65 => X"0000005b000000000000007b000000000000009b00000000000000c200000000",
            INIT_66 => X"00000056000000000000005f0000000000000054000000000000005400000000",
            INIT_67 => X"00000049000000000000004f0000000000000049000000000000005400000000",
            INIT_68 => X"000000b90000000000000098000000000000005d00000000000000bd00000000",
            INIT_69 => X"000000a700000000000000ad0000000000000088000000000000007700000000",
            INIT_6A => X"000000a700000000000000910000000000000093000000000000006700000000",
            INIT_6B => X"0000008d00000000000000b400000000000000e200000000000000bd00000000",
            INIT_6C => X"0000009a00000000000000470000000000000075000000000000007e00000000",
            INIT_6D => X"000000570000000000000072000000000000009500000000000000ba00000000",
            INIT_6E => X"0000006300000000000000500000000000000048000000000000005000000000",
            INIT_6F => X"0000005e0000000000000061000000000000005a000000000000006400000000",
            INIT_70 => X"000000ba00000000000000a8000000000000006c00000000000000c200000000",
            INIT_71 => X"000000a7000000000000009c0000000000000063000000000000006900000000",
            INIT_72 => X"000000c6000000000000008a0000000000000073000000000000006400000000",
            INIT_73 => X"0000009a000000000000009100000000000000ac00000000000000be00000000",
            INIT_74 => X"0000009800000000000000470000000000000067000000000000009200000000",
            INIT_75 => X"0000006e0000000000000082000000000000008900000000000000b300000000",
            INIT_76 => X"0000006d000000000000005f000000000000005b000000000000005500000000",
            INIT_77 => X"0000007500000000000000610000000000000064000000000000007300000000",
            INIT_78 => X"000000b800000000000000ac000000000000008400000000000000c500000000",
            INIT_79 => X"0000009b000000000000008c000000000000004e000000000000008200000000",
            INIT_7A => X"000000e6000000000000008f0000000000000082000000000000007300000000",
            INIT_7B => X"000000830000000000000087000000000000009100000000000000f200000000",
            INIT_7C => X"00000090000000000000005f000000000000006c000000000000007900000000",
            INIT_7D => X"000000570000000000000070000000000000009800000000000000a800000000",
            INIT_7E => X"0000007000000000000000690000000000000057000000000000004700000000",
            INIT_7F => X"0000008800000000000000790000000000000067000000000000007800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE0;


    MEM_IFMAP_LAYER0_INSTANCE1 : if BRAM_NAME = "ifmap_layer0_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bf00000000000000a8000000000000009200000000000000cb00000000",
            INIT_01 => X"0000008a000000000000007e000000000000004e00000000000000a800000000",
            INIT_02 => X"000000ad000000000000009a0000000000000060000000000000008a00000000",
            INIT_03 => X"000000710000000000000071000000000000008c00000000000000a200000000",
            INIT_04 => X"000000ab00000000000000700000000000000069000000000000006500000000",
            INIT_05 => X"0000006d00000000000000870000000000000094000000000000009c00000000",
            INIT_06 => X"00000065000000000000005e000000000000004f000000000000004e00000000",
            INIT_07 => X"000000900000000000000097000000000000007d000000000000006b00000000",
            INIT_08 => X"000000b700000000000000a400000000000000a300000000000000d600000000",
            INIT_09 => X"0000009c0000000000000060000000000000005e00000000000000b000000000",
            INIT_0A => X"000000760000000000000081000000000000006a000000000000009400000000",
            INIT_0B => X"0000007300000000000000660000000000000074000000000000007200000000",
            INIT_0C => X"0000007600000000000000900000000000000065000000000000005600000000",
            INIT_0D => X"0000004b00000000000000850000000000000080000000000000004400000000",
            INIT_0E => X"000000660000000000000047000000000000003a000000000000003c00000000",
            INIT_0F => X"0000008c0000000000000096000000000000008f000000000000007400000000",
            INIT_10 => X"000000ad00000000000000a700000000000000b200000000000000d400000000",
            INIT_11 => X"0000008d0000000000000056000000000000007c00000000000000b000000000",
            INIT_12 => X"0000004d00000000000000680000000000000087000000000000009900000000",
            INIT_13 => X"000000930000000000000081000000000000007c000000000000008600000000",
            INIT_14 => X"000000840000000000000096000000000000005c000000000000005500000000",
            INIT_15 => X"00000040000000000000004b000000000000006b000000000000007500000000",
            INIT_16 => X"0000008500000000000000560000000000000041000000000000002c00000000",
            INIT_17 => X"00000097000000000000009a00000000000000a0000000000000009b00000000",
            INIT_18 => X"000000ae00000000000000ab00000000000000bb00000000000000c700000000",
            INIT_19 => X"000000770000000000000056000000000000009000000000000000b100000000",
            INIT_1A => X"0000004600000000000000900000000000000089000000000000007a00000000",
            INIT_1B => X"000000b80000000000000091000000000000006c000000000000008100000000",
            INIT_1C => X"0000008900000000000000830000000000000049000000000000007400000000",
            INIT_1D => X"0000003400000000000000330000000000000059000000000000008600000000",
            INIT_1E => X"000000a30000000000000079000000000000005a000000000000002f00000000",
            INIT_1F => X"00000095000000000000009e00000000000000a400000000000000ab00000000",
            INIT_20 => X"000000b100000000000000b300000000000000c300000000000000a500000000",
            INIT_21 => X"000000830000000000000063000000000000009800000000000000b500000000",
            INIT_22 => X"00000050000000000000005d000000000000006700000000000000ab00000000",
            INIT_23 => X"000000bf00000000000000b2000000000000007a000000000000005d00000000",
            INIT_24 => X"0000005700000000000000590000000000000064000000000000009600000000",
            INIT_25 => X"000000180000000000000026000000000000002e000000000000003c00000000",
            INIT_26 => X"00000090000000000000006c000000000000003c000000000000002e00000000",
            INIT_27 => X"00000078000000000000007f0000000000000080000000000000009000000000",
            INIT_28 => X"000000b200000000000000b100000000000000c3000000000000007500000000",
            INIT_29 => X"000000960000000000000053000000000000008a00000000000000b500000000",
            INIT_2A => X"00000086000000000000008500000000000000db00000000000000f500000000",
            INIT_2B => X"000000c200000000000000be00000000000000b0000000000000009500000000",
            INIT_2C => X"0000003d000000000000006e000000000000007d00000000000000a800000000",
            INIT_2D => X"0000003a00000000000000310000000000000022000000000000002300000000",
            INIT_2E => X"000000480000000000000045000000000000003a000000000000003d00000000",
            INIT_2F => X"00000037000000000000003b0000000000000045000000000000004e00000000",
            INIT_30 => X"000000b000000000000000ae00000000000000af000000000000004f00000000",
            INIT_31 => X"000000d3000000000000006d000000000000008c00000000000000b100000000",
            INIT_32 => X"0000007c00000000000000d000000000000000fc00000000000000fd00000000",
            INIT_33 => X"0000007a0000000000000074000000000000007c000000000000007200000000",
            INIT_34 => X"0000003c00000000000000440000000000000044000000000000006800000000",
            INIT_35 => X"0000003800000000000000330000000000000032000000000000003400000000",
            INIT_36 => X"00000033000000000000002b0000000000000033000000000000003800000000",
            INIT_37 => X"0000002a000000000000002b0000000000000030000000000000003b00000000",
            INIT_38 => X"000000a800000000000000900000000000000060000000000000002900000000",
            INIT_39 => X"000000f600000000000000a500000000000000a500000000000000b200000000",
            INIT_3A => X"0000003c000000000000006e00000000000000e300000000000000fd00000000",
            INIT_3B => X"0000003000000000000000310000000000000031000000000000003500000000",
            INIT_3C => X"0000002a000000000000002e000000000000002a000000000000002d00000000",
            INIT_3D => X"0000002b000000000000002e000000000000002e000000000000002600000000",
            INIT_3E => X"00000032000000000000002e000000000000002e000000000000002a00000000",
            INIT_3F => X"0000002d00000000000000330000000000000035000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000083000000000000003b000000000000001d000000000000001d00000000",
            INIT_41 => X"000000fe00000000000000c2000000000000008400000000000000a600000000",
            INIT_42 => X"00000032000000000000003d000000000000008d00000000000000f100000000",
            INIT_43 => X"0000003200000000000000310000000000000033000000000000003200000000",
            INIT_44 => X"000000220000000000000027000000000000002a000000000000002f00000000",
            INIT_45 => X"0000002a00000000000000260000000000000027000000000000002300000000",
            INIT_46 => X"0000003b000000000000003e0000000000000038000000000000002d00000000",
            INIT_47 => X"00000033000000000000002e0000000000000032000000000000003800000000",
            INIT_48 => X"000000490000000000000022000000000000001e000000000000003000000000",
            INIT_49 => X"0000010000000000000000d70000000000000080000000000000008000000000",
            INIT_4A => X"000000320000000000000036000000000000004200000000000000bb00000000",
            INIT_4B => X"0000002d000000000000002e0000000000000034000000000000003400000000",
            INIT_4C => X"0000002700000000000000240000000000000029000000000000002b00000000",
            INIT_4D => X"0000002e000000000000002b0000000000000028000000000000002800000000",
            INIT_4E => X"0000003b0000000000000040000000000000003e000000000000003b00000000",
            INIT_4F => X"0000005300000000000000460000000000000032000000000000003600000000",
            INIT_50 => X"00000029000000000000001f0000000000000023000000000000003400000000",
            INIT_51 => X"000000f000000000000000e00000000000000080000000000000004200000000",
            INIT_52 => X"000000380000000000000031000000000000003a000000000000007c00000000",
            INIT_53 => X"0000002f000000000000002c000000000000002c000000000000003600000000",
            INIT_54 => X"0000002c000000000000002b000000000000002b000000000000002e00000000",
            INIT_55 => X"0000003a0000000000000036000000000000002d000000000000002c00000000",
            INIT_56 => X"00000024000000000000002b000000000000002e000000000000003600000000",
            INIT_57 => X"0000004c00000000000000550000000000000049000000000000003300000000",
            INIT_58 => X"00000023000000000000001d0000000000000023000000000000003200000000",
            INIT_59 => X"000000d300000000000000ca000000000000004e000000000000002c00000000",
            INIT_5A => X"0000003000000000000000360000000000000041000000000000006100000000",
            INIT_5B => X"0000002d00000000000000280000000000000030000000000000003a00000000",
            INIT_5C => X"0000002e000000000000002f0000000000000030000000000000002f00000000",
            INIT_5D => X"0000003000000000000000270000000000000027000000000000003300000000",
            INIT_5E => X"00000028000000000000001c0000000000000027000000000000002f00000000",
            INIT_5F => X"00000033000000000000002e0000000000000043000000000000004300000000",
            INIT_60 => X"0000002100000000000000200000000000000023000000000000003200000000",
            INIT_61 => X"000000aa0000000000000068000000000000002e000000000000002900000000",
            INIT_62 => X"0000003500000000000000340000000000000036000000000000004000000000",
            INIT_63 => X"0000002d0000000000000036000000000000003a000000000000003d00000000",
            INIT_64 => X"00000031000000000000002e0000000000000029000000000000002a00000000",
            INIT_65 => X"000000270000000000000028000000000000002a000000000000002e00000000",
            INIT_66 => X"0000003f000000000000002c0000000000000028000000000000002500000000",
            INIT_67 => X"00000033000000000000000f000000000000001f000000000000002f00000000",
            INIT_68 => X"00000026000000000000001f000000000000002a000000000000004400000000",
            INIT_69 => X"00000047000000000000002a000000000000002b000000000000002500000000",
            INIT_6A => X"00000026000000000000001b000000000000001f000000000000003100000000",
            INIT_6B => X"00000035000000000000003a0000000000000038000000000000003100000000",
            INIT_6C => X"000000350000000000000039000000000000003c000000000000003800000000",
            INIT_6D => X"000000210000000000000027000000000000002d000000000000003200000000",
            INIT_6E => X"00000049000000000000004f000000000000003e000000000000002a00000000",
            INIT_6F => X"00000028000000000000000d0000000000000026000000000000003800000000",
            INIT_70 => X"0000002b00000000000000230000000000000031000000000000003d00000000",
            INIT_71 => X"00000028000000000000002c000000000000002a000000000000002700000000",
            INIT_72 => X"0000001e0000000000000017000000000000001b000000000000002a00000000",
            INIT_73 => X"0000002f0000000000000024000000000000001d000000000000001b00000000",
            INIT_74 => X"0000004b0000000000000042000000000000003e000000000000003800000000",
            INIT_75 => X"0000002b000000000000002b0000000000000031000000000000004500000000",
            INIT_76 => X"0000005d000000000000006d0000000000000055000000000000003c00000000",
            INIT_77 => X"00000014000000000000001d000000000000001a000000000000003c00000000",
            INIT_78 => X"0000002b000000000000002d0000000000000038000000000000003600000000",
            INIT_79 => X"0000002600000000000000280000000000000028000000000000002800000000",
            INIT_7A => X"0000001d0000000000000016000000000000001a000000000000002400000000",
            INIT_7B => X"000000120000000000000013000000000000001d000000000000001900000000",
            INIT_7C => X"0000004a000000000000003d000000000000002f000000000000002000000000",
            INIT_7D => X"0000002d00000000000000340000000000000035000000000000004200000000",
            INIT_7E => X"0000005900000000000000690000000000000059000000000000004300000000",
            INIT_7F => X"0000001500000000000000220000000000000018000000000000003000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE1;


    MEM_IFMAP_LAYER0_INSTANCE2 : if BRAM_NAME = "ifmap_layer0_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000760000000000000074000000000000006f000000000000007000000000",
            INIT_01 => X"000000710000000000000073000000000000006d000000000000007000000000",
            INIT_02 => X"0000006f00000000000000740000000000000071000000000000006f00000000",
            INIT_03 => X"0000007700000000000000750000000000000075000000000000006f00000000",
            INIT_04 => X"00000070000000000000006f0000000000000071000000000000007500000000",
            INIT_05 => X"0000006a000000000000006b000000000000006b000000000000006d00000000",
            INIT_06 => X"0000006100000000000000620000000000000065000000000000006b00000000",
            INIT_07 => X"00000055000000000000005b000000000000005f000000000000006100000000",
            INIT_08 => X"000000740000000000000072000000000000006e000000000000007000000000",
            INIT_09 => X"0000007200000000000000750000000000000071000000000000007000000000",
            INIT_0A => X"0000006e000000000000006f000000000000006e000000000000007400000000",
            INIT_0B => X"0000007300000000000000750000000000000077000000000000007100000000",
            INIT_0C => X"000000730000000000000070000000000000006f000000000000007300000000",
            INIT_0D => X"0000006400000000000000660000000000000068000000000000006e00000000",
            INIT_0E => X"0000006100000000000000660000000000000066000000000000006900000000",
            INIT_0F => X"00000058000000000000005b000000000000005f000000000000006200000000",
            INIT_10 => X"0000006f000000000000006f000000000000006d000000000000006e00000000",
            INIT_11 => X"0000007500000000000000750000000000000073000000000000006a00000000",
            INIT_12 => X"0000006d00000000000000720000000000000073000000000000007300000000",
            INIT_13 => X"0000007100000000000000720000000000000073000000000000006f00000000",
            INIT_14 => X"00000060000000000000006f0000000000000072000000000000007400000000",
            INIT_15 => X"00000055000000000000004d000000000000004e000000000000005a00000000",
            INIT_16 => X"0000006300000000000000670000000000000060000000000000005600000000",
            INIT_17 => X"00000059000000000000005f0000000000000062000000000000006300000000",
            INIT_18 => X"00000070000000000000006d000000000000006e000000000000006b00000000",
            INIT_19 => X"0000007700000000000000780000000000000075000000000000006e00000000",
            INIT_1A => X"00000092000000000000007b0000000000000075000000000000007300000000",
            INIT_1B => X"000000720000000000000073000000000000006f000000000000008200000000",
            INIT_1C => X"000000570000000000000050000000000000006f000000000000007000000000",
            INIT_1D => X"0000003f000000000000004b000000000000005a000000000000005a00000000",
            INIT_1E => X"000000620000000000000055000000000000003e000000000000004600000000",
            INIT_1F => X"0000005e00000000000000630000000000000065000000000000006600000000",
            INIT_20 => X"0000007200000000000000730000000000000072000000000000006b00000000",
            INIT_21 => X"0000007400000000000000780000000000000071000000000000007200000000",
            INIT_22 => X"000000d600000000000000800000000000000074000000000000007100000000",
            INIT_23 => X"0000006c000000000000006f0000000000000072000000000000009c00000000",
            INIT_24 => X"0000006700000000000000450000000000000035000000000000005000000000",
            INIT_25 => X"0000005e00000000000000660000000000000072000000000000006e00000000",
            INIT_26 => X"000000530000000000000049000000000000004e000000000000004800000000",
            INIT_27 => X"0000005d000000000000005e0000000000000065000000000000006000000000",
            INIT_28 => X"0000007000000000000000640000000000000068000000000000006d00000000",
            INIT_29 => X"0000007300000000000000740000000000000071000000000000007300000000",
            INIT_2A => X"0000008a00000000000000760000000000000074000000000000006f00000000",
            INIT_2B => X"00000032000000000000004b0000000000000066000000000000007a00000000",
            INIT_2C => X"0000007100000000000000530000000000000038000000000000003a00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007900000000",
            INIT_2E => X"0000003a000000000000003a000000000000005b000000000000006400000000",
            INIT_2F => X"0000005f00000000000000620000000000000069000000000000005400000000",
            INIT_30 => X"0000004a0000000000000025000000000000005f000000000000006400000000",
            INIT_31 => X"0000007600000000000000730000000000000076000000000000007500000000",
            INIT_32 => X"0000006b00000000000000780000000000000074000000000000007500000000",
            INIT_33 => X"000000430000000000000057000000000000006c000000000000006200000000",
            INIT_34 => X"000000820000000000000054000000000000004b000000000000005300000000",
            INIT_35 => X"0000006600000000000000630000000000000076000000000000008e00000000",
            INIT_36 => X"0000002f00000000000000470000000000000053000000000000006f00000000",
            INIT_37 => X"0000005d00000000000000630000000000000062000000000000003d00000000",
            INIT_38 => X"00000040000000000000002b0000000000000060000000000000007300000000",
            INIT_39 => X"0000007400000000000000720000000000000075000000000000006f00000000",
            INIT_3A => X"0000005e000000000000006d0000000000000071000000000000007700000000",
            INIT_3B => X"00000057000000000000006a0000000000000083000000000000006e00000000",
            INIT_3C => X"00000076000000000000004d0000000000000058000000000000005f00000000",
            INIT_3D => X"00000062000000000000005d000000000000007c000000000000009900000000",
            INIT_3E => X"00000035000000000000003c0000000000000051000000000000005d00000000",
            INIT_3F => X"0000006100000000000000670000000000000053000000000000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000079000000000000003a000000000000006900000000000000a100000000",
            INIT_41 => X"0000007a00000000000000750000000000000071000000000000007c00000000",
            INIT_42 => X"0000006900000000000000590000000000000087000000000000007900000000",
            INIT_43 => X"00000050000000000000006f000000000000008f000000000000008d00000000",
            INIT_44 => X"00000047000000000000004e0000000000000055000000000000005100000000",
            INIT_45 => X"0000004f00000000000000670000000000000087000000000000007d00000000",
            INIT_46 => X"0000003900000000000000490000000000000052000000000000004d00000000",
            INIT_47 => X"00000067000000000000006a000000000000003b000000000000002300000000",
            INIT_48 => X"0000009a0000000000000064000000000000008b00000000000000b000000000",
            INIT_49 => X"0000007600000000000000740000000000000074000000000000009500000000",
            INIT_4A => X"0000008300000000000000b400000000000000d600000000000000b400000000",
            INIT_4B => X"00000055000000000000006e0000000000000083000000000000009900000000",
            INIT_4C => X"000000440000000000000039000000000000004a000000000000005400000000",
            INIT_4D => X"00000062000000000000007c0000000000000085000000000000007d00000000",
            INIT_4E => X"0000004c00000000000000550000000000000055000000000000005100000000",
            INIT_4F => X"00000067000000000000004b000000000000001e000000000000003100000000",
            INIT_50 => X"000000a90000000000000097000000000000007400000000000000b700000000",
            INIT_51 => X"0000005900000000000000760000000000000070000000000000009c00000000",
            INIT_52 => X"0000008700000000000000bf00000000000000e000000000000000c500000000",
            INIT_53 => X"0000006f000000000000006c0000000000000089000000000000009f00000000",
            INIT_54 => X"00000055000000000000002c0000000000000050000000000000004c00000000",
            INIT_55 => X"000000640000000000000093000000000000009300000000000000a500000000",
            INIT_56 => X"0000004f00000000000000580000000000000066000000000000005300000000",
            INIT_57 => X"00000051000000000000002e0000000000000024000000000000003b00000000",
            INIT_58 => X"000000af0000000000000090000000000000006c00000000000000bf00000000",
            INIT_59 => X"0000005d000000000000007b000000000000007800000000000000a700000000",
            INIT_5A => X"0000008e00000000000000ab00000000000000b6000000000000005f00000000",
            INIT_5B => X"0000006b000000000000007700000000000000ab00000000000000a100000000",
            INIT_5C => X"0000007900000000000000260000000000000054000000000000006200000000",
            INIT_5D => X"00000059000000000000008b000000000000009800000000000000c900000000",
            INIT_5E => X"000000570000000000000068000000000000005d000000000000005000000000",
            INIT_5F => X"0000003800000000000000370000000000000035000000000000004b00000000",
            INIT_60 => X"000000b40000000000000086000000000000006000000000000000c200000000",
            INIT_61 => X"0000006d000000000000007b000000000000007b000000000000009c00000000",
            INIT_62 => X"000000720000000000000090000000000000009a000000000000004400000000",
            INIT_63 => X"00000071000000000000009500000000000000ca00000000000000a600000000",
            INIT_64 => X"0000009300000000000000320000000000000072000000000000007200000000",
            INIT_65 => X"000000580000000000000076000000000000009500000000000000bb00000000",
            INIT_66 => X"00000057000000000000005f0000000000000054000000000000005300000000",
            INIT_67 => X"00000037000000000000004a0000000000000049000000000000005700000000",
            INIT_68 => X"000000bc000000000000009a000000000000005f00000000000000c000000000",
            INIT_69 => X"00000074000000000000007c000000000000006a000000000000006e00000000",
            INIT_6A => X"00000095000000000000007d0000000000000084000000000000004800000000",
            INIT_6B => X"0000008300000000000000ac00000000000000d800000000000000ae00000000",
            INIT_6C => X"0000009800000000000000470000000000000072000000000000007500000000",
            INIT_6D => X"00000055000000000000006e000000000000009000000000000000b500000000",
            INIT_6E => X"0000006400000000000000500000000000000049000000000000005000000000",
            INIT_6F => X"0000004900000000000000590000000000000058000000000000006500000000",
            INIT_70 => X"000000ba00000000000000a7000000000000006b00000000000000c400000000",
            INIT_71 => X"0000007a00000000000000770000000000000059000000000000006d00000000",
            INIT_72 => X"000000b9000000000000007b000000000000006a000000000000004a00000000",
            INIT_73 => X"0000008f000000000000008c00000000000000a500000000000000b400000000",
            INIT_74 => X"0000009800000000000000470000000000000064000000000000008800000000",
            INIT_75 => X"0000006d0000000000000080000000000000008500000000000000af00000000",
            INIT_76 => X"0000006e0000000000000060000000000000005d000000000000005600000000",
            INIT_77 => X"0000005f00000000000000550000000000000060000000000000007400000000",
            INIT_78 => X"000000b200000000000000a7000000000000008100000000000000c500000000",
            INIT_79 => X"0000007d00000000000000780000000000000053000000000000008900000000",
            INIT_7A => X"000000dd00000000000000830000000000000078000000000000005e00000000",
            INIT_7B => X"000000790000000000000082000000000000008a00000000000000ec00000000",
            INIT_7C => X"0000008600000000000000580000000000000068000000000000007000000000",
            INIT_7D => X"00000055000000000000006c0000000000000093000000000000009f00000000",
            INIT_7E => X"0000006d00000000000000680000000000000058000000000000004800000000",
            INIT_7F => X"0000006800000000000000600000000000000056000000000000006e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE2;


    MEM_IFMAP_LAYER0_INSTANCE3 : if BRAM_NAME = "ifmap_layer0_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b600000000000000a4000000000000009200000000000000cb00000000",
            INIT_01 => X"0000007e000000000000007d000000000000005600000000000000aa00000000",
            INIT_02 => X"000000a3000000000000008f0000000000000050000000000000007900000000",
            INIT_03 => X"0000006a000000000000006a0000000000000084000000000000009800000000",
            INIT_04 => X"0000008f000000000000005a0000000000000065000000000000006500000000",
            INIT_05 => X"000000690000000000000082000000000000008d000000000000008a00000000",
            INIT_06 => X"0000005b000000000000005d000000000000004f000000000000004c00000000",
            INIT_07 => X"00000068000000000000006c0000000000000058000000000000005300000000",
            INIT_08 => X"000000b800000000000000a700000000000000a600000000000000d700000000",
            INIT_09 => X"000000950000000000000060000000000000006600000000000000b600000000",
            INIT_0A => X"000000690000000000000074000000000000005d000000000000008900000000",
            INIT_0B => X"0000006e000000000000005b0000000000000069000000000000006600000000",
            INIT_0C => X"0000006000000000000000800000000000000067000000000000005b00000000",
            INIT_0D => X"00000045000000000000007e0000000000000078000000000000003800000000",
            INIT_0E => X"0000005d00000000000000460000000000000038000000000000003800000000",
            INIT_0F => X"0000006e00000000000000740000000000000070000000000000005e00000000",
            INIT_10 => X"000000b500000000000000af00000000000000b800000000000000d300000000",
            INIT_11 => X"0000008b0000000000000058000000000000008300000000000000b800000000",
            INIT_12 => X"00000040000000000000005a0000000000000080000000000000009400000000",
            INIT_13 => X"0000008f0000000000000075000000000000006f000000000000007900000000",
            INIT_14 => X"00000075000000000000008b0000000000000060000000000000005c00000000",
            INIT_15 => X"0000003b00000000000000440000000000000063000000000000006d00000000",
            INIT_16 => X"000000690000000000000045000000000000003e000000000000002900000000",
            INIT_17 => X"0000006f00000000000000730000000000000078000000000000007700000000",
            INIT_18 => X"000000b300000000000000b000000000000000bd00000000000000c000000000",
            INIT_19 => X"00000079000000000000005a000000000000009500000000000000b600000000",
            INIT_1A => X"0000003b00000000000000860000000000000088000000000000007c00000000",
            INIT_1B => X"000000b000000000000000860000000000000061000000000000007600000000",
            INIT_1C => X"0000007c0000000000000077000000000000004b000000000000007600000000",
            INIT_1D => X"0000003300000000000000310000000000000056000000000000008100000000",
            INIT_1E => X"00000076000000000000005b000000000000005a000000000000003100000000",
            INIT_1F => X"0000006b000000000000006f0000000000000071000000000000007900000000",
            INIT_20 => X"000000ad00000000000000b200000000000000c1000000000000009c00000000",
            INIT_21 => X"000000870000000000000067000000000000009d00000000000000b500000000",
            INIT_22 => X"0000004d000000000000005a000000000000006900000000000000af00000000",
            INIT_23 => X"000000b600000000000000ad0000000000000076000000000000005a00000000",
            INIT_24 => X"0000004d000000000000004e0000000000000064000000000000009400000000",
            INIT_25 => X"00000021000000000000002e0000000000000034000000000000003d00000000",
            INIT_26 => X"0000007d00000000000000640000000000000047000000000000003900000000",
            INIT_27 => X"000000690000000000000071000000000000006d000000000000007b00000000",
            INIT_28 => X"000000a900000000000000b200000000000000c8000000000000007800000000",
            INIT_29 => X"000000990000000000000057000000000000009000000000000000b300000000",
            INIT_2A => X"0000008d000000000000008c00000000000000de00000000000000f700000000",
            INIT_2B => X"000000c000000000000000c400000000000000b6000000000000009c00000000",
            INIT_2C => X"0000003e000000000000006d000000000000008500000000000000ac00000000",
            INIT_2D => X"0000005100000000000000460000000000000036000000000000003100000000",
            INIT_2E => X"0000006500000000000000630000000000000054000000000000005500000000",
            INIT_2F => X"0000005a000000000000005c0000000000000060000000000000006800000000",
            INIT_30 => X"000000ac00000000000000b700000000000000c5000000000000006900000000",
            INIT_31 => X"000000d30000000000000070000000000000009200000000000000b100000000",
            INIT_32 => X"0000008f00000000000000e000000000000000fd00000000000000fc00000000",
            INIT_33 => X"000000850000000000000085000000000000008d000000000000008400000000",
            INIT_34 => X"000000520000000000000057000000000000005d000000000000007c00000000",
            INIT_35 => X"0000005d00000000000000550000000000000054000000000000005400000000",
            INIT_36 => X"000000680000000000000060000000000000005b000000000000005e00000000",
            INIT_37 => X"0000005f00000000000000610000000000000061000000000000006c00000000",
            INIT_38 => X"000000ae00000000000000a80000000000000089000000000000005900000000",
            INIT_39 => X"000000f500000000000000a600000000000000aa00000000000000b600000000",
            INIT_3A => X"00000058000000000000008800000000000000e700000000000000fb00000000",
            INIT_3B => X"00000048000000000000004b000000000000004c000000000000005000000000",
            INIT_3C => X"0000005200000000000000510000000000000051000000000000004f00000000",
            INIT_3D => X"000000570000000000000059000000000000005a000000000000005600000000",
            INIT_3E => X"00000060000000000000005e000000000000005d000000000000005900000000",
            INIT_3F => X"0000005a000000000000005f000000000000005e000000000000006000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009900000000000000660000000000000057000000000000005b00000000",
            INIT_41 => X"000000fa00000000000000bd000000000000008800000000000000b300000000",
            INIT_42 => X"00000054000000000000005e000000000000009f00000000000000f500000000",
            INIT_43 => X"0000005400000000000000530000000000000055000000000000005400000000",
            INIT_44 => X"0000004f00000000000000520000000000000054000000000000005600000000",
            INIT_45 => X"0000005900000000000000550000000000000056000000000000005300000000",
            INIT_46 => X"0000006500000000000000670000000000000067000000000000005c00000000",
            INIT_47 => X"00000067000000000000005e0000000000000063000000000000006600000000",
            INIT_48 => X"0000006a0000000000000055000000000000005e000000000000006f00000000",
            INIT_49 => X"000000fd00000000000000d50000000000000088000000000000009400000000",
            INIT_4A => X"00000058000000000000005b000000000000005d00000000000000c600000000",
            INIT_4B => X"000000520000000000000053000000000000005a000000000000005a00000000",
            INIT_4C => X"0000005300000000000000500000000000000051000000000000005200000000",
            INIT_4D => X"0000005f000000000000005c0000000000000059000000000000005600000000",
            INIT_4E => X"0000006c000000000000006d000000000000006e000000000000006c00000000",
            INIT_4F => X"00000089000000000000007b0000000000000069000000000000006c00000000",
            INIT_50 => X"0000005300000000000000560000000000000063000000000000007200000000",
            INIT_51 => X"000000f500000000000000e50000000000000091000000000000005f00000000",
            INIT_52 => X"0000005e0000000000000057000000000000005c000000000000008f00000000",
            INIT_53 => X"0000005300000000000000520000000000000052000000000000005c00000000",
            INIT_54 => X"0000005800000000000000560000000000000053000000000000005400000000",
            INIT_55 => X"0000006e000000000000006a0000000000000061000000000000005a00000000",
            INIT_56 => X"0000005b000000000000005f0000000000000061000000000000006900000000",
            INIT_57 => X"0000007d000000000000008a0000000000000082000000000000006c00000000",
            INIT_58 => X"0000005600000000000000590000000000000062000000000000006e00000000",
            INIT_59 => X"000000e400000000000000db000000000000006a000000000000005300000000",
            INIT_5A => X"00000057000000000000005e0000000000000068000000000000007e00000000",
            INIT_5B => X"0000005200000000000000500000000000000057000000000000006100000000",
            INIT_5C => X"0000005900000000000000590000000000000057000000000000005400000000",
            INIT_5D => X"00000066000000000000005d000000000000005c000000000000006100000000",
            INIT_5E => X"000000650000000000000055000000000000005d000000000000006500000000",
            INIT_5F => X"000000600000000000000062000000000000007e000000000000008100000000",
            INIT_60 => X"00000058000000000000005c0000000000000061000000000000006c00000000",
            INIT_61 => X"000000c500000000000000850000000000000054000000000000005800000000",
            INIT_62 => X"0000005f000000000000005e0000000000000061000000000000006400000000",
            INIT_63 => X"0000005300000000000000600000000000000064000000000000006700000000",
            INIT_64 => X"0000005c00000000000000580000000000000050000000000000004f00000000",
            INIT_65 => X"0000005c000000000000005d000000000000005f000000000000005c00000000",
            INIT_66 => X"0000007d0000000000000066000000000000005d000000000000005a00000000",
            INIT_67 => X"0000005d000000000000003c000000000000005a000000000000006e00000000",
            INIT_68 => X"0000005b00000000000000580000000000000064000000000000007c00000000",
            INIT_69 => X"0000006b000000000000004f0000000000000059000000000000005700000000",
            INIT_6A => X"000000520000000000000047000000000000004d000000000000005900000000",
            INIT_6B => X"0000005c00000000000000660000000000000064000000000000005d00000000",
            INIT_6C => X"0000006100000000000000630000000000000063000000000000005e00000000",
            INIT_6D => X"000000530000000000000058000000000000005e000000000000005f00000000",
            INIT_6E => X"0000008300000000000000840000000000000070000000000000005b00000000",
            INIT_6F => X"0000005500000000000000400000000000000061000000000000007400000000",
            INIT_70 => X"0000005b00000000000000550000000000000066000000000000007400000000",
            INIT_71 => X"000000510000000000000058000000000000005c000000000000005a00000000",
            INIT_72 => X"0000004a00000000000000430000000000000048000000000000005500000000",
            INIT_73 => X"0000005600000000000000500000000000000049000000000000004700000000",
            INIT_74 => X"00000077000000000000006d0000000000000065000000000000005f00000000",
            INIT_75 => X"000000580000000000000058000000000000005f000000000000007100000000",
            INIT_76 => X"00000091000000000000009c0000000000000082000000000000006900000000",
            INIT_77 => X"0000004000000000000000520000000000000052000000000000007300000000",
            INIT_78 => X"0000005600000000000000590000000000000069000000000000006b00000000",
            INIT_79 => X"000000510000000000000057000000000000005c000000000000005900000000",
            INIT_7A => X"0000004900000000000000420000000000000045000000000000004f00000000",
            INIT_7B => X"0000003a000000000000003f0000000000000049000000000000004500000000",
            INIT_7C => X"0000007700000000000000680000000000000057000000000000004600000000",
            INIT_7D => X"00000057000000000000005f0000000000000060000000000000006f00000000",
            INIT_7E => X"0000008700000000000000920000000000000083000000000000006d00000000",
            INIT_7F => X"000000430000000000000054000000000000004d000000000000006300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE3;


    MEM_IFMAP_LAYER0_INSTANCE4 : if BRAM_NAME = "ifmap_layer0_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000350000000000000033000000000000002f000000000000003100000000",
            INIT_01 => X"0000002d000000000000002f0000000000000029000000000000002e00000000",
            INIT_02 => X"0000003400000000000000290000000000000029000000000000002c00000000",
            INIT_03 => X"0000002c000000000000002d0000000000000029000000000000003100000000",
            INIT_04 => X"0000002b00000000000000270000000000000026000000000000002800000000",
            INIT_05 => X"0000002b000000000000002d000000000000002d000000000000002c00000000",
            INIT_06 => X"00000029000000000000002b0000000000000027000000000000002c00000000",
            INIT_07 => X"0000002100000000000000240000000000000024000000000000002600000000",
            INIT_08 => X"00000038000000000000002d0000000000000028000000000000003300000000",
            INIT_09 => X"0000002d000000000000002f000000000000002b000000000000003100000000",
            INIT_0A => X"0000003600000000000000290000000000000026000000000000002e00000000",
            INIT_0B => X"0000002100000000000000280000000000000029000000000000003400000000",
            INIT_0C => X"0000003200000000000000290000000000000021000000000000001e00000000",
            INIT_0D => X"0000003000000000000000340000000000000037000000000000003500000000",
            INIT_0E => X"00000026000000000000002d000000000000002e000000000000003200000000",
            INIT_0F => X"000000220000000000000020000000000000001f000000000000002200000000",
            INIT_10 => X"0000003000000000000000240000000000000021000000000000002f00000000",
            INIT_11 => X"0000002d000000000000002d000000000000002c000000000000002a00000000",
            INIT_12 => X"000000390000000000000030000000000000002b000000000000002b00000000",
            INIT_13 => X"0000002300000000000000250000000000000026000000000000003300000000",
            INIT_14 => X"000000310000000000000036000000000000002f000000000000002700000000",
            INIT_15 => X"00000032000000000000002f0000000000000032000000000000003400000000",
            INIT_16 => X"0000002700000000000000330000000000000037000000000000003000000000",
            INIT_17 => X"0000002100000000000000220000000000000022000000000000002300000000",
            INIT_18 => X"0000002c000000000000001f0000000000000020000000000000002800000000",
            INIT_19 => X"000000300000000000000030000000000000002e000000000000002b00000000",
            INIT_1A => X"0000005f0000000000000039000000000000002d000000000000002c00000000",
            INIT_1B => X"00000036000000000000002f0000000000000029000000000000004b00000000",
            INIT_1C => X"00000041000000000000002f0000000000000043000000000000003a00000000",
            INIT_1D => X"0000003200000000000000420000000000000054000000000000004c00000000",
            INIT_1E => X"0000002e000000000000002d0000000000000027000000000000003400000000",
            INIT_1F => X"0000002400000000000000270000000000000027000000000000002b00000000",
            INIT_20 => X"0000002f00000000000000310000000000000030000000000000002900000000",
            INIT_21 => X"0000002c000000000000002f0000000000000028000000000000002b00000000",
            INIT_22 => X"000000a4000000000000003b000000000000002a000000000000002900000000",
            INIT_23 => X"00000047000000000000003c0000000000000038000000000000006b00000000",
            INIT_24 => X"000000620000000000000038000000000000001f000000000000003200000000",
            INIT_25 => X"0000005d00000000000000690000000000000076000000000000006f00000000",
            INIT_26 => X"0000002d000000000000002f0000000000000046000000000000004300000000",
            INIT_27 => X"000000240000000000000024000000000000002e000000000000003000000000",
            INIT_28 => X"0000003500000000000000390000000000000040000000000000003600000000",
            INIT_29 => X"0000002900000000000000290000000000000027000000000000002c00000000",
            INIT_2A => X"00000055000000000000002a0000000000000027000000000000002500000000",
            INIT_2B => X"0000001f000000000000002b000000000000003a000000000000004e00000000",
            INIT_2C => X"0000006e000000000000004c000000000000002d000000000000002b00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007800000000",
            INIT_2E => X"00000025000000000000002f0000000000000056000000000000006100000000",
            INIT_2F => X"00000028000000000000002c000000000000003a000000000000003100000000",
            INIT_30 => X"0000001c00000000000000110000000000000050000000000000003900000000",
            INIT_31 => X"0000002b0000000000000028000000000000002b000000000000003000000000",
            INIT_32 => X"0000003400000000000000270000000000000025000000000000002a00000000",
            INIT_33 => X"000000390000000000000046000000000000004b000000000000003b00000000",
            INIT_34 => X"00000079000000000000004a0000000000000040000000000000004800000000",
            INIT_35 => X"0000005e000000000000005a000000000000006c000000000000008400000000",
            INIT_36 => X"000000270000000000000045000000000000004d000000000000006700000000",
            INIT_37 => X"000000270000000000000030000000000000003a000000000000002400000000",
            INIT_38 => X"000000290000000000000026000000000000005c000000000000005a00000000",
            INIT_39 => X"000000270000000000000024000000000000002a000000000000003800000000",
            INIT_3A => X"0000003100000000000000330000000000000033000000000000003100000000",
            INIT_3B => X"0000004f000000000000005d000000000000006b000000000000004d00000000",
            INIT_3C => X"0000006b00000000000000450000000000000052000000000000005800000000",
            INIT_3D => X"0000005800000000000000510000000000000070000000000000008c00000000",
            INIT_3E => X"00000031000000000000003a000000000000004a000000000000005400000000",
            INIT_3F => X"0000002700000000000000330000000000000032000000000000002000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000071000000000000003b0000000000000069000000000000009000000000",
            INIT_41 => X"000000320000000000000029000000000000002b000000000000005200000000",
            INIT_42 => X"0000004e000000000000003b000000000000005f000000000000004200000000",
            INIT_43 => X"0000004a00000000000000650000000000000080000000000000007900000000",
            INIT_44 => X"0000003d00000000000000490000000000000052000000000000004d00000000",
            INIT_45 => X"00000046000000000000005d000000000000007b000000000000007000000000",
            INIT_46 => X"000000350000000000000043000000000000004c000000000000004500000000",
            INIT_47 => X"0000002d000000000000003b0000000000000023000000000000001b00000000",
            INIT_48 => X"000000950000000000000069000000000000008f00000000000000a300000000",
            INIT_49 => X"0000003c000000000000002f0000000000000033000000000000007000000000",
            INIT_4A => X"0000007700000000000000a600000000000000c6000000000000009200000000",
            INIT_4B => X"0000004f000000000000006b000000000000007d000000000000009100000000",
            INIT_4C => X"0000003a00000000000000350000000000000047000000000000004f00000000",
            INIT_4D => X"000000590000000000000072000000000000007a000000000000007000000000",
            INIT_4E => X"00000047000000000000004e000000000000004e000000000000004a00000000",
            INIT_4F => X"00000039000000000000002c000000000000000f000000000000002b00000000",
            INIT_50 => X"000000a8000000000000009e000000000000007a00000000000000af00000000",
            INIT_51 => X"0000002f00000000000000330000000000000032000000000000007a00000000",
            INIT_52 => X"0000008300000000000000bc00000000000000e200000000000000b300000000",
            INIT_53 => X"0000006800000000000000680000000000000084000000000000009b00000000",
            INIT_54 => X"0000004d0000000000000028000000000000004d000000000000004500000000",
            INIT_55 => X"0000005c000000000000008a0000000000000089000000000000009a00000000",
            INIT_56 => X"00000049000000000000004f0000000000000060000000000000004d00000000",
            INIT_57 => X"0000002e000000000000001f0000000000000021000000000000003b00000000",
            INIT_58 => X"000000b20000000000000099000000000000007400000000000000bd00000000",
            INIT_59 => X"0000002c0000000000000037000000000000003b000000000000008800000000",
            INIT_5A => X"0000008500000000000000a400000000000000bc000000000000005000000000",
            INIT_5B => X"0000005f000000000000006a000000000000009f000000000000009700000000",
            INIT_5C => X"000000710000000000000022000000000000004f000000000000005900000000",
            INIT_5D => X"000000520000000000000082000000000000008e00000000000000c000000000",
            INIT_5E => X"00000051000000000000005e0000000000000058000000000000004b00000000",
            INIT_5F => X"0000001a00000000000000300000000000000037000000000000004e00000000",
            INIT_60 => X"000000b90000000000000090000000000000006900000000000000c200000000",
            INIT_61 => X"0000002f00000000000000350000000000000044000000000000008500000000",
            INIT_62 => X"0000005e000000000000007e0000000000000098000000000000002c00000000",
            INIT_63 => X"00000062000000000000008100000000000000b7000000000000009400000000",
            INIT_64 => X"0000008c000000000000002f000000000000006d000000000000006900000000",
            INIT_65 => X"00000053000000000000006f000000000000008c00000000000000b200000000",
            INIT_66 => X"0000005100000000000000550000000000000050000000000000004f00000000",
            INIT_67 => X"0000001800000000000000400000000000000049000000000000005900000000",
            INIT_68 => X"000000c000000000000000a3000000000000006700000000000000c100000000",
            INIT_69 => X"00000032000000000000003a0000000000000042000000000000006200000000",
            INIT_6A => X"0000007f00000000000000670000000000000078000000000000002700000000",
            INIT_6B => X"00000075000000000000009d00000000000000c8000000000000009b00000000",
            INIT_6C => X"000000930000000000000044000000000000006d000000000000006b00000000",
            INIT_6D => X"000000500000000000000068000000000000008800000000000000ae00000000",
            INIT_6E => X"0000005e00000000000000480000000000000046000000000000004c00000000",
            INIT_6F => X"0000002200000000000000450000000000000051000000000000006300000000",
            INIT_70 => X"000000bc00000000000000ac000000000000007000000000000000c400000000",
            INIT_71 => X"00000037000000000000003e0000000000000043000000000000006d00000000",
            INIT_72 => X"000000a900000000000000670000000000000058000000000000002200000000",
            INIT_73 => X"00000086000000000000008c000000000000009f00000000000000a900000000",
            INIT_74 => X"000000950000000000000046000000000000005f000000000000007d00000000",
            INIT_75 => X"00000069000000000000007a000000000000007f00000000000000aa00000000",
            INIT_76 => X"00000068000000000000005a000000000000005b000000000000005300000000",
            INIT_77 => X"0000002f00000000000000350000000000000050000000000000006f00000000",
            INIT_78 => X"000000b500000000000000ae000000000000008800000000000000c500000000",
            INIT_79 => X"0000004d0000000000000058000000000000004d000000000000008e00000000",
            INIT_7A => X"000000d30000000000000074000000000000005d000000000000003400000000",
            INIT_7B => X"000000700000000000000082000000000000008900000000000000e600000000",
            INIT_7C => X"00000076000000000000004b000000000000005f000000000000006500000000",
            INIT_7D => X"000000500000000000000065000000000000008a000000000000009200000000",
            INIT_7E => X"0000006300000000000000630000000000000057000000000000004400000000",
            INIT_7F => X"0000003000000000000000300000000000000036000000000000005d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE4;


    MEM_IFMAP_LAYER0_INSTANCE5 : if BRAM_NAME = "ifmap_layer0_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bc00000000000000b200000000000000a000000000000000cc00000000",
            INIT_01 => X"00000071000000000000007e000000000000005a00000000000000ac00000000",
            INIT_02 => X"0000009b00000000000000850000000000000025000000000000005200000000",
            INIT_03 => X"0000005a00000000000000580000000000000075000000000000008d00000000",
            INIT_04 => X"00000068000000000000003a0000000000000057000000000000005c00000000",
            INIT_05 => X"000000610000000000000076000000000000007e000000000000006d00000000",
            INIT_06 => X"00000052000000000000005e000000000000004d000000000000004800000000",
            INIT_07 => X"0000002e0000000000000037000000000000002d000000000000003700000000",
            INIT_08 => X"000000c200000000000000b800000000000000b400000000000000d700000000",
            INIT_09 => X"000000910000000000000066000000000000006900000000000000ba00000000",
            INIT_0A => X"0000005f0000000000000069000000000000003d000000000000006f00000000",
            INIT_0B => X"0000006200000000000000490000000000000059000000000000005900000000",
            INIT_0C => X"000000400000000000000066000000000000005f000000000000005800000000",
            INIT_0D => X"0000003d00000000000000730000000000000069000000000000002000000000",
            INIT_0E => X"0000004e00000000000000410000000000000035000000000000003300000000",
            INIT_0F => X"0000003600000000000000400000000000000044000000000000004000000000",
            INIT_10 => X"000000c100000000000000bd00000000000000c000000000000000cd00000000",
            INIT_11 => X"0000008f0000000000000060000000000000008500000000000000bc00000000",
            INIT_12 => X"000000370000000000000050000000000000006f000000000000008d00000000",
            INIT_13 => X"0000008500000000000000640000000000000060000000000000006c00000000",
            INIT_14 => X"0000005d0000000000000078000000000000005d000000000000005d00000000",
            INIT_15 => X"00000034000000000000003a0000000000000056000000000000005c00000000",
            INIT_16 => X"0000003b0000000000000028000000000000003c000000000000002700000000",
            INIT_17 => X"0000002e000000000000002d0000000000000036000000000000003e00000000",
            INIT_18 => X"000000b900000000000000b500000000000000bb00000000000000b400000000",
            INIT_19 => X"000000840000000000000063000000000000009800000000000000b800000000",
            INIT_1A => X"00000033000000000000007e0000000000000087000000000000008200000000",
            INIT_1B => X"000000a8000000000000007b0000000000000056000000000000006c00000000",
            INIT_1C => X"0000006900000000000000670000000000000049000000000000007600000000",
            INIT_1D => X"00000032000000000000002c000000000000004e000000000000007600000000",
            INIT_1E => X"00000044000000000000003c000000000000005d000000000000003400000000",
            INIT_1F => X"0000002e00000000000000320000000000000034000000000000004000000000",
            INIT_20 => X"000000ac00000000000000af00000000000000bb000000000000009200000000",
            INIT_21 => X"00000092000000000000006f00000000000000a000000000000000b400000000",
            INIT_22 => X"000000490000000000000057000000000000006f00000000000000b900000000",
            INIT_23 => X"000000b100000000000000ad0000000000000074000000000000005600000000",
            INIT_24 => X"0000003f00000000000000420000000000000065000000000000009400000000",
            INIT_25 => X"0000002900000000000000330000000000000036000000000000003900000000",
            INIT_26 => X"00000052000000000000004b0000000000000053000000000000004500000000",
            INIT_27 => X"0000003f0000000000000045000000000000003d000000000000004c00000000",
            INIT_28 => X"000000a800000000000000b000000000000000c8000000000000007c00000000",
            INIT_29 => X"0000009f000000000000005b000000000000009300000000000000b300000000",
            INIT_2A => X"00000093000000000000009000000000000000e100000000000000fa00000000",
            INIT_2B => X"000000c500000000000000d000000000000000c000000000000000a400000000",
            INIT_2C => X"0000003e000000000000006d000000000000008f00000000000000b500000000",
            INIT_2D => X"0000006600000000000000570000000000000044000000000000003a00000000",
            INIT_2E => X"00000077000000000000007a000000000000006f000000000000006e00000000",
            INIT_2F => X"0000007300000000000000700000000000000070000000000000007800000000",
            INIT_30 => X"000000b100000000000000c000000000000000d5000000000000008500000000",
            INIT_31 => X"000000d10000000000000071000000000000009600000000000000b600000000",
            INIT_32 => X"0000009d00000000000000e800000000000000fc00000000000000f700000000",
            INIT_33 => X"00000098000000000000009c00000000000000a2000000000000009500000000",
            INIT_34 => X"0000006500000000000000680000000000000077000000000000009400000000",
            INIT_35 => X"0000007d0000000000000073000000000000006e000000000000006f00000000",
            INIT_36 => X"0000008d00000000000000870000000000000082000000000000008300000000",
            INIT_37 => X"0000008400000000000000890000000000000084000000000000008e00000000",
            INIT_38 => X"000000bc00000000000000bc00000000000000a8000000000000008700000000",
            INIT_39 => X"000000ed00000000000000a400000000000000ae00000000000000c000000000",
            INIT_3A => X"0000006f000000000000009900000000000000e400000000000000f100000000",
            INIT_3B => X"00000065000000000000006b0000000000000069000000000000006900000000",
            INIT_3C => X"0000007400000000000000710000000000000078000000000000007300000000",
            INIT_3D => X"00000080000000000000007e000000000000007d000000000000007d00000000",
            INIT_3E => X"000000890000000000000089000000000000008b000000000000008400000000",
            INIT_3F => X"00000085000000000000008b0000000000000086000000000000008700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b000000000000000860000000000000082000000000000008d00000000",
            INIT_41 => X"000000f200000000000000b5000000000000008900000000000000bf00000000",
            INIT_42 => X"00000076000000000000007f00000000000000af00000000000000f500000000",
            INIT_43 => X"0000007400000000000000780000000000000079000000000000007700000000",
            INIT_44 => X"0000007100000000000000730000000000000075000000000000007500000000",
            INIT_45 => X"00000082000000000000007d000000000000007d000000000000007800000000",
            INIT_46 => X"0000008e000000000000008e0000000000000091000000000000008600000000",
            INIT_47 => X"00000095000000000000008c0000000000000090000000000000009200000000",
            INIT_48 => X"00000088000000000000007c000000000000008c00000000000000a200000000",
            INIT_49 => X"000000f900000000000000d1000000000000008f00000000000000a700000000",
            INIT_4A => X"0000007d0000000000000080000000000000007600000000000000cd00000000",
            INIT_4B => X"000000730000000000000079000000000000007f000000000000007f00000000",
            INIT_4C => X"0000007500000000000000710000000000000070000000000000007100000000",
            INIT_4D => X"0000008a00000000000000860000000000000083000000000000007b00000000",
            INIT_4E => X"0000009500000000000000930000000000000098000000000000009600000000",
            INIT_4F => X"000000b600000000000000a70000000000000098000000000000009a00000000",
            INIT_50 => X"0000007a0000000000000082000000000000009300000000000000a500000000",
            INIT_51 => X"000000f700000000000000ea00000000000000a4000000000000007e00000000",
            INIT_52 => X"00000083000000000000007b0000000000000072000000000000009900000000",
            INIT_53 => X"0000007700000000000000770000000000000077000000000000008100000000",
            INIT_54 => X"0000007f000000000000007b0000000000000077000000000000007700000000",
            INIT_55 => X"0000009a0000000000000096000000000000008d000000000000008300000000",
            INIT_56 => X"0000008a000000000000008c000000000000008d000000000000009600000000",
            INIT_57 => X"000000a900000000000000b600000000000000b2000000000000009e00000000",
            INIT_58 => X"00000085000000000000008a000000000000009500000000000000a200000000",
            INIT_59 => X"000000ea00000000000000e9000000000000008a000000000000007e00000000",
            INIT_5A => X"0000007c0000000000000081000000000000007e000000000000008c00000000",
            INIT_5B => X"000000770000000000000074000000000000007b000000000000008500000000",
            INIT_5C => X"000000840000000000000082000000000000007e000000000000007a00000000",
            INIT_5D => X"00000094000000000000008b000000000000008a000000000000008c00000000",
            INIT_5E => X"000000990000000000000085000000000000008b000000000000009300000000",
            INIT_5F => X"0000008b000000000000008e00000000000000b000000000000000b600000000",
            INIT_60 => X"0000008d000000000000008f000000000000009300000000000000a100000000",
            INIT_61 => X"000000d3000000000000009f000000000000007d000000000000008a00000000",
            INIT_62 => X"0000008200000000000000800000000000000079000000000000007700000000",
            INIT_63 => X"0000007800000000000000830000000000000087000000000000008b00000000",
            INIT_64 => X"0000008700000000000000820000000000000078000000000000007600000000",
            INIT_65 => X"00000088000000000000008a000000000000008b000000000000008800000000",
            INIT_66 => X"000000b20000000000000097000000000000008a000000000000008700000000",
            INIT_67 => X"000000880000000000000067000000000000008c00000000000000a400000000",
            INIT_68 => X"000000920000000000000089000000000000009400000000000000b100000000",
            INIT_69 => X"0000008500000000000000710000000000000084000000000000008b00000000",
            INIT_6A => X"0000007500000000000000690000000000000069000000000000007200000000",
            INIT_6B => X"0000008000000000000000890000000000000087000000000000008000000000",
            INIT_6C => X"0000008a000000000000008b0000000000000089000000000000008300000000",
            INIT_6D => X"0000007d00000000000000830000000000000088000000000000008900000000",
            INIT_6E => X"000000b500000000000000b3000000000000009a000000000000008500000000",
            INIT_6F => X"0000007f000000000000006c000000000000009200000000000000a800000000",
            INIT_70 => X"0000008f0000000000000084000000000000009400000000000000a800000000",
            INIT_71 => X"00000070000000000000007d0000000000000086000000000000008b00000000",
            INIT_72 => X"0000006d00000000000000660000000000000068000000000000007300000000",
            INIT_73 => X"000000780000000000000073000000000000006c000000000000006a00000000",
            INIT_74 => X"0000009c00000000000000900000000000000087000000000000008000000000",
            INIT_75 => X"0000007f000000000000007f0000000000000086000000000000009800000000",
            INIT_76 => X"000000be00000000000000c500000000000000aa000000000000009000000000",
            INIT_77 => X"0000006b000000000000007e000000000000008200000000000000a400000000",
            INIT_78 => X"000000860000000000000084000000000000009500000000000000a000000000",
            INIT_79 => X"00000073000000000000007b0000000000000084000000000000008600000000",
            INIT_7A => X"0000006c00000000000000650000000000000069000000000000007200000000",
            INIT_7B => X"000000590000000000000062000000000000006c000000000000006800000000",
            INIT_7C => X"0000009800000000000000890000000000000076000000000000006400000000",
            INIT_7D => X"0000007b00000000000000820000000000000083000000000000009100000000",
            INIT_7E => X"000000af00000000000000b600000000000000a7000000000000009100000000",
            INIT_7F => X"0000006e0000000000000081000000000000007c000000000000009100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE5;


    MEM_IFMAP_LAYER1_INSTANCE0 : if BRAM_NAME = "ifmap_layer1_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000200000000000000000000000000000000000000000000000500000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000005400000000",
            INIT_06 => X"0000000200000000000000000000000000000002000000000000001b00000000",
            INIT_07 => X"0000000400000000000000000000000000000000000000000000000500000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000004a00000000000000070000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000750000000000000000000000000000001c00000000",
            INIT_0C => X"0000000d000000000000000c0000000000000001000000000000000900000000",
            INIT_0D => X"0000000000000000000000310000000000000000000000000000000000000000",
            INIT_0E => X"0000003600000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000002800000000000000000000000000000054000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000003400000000",
            INIT_11 => X"0000000000000000000000000000000000000058000000000000000000000000",
            INIT_12 => X"0000000000000000000000060000000000000000000000000000000a00000000",
            INIT_13 => X"0000004200000000000000000000000000000000000000000000001f00000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"000000070000000000000000000000000000000000000000000000d900000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000004d00000000000000440000000000000000000000000000000000000000",
            INIT_18 => X"000000a800000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000001b00000000000000040000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000510000000000000016000000000000000000000000",
            INIT_1C => X"0000000000000000000000620000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_1E => X"0000003800000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000120000000000000000000000000000001700000000",
            INIT_21 => X"000000000000000000000012000000000000001d000000000000000600000000",
            INIT_22 => X"0000000000000000000000470000000000000000000000000000000000000000",
            INIT_23 => X"00000000000000000000000e000000000000001a000000000000000000000000",
            INIT_24 => X"0000003400000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000610000000000000000000000000000003700000000",
            INIT_26 => X"00000000000000000000000000000000000000cb000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_28 => X"0000000500000000000000100000000000000024000000000000001700000000",
            INIT_29 => X"00000000000000000000000e000000000000001d000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000009200000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_2D => X"000000000000000000000038000000000000001f000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000d00000000000000090000000000000004000000000000000000000000",
            INIT_30 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_31 => X"000000000000000000000000000000000000004f000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000002900000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000500000000000000080000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000380000000000000000000000000000000000000000",
            INIT_38 => X"000000ab00000000000000ab00000000000000a4000000000000000000000000",
            INIT_39 => X"000000ae00000000000000ac00000000000000a800000000000000ac00000000",
            INIT_3A => X"00000083000000000000009500000000000000a300000000000000ab00000000",
            INIT_3B => X"0000007a000000000000008a0000000000000093000000000000008b00000000",
            INIT_3C => X"000000af00000000000000b000000000000000ab00000000000000a400000000",
            INIT_3D => X"0000009e00000000000000b3000000000000011100000000000000b700000000",
            INIT_3E => X"0000007400000000000000940000000000000095000000000000007000000000",
            INIT_3F => X"0000007800000000000000860000000000000084000000000000006f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ae00000000000000ac00000000000000ad000000000000009a00000000",
            INIT_41 => X"00000054000000000000005e000000000000008e00000000000000ee00000000",
            INIT_42 => X"0000007400000000000000ae00000000000000cd00000000000000e400000000",
            INIT_43 => X"000000aa000000000000006b0000000000000093000000000000005300000000",
            INIT_44 => X"000000b500000000000000ae00000000000000b900000000000000b400000000",
            INIT_45 => X"000000df000000000000007c000000000000007a00000000000000cc00000000",
            INIT_46 => X"000000280000000000000067000000000000009200000000000000d100000000",
            INIT_47 => X"000000bf000000000000013100000000000000e0000000000000008500000000",
            INIT_48 => X"000000f20000000000000123000000000000017d00000000000000fc00000000",
            INIT_49 => X"0000010800000000000000bf000000000000005c000000000000008800000000",
            INIT_4A => X"00000039000000000000004c0000000000000089000000000000008f00000000",
            INIT_4B => X"0000009500000000000000d0000000000000015f00000000000000f400000000",
            INIT_4C => X"000000bc000000000000012e000000000000011f000000000000015c00000000",
            INIT_4D => X"0000008c000000000000011d000000000000012b000000000000006600000000",
            INIT_4E => X"0000010000000000000000480000000000000080000000000000009b00000000",
            INIT_4F => X"000000ee000000000000008000000000000000bb000000000000014400000000",
            INIT_50 => X"0000009100000000000000f70000000000000167000000000000014100000000",
            INIT_51 => X"0000008c00000000000000920000000000000100000000000000015600000000",
            INIT_52 => X"000001610000000000000134000000000000008500000000000000ae00000000",
            INIT_53 => X"0000018300000000000000cd00000000000000be00000000000000c400000000",
            INIT_54 => X"00000123000000000000009200000000000000d8000000000000010f00000000",
            INIT_55 => X"000000ad0000000000000096000000000000009000000000000000f800000000",
            INIT_56 => X"000000c1000000000000018a000000000000016d000000000000009300000000",
            INIT_57 => X"000000bf00000000000000d200000000000000b4000000000000010b00000000",
            INIT_58 => X"000000ad00000000000000c700000000000000c900000000000000b800000000",
            INIT_59 => X"000000ad000000000000009e0000000000000059000000000000005600000000",
            INIT_5A => X"0000012800000000000000ef0000000000000184000000000000018200000000",
            INIT_5B => X"0000012b00000000000000f9000000000000009100000000000000cf00000000",
            INIT_5C => X"000000290000000000000057000000000000009c00000000000000b100000000",
            INIT_5D => X"0000018f00000000000000b300000000000000ce000000000000007d00000000",
            INIT_5E => X"0000019500000000000001b000000000000000fa000000000000017a00000000",
            INIT_5F => X"000000ba000000000000014c000000000000014700000000000000fd00000000",
            INIT_60 => X"000000a7000000000000007e0000000000000061000000000000007000000000",
            INIT_61 => X"00000175000000000000012500000000000000a900000000000000cd00000000",
            INIT_62 => X"000000ae00000000000001770000000000000225000000000000014800000000",
            INIT_63 => X"0000008b000000000000008d00000000000000a900000000000000b200000000",
            INIT_64 => X"000000c900000000000000bb00000000000000ab000000000000009c00000000",
            INIT_65 => X"0000017900000000000000fc00000000000000b600000000000000b900000000",
            INIT_66 => X"0000009b00000000000000a600000000000000ba00000000000001e100000000",
            INIT_67 => X"000000b5000000000000009a0000000000000093000000000000009600000000",
            INIT_68 => X"000000f600000000000000cd00000000000000ce00000000000000c900000000",
            INIT_69 => X"0000016b000000000000013400000000000000ad00000000000000b900000000",
            INIT_6A => X"0000009700000000000000a800000000000000b900000000000000a500000000",
            INIT_6B => X"000000c100000000000000b900000000000000af000000000000009d00000000",
            INIT_6C => X"000000bd00000000000000d200000000000000e000000000000000b900000000",
            INIT_6D => X"0000008100000000000000ce00000000000000b200000000000000b100000000",
            INIT_6E => X"000000bc00000000000000a800000000000000a3000000000000009200000000",
            INIT_6F => X"0000010300000000000000b200000000000000b000000000000000cf00000000",
            INIT_70 => X"000000000000000000000000000000000000009c000000000000010e00000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000033000000000000000000000000",
            INIT_7A => X"00000000000000000000000a0000000000000023000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000090000000000000000000000000000004700000000",
            INIT_7F => X"0000001e00000000000000000000000000000013000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE0;


    MEM_IFMAP_LAYER1_INSTANCE1 : if BRAM_NAME = "ifmap_layer1_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000050000000000000012000000000000000000000000",
            INIT_01 => X"0000002700000000000000000000000000000000000000000000000600000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_03 => X"0000000000000000000000470000000000000011000000000000000000000000",
            INIT_04 => X"0000000a000000000000003a000000000000009c000000000000000400000000",
            INIT_05 => X"0000001200000000000000620000000000000000000000000000000000000000",
            INIT_06 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_07 => X"00000000000000000000000c000000000000002c000000000000000800000000",
            INIT_08 => X"00000000000000000000003f0000000000000038000000000000004800000000",
            INIT_09 => X"0000000000000000000000050000000000000073000000000000000000000000",
            INIT_0A => X"0000001f00000000000000000000000000000004000000000000000000000000",
            INIT_0B => X"0000001000000000000000000000000000000000000000000000002a00000000",
            INIT_0C => X"0000000000000000000000260000000000000018000000000000007a00000000",
            INIT_0D => X"000000110000000000000000000000000000000f000000000000005700000000",
            INIT_0E => X"0000005900000000000000300000000000000000000000000000001700000000",
            INIT_0F => X"000000390000000000000000000000000000002b000000000000000000000000",
            INIT_10 => X"00000000000000000000000e0000000000000000000000000000000700000000",
            INIT_11 => X"00000004000000000000000c0000000000000000000000000000003400000000",
            INIT_12 => X"0000000000000000000000560000000000000052000000000000000000000000",
            INIT_13 => X"0000001c00000000000000000000000000000009000000000000004200000000",
            INIT_14 => X"0000000000000000000000190000000000000008000000000000000600000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"000000800000000000000000000000000000004d000000000000007500000000",
            INIT_17 => X"0000004e00000000000000500000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000008d0000000000000001000000000000001a000000000000000900000000",
            INIT_1A => X"0000005000000000000000940000000000000022000000000000007200000000",
            INIT_1B => X"000000150000000000000038000000000000003b000000000000002900000000",
            INIT_1C => X"0000001e000000000000001d0000000000000013000000000000001000000000",
            INIT_1D => X"00000073000000000000000e000000000000001a000000000000002000000000",
            INIT_1E => X"000000140000000000000009000000000000007a000000000000006d00000000",
            INIT_1F => X"0000000e000000000000000b0000000000000010000000000000001200000000",
            INIT_20 => X"000000290000000000000026000000000000001e000000000000001600000000",
            INIT_21 => X"0000009e000000000000001b0000000000000014000000000000002800000000",
            INIT_22 => X"00000009000000000000001c0000000000000007000000000000004d00000000",
            INIT_23 => X"00000022000000000000001c0000000000000017000000000000001200000000",
            INIT_24 => X"0000003b0000000000000034000000000000001c000000000000002f00000000",
            INIT_25 => X"0000004300000000000000270000000000000023000000000000001100000000",
            INIT_26 => X"0000001500000000000000280000000000000029000000000000000d00000000",
            INIT_27 => X"0000001b00000000000000150000000000000018000000000000001800000000",
            INIT_28 => X"0000000000000000000000000000000000000025000000000000003000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000d00000000000000060000000000000009000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000004000000000000001700000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000300000000000000060000000000000003000000000000000b00000000",
            INIT_37 => X"000000240000000000000000000000000000000a000000000000001100000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"00000008000000000000000e0000000000000005000000000000000000000000",
            INIT_3A => X"0000000a000000000000000a0000000000000006000000000000001500000000",
            INIT_3B => X"00000005000000000000002d0000000000000000000000000000000f00000000",
            INIT_3C => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000400000000000000060000000000000008000000000000000000000000",
            INIT_3E => X"00000014000000000000000b0000000000000017000000000000000600000000",
            INIT_3F => X"000000000000000000000000000000000000003a000000000000001500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"000000140000000000000000000000000000000b000000000000000e00000000",
            INIT_42 => X"000000080000000000000011000000000000000f000000000000001300000000",
            INIT_43 => X"000000000000000000000011000000000000001c000000000000002d00000000",
            INIT_44 => X"00000004000000000000000c0000000000000000000000000000000000000000",
            INIT_45 => X"0000001000000000000000060000000000000000000000000000000d00000000",
            INIT_46 => X"0000002600000000000000000000000000000003000000000000001100000000",
            INIT_47 => X"0000000000000000000000090000000000000025000000000000001d00000000",
            INIT_48 => X"0000000e00000000000000000000000000000008000000000000000700000000",
            INIT_49 => X"0000000b00000000000000110000000000000000000000000000000000000000",
            INIT_4A => X"0000001800000000000000150000000000000000000000000000000000000000",
            INIT_4B => X"0000001100000000000000140000000000000018000000000000001f00000000",
            INIT_4C => X"0000000100000000000000080000000000000005000000000000001800000000",
            INIT_4D => X"000000000000000000000005000000000000001c000000000000000d00000000",
            INIT_4E => X"0000001c00000000000000180000000000000013000000000000000000000000",
            INIT_4F => X"00000010000000000000001b000000000000001e000000000000001d00000000",
            INIT_50 => X"0000003300000000000000230000000000000028000000000000001f00000000",
            INIT_51 => X"0000002600000000000000240000000000000030000000000000003500000000",
            INIT_52 => X"00000000000000000000002a0000000000000031000000000000003400000000",
            INIT_53 => X"00000043000000000000003f000000000000004d000000000000000b00000000",
            INIT_54 => X"0000004d00000000000000490000000000000045000000000000004800000000",
            INIT_55 => X"000000570000000000000053000000000000004e000000000000005300000000",
            INIT_56 => X"000000500000000000000000000000000000003b000000000000003900000000",
            INIT_57 => X"0000004900000000000000480000000000000049000000000000004c00000000",
            INIT_58 => X"0000004f00000000000000540000000000000053000000000000004d00000000",
            INIT_59 => X"0000005800000000000000640000000000000060000000000000005700000000",
            INIT_5A => X"0000004b0000000000000046000000000000001d000000000000003800000000",
            INIT_5B => X"00000051000000000000004e000000000000004a000000000000004c00000000",
            INIT_5C => X"0000005f000000000000005d0000000000000057000000000000005400000000",
            INIT_5D => X"0000004b000000000000005e0000000000000061000000000000005000000000",
            INIT_5E => X"0000004a00000000000000480000000000000044000000000000003e00000000",
            INIT_5F => X"00000051000000000000004f000000000000004a000000000000004e00000000",
            INIT_60 => X"000000610000000000000055000000000000005a000000000000005800000000",
            INIT_61 => X"0000008600000000000000850000000000000086000000000000008100000000",
            INIT_62 => X"00000092000000000000008b0000000000000080000000000000008400000000",
            INIT_63 => X"0000006900000000000000640000000000000072000000000000008600000000",
            INIT_64 => X"0000008000000000000000720000000000000075000000000000006c00000000",
            INIT_65 => X"000000880000000000000088000000000000008d000000000000008b00000000",
            INIT_66 => X"0000005900000000000000780000000000000078000000000000007800000000",
            INIT_67 => X"00000046000000000000002c000000000000001c000000000000003600000000",
            INIT_68 => X"000000710000000000000062000000000000006e000000000000005f00000000",
            INIT_69 => X"00000094000000000000008c000000000000008a000000000000008800000000",
            INIT_6A => X"0000003600000000000000270000000000000035000000000000004100000000",
            INIT_6B => X"000000390000000000000019000000000000001e000000000000002000000000",
            INIT_6C => X"0000007c00000000000000490000000000000015000000000000006100000000",
            INIT_6D => X"0000003900000000000000570000000000000072000000000000008c00000000",
            INIT_6E => X"0000002000000000000000480000000000000018000000000000001f00000000",
            INIT_6F => X"0000005c0000000000000011000000000000000e000000000000002900000000",
            INIT_70 => X"000000850000000000000066000000000000003f000000000000000000000000",
            INIT_71 => X"0000001a000000000000002f0000000000000049000000000000005100000000",
            INIT_72 => X"00000019000000000000002e0000000000000033000000000000001900000000",
            INIT_73 => X"000000030000000000000039000000000000000f000000000000002100000000",
            INIT_74 => X"0000005400000000000000630000000000000059000000000000002d00000000",
            INIT_75 => X"000000100000000000000028000000000000002a000000000000003c00000000",
            INIT_76 => X"0000002900000000000000100000000000000027000000000000005100000000",
            INIT_77 => X"0000001f00000000000000000000000000000010000000000000001700000000",
            INIT_78 => X"0000004000000000000000670000000000000065000000000000004800000000",
            INIT_79 => X"0000005500000000000000170000000000000020000000000000004100000000",
            INIT_7A => X"0000001b0000000000000019000000000000000f000000000000001100000000",
            INIT_7B => X"0000002000000000000000180000000000000006000000000000001e00000000",
            INIT_7C => X"0000002e00000000000000610000000000000055000000000000004000000000",
            INIT_7D => X"0000001b0000000000000062000000000000001a000000000000003000000000",
            INIT_7E => X"00000041000000000000002e0000000000000023000000000000001100000000",
            INIT_7F => X"000000280000000000000000000000000000001f000000000000000b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE1;


    MEM_IFMAP_LAYER1_INSTANCE2 : if BRAM_NAME = "ifmap_layer1_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002100000000000000220000000000000037000000000000002b00000000",
            INIT_01 => X"0000001a0000000000000035000000000000003e000000000000002e00000000",
            INIT_02 => X"00000020000000000000006c0000000000000041000000000000002200000000",
            INIT_03 => X"0000001900000000000000240000000000000000000000000000002100000000",
            INIT_04 => X"0000002700000000000000200000000000000031000000000000003000000000",
            INIT_05 => X"00000029000000000000000f0000000000000018000000000000003600000000",
            INIT_06 => X"000000220000000000000022000000000000006b000000000000006900000000",
            INIT_07 => X"0000000e00000000000000000000000000000044000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000020000000000000002d00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"00000010000000000000000f0000000000000009000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000005900000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000003000000000000000160000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"000000250000000000000024000000000000002a000000000000000000000000",
            INIT_1A => X"0000002a00000000000000230000000000000027000000000000002500000000",
            INIT_1B => X"0000002000000000000000210000000000000023000000000000002a00000000",
            INIT_1C => X"000000210000000000000025000000000000001f000000000000002600000000",
            INIT_1D => X"0000002500000000000000260000000000000027000000000000002a00000000",
            INIT_1E => X"00000022000000000000001b0000000000000020000000000000002300000000",
            INIT_1F => X"00000021000000000000000a000000000000000f000000000000000900000000",
            INIT_20 => X"000000270000000000000026000000000000002b000000000000003100000000",
            INIT_21 => X"0000002c0000000000000025000000000000002c000000000000003100000000",
            INIT_22 => X"0000001200000000000000110000000000000001000000000000003a00000000",
            INIT_23 => X"0000000e0000000000000007000000000000000b000000000000002100000000",
            INIT_24 => X"000000570000000000000000000000000000002d000000000000003600000000",
            INIT_25 => X"0000001000000000000000200000000000000027000000000000003000000000",
            INIT_26 => X"0000003500000000000000150000000000000006000000000000000a00000000",
            INIT_27 => X"0000001e00000000000000020000000000000016000000000000000000000000",
            INIT_28 => X"0000001b000000000000003d0000000000000000000000000000004300000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_2A => X"000000040000000000000028000000000000001a000000000000000100000000",
            INIT_2B => X"0000004300000000000000070000000000000018000000000000000000000000",
            INIT_2C => X"0000001900000000000000100000000000000027000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_2E => X"000000000000000000000000000000000000004f000000000000000900000000",
            INIT_2F => X"00000000000000000000000e0000000000000005000000000000001f00000000",
            INIT_30 => X"0000003b00000000000000020000000000000023000000000000001900000000",
            INIT_31 => X"0000000000000000000000000000000000000004000000000000001200000000",
            INIT_32 => X"0000001c00000000000000020000000000000000000000000000005100000000",
            INIT_33 => X"0000000000000000000000000000000000000015000000000000001300000000",
            INIT_34 => X"0000002c000000000000001c000000000000000c000000000000000e00000000",
            INIT_35 => X"0000004a00000000000000010000000000000011000000000000000000000000",
            INIT_36 => X"00000024000000000000001e0000000000000004000000000000000000000000",
            INIT_37 => X"0000000000000000000000020000000000000000000000000000001c00000000",
            INIT_38 => X"000000070000000000000013000000000000000f000000000000001b00000000",
            INIT_39 => X"00000029000000000000001c0000000000000020000000000000001300000000",
            INIT_3A => X"0000002b00000000000000270000000000000028000000000000000200000000",
            INIT_3B => X"0000002100000000000000000000000000000006000000000000000000000000",
            INIT_3C => X"00000000000000000000000c0000000000000013000000000000000000000000",
            INIT_3D => X"0000000e0000000000000000000000000000000e000000000000002800000000",
            INIT_3E => X"000000230000000000000021000000000000003f000000000000003100000000",
            INIT_3F => X"0000000000000000000000370000000000000000000000000000000400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000019000000000000000000000000",
            INIT_41 => X"0000001d00000000000000090000000000000011000000000000000000000000",
            INIT_42 => X"0000000c00000000000000480000000000000006000000000000001d00000000",
            INIT_43 => X"0000000000000000000000000000000000000039000000000000000000000000",
            INIT_44 => X"0000000900000000000000040000000000000011000000000000001700000000",
            INIT_45 => X"00000013000000000000000a000000000000000f000000000000000f00000000",
            INIT_46 => X"0000001300000000000000440000000000000011000000000000000800000000",
            INIT_47 => X"0000000900000000000000080000000000000000000000000000001700000000",
            INIT_48 => X"0000000e0000000000000010000000000000000f000000000000000e00000000",
            INIT_49 => X"0000000900000000000000040000000000000010000000000000001100000000",
            INIT_4A => X"0000000000000000000000520000000000000013000000000000000200000000",
            INIT_4B => X"0000000f00000000000000050000000000000010000000000000000000000000",
            INIT_4C => X"00000011000000000000000f000000000000000d000000000000000a00000000",
            INIT_4D => X"0000000000000000000000160000000000000015000000000000000500000000",
            INIT_4E => X"0000001100000000000000200000000000000019000000000000000c00000000",
            INIT_4F => X"0000000900000000000000080000000000000011000000000000001d00000000",
            INIT_50 => X"0000000d000000000000000d000000000000000a000000000000000900000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000001200000000000000020000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000005000000000000001200000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"000000010000000000000000000000000000000c000000000000000000000000",
            INIT_5B => X"0000002e000000000000003f000000000000003b000000000000000500000000",
            INIT_5C => X"000000060000000000000000000000000000000b000000000000001c00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_5E => X"0000002600000000000000140000000000000010000000000000000000000000",
            INIT_5F => X"000000210000000000000029000000000000002b000000000000004200000000",
            INIT_60 => X"0000004400000000000000210000000000000004000000000000001300000000",
            INIT_61 => X"0000001200000000000000140000000000000000000000000000000000000000",
            INIT_62 => X"00000029000000000000002b000000000000001e000000000000002c00000000",
            INIT_63 => X"0000001300000000000000270000000000000015000000000000003100000000",
            INIT_64 => X"0000000000000000000000680000000000000046000000000000000f00000000",
            INIT_65 => X"000000310000000000000026000000000000006e000000000000000000000000",
            INIT_66 => X"00000041000000000000004e0000000000000020000000000000001f00000000",
            INIT_67 => X"0000000d00000000000000220000000000000031000000000000002100000000",
            INIT_68 => X"000000000000000000000002000000000000006f000000000000003900000000",
            INIT_69 => X"0000002a00000000000000510000000000000033000000000000003300000000",
            INIT_6A => X"00000028000000000000003b000000000000006c000000000000002300000000",
            INIT_6B => X"00000048000000000000001f0000000000000031000000000000002f00000000",
            INIT_6C => X"0000000b0000000000000000000000000000001e000000000000006200000000",
            INIT_6D => X"0000002000000000000000440000000000000048000000000000006100000000",
            INIT_6E => X"0000003500000000000000300000000000000038000000000000005600000000",
            INIT_6F => X"0000007c00000000000000630000000000000004000000000000003600000000",
            INIT_70 => X"0000003d00000000000000150000000000000042000000000000003b00000000",
            INIT_71 => X"0000002000000000000000290000000000000031000000000000002900000000",
            INIT_72 => X"00000015000000000000002a0000000000000022000000000000003900000000",
            INIT_73 => X"00000048000000000000007a000000000000006f000000000000000000000000",
            INIT_74 => X"0000002d000000000000001b0000000000000036000000000000006300000000",
            INIT_75 => X"0000001f0000000000000026000000000000003a000000000000004000000000",
            INIT_76 => X"000000000000000000000000000000000000001e000000000000001600000000",
            INIT_77 => X"0000007a000000000000004f000000000000006b000000000000008900000000",
            INIT_78 => X"0000007200000000000000680000000000000038000000000000004000000000",
            INIT_79 => X"00000045000000000000003c000000000000002b000000000000003a00000000",
            INIT_7A => X"000000c5000000000000004e0000000000000063000000000000005e00000000",
            INIT_7B => X"000000930000000000000099000000000000004e000000000000008f00000000",
            INIT_7C => X"000000770000000000000087000000000000008b000000000000007c00000000",
            INIT_7D => X"00000096000000000000008e0000000000000085000000000000007600000000",
            INIT_7E => X"000000b100000000000000a70000000000000096000000000000009d00000000",
            INIT_7F => X"00000080000000000000006c00000000000000a5000000000000007700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE2;


    MEM_IFMAP_LAYER1_INSTANCE3 : if BRAM_NAME = "ifmap_layer1_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000087000000000000007f000000000000007f000000000000007f00000000",
            INIT_01 => X"0000009d00000000000000a0000000000000009c000000000000009300000000",
            INIT_02 => X"000000b1000000000000009c00000000000000ac00000000000000a900000000",
            INIT_03 => X"00000082000000000000008a000000000000006e00000000000000a600000000",
            INIT_04 => X"000000a100000000000000910000000000000084000000000000008200000000",
            INIT_05 => X"000000c200000000000000b700000000000000a300000000000000ac00000000",
            INIT_06 => X"000000a5000000000000009b00000000000000a700000000000000aa00000000",
            INIT_07 => X"00000083000000000000008f0000000000000091000000000000008200000000",
            INIT_08 => X"0000009900000000000000970000000000000095000000000000008600000000",
            INIT_09 => X"00000078000000000000009900000000000000bd00000000000000a400000000",
            INIT_0A => X"0000007e000000000000007f000000000000007b000000000000007b00000000",
            INIT_0B => X"00000082000000000000008b000000000000007c000000000000007600000000",
            INIT_0C => X"0000006100000000000000560000000000000053000000000000006500000000",
            INIT_0D => X"00000081000000000000007a0000000000000073000000000000006e00000000",
            INIT_0E => X"00000061000000000000007f0000000000000081000000000000007e00000000",
            INIT_0F => X"0000003200000000000000500000000000000063000000000000006f00000000",
            INIT_10 => X"00000050000000000000002f0000000000000020000000000000001d00000000",
            INIT_11 => X"0000008100000000000000500000000000000047000000000000006900000000",
            INIT_12 => X"0000004e00000000000000670000000000000083000000000000008500000000",
            INIT_13 => X"0000001d0000000000000013000000000000002a000000000000003900000000",
            INIT_14 => X"0000004d0000000000000029000000000000001d000000000000001e00000000",
            INIT_15 => X"0000007f00000000000000730000000000000021000000000000003100000000",
            INIT_16 => X"0000002900000000000000320000000000000053000000000000006700000000",
            INIT_17 => X"000000230000000000000029000000000000001a000000000000001a00000000",
            INIT_18 => X"000000280000000000000031000000000000001f000000000000002200000000",
            INIT_19 => X"0000002b00000000000000690000000000000067000000000000000c00000000",
            INIT_1A => X"0000001800000000000000250000000000000029000000000000003100000000",
            INIT_1B => X"0000001c000000000000002a0000000000000028000000000000001d00000000",
            INIT_1C => X"0000000600000000000000220000000000000022000000000000002000000000",
            INIT_1D => X"0000003600000000000000150000000000000068000000000000006600000000",
            INIT_1E => X"00000004000000000000001e000000000000002f000000000000002700000000",
            INIT_1F => X"0000001e00000000000000190000000000000029000000000000002400000000",
            INIT_20 => X"0000003e0000000000000000000000000000002b000000000000001d00000000",
            INIT_21 => X"0000001c00000000000000270000000000000028000000000000006d00000000",
            INIT_22 => X"0000002700000000000000000000000000000025000000000000002800000000",
            INIT_23 => X"00000026000000000000001a0000000000000019000000000000002200000000",
            INIT_24 => X"0000003b0000000000000022000000000000000c000000000000001d00000000",
            INIT_25 => X"0000001e0000000000000026000000000000000e000000000000004300000000",
            INIT_26 => X"00000026000000000000002b0000000000000022000000000000002d00000000",
            INIT_27 => X"00000012000000000000004f000000000000001e000000000000001600000000",
            INIT_28 => X"00000031000000000000000c000000000000001c000000000000000000000000",
            INIT_29 => X"0000001d000000000000001f0000000000000032000000000000002900000000",
            INIT_2A => X"0000001c00000000000000280000000000000029000000000000003400000000",
            INIT_2B => X"0000000c0000000000000016000000000000005c000000000000003b00000000",
            INIT_2C => X"0000002300000000000000180000000000000000000000000000001600000000",
            INIT_2D => X"00000025000000000000001d0000000000000018000000000000002100000000",
            INIT_2E => X"00000040000000000000000c0000000000000014000000000000001b00000000",
            INIT_2F => X"00000016000000000000000f0000000000000000000000000000005e00000000",
            INIT_30 => X"00000000000000000000000a0000000000000014000000000000000000000000",
            INIT_31 => X"0000000000000000000000040000000000000001000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000040000000000000000000000000000000500000000",
            INIT_43 => X"0000000000000000000000030000000000000001000000000000000000000000",
            INIT_44 => X"0000001100000000000000020000000000000000000000000000000000000000",
            INIT_45 => X"0000000200000000000000000000000000000000000000000000000400000000",
            INIT_46 => X"0000000800000000000000000000000000000005000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000001600000000000000000000000000000000000000000000001500000000",
            INIT_49 => X"0000004400000000000000000000000000000000000000000000001c00000000",
            INIT_4A => X"0000001c00000000000000080000000000000000000000000000000400000000",
            INIT_4B => X"0000003d00000000000000090000000000000000000000000000000000000000",
            INIT_4C => X"0000002400000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"00000000000000000000005f0000000000000000000000000000002200000000",
            INIT_4E => X"0000000000000000000000160000000000000000000000000000000800000000",
            INIT_4F => X"00000000000000000000006d0000000000000000000000000000000000000000",
            INIT_50 => X"0000005f00000000000000000000000000000000000000000000000200000000",
            INIT_51 => X"000000520000000000000000000000000000001c000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000086000000000000000000000000",
            INIT_54 => X"0000000000000000000000330000000000000000000000000000000000000000",
            INIT_55 => X"0000007600000000000000190000000000000000000000000000001800000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_57 => X"000000130000000000000000000000000000000000000000000000d200000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"00000040000000000000005f0000000000000000000000000000000f00000000",
            INIT_5A => X"000000b100000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"00000010000000000000000b0000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"000000000000000000000054000000000000003d000000000000000000000000",
            INIT_5E => X"0000000000000000000000740000000000000000000000000000000500000000",
            INIT_5F => X"00000000000000000000000f0000000000000025000000000000000000000000",
            INIT_60 => X"0000003100000000000000000000000000000007000000000000000000000000",
            INIT_61 => X"000000000000000000000000000000000000002e000000000000000000000000",
            INIT_62 => X"0000000000000000000000200000000000000000000000000000002700000000",
            INIT_63 => X"00000000000000000000000b0000000000000025000000000000002b00000000",
            INIT_64 => X"0000000000000000000000550000000000000000000000000000000d00000000",
            INIT_65 => X"0000000000000000000000000000000000000034000000000000000c00000000",
            INIT_66 => X"0000002f00000000000000040000000000000000000000000000000300000000",
            INIT_67 => X"00000005000000000000005a0000000000000000000000000000002900000000",
            INIT_68 => X"00000000000000000000000000000000000000aa000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000003e00000000",
            INIT_6A => X"0000001f00000000000000160000000000000006000000000000000000000000",
            INIT_6B => X"00000000000000000000004c0000000000000075000000000000000000000000",
            INIT_6C => X"0000001f00000000000000000000000000000000000000000000007a00000000",
            INIT_6D => X"0000000c00000000000000080000000000000000000000000000001a00000000",
            INIT_6E => X"00000000000000000000000d000000000000000c000000000000001000000000",
            INIT_6F => X"0000000000000000000000840000000000000071000000000000000000000000",
            INIT_70 => X"0000000600000000000000000000000000000002000000000000000000000000",
            INIT_71 => X"00000008000000000000000d0000000000000009000000000000000200000000",
            INIT_72 => X"00000000000000000000000e000000000000000f000000000000000600000000",
            INIT_73 => X"00000000000000000000000000000000000000bd000000000000001100000000",
            INIT_74 => X"0000000e00000000000000010000000000000000000000000000000c00000000",
            INIT_75 => X"000000040000000000000010000000000000000b000000000000000b00000000",
            INIT_76 => X"0000000c00000000000000000000000000000000000000000000002000000000",
            INIT_77 => X"0000002500000000000000000000000000000007000000000000002300000000",
            INIT_78 => X"00000000000000000000000b0000000000000006000000000000001800000000",
            INIT_79 => X"00000000000000000000002d000000000000000f000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000002500000000000000160000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000004000000000000001c00000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000e00000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE3;


    MEM_IFMAP_LAYER1_INSTANCE4 : if BRAM_NAME = "ifmap_layer1_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000000000000c000000000000004500000000",
            INIT_01 => X"0000002700000000000000000000000000000018000000000000001d00000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_03 => X"00000001000000000000002b0000000000000025000000000000004e00000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000006000000000000001e00000000",
            INIT_06 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"00000000000000000000000a0000000000000010000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_0B => X"0000000000000000000000070000000000000009000000000000000000000000",
            INIT_0C => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000002900000000000000000000000000000000000000000000000a00000000",
            INIT_0E => X"0000000000000000000000000000000000000022000000000000006400000000",
            INIT_0F => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_11 => X"000000280000000000000000000000000000001a000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000600000000000000050000000000000000000000000000000000000000",
            INIT_16 => X"000000050000000000000000000000000000002b000000000000002000000000",
            INIT_17 => X"00000007000000000000000b0000000000000000000000000000000100000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000600000000000000540000000000000000000000000000000000000000",
            INIT_1A => X"0000003100000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"000000000000000000000000000000000000001f000000000000003a00000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_1D => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_1E => X"0000001a0000000000000037000000000000003f000000000000000000000000",
            INIT_1F => X"0000001000000000000000050000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"00000008000000000000002f0000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"000000320000000000000065000000000000002b000000000000002700000000",
            INIT_24 => X"0000006800000000000000500000000000000000000000000000000000000000",
            INIT_25 => X"00000013000000000000001e0000000000000043000000000000004600000000",
            INIT_26 => X"0000000000000000000000000000000000000009000000000000000500000000",
            INIT_27 => X"0000001900000000000000490000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000056000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_2B => X"0000004100000000000000510000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_2D => X"0000001300000000000000060000000000000000000000000000000200000000",
            INIT_2E => X"0000000000000000000000260000000000000000000000000000000800000000",
            INIT_2F => X"0000001f000000000000004e000000000000000b000000000000000000000000",
            INIT_30 => X"0000000000000000000000010000000000000024000000000000002400000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"000000a600000000000000a80000000000000000000000000000000000000000",
            INIT_33 => X"000000a400000000000000ad00000000000000ad00000000000000af00000000",
            INIT_34 => X"0000009100000000000000aa00000000000000b700000000000000b800000000",
            INIT_35 => X"00000096000000000000008f0000000000000086000000000000007b00000000",
            INIT_36 => X"000000b500000000000000b300000000000000ab000000000000008a00000000",
            INIT_37 => X"000000b300000000000000c400000000000000b400000000000000b200000000",
            INIT_38 => X"0000004f0000000000000057000000000000006400000000000000a000000000",
            INIT_39 => X"000000920000000000000080000000000000005d000000000000005200000000",
            INIT_3A => X"000000b100000000000000b6000000000000008d000000000000007200000000",
            INIT_3B => X"000000350000000000000054000000000000008b00000000000000b600000000",
            INIT_3C => X"0000003b00000000000000460000000000000065000000000000004100000000",
            INIT_3D => X"0000002a00000000000000850000000000000051000000000000003500000000",
            INIT_3E => X"000000a200000000000000b700000000000000b9000000000000009400000000",
            INIT_3F => X"00000034000000000000003f0000000000000071000000000000007f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000014000000000000003d0000000000000043000000000000006900000000",
            INIT_41 => X"000000a3000000000000002f0000000000000076000000000000001e00000000",
            INIT_42 => X"000000ac00000000000000c600000000000000bf00000000000000ad00000000",
            INIT_43 => X"00000063000000000000001c0000000000000036000000000000005a00000000",
            INIT_44 => X"0000001f000000000000003b0000000000000040000000000000006900000000",
            INIT_45 => X"000000a400000000000000770000000000000039000000000000004f00000000",
            INIT_46 => X"0000006800000000000000670000000000000057000000000000008400000000",
            INIT_47 => X"0000006200000000000000ac0000000000000021000000000000004900000000",
            INIT_48 => X"0000002f000000000000002c000000000000003e000000000000001f00000000",
            INIT_49 => X"00000077000000000000007c000000000000005a000000000000004400000000",
            INIT_4A => X"0000005d000000000000007b0000000000000095000000000000006e00000000",
            INIT_4B => X"0000002e000000000000003d000000000000009e000000000000002400000000",
            INIT_4C => X"0000005c00000000000000420000000000000043000000000000003500000000",
            INIT_4D => X"00000080000000000000007c0000000000000069000000000000005400000000",
            INIT_4E => X"0000002a0000000000000041000000000000004700000000000000ae00000000",
            INIT_4F => X"000000380000000000000022000000000000003e000000000000008f00000000",
            INIT_50 => X"0000006d000000000000005a0000000000000058000000000000004b00000000",
            INIT_51 => X"0000003600000000000000740000000000000065000000000000002b00000000",
            INIT_52 => X"00000064000000000000005f0000000000000048000000000000003b00000000",
            INIT_53 => X"0000005e00000000000000220000000000000004000000000000004400000000",
            INIT_54 => X"000000220000000000000069000000000000005a00000000000000a300000000",
            INIT_55 => X"000000630000000000000053000000000000004b000000000000005e00000000",
            INIT_56 => X"0000000800000000000000400000000000000059000000000000006a00000000",
            INIT_57 => X"0000009400000000000000a7000000000000004c000000000000000800000000",
            INIT_58 => X"000000b3000000000000001f0000000000000074000000000000006d00000000",
            INIT_59 => X"0000004d00000000000000850000000000000077000000000000007c00000000",
            INIT_5A => X"0000002000000000000000110000000000000015000000000000001f00000000",
            INIT_5B => X"00000024000000000000002d000000000000003c000000000000002900000000",
            INIT_5C => X"0000002200000000000000de0000000000000059000000000000004f00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"000000000000000000000000000000000000008d000000000000006f00000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000005a00000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000c00000000000000000000000000000000000000000000000900000000",
            INIT_6B => X"0000000e0000000000000011000000000000000b000000000000001100000000",
            INIT_6C => X"0000000d0000000000000011000000000000000d000000000000000900000000",
            INIT_6D => X"000000090000000000000003000000000000000e000000000000000d00000000",
            INIT_6E => X"0000000900000000000000060000000000000013000000000000000f00000000",
            INIT_6F => X"0000000000000000000000070000000000000014000000000000000800000000",
            INIT_70 => X"0000000000000000000000270000000000000009000000000000002100000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_72 => X"0000000900000000000000000000000000000013000000000000000b00000000",
            INIT_73 => X"0000003a000000000000000e0000000000000007000000000000001200000000",
            INIT_74 => X"0000003100000000000000000000000000000000000000000000001000000000",
            INIT_75 => X"000000000000000000000000000000000000002e000000000000002600000000",
            INIT_76 => X"00000001000000000000000a0000000000000000000000000000005e00000000",
            INIT_77 => X"0000002700000000000000140000000000000000000000000000000f00000000",
            INIT_78 => X"0000001a00000000000000540000000000000000000000000000001500000000",
            INIT_79 => X"0000007d00000000000000000000000000000013000000000000003500000000",
            INIT_7A => X"0000001800000000000000000000000000000037000000000000000000000000",
            INIT_7B => X"0000002200000000000000390000000000000052000000000000002800000000",
            INIT_7C => X"0000000700000000000000490000000000000023000000000000000000000000",
            INIT_7D => X"00000009000000000000006c0000000000000000000000000000002d00000000",
            INIT_7E => X"0000004c0000000000000000000000000000001b000000000000004e00000000",
            INIT_7F => X"000000000000000000000040000000000000003b000000000000005100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE4;


    MEM_IFMAP_LAYER1_INSTANCE5 : if BRAM_NAME = "ifmap_layer1_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000270000000000000000000000000000005f000000000000006b00000000",
            INIT_01 => X"00000013000000000000003f0000000000000068000000000000001400000000",
            INIT_02 => X"0000004100000000000000000000000000000000000000000000004700000000",
            INIT_03 => X"0000007900000000000000000000000000000059000000000000004a00000000",
            INIT_04 => X"0000002800000000000000000000000000000002000000000000003900000000",
            INIT_05 => X"000000210000000000000023000000000000004e000000000000005700000000",
            INIT_06 => X"0000003200000000000000900000000000000000000000000000000000000000",
            INIT_07 => X"00000045000000000000005a0000000000000000000000000000004200000000",
            INIT_08 => X"00000065000000000000002c0000000000000013000000000000000000000000",
            INIT_09 => X"0000001d0000000000000000000000000000007d000000000000002400000000",
            INIT_0A => X"00000000000000000000000f0000000000000031000000000000002600000000",
            INIT_0B => X"00000000000000000000005b0000000000000000000000000000002800000000",
            INIT_0C => X"0000003000000000000000460000000000000000000000000000000000000000",
            INIT_0D => X"0000001500000000000000440000000000000000000000000000008f00000000",
            INIT_0E => X"0000002d0000000000000015000000000000002f000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000007000000000000005400000000",
            INIT_10 => X"00000089000000000000002c0000000000000000000000000000001700000000",
            INIT_11 => X"000000000000000000000023000000000000008d000000000000000000000000",
            INIT_12 => X"0000000000000000000000280000000000000069000000000000004e00000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"000000000000000000000054000000000000000c000000000000000000000000",
            INIT_15 => X"000000110000000000000010000000000000006400000000000000c200000000",
            INIT_16 => X"0000000800000000000000080000000000000009000000000000001c00000000",
            INIT_17 => X"00000021000000000000001b000000000000000f000000000000000c00000000",
            INIT_18 => X"000000b600000000000000410000000000000000000000000000000000000000",
            INIT_19 => X"000000110000000000000011000000000000001a000000000000001400000000",
            INIT_1A => X"0000001500000000000000030000000000000004000000000000000800000000",
            INIT_1B => X"0000000600000000000000310000000000000003000000000000001700000000",
            INIT_1C => X"0000000b00000000000000410000000000000091000000000000000000000000",
            INIT_1D => X"0000000c000000000000000e0000000000000010000000000000002000000000",
            INIT_1E => X"00000000000000000000001f0000000000000014000000000000001200000000",
            INIT_1F => X"0000000700000000000000110000000000000040000000000000003700000000",
            INIT_20 => X"000000150000000000000000000000000000001f000000000000001d00000000",
            INIT_21 => X"000000220000000000000011000000000000000b000000000000001a00000000",
            INIT_22 => X"00000050000000000000002f0000000000000000000000000000001000000000",
            INIT_23 => X"00000053000000000000004b0000000000000053000000000000004d00000000",
            INIT_24 => X"000000550000000000000054000000000000004a000000000000004f00000000",
            INIT_25 => X"000000400000000000000047000000000000004a000000000000004e00000000",
            INIT_26 => X"0000004a0000000000000049000000000000004b000000000000004800000000",
            INIT_27 => X"000000490000000000000058000000000000004a000000000000004f00000000",
            INIT_28 => X"00000054000000000000004f0000000000000068000000000000004c00000000",
            INIT_29 => X"0000002600000000000000340000000000000041000000000000002c00000000",
            INIT_2A => X"00000032000000000000004f0000000000000048000000000000003a00000000",
            INIT_2B => X"00000049000000000000004b0000000000000057000000000000005200000000",
            INIT_2C => X"00000009000000000000001f0000000000000040000000000000007c00000000",
            INIT_2D => X"0000001700000000000000530000000000000050000000000000006200000000",
            INIT_2E => X"0000005b0000000000000000000000000000008e000000000000003600000000",
            INIT_2F => X"00000056000000000000002f0000000000000059000000000000004700000000",
            INIT_30 => X"0000008e0000000000000000000000000000003a000000000000004500000000",
            INIT_31 => X"000000000000000000000036000000000000005c000000000000004300000000",
            INIT_32 => X"000000040000000000000082000000000000002500000000000000b200000000",
            INIT_33 => X"00000065000000000000008f0000000000000053000000000000007a00000000",
            INIT_34 => X"00000075000000000000006a0000000000000000000000000000004500000000",
            INIT_35 => X"0000009400000000000000000000000000000050000000000000003200000000",
            INIT_36 => X"00000044000000000000003b00000000000000a1000000000000006800000000",
            INIT_37 => X"0000006c000000000000006d00000000000000aa000000000000008900000000",
            INIT_38 => X"00000029000000000000008b00000000000000a9000000000000000000000000",
            INIT_39 => X"0000009500000000000000950000000000000036000000000000004a00000000",
            INIT_3A => X"0000003800000000000000000000000000000086000000000000006f00000000",
            INIT_3B => X"00000000000000000000008a0000000000000089000000000000009700000000",
            INIT_3C => X"0000002f000000000000002b000000000000006b00000000000000be00000000",
            INIT_3D => X"0000005600000000000000a40000000000000095000000000000005600000000",
            INIT_3E => X"000000be000000000000002a0000000000000009000000000000007700000000",
            INIT_3F => X"000000990000000000000000000000000000007b000000000000006700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005a0000000000000041000000000000001c000000000000007700000000",
            INIT_41 => X"0000004200000000000000b2000000000000007900000000000000ad00000000",
            INIT_42 => X"0000004d00000000000000740000000000000050000000000000005600000000",
            INIT_43 => X"00000077000000000000003e000000000000005c000000000000002900000000",
            INIT_44 => X"00000097000000000000003b0000000000000032000000000000001600000000",
            INIT_45 => X"0000008d000000000000000e00000000000000d6000000000000007a00000000",
            INIT_46 => X"0000003f0000000000000080000000000000002b000000000000002c00000000",
            INIT_47 => X"000000030000000000000021000000000000006d000000000000005d00000000",
            INIT_48 => X"0000007f0000000000000042000000000000005f000000000000002600000000",
            INIT_49 => X"0000006000000000000000ec000000000000000000000000000000ce00000000",
            INIT_4A => X"0000004a000000000000009d0000000000000092000000000000002300000000",
            INIT_4B => X"00000028000000000000000f000000000000000d000000000000001500000000",
            INIT_4C => X"0000009d00000000000000600000000000000006000000000000004300000000",
            INIT_4D => X"0000003f000000000000009e0000000000000111000000000000001600000000",
            INIT_4E => X"00000029000000000000002a000000000000004a000000000000004300000000",
            INIT_4F => X"0000004000000000000000300000000000000030000000000000002700000000",
            INIT_50 => X"000000ac00000000000000270000000000000001000000000000004300000000",
            INIT_51 => X"0000002f0000000000000036000000000000003600000000000000e100000000",
            INIT_52 => X"0000002800000000000000230000000000000025000000000000002e00000000",
            INIT_53 => X"0000005400000000000000300000000000000036000000000000003700000000",
            INIT_54 => X"0000006600000000000000f30000000000000000000000000000002a00000000",
            INIT_55 => X"00000028000000000000002f0000000000000042000000000000002b00000000",
            INIT_56 => X"0000003e0000000000000037000000000000002d000000000000002900000000",
            INIT_57 => X"0000002f000000000000005e0000000000000057000000000000001800000000",
            INIT_58 => X"0000001e000000000000003a0000000000000055000000000000002b00000000",
            INIT_59 => X"0000003600000000000000290000000000000038000000000000003200000000",
            INIT_5A => X"000000570000000000000014000000000000002b000000000000004100000000",
            INIT_5B => X"0000003b0000000000000034000000000000003a000000000000006f00000000",
            INIT_5C => X"0000004200000000000000340000000000000039000000000000003800000000",
            INIT_5D => X"0000002f000000000000002f0000000000000039000000000000004600000000",
            INIT_5E => X"0000002c00000000000000320000000000000032000000000000003400000000",
            INIT_5F => X"0000003b000000000000003a000000000000003b000000000000004000000000",
            INIT_60 => X"000000370000000000000039000000000000001f000000000000003700000000",
            INIT_61 => X"000000080000000000000000000000000000000c000000000000002700000000",
            INIT_62 => X"0000002400000000000000300000000000000037000000000000002300000000",
            INIT_63 => X"0000003c00000000000000400000000000000041000000000000004f00000000",
            INIT_64 => X"0000000100000000000000130000000000000025000000000000001100000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000001c0000000000000000000000000000002e000000000000001a00000000",
            INIT_67 => X"0000001f000000000000002e000000000000003d000000000000004400000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000003800000000000000000000000000000000000000000000002500000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"00000002000000000000003d0000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"00000000000000000000001c0000000000000047000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000022000000000000000400000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000001a00000000000000030000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE5;


    MEM_IFMAP_LAYER1_INSTANCE6 : if BRAM_NAME = "ifmap_layer1_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000031000000000000001b000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000002400000000000000240000000000000000000000000000000000000000",
            INIT_14 => X"0000001c000000000000001f000000000000001e000000000000002000000000",
            INIT_15 => X"0000002400000000000000200000000000000029000000000000002700000000",
            INIT_16 => X"00000021000000000000001e0000000000000029000000000000002d00000000",
            INIT_17 => X"00000021000000000000001d000000000000001f000000000000001e00000000",
            INIT_18 => X"0000001d00000000000000000000000000000017000000000000002100000000",
            INIT_19 => X"000000000000000000000000000000000000003d000000000000002800000000",
            INIT_1A => X"00000019000000000000001d0000000000000023000000000000000700000000",
            INIT_1B => X"00000023000000000000001f0000000000000031000000000000003b00000000",
            INIT_1C => X"0000002200000000000000330000000000000042000000000000002400000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"000000000000000000000014000000000000001e000000000000000000000000",
            INIT_1F => X"0000001b000000000000001a0000000000000019000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000d0000000000000015000000000000000a000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000014000000000000001100000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_24 => X"0000000000000000000000180000000000000006000000000000000900000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000001e00000000000000000000000000000008000000000000002200000000",
            INIT_27 => X"00000000000000000000001f000000000000002b000000000000004400000000",
            INIT_28 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_2A => X"00000020000000000000002b0000000000000002000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_2C => X"00000000000000000000000c0000000000000000000000000000000100000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000a00000000000000250000000000000032000000000000000000000000",
            INIT_30 => X"00000000000000000000000d000000000000000d000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000013000000000000001000000000",
            INIT_32 => X"0000003800000000000000080000000000000000000000000000000c00000000",
            INIT_33 => X"0000001e00000000000000000000000000000000000000000000000d00000000",
            INIT_34 => X"000000000000000000000018000000000000003d000000000000001500000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_36 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_37 => X"000000330000000000000028000000000000000e000000000000000000000000",
            INIT_38 => X"0000001e00000000000000000000000000000000000000000000000700000000",
            INIT_39 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_3A => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_3C => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000004700000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"00000000000000000000000d0000000000000012000000000000002e00000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000100000000000000120000000000000017000000000000000700000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"00000000000000000000001c000000000000000e000000000000000000000000",
            INIT_52 => X"0000000c000000000000000d0000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000290000000000000022000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"00000004000000000000000e0000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_5A => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_5F => X"0000000900000000000000150000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_62 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"000000060000000000000014000000000000001d000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_6A => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"00000000000000000000000c0000000000000005000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000001400000000000000040000000000000000000000000000000000000000",
            INIT_6F => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000070000000000000000000000000000001600000000",
            INIT_71 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_72 => X"0000002f00000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000023000000000000002e00000000",
            INIT_74 => X"0000001b00000000000000190000000000000005000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000021000000000000002d00000000",
            INIT_76 => X"000000000000000000000000000000000000000e000000000000001500000000",
            INIT_77 => X"0000000000000000000000010000000000000002000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"00000003000000000000000b000000000000000b000000000000001c00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"000000000000000000000003000000000000001f000000000000003100000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE6;


    MEM_IFMAP_LAYER1_INSTANCE7 : if BRAM_NAME = "ifmap_layer1_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_01 => X"0000000a00000000000000030000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE7;


    MEM_IFMAP_LAYER2_INSTANCE0 : if BRAM_NAME = "ifmap_layer2_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_01 => X"000000d500000000000000040000000000000000000000000000002000000000",
            INIT_02 => X"0000006100000000000000080000000000000000000000000000002c00000000",
            INIT_03 => X"0000002a0000000000000042000000000000002a000000000000000700000000",
            INIT_04 => X"0000001e00000000000001540000000000000000000000000000000000000000",
            INIT_05 => X"00000000000000000000004e0000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000042000000000000002800000000",
            INIT_07 => X"00000000000000000000001e0000000000000140000000000000000000000000",
            INIT_08 => X"000000000000000000000000000000000000004c000000000000000000000000",
            INIT_09 => X"0000004200000000000000000000000000000032000000000000000000000000",
            INIT_0A => X"0000000000000000000000180000000000000000000000000000000f00000000",
            INIT_0B => X"000000040000000000000004000000000000000c000000000000003c00000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"000000020000000000000000000000000000007a000000000000007b00000000",
            INIT_0E => X"0000002900000000000000000000000000000000000000000000003b00000000",
            INIT_0F => X"0000000000000000000000760000000000000010000000000000000000000000",
            INIT_10 => X"0000007400000000000000000000000000000000000000000000007a00000000",
            INIT_11 => X"0000003000000000000000000000000000000000000000000000008400000000",
            INIT_12 => X"000000c700000000000000000000000000000067000000000000000000000000",
            INIT_13 => X"0000000f00000000000000a20000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000af000000000000005f000000000000000000000000",
            INIT_15 => X"00000021000000000000016d0000000000000000000000000000000000000000",
            INIT_16 => X"0000008b00000000000000000000000000000000000000000000004900000000",
            INIT_17 => X"0000000000000000000000190000000000000078000000000000000000000000",
            INIT_18 => X"0000003e00000000000000470000000000000000000000000000000400000000",
            INIT_19 => X"0000005d0000000000000044000000000000003c000000000000004a00000000",
            INIT_1A => X"00000067000000000000005b0000000000000068000000000000007500000000",
            INIT_1B => X"000000700000000000000067000000000000002d000000000000005a00000000",
            INIT_1C => X"0000005d000000000000004d000000000000003c000000000000004200000000",
            INIT_1D => X"000000000000000000000056000000000000004c000000000000000000000000",
            INIT_1E => X"00000035000000000000005c0000000000000012000000000000002800000000",
            INIT_1F => X"0000001000000000000000000000000000000092000000000000007300000000",
            INIT_20 => X"0000002800000000000000260000000000000032000000000000003c00000000",
            INIT_21 => X"0000000000000000000000000000000000000002000000000000007000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"000000000000000000000000000000000000001b000000000000000000000000",
            INIT_24 => X"0000003600000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000045000000000000007100000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000002a0000000000000000000000000000001f000000000000001200000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000001b00000000000000000000000000000000000000000000000e00000000",
            INIT_2A => X"0000001a00000000000000010000000000000000000000000000000000000000",
            INIT_2B => X"00000000000000000000004d0000000000000036000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"00000103000000000000000000000000000000b0000000000000000000000000",
            INIT_33 => X"0000000e00000000000000420000000000000077000000000000000000000000",
            INIT_34 => X"0000015000000000000000b50000000000000135000000000000004700000000",
            INIT_35 => X"0000005d0000000000000064000000000000003c000000000000000000000000",
            INIT_36 => X"0000000000000000000000390000000000000029000000000000000000000000",
            INIT_37 => X"000000000000000000000027000000000000013a000000000000000000000000",
            INIT_38 => X"00000000000000000000010f0000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000180000000000000010000000000000005300000000",
            INIT_3A => X"0000000000000000000000000000000000000062000000000000014500000000",
            INIT_3B => X"0000000000000000000001d40000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_3D => X"000000460000000000000086000000000000003c000000000000001c00000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_3F => X"0000001d00000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000700000000000000000000000000000032000000000000000000000000",
            INIT_41 => X"000000000000000000000040000000000000000e000000000000000000000000",
            INIT_42 => X"00000000000000000000001b0000000000000000000000000000004e00000000",
            INIT_43 => X"0000003400000000000000000000000000000069000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000031000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_4D => X"0000005500000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000005500000000000000000000000000000044000000000000000000000000",
            INIT_4F => X"0000000000000000000000270000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000540000000000000000000000000000002e00000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000003600000000",
            INIT_52 => X"000000c000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000039000000000000000000000000",
            INIT_54 => X"0000003800000000000000620000000000000000000000000000005d00000000",
            INIT_55 => X"0000000000000000000000450000000000000003000000000000002b00000000",
            INIT_56 => X"0000004400000000000000010000000000000025000000000000000000000000",
            INIT_57 => X"0000007500000000000000030000000000000000000000000000004600000000",
            INIT_58 => X"0000001000000000000000000000000000000030000000000000007300000000",
            INIT_59 => X"0000004d00000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000004400000000000000040000000000000000000000000000008600000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000008400000000",
            INIT_5C => X"0000005800000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"000000000000000000000092000000000000000c000000000000007400000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000006900000000000000100000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000005300000000",
            INIT_61 => X"0000000000000000000000000000000000000015000000000000000900000000",
            INIT_62 => X"0000008d00000000000000000000000000000005000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000200000000000000029000000000000000000000000",
            INIT_65 => X"0000000000000000000000010000000000000000000000000000004900000000",
            INIT_66 => X"0000006900000000000000000000000000000061000000000000000000000000",
            INIT_67 => X"0000004f00000000000000000000000000000048000000000000000000000000",
            INIT_68 => X"0000000000000000000000140000000000000000000000000000006700000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000005c00000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000006a00000000",
            INIT_6B => X"0000000000000000000000000000000000000023000000000000000000000000",
            INIT_6C => X"0000008d00000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000200000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000230000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000048000000000000003900000000",
            INIT_74 => X"0000004100000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"00000000000000000000002e0000000000000014000000000000001700000000",
            INIT_77 => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"000000000000000000000000000000000000000000000000000000ca00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000003400000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"000000450000000000000000000000000000000300000000000000a600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE0;


    MEM_IFMAP_LAYER2_INSTANCE1 : if BRAM_NAME = "ifmap_layer2_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"00000107000000000000000c0000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000004f00000000",
            INIT_03 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_04 => X"00000027000000000000002e0000000000000022000000000000000000000000",
            INIT_05 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"00000000000000000000001e000000000000004b000000000000002800000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000970000000000000000000000000000000000000000",
            INIT_0A => X"00000000000000000000004e0000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000106000000000000000000000000",
            INIT_0C => X"00000000000000000000002e0000000000000000000000000000000000000000",
            INIT_0D => X"000000000000000000000000000000000000000000000000000000d800000000",
            INIT_0E => X"0000000000000000000000000000000000000028000000000000006500000000",
            INIT_0F => X"0000007100000000000000b80000000000000000000000000000000000000000",
            INIT_10 => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"000000000000000000000000000000000000014a000000000000002a00000000",
            INIT_12 => X"0000000f000000000000007f000000000000000e000000000000001000000000",
            INIT_13 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_17 => X"0000000000000000000000000000000000000051000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000900000000000000120000000000000000000000000000000000000000",
            INIT_1A => X"0000005a00000000000000060000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000001200000000000000000000000000000000000000000000004f00000000",
            INIT_1D => X"0000000000000000000000000000000000000003000000000000002200000000",
            INIT_1E => X"0000000200000000000000290000000000000023000000000000003c00000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000004900000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"00000000000000000000005c0000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000006100000000",
            INIT_24 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000009500000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000009500000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000001c00000000000000000000000000000038000000000000008300000000",
            INIT_36 => X"0000004d00000000000000830000000000000063000000000000001b00000000",
            INIT_37 => X"0000000000000000000000150000000000000046000000000000004300000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"000000000000000000000000000000000000000a000000000000006b00000000",
            INIT_4F => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000890000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000310000000000000000000000000000000000000000",
            INIT_52 => X"0000007200000000000000340000000000000014000000000000000000000000",
            INIT_53 => X"00000000000000000000000000000000000000a1000000000000000000000000",
            INIT_54 => X"0000000000000000000000c80000000000000000000000000000000000000000",
            INIT_55 => X"000000000000000000000080000000000000005f000000000000009000000000",
            INIT_56 => X"000000000000000000000000000000000000003b000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"00000000000000000000000f0000000000000013000000000000005600000000",
            INIT_5B => X"000000650000000000000069000000000000002b000000000000000000000000",
            INIT_5C => X"0000000000000000000000200000000000000000000000000000001f00000000",
            INIT_5D => X"0000005d00000000000000200000000000000028000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000006c00000000",
            INIT_5F => X"0000007300000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_61 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_63 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_64 => X"00000036000000000000001e0000000000000000000000000000000000000000",
            INIT_65 => X"00000039000000000000000000000000000000d8000000000000009500000000",
            INIT_66 => X"000000a300000000000000910000000000000065000000000000008500000000",
            INIT_67 => X"00000060000000000000005a0000000000000070000000000000010e00000000",
            INIT_68 => X"00000000000000000000004b000000000000007b000000000000006a00000000",
            INIT_69 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000350000000000000000000000000000002300000000",
            INIT_6B => X"000000180000000000000000000000000000001a000000000000005d00000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000b00000000000000000000000000000000000000000000001700000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000001000000000000000000000000000000023000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000007500000000",
            INIT_72 => X"0000002e00000000000000360000000000000052000000000000002700000000",
            INIT_73 => X"0000000000000000000000000000000000000027000000000000002500000000",
            INIT_74 => X"0000002600000000000000000000000000000020000000000000000000000000",
            INIT_75 => X"0000005200000000000000a70000000000000059000000000000004e00000000",
            INIT_76 => X"000000f100000000000000450000000000000059000000000000004b00000000",
            INIT_77 => X"000000d800000000000000800000000000000077000000000000006d00000000",
            INIT_78 => X"0000009c00000000000000bc0000000000000055000000000000009100000000",
            INIT_79 => X"00000078000000000000019a000000000000009d000000000000003e00000000",
            INIT_7A => X"000000da000000000000004e0000000000000037000000000000002400000000",
            INIT_7B => X"0000006e00000000000000640000000000000133000000000000008200000000",
            INIT_7C => X"00000053000000000000007b0000000000000112000000000000004a00000000",
            INIT_7D => X"0000000000000000000000530000000000000000000000000000002e00000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000014000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE1;


    MEM_IFMAP_LAYER2_INSTANCE2 : if BRAM_NAME = "ifmap_layer2_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"00000039000000000000002c0000000000000036000000000000000000000000",
            INIT_02 => X"000000080000000000000000000000000000001f000000000000002b00000000",
            INIT_03 => X"000000000000000000000000000000000000000b000000000000006a00000000",
            INIT_04 => X"0000009100000000000000270000000000000000000000000000002600000000",
            INIT_05 => X"0000005200000000000000000000000000000034000000000000001400000000",
            INIT_06 => X"000000000000000000000035000000000000000c000000000000001900000000",
            INIT_07 => X"00000034000000000000005a0000000000000027000000000000000000000000",
            INIT_08 => X"0000000000000000000000770000000000000018000000000000004d00000000",
            INIT_09 => X"000000080000000000000032000000000000002c000000000000001400000000",
            INIT_0A => X"0000002e000000000000007d0000000000000085000000000000000000000000",
            INIT_0B => X"00000031000000000000004d0000000000000050000000000000003500000000",
            INIT_0C => X"0000003e000000000000004c0000000000000017000000000000003f00000000",
            INIT_0D => X"0000009100000000000000840000000000000065000000000000004800000000",
            INIT_0E => X"000000430000000000000051000000000000002e000000000000009300000000",
            INIT_0F => X"0000007400000000000000ca0000000000000078000000000000005a00000000",
            INIT_10 => X"0000005e0000000000000059000000000000008a000000000000006000000000",
            INIT_11 => X"0000005d000000000000006f000000000000006c000000000000008900000000",
            INIT_12 => X"0000003700000000000000600000000000000055000000000000009c00000000",
            INIT_13 => X"0000006b00000000000000220000000000000020000000000000007800000000",
            INIT_14 => X"000000cf0000000000000022000000000000008b000000000000005900000000",
            INIT_15 => X"0000000000000000000000000000000000000075000000000000005d00000000",
            INIT_16 => X"0000000000000000000000090000000000000000000000000000006e00000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000005700000000000000000000000000000059000000000000000000000000",
            INIT_1B => X"0000004000000000000000900000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000e50000000000000000000000000000000700000000",
            INIT_1D => X"0000002f00000000000000080000000000000025000000000000000000000000",
            INIT_1E => X"00000000000000000000000000000000000001e8000000000000000000000000",
            INIT_1F => X"0000000000000000000000bd0000000000000000000000000000000000000000",
            INIT_20 => X"00000000000000000000002b0000000000000000000000000000010a00000000",
            INIT_21 => X"000000000000000000000000000000000000000000000000000000ec00000000",
            INIT_22 => X"0000018a0000000000000057000000000000009b000000000000000000000000",
            INIT_23 => X"0000006b00000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000e0000000000000000000000000000008a000000000000003300000000",
            INIT_25 => X"0000009300000000000000570000000000000050000000000000001700000000",
            INIT_26 => X"0000005300000000000000000000000000000019000000000000000000000000",
            INIT_27 => X"000000000000000000000000000000000000004d000000000000000000000000",
            INIT_28 => X"0000000000000000000000a5000000000000000d000000000000000000000000",
            INIT_29 => X"00000000000000000000009e000000000000003b00000000000000bd00000000",
            INIT_2A => X"000000f300000000000000000000000000000131000000000000000000000000",
            INIT_2B => X"00000000000000000000000d0000000000000124000000000000004800000000",
            INIT_2C => X"0000000000000000000000b60000000000000000000000000000008900000000",
            INIT_2D => X"00000033000000000000001b000000000000000000000000000000cb00000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000006700000000",
            INIT_2F => X"0000002f000000000000000000000000000000e5000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000031000000000000003500000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000b0000000000000000000000000000002a000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000002e00000000",
            INIT_3A => X"0000000000000000000000720000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000007400000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_3E => X"0000000000000000000000260000000000000000000000000000000000000000",
            INIT_3F => X"000000420000000000000075000000000000009d000000000000000e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002300000000000000000000000000000000000000000000005900000000",
            INIT_41 => X"0000001800000000000000000000000000000000000000000000001a00000000",
            INIT_42 => X"000000000000000000000079000000000000006b000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_44 => X"0000000000000000000000350000000000000053000000000000001e00000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_46 => X"00000062000000000000009a0000000000000021000000000000000c00000000",
            INIT_47 => X"000000e4000000000000002300000000000000c0000000000000003f00000000",
            INIT_48 => X"0000001000000000000000000000000000000018000000000000008400000000",
            INIT_49 => X"0000000000000000000000370000000000000102000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000001700000000000000180000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"000000400000000000000009000000000000003d000000000000001e00000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000007a00000000",
            INIT_51 => X"0000009d00000000000000000000000000000024000000000000000000000000",
            INIT_52 => X"00000010000000000000005a0000000000000016000000000000008900000000",
            INIT_53 => X"000000a700000000000000fe0000000000000000000000000000004800000000",
            INIT_54 => X"0000011600000000000000f500000000000000f800000000000000b900000000",
            INIT_55 => X"00000117000000000000013c0000000000000122000000000000013c00000000",
            INIT_56 => X"000001530000000000000127000000000000011e000000000000010e00000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000004300000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"000000000000000000000087000000000000003c000000000000003200000000",
            INIT_5B => X"0000001f00000000000000a1000000000000001b000000000000000000000000",
            INIT_5C => X"00000000000000000000000b0000000000000057000000000000004100000000",
            INIT_5D => X"0000002e000000000000000000000000000000be000000000000000000000000",
            INIT_5E => X"0000001a0000000000000000000000000000005f000000000000005900000000",
            INIT_5F => X"0000000000000000000000480000000000000000000000000000000000000000",
            INIT_60 => X"0000007c0000000000000000000000000000000000000000000000b900000000",
            INIT_61 => X"0000000000000000000000f2000000000000005400000000000000ac00000000",
            INIT_62 => X"000000b200000000000000c900000000000000ab000000000000005d00000000",
            INIT_63 => X"000000b900000000000000aa000000000000008300000000000000c000000000",
            INIT_64 => X"0000006200000000000000600000000000000062000000000000007300000000",
            INIT_65 => X"0000005800000000000000a300000000000000b800000000000000a900000000",
            INIT_66 => X"000000000000000000000061000000000000001e000000000000006100000000",
            INIT_67 => X"0000007e000000000000000e0000000000000000000000000000008800000000",
            INIT_68 => X"0000006c00000000000000000000000000000039000000000000000400000000",
            INIT_69 => X"0000000000000000000000620000000000000000000000000000006500000000",
            INIT_6A => X"0000002b00000000000000110000000000000000000000000000003d00000000",
            INIT_6B => X"0000006c000000000000001f000000000000000b000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"000000e300000000000000fc0000000000000000000000000000000000000000",
            INIT_70 => X"0000005c000000000000008d00000000000000f0000000000000006b00000000",
            INIT_71 => X"0000007600000000000000c9000000000000004b00000000000000c700000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_77 => X"0000002000000000000000380000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE2;


    MEM_IFMAP_LAYER2_INSTANCE3 : if BRAM_NAME = "ifmap_layer2_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_04 => X"0000001e00000000000001170000000000000000000000000000000000000000",
            INIT_05 => X"0000008c000000000000006500000000000000bd000000000000007a00000000",
            INIT_06 => X"0000008d000000000000011200000000000000c7000000000000009900000000",
            INIT_07 => X"000000cd00000000000000ce000000000000009b000000000000008800000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE3;


    MEM_GOLD_LAYER0_INSTANCE0 : if BRAM_NAME = "gold_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000200000000000000000000000000000000000000000000000500000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000005400000000",
            INIT_06 => X"0000000200000000000000000000000000000002000000000000001b00000000",
            INIT_07 => X"0000000400000000000000000000000000000000000000000000000500000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000004a00000000000000070000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000750000000000000000000000000000001c00000000",
            INIT_0C => X"0000000d000000000000000c0000000000000001000000000000000900000000",
            INIT_0D => X"0000000000000000000000310000000000000000000000000000000000000000",
            INIT_0E => X"0000003600000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000002800000000000000000000000000000054000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000003400000000",
            INIT_11 => X"0000000000000000000000000000000000000058000000000000000000000000",
            INIT_12 => X"0000000000000000000000060000000000000000000000000000000a00000000",
            INIT_13 => X"0000004200000000000000000000000000000000000000000000001f00000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"000000070000000000000000000000000000000000000000000000d900000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000004d00000000000000440000000000000000000000000000000000000000",
            INIT_18 => X"000000a800000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000001b00000000000000040000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000510000000000000016000000000000000000000000",
            INIT_1C => X"0000000000000000000000620000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_1E => X"0000003800000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000120000000000000000000000000000001700000000",
            INIT_21 => X"000000000000000000000012000000000000001d000000000000000600000000",
            INIT_22 => X"0000000000000000000000470000000000000000000000000000000000000000",
            INIT_23 => X"00000000000000000000000e000000000000001a000000000000000000000000",
            INIT_24 => X"0000003400000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000610000000000000000000000000000003700000000",
            INIT_26 => X"00000000000000000000000000000000000000cb000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_28 => X"0000000500000000000000100000000000000024000000000000001700000000",
            INIT_29 => X"00000000000000000000000e000000000000001d000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000009200000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_2D => X"000000000000000000000038000000000000001f000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000d00000000000000090000000000000004000000000000000000000000",
            INIT_30 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_31 => X"000000000000000000000000000000000000004f000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000002900000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000500000000000000080000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000380000000000000000000000000000000000000000",
            INIT_38 => X"000000ab00000000000000ab00000000000000a4000000000000000000000000",
            INIT_39 => X"000000ae00000000000000ac00000000000000a800000000000000ac00000000",
            INIT_3A => X"00000083000000000000009500000000000000a300000000000000ab00000000",
            INIT_3B => X"0000007a000000000000008a0000000000000093000000000000008b00000000",
            INIT_3C => X"000000af00000000000000b000000000000000ab00000000000000a400000000",
            INIT_3D => X"0000009e00000000000000b3000000000000011100000000000000b700000000",
            INIT_3E => X"0000007400000000000000940000000000000095000000000000007000000000",
            INIT_3F => X"0000007800000000000000860000000000000084000000000000006f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ae00000000000000ac00000000000000ad000000000000009a00000000",
            INIT_41 => X"00000054000000000000005e000000000000008e00000000000000ee00000000",
            INIT_42 => X"0000007400000000000000ae00000000000000cd00000000000000e400000000",
            INIT_43 => X"000000aa000000000000006b0000000000000093000000000000005300000000",
            INIT_44 => X"000000b500000000000000ae00000000000000b900000000000000b400000000",
            INIT_45 => X"000000df000000000000007c000000000000007a00000000000000cc00000000",
            INIT_46 => X"000000280000000000000067000000000000009200000000000000d100000000",
            INIT_47 => X"000000bf000000000000013100000000000000e0000000000000008500000000",
            INIT_48 => X"000000f20000000000000123000000000000017d00000000000000fc00000000",
            INIT_49 => X"0000010800000000000000bf000000000000005c000000000000008800000000",
            INIT_4A => X"00000039000000000000004c0000000000000089000000000000008f00000000",
            INIT_4B => X"0000009500000000000000d0000000000000015f00000000000000f400000000",
            INIT_4C => X"000000bc000000000000012e000000000000011f000000000000015c00000000",
            INIT_4D => X"0000008c000000000000011d000000000000012b000000000000006600000000",
            INIT_4E => X"0000010000000000000000480000000000000080000000000000009b00000000",
            INIT_4F => X"000000ee000000000000008000000000000000bb000000000000014400000000",
            INIT_50 => X"0000009100000000000000f70000000000000167000000000000014100000000",
            INIT_51 => X"0000008c00000000000000920000000000000100000000000000015600000000",
            INIT_52 => X"000001610000000000000134000000000000008500000000000000ae00000000",
            INIT_53 => X"0000018300000000000000cd00000000000000be00000000000000c400000000",
            INIT_54 => X"00000123000000000000009200000000000000d8000000000000010f00000000",
            INIT_55 => X"000000ad0000000000000096000000000000009000000000000000f800000000",
            INIT_56 => X"000000c1000000000000018a000000000000016d000000000000009300000000",
            INIT_57 => X"000000bf00000000000000d200000000000000b4000000000000010b00000000",
            INIT_58 => X"000000ad00000000000000c700000000000000c900000000000000b800000000",
            INIT_59 => X"000000ad000000000000009e0000000000000059000000000000005600000000",
            INIT_5A => X"0000012800000000000000ef0000000000000184000000000000018200000000",
            INIT_5B => X"0000012b00000000000000f9000000000000009100000000000000cf00000000",
            INIT_5C => X"000000290000000000000057000000000000009c00000000000000b100000000",
            INIT_5D => X"0000018f00000000000000b300000000000000ce000000000000007d00000000",
            INIT_5E => X"0000019500000000000001b000000000000000fa000000000000017a00000000",
            INIT_5F => X"000000ba000000000000014c000000000000014700000000000000fd00000000",
            INIT_60 => X"000000a7000000000000007e0000000000000061000000000000007000000000",
            INIT_61 => X"00000175000000000000012500000000000000a900000000000000cd00000000",
            INIT_62 => X"000000ae00000000000001770000000000000225000000000000014800000000",
            INIT_63 => X"0000008b000000000000008d00000000000000a900000000000000b200000000",
            INIT_64 => X"000000c900000000000000bb00000000000000ab000000000000009c00000000",
            INIT_65 => X"0000017900000000000000fc00000000000000b600000000000000b900000000",
            INIT_66 => X"0000009b00000000000000a600000000000000ba00000000000001e100000000",
            INIT_67 => X"000000b5000000000000009a0000000000000093000000000000009600000000",
            INIT_68 => X"000000f600000000000000cd00000000000000ce00000000000000c900000000",
            INIT_69 => X"0000016b000000000000013400000000000000ad00000000000000b900000000",
            INIT_6A => X"0000009700000000000000a800000000000000b900000000000000a500000000",
            INIT_6B => X"000000c100000000000000b900000000000000af000000000000009d00000000",
            INIT_6C => X"000000bd00000000000000d200000000000000e000000000000000b900000000",
            INIT_6D => X"0000008100000000000000ce00000000000000b200000000000000b100000000",
            INIT_6E => X"000000bc00000000000000a800000000000000a3000000000000009200000000",
            INIT_6F => X"0000010300000000000000b200000000000000b000000000000000cf00000000",
            INIT_70 => X"000000000000000000000000000000000000009c000000000000010e00000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000033000000000000000000000000",
            INIT_7A => X"00000000000000000000000a0000000000000023000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000090000000000000000000000000000004700000000",
            INIT_7F => X"0000001e00000000000000000000000000000013000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE0;


    MEM_GOLD_LAYER0_INSTANCE1 : if BRAM_NAME = "gold_layer0_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000050000000000000012000000000000000000000000",
            INIT_01 => X"0000002700000000000000000000000000000000000000000000000600000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_03 => X"0000000000000000000000470000000000000011000000000000000000000000",
            INIT_04 => X"0000000a000000000000003a000000000000009c000000000000000400000000",
            INIT_05 => X"0000001200000000000000620000000000000000000000000000000000000000",
            INIT_06 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_07 => X"00000000000000000000000c000000000000002c000000000000000800000000",
            INIT_08 => X"00000000000000000000003f0000000000000038000000000000004800000000",
            INIT_09 => X"0000000000000000000000050000000000000073000000000000000000000000",
            INIT_0A => X"0000001f00000000000000000000000000000004000000000000000000000000",
            INIT_0B => X"0000001000000000000000000000000000000000000000000000002a00000000",
            INIT_0C => X"0000000000000000000000260000000000000018000000000000007a00000000",
            INIT_0D => X"000000110000000000000000000000000000000f000000000000005700000000",
            INIT_0E => X"0000005900000000000000300000000000000000000000000000001700000000",
            INIT_0F => X"000000390000000000000000000000000000002b000000000000000000000000",
            INIT_10 => X"00000000000000000000000e0000000000000000000000000000000700000000",
            INIT_11 => X"00000004000000000000000c0000000000000000000000000000003400000000",
            INIT_12 => X"0000000000000000000000560000000000000052000000000000000000000000",
            INIT_13 => X"0000001c00000000000000000000000000000009000000000000004200000000",
            INIT_14 => X"0000000000000000000000190000000000000008000000000000000600000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"000000800000000000000000000000000000004d000000000000007500000000",
            INIT_17 => X"0000004e00000000000000500000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000008d0000000000000001000000000000001a000000000000000900000000",
            INIT_1A => X"0000005000000000000000940000000000000022000000000000007200000000",
            INIT_1B => X"000000150000000000000038000000000000003b000000000000002900000000",
            INIT_1C => X"0000001e000000000000001d0000000000000013000000000000001000000000",
            INIT_1D => X"00000073000000000000000e000000000000001a000000000000002000000000",
            INIT_1E => X"000000140000000000000009000000000000007a000000000000006d00000000",
            INIT_1F => X"0000000e000000000000000b0000000000000010000000000000001200000000",
            INIT_20 => X"000000290000000000000026000000000000001e000000000000001600000000",
            INIT_21 => X"0000009e000000000000001b0000000000000014000000000000002800000000",
            INIT_22 => X"00000009000000000000001c0000000000000007000000000000004d00000000",
            INIT_23 => X"00000022000000000000001c0000000000000017000000000000001200000000",
            INIT_24 => X"0000003b0000000000000034000000000000001c000000000000002f00000000",
            INIT_25 => X"0000004300000000000000270000000000000023000000000000001100000000",
            INIT_26 => X"0000001500000000000000280000000000000029000000000000000d00000000",
            INIT_27 => X"0000001b00000000000000150000000000000018000000000000001800000000",
            INIT_28 => X"0000000000000000000000000000000000000025000000000000003000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000d00000000000000060000000000000009000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000004000000000000001700000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000300000000000000060000000000000003000000000000000b00000000",
            INIT_37 => X"000000240000000000000000000000000000000a000000000000001100000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"00000008000000000000000e0000000000000005000000000000000000000000",
            INIT_3A => X"0000000a000000000000000a0000000000000006000000000000001500000000",
            INIT_3B => X"00000005000000000000002d0000000000000000000000000000000f00000000",
            INIT_3C => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000400000000000000060000000000000008000000000000000000000000",
            INIT_3E => X"00000014000000000000000b0000000000000017000000000000000600000000",
            INIT_3F => X"000000000000000000000000000000000000003a000000000000001500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"000000140000000000000000000000000000000b000000000000000e00000000",
            INIT_42 => X"000000080000000000000011000000000000000f000000000000001300000000",
            INIT_43 => X"000000000000000000000011000000000000001c000000000000002d00000000",
            INIT_44 => X"00000004000000000000000c0000000000000000000000000000000000000000",
            INIT_45 => X"0000001000000000000000060000000000000000000000000000000d00000000",
            INIT_46 => X"0000002600000000000000000000000000000003000000000000001100000000",
            INIT_47 => X"0000000000000000000000090000000000000025000000000000001d00000000",
            INIT_48 => X"0000000e00000000000000000000000000000008000000000000000700000000",
            INIT_49 => X"0000000b00000000000000110000000000000000000000000000000000000000",
            INIT_4A => X"0000001800000000000000150000000000000000000000000000000000000000",
            INIT_4B => X"0000001100000000000000140000000000000018000000000000001f00000000",
            INIT_4C => X"0000000100000000000000080000000000000005000000000000001800000000",
            INIT_4D => X"000000000000000000000005000000000000001c000000000000000d00000000",
            INIT_4E => X"0000001c00000000000000180000000000000013000000000000000000000000",
            INIT_4F => X"00000010000000000000001b000000000000001e000000000000001d00000000",
            INIT_50 => X"0000003300000000000000230000000000000028000000000000001f00000000",
            INIT_51 => X"0000002600000000000000240000000000000030000000000000003500000000",
            INIT_52 => X"00000000000000000000002a0000000000000031000000000000003400000000",
            INIT_53 => X"00000043000000000000003f000000000000004d000000000000000b00000000",
            INIT_54 => X"0000004d00000000000000490000000000000045000000000000004800000000",
            INIT_55 => X"000000570000000000000053000000000000004e000000000000005300000000",
            INIT_56 => X"000000500000000000000000000000000000003b000000000000003900000000",
            INIT_57 => X"0000004900000000000000480000000000000049000000000000004c00000000",
            INIT_58 => X"0000004f00000000000000540000000000000053000000000000004d00000000",
            INIT_59 => X"0000005800000000000000640000000000000060000000000000005700000000",
            INIT_5A => X"0000004b0000000000000046000000000000001d000000000000003800000000",
            INIT_5B => X"00000051000000000000004e000000000000004a000000000000004c00000000",
            INIT_5C => X"0000005f000000000000005d0000000000000057000000000000005400000000",
            INIT_5D => X"0000004b000000000000005e0000000000000061000000000000005000000000",
            INIT_5E => X"0000004a00000000000000480000000000000044000000000000003e00000000",
            INIT_5F => X"00000051000000000000004f000000000000004a000000000000004e00000000",
            INIT_60 => X"000000610000000000000055000000000000005a000000000000005800000000",
            INIT_61 => X"0000008600000000000000850000000000000086000000000000008100000000",
            INIT_62 => X"00000092000000000000008b0000000000000080000000000000008400000000",
            INIT_63 => X"0000006900000000000000640000000000000072000000000000008600000000",
            INIT_64 => X"0000008000000000000000720000000000000075000000000000006c00000000",
            INIT_65 => X"000000880000000000000088000000000000008d000000000000008b00000000",
            INIT_66 => X"0000005900000000000000780000000000000078000000000000007800000000",
            INIT_67 => X"00000046000000000000002c000000000000001c000000000000003600000000",
            INIT_68 => X"000000710000000000000062000000000000006e000000000000005f00000000",
            INIT_69 => X"00000094000000000000008c000000000000008a000000000000008800000000",
            INIT_6A => X"0000003600000000000000270000000000000035000000000000004100000000",
            INIT_6B => X"000000390000000000000019000000000000001e000000000000002000000000",
            INIT_6C => X"0000007c00000000000000490000000000000015000000000000006100000000",
            INIT_6D => X"0000003900000000000000570000000000000072000000000000008c00000000",
            INIT_6E => X"0000002000000000000000480000000000000018000000000000001f00000000",
            INIT_6F => X"0000005c0000000000000011000000000000000e000000000000002900000000",
            INIT_70 => X"000000850000000000000066000000000000003f000000000000000000000000",
            INIT_71 => X"0000001a000000000000002f0000000000000049000000000000005100000000",
            INIT_72 => X"00000019000000000000002e0000000000000033000000000000001900000000",
            INIT_73 => X"000000030000000000000039000000000000000f000000000000002100000000",
            INIT_74 => X"0000005400000000000000630000000000000059000000000000002d00000000",
            INIT_75 => X"000000100000000000000028000000000000002a000000000000003c00000000",
            INIT_76 => X"0000002900000000000000100000000000000027000000000000005100000000",
            INIT_77 => X"0000001f00000000000000000000000000000010000000000000001700000000",
            INIT_78 => X"0000004000000000000000670000000000000065000000000000004800000000",
            INIT_79 => X"0000005500000000000000170000000000000020000000000000004100000000",
            INIT_7A => X"0000001b0000000000000019000000000000000f000000000000001100000000",
            INIT_7B => X"0000002000000000000000180000000000000006000000000000001e00000000",
            INIT_7C => X"0000002e00000000000000610000000000000055000000000000004000000000",
            INIT_7D => X"0000001b0000000000000062000000000000001a000000000000003000000000",
            INIT_7E => X"00000041000000000000002e0000000000000023000000000000001100000000",
            INIT_7F => X"000000280000000000000000000000000000001f000000000000000b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE1;


    MEM_GOLD_LAYER0_INSTANCE2 : if BRAM_NAME = "gold_layer0_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002100000000000000220000000000000037000000000000002b00000000",
            INIT_01 => X"0000001a0000000000000035000000000000003e000000000000002e00000000",
            INIT_02 => X"00000020000000000000006c0000000000000041000000000000002200000000",
            INIT_03 => X"0000001900000000000000240000000000000000000000000000002100000000",
            INIT_04 => X"0000002700000000000000200000000000000031000000000000003000000000",
            INIT_05 => X"00000029000000000000000f0000000000000018000000000000003600000000",
            INIT_06 => X"000000220000000000000022000000000000006b000000000000006900000000",
            INIT_07 => X"0000000e00000000000000000000000000000044000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000020000000000000002d00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"00000010000000000000000f0000000000000009000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000005900000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000003000000000000000160000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"000000250000000000000024000000000000002a000000000000000000000000",
            INIT_1A => X"0000002a00000000000000230000000000000027000000000000002500000000",
            INIT_1B => X"0000002000000000000000210000000000000023000000000000002a00000000",
            INIT_1C => X"000000210000000000000025000000000000001f000000000000002600000000",
            INIT_1D => X"0000002500000000000000260000000000000027000000000000002a00000000",
            INIT_1E => X"00000022000000000000001b0000000000000020000000000000002300000000",
            INIT_1F => X"00000021000000000000000a000000000000000f000000000000000900000000",
            INIT_20 => X"000000270000000000000026000000000000002b000000000000003100000000",
            INIT_21 => X"0000002c0000000000000025000000000000002c000000000000003100000000",
            INIT_22 => X"0000001200000000000000110000000000000001000000000000003a00000000",
            INIT_23 => X"0000000e0000000000000007000000000000000b000000000000002100000000",
            INIT_24 => X"000000570000000000000000000000000000002d000000000000003600000000",
            INIT_25 => X"0000001000000000000000200000000000000027000000000000003000000000",
            INIT_26 => X"0000003500000000000000150000000000000006000000000000000a00000000",
            INIT_27 => X"0000001e00000000000000020000000000000016000000000000000000000000",
            INIT_28 => X"0000001b000000000000003d0000000000000000000000000000004300000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_2A => X"000000040000000000000028000000000000001a000000000000000100000000",
            INIT_2B => X"0000004300000000000000070000000000000018000000000000000000000000",
            INIT_2C => X"0000001900000000000000100000000000000027000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_2E => X"000000000000000000000000000000000000004f000000000000000900000000",
            INIT_2F => X"00000000000000000000000e0000000000000005000000000000001f00000000",
            INIT_30 => X"0000003b00000000000000020000000000000023000000000000001900000000",
            INIT_31 => X"0000000000000000000000000000000000000004000000000000001200000000",
            INIT_32 => X"0000001c00000000000000020000000000000000000000000000005100000000",
            INIT_33 => X"0000000000000000000000000000000000000015000000000000001300000000",
            INIT_34 => X"0000002c000000000000001c000000000000000c000000000000000e00000000",
            INIT_35 => X"0000004a00000000000000010000000000000011000000000000000000000000",
            INIT_36 => X"00000024000000000000001e0000000000000004000000000000000000000000",
            INIT_37 => X"0000000000000000000000020000000000000000000000000000001c00000000",
            INIT_38 => X"000000070000000000000013000000000000000f000000000000001b00000000",
            INIT_39 => X"00000029000000000000001c0000000000000020000000000000001300000000",
            INIT_3A => X"0000002b00000000000000270000000000000028000000000000000200000000",
            INIT_3B => X"0000002100000000000000000000000000000006000000000000000000000000",
            INIT_3C => X"00000000000000000000000c0000000000000013000000000000000000000000",
            INIT_3D => X"0000000e0000000000000000000000000000000e000000000000002800000000",
            INIT_3E => X"000000230000000000000021000000000000003f000000000000003100000000",
            INIT_3F => X"0000000000000000000000370000000000000000000000000000000400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000019000000000000000000000000",
            INIT_41 => X"0000001d00000000000000090000000000000011000000000000000000000000",
            INIT_42 => X"0000000c00000000000000480000000000000006000000000000001d00000000",
            INIT_43 => X"0000000000000000000000000000000000000039000000000000000000000000",
            INIT_44 => X"0000000900000000000000040000000000000011000000000000001700000000",
            INIT_45 => X"00000013000000000000000a000000000000000f000000000000000f00000000",
            INIT_46 => X"0000001300000000000000440000000000000011000000000000000800000000",
            INIT_47 => X"0000000900000000000000080000000000000000000000000000001700000000",
            INIT_48 => X"0000000e0000000000000010000000000000000f000000000000000e00000000",
            INIT_49 => X"0000000900000000000000040000000000000010000000000000001100000000",
            INIT_4A => X"0000000000000000000000520000000000000013000000000000000200000000",
            INIT_4B => X"0000000f00000000000000050000000000000010000000000000000000000000",
            INIT_4C => X"00000011000000000000000f000000000000000d000000000000000a00000000",
            INIT_4D => X"0000000000000000000000160000000000000015000000000000000500000000",
            INIT_4E => X"0000001100000000000000200000000000000019000000000000000c00000000",
            INIT_4F => X"0000000900000000000000080000000000000011000000000000001d00000000",
            INIT_50 => X"0000000d000000000000000d000000000000000a000000000000000900000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000001200000000000000020000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000005000000000000001200000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"000000010000000000000000000000000000000c000000000000000000000000",
            INIT_5B => X"0000002e000000000000003f000000000000003b000000000000000500000000",
            INIT_5C => X"000000060000000000000000000000000000000b000000000000001c00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_5E => X"0000002600000000000000140000000000000010000000000000000000000000",
            INIT_5F => X"000000210000000000000029000000000000002b000000000000004200000000",
            INIT_60 => X"0000004400000000000000210000000000000004000000000000001300000000",
            INIT_61 => X"0000001200000000000000140000000000000000000000000000000000000000",
            INIT_62 => X"00000029000000000000002b000000000000001e000000000000002c00000000",
            INIT_63 => X"0000001300000000000000270000000000000015000000000000003100000000",
            INIT_64 => X"0000000000000000000000680000000000000046000000000000000f00000000",
            INIT_65 => X"000000310000000000000026000000000000006e000000000000000000000000",
            INIT_66 => X"00000041000000000000004e0000000000000020000000000000001f00000000",
            INIT_67 => X"0000000d00000000000000220000000000000031000000000000002100000000",
            INIT_68 => X"000000000000000000000002000000000000006f000000000000003900000000",
            INIT_69 => X"0000002a00000000000000510000000000000033000000000000003300000000",
            INIT_6A => X"00000028000000000000003b000000000000006c000000000000002300000000",
            INIT_6B => X"00000048000000000000001f0000000000000031000000000000002f00000000",
            INIT_6C => X"0000000b0000000000000000000000000000001e000000000000006200000000",
            INIT_6D => X"0000002000000000000000440000000000000048000000000000006100000000",
            INIT_6E => X"0000003500000000000000300000000000000038000000000000005600000000",
            INIT_6F => X"0000007c00000000000000630000000000000004000000000000003600000000",
            INIT_70 => X"0000003d00000000000000150000000000000042000000000000003b00000000",
            INIT_71 => X"0000002000000000000000290000000000000031000000000000002900000000",
            INIT_72 => X"00000015000000000000002a0000000000000022000000000000003900000000",
            INIT_73 => X"00000048000000000000007a000000000000006f000000000000000000000000",
            INIT_74 => X"0000002d000000000000001b0000000000000036000000000000006300000000",
            INIT_75 => X"0000001f0000000000000026000000000000003a000000000000004000000000",
            INIT_76 => X"000000000000000000000000000000000000001e000000000000001600000000",
            INIT_77 => X"0000007a000000000000004f000000000000006b000000000000008900000000",
            INIT_78 => X"0000007200000000000000680000000000000038000000000000004000000000",
            INIT_79 => X"00000045000000000000003c000000000000002b000000000000003a00000000",
            INIT_7A => X"000000c5000000000000004e0000000000000063000000000000005e00000000",
            INIT_7B => X"000000930000000000000099000000000000004e000000000000008f00000000",
            INIT_7C => X"000000770000000000000087000000000000008b000000000000007c00000000",
            INIT_7D => X"00000096000000000000008e0000000000000085000000000000007600000000",
            INIT_7E => X"000000b100000000000000a70000000000000096000000000000009d00000000",
            INIT_7F => X"00000080000000000000006c00000000000000a5000000000000007700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE2;


    MEM_GOLD_LAYER0_INSTANCE3 : if BRAM_NAME = "gold_layer0_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000087000000000000007f000000000000007f000000000000007f00000000",
            INIT_01 => X"0000009d00000000000000a0000000000000009c000000000000009300000000",
            INIT_02 => X"000000b1000000000000009c00000000000000ac00000000000000a900000000",
            INIT_03 => X"00000082000000000000008a000000000000006e00000000000000a600000000",
            INIT_04 => X"000000a100000000000000910000000000000084000000000000008200000000",
            INIT_05 => X"000000c200000000000000b700000000000000a300000000000000ac00000000",
            INIT_06 => X"000000a5000000000000009b00000000000000a700000000000000aa00000000",
            INIT_07 => X"00000083000000000000008f0000000000000091000000000000008200000000",
            INIT_08 => X"0000009900000000000000970000000000000095000000000000008600000000",
            INIT_09 => X"00000078000000000000009900000000000000bd00000000000000a400000000",
            INIT_0A => X"0000007e000000000000007f000000000000007b000000000000007b00000000",
            INIT_0B => X"00000082000000000000008b000000000000007c000000000000007600000000",
            INIT_0C => X"0000006100000000000000560000000000000053000000000000006500000000",
            INIT_0D => X"00000081000000000000007a0000000000000073000000000000006e00000000",
            INIT_0E => X"00000061000000000000007f0000000000000081000000000000007e00000000",
            INIT_0F => X"0000003200000000000000500000000000000063000000000000006f00000000",
            INIT_10 => X"00000050000000000000002f0000000000000020000000000000001d00000000",
            INIT_11 => X"0000008100000000000000500000000000000047000000000000006900000000",
            INIT_12 => X"0000004e00000000000000670000000000000083000000000000008500000000",
            INIT_13 => X"0000001d0000000000000013000000000000002a000000000000003900000000",
            INIT_14 => X"0000004d0000000000000029000000000000001d000000000000001e00000000",
            INIT_15 => X"0000007f00000000000000730000000000000021000000000000003100000000",
            INIT_16 => X"0000002900000000000000320000000000000053000000000000006700000000",
            INIT_17 => X"000000230000000000000029000000000000001a000000000000001a00000000",
            INIT_18 => X"000000280000000000000031000000000000001f000000000000002200000000",
            INIT_19 => X"0000002b00000000000000690000000000000067000000000000000c00000000",
            INIT_1A => X"0000001800000000000000250000000000000029000000000000003100000000",
            INIT_1B => X"0000001c000000000000002a0000000000000028000000000000001d00000000",
            INIT_1C => X"0000000600000000000000220000000000000022000000000000002000000000",
            INIT_1D => X"0000003600000000000000150000000000000068000000000000006600000000",
            INIT_1E => X"00000004000000000000001e000000000000002f000000000000002700000000",
            INIT_1F => X"0000001e00000000000000190000000000000029000000000000002400000000",
            INIT_20 => X"0000003e0000000000000000000000000000002b000000000000001d00000000",
            INIT_21 => X"0000001c00000000000000270000000000000028000000000000006d00000000",
            INIT_22 => X"0000002700000000000000000000000000000025000000000000002800000000",
            INIT_23 => X"00000026000000000000001a0000000000000019000000000000002200000000",
            INIT_24 => X"0000003b0000000000000022000000000000000c000000000000001d00000000",
            INIT_25 => X"0000001e0000000000000026000000000000000e000000000000004300000000",
            INIT_26 => X"00000026000000000000002b0000000000000022000000000000002d00000000",
            INIT_27 => X"00000012000000000000004f000000000000001e000000000000001600000000",
            INIT_28 => X"00000031000000000000000c000000000000001c000000000000000000000000",
            INIT_29 => X"0000001d000000000000001f0000000000000032000000000000002900000000",
            INIT_2A => X"0000001c00000000000000280000000000000029000000000000003400000000",
            INIT_2B => X"0000000c0000000000000016000000000000005c000000000000003b00000000",
            INIT_2C => X"0000002300000000000000180000000000000000000000000000001600000000",
            INIT_2D => X"00000025000000000000001d0000000000000018000000000000002100000000",
            INIT_2E => X"00000040000000000000000c0000000000000014000000000000001b00000000",
            INIT_2F => X"00000016000000000000000f0000000000000000000000000000005e00000000",
            INIT_30 => X"00000000000000000000000a0000000000000014000000000000000000000000",
            INIT_31 => X"0000000000000000000000040000000000000001000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000040000000000000000000000000000000500000000",
            INIT_43 => X"0000000000000000000000030000000000000001000000000000000000000000",
            INIT_44 => X"0000001100000000000000020000000000000000000000000000000000000000",
            INIT_45 => X"0000000200000000000000000000000000000000000000000000000400000000",
            INIT_46 => X"0000000800000000000000000000000000000005000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000001600000000000000000000000000000000000000000000001500000000",
            INIT_49 => X"0000004400000000000000000000000000000000000000000000001c00000000",
            INIT_4A => X"0000001c00000000000000080000000000000000000000000000000400000000",
            INIT_4B => X"0000003d00000000000000090000000000000000000000000000000000000000",
            INIT_4C => X"0000002400000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"00000000000000000000005f0000000000000000000000000000002200000000",
            INIT_4E => X"0000000000000000000000160000000000000000000000000000000800000000",
            INIT_4F => X"00000000000000000000006d0000000000000000000000000000000000000000",
            INIT_50 => X"0000005f00000000000000000000000000000000000000000000000200000000",
            INIT_51 => X"000000520000000000000000000000000000001c000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000086000000000000000000000000",
            INIT_54 => X"0000000000000000000000330000000000000000000000000000000000000000",
            INIT_55 => X"0000007600000000000000190000000000000000000000000000001800000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_57 => X"000000130000000000000000000000000000000000000000000000d200000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"00000040000000000000005f0000000000000000000000000000000f00000000",
            INIT_5A => X"000000b100000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"00000010000000000000000b0000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"000000000000000000000054000000000000003d000000000000000000000000",
            INIT_5E => X"0000000000000000000000740000000000000000000000000000000500000000",
            INIT_5F => X"00000000000000000000000f0000000000000025000000000000000000000000",
            INIT_60 => X"0000003100000000000000000000000000000007000000000000000000000000",
            INIT_61 => X"000000000000000000000000000000000000002e000000000000000000000000",
            INIT_62 => X"0000000000000000000000200000000000000000000000000000002700000000",
            INIT_63 => X"00000000000000000000000b0000000000000025000000000000002b00000000",
            INIT_64 => X"0000000000000000000000550000000000000000000000000000000d00000000",
            INIT_65 => X"0000000000000000000000000000000000000034000000000000000c00000000",
            INIT_66 => X"0000002f00000000000000040000000000000000000000000000000300000000",
            INIT_67 => X"00000005000000000000005a0000000000000000000000000000002900000000",
            INIT_68 => X"00000000000000000000000000000000000000aa000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000003e00000000",
            INIT_6A => X"0000001f00000000000000160000000000000006000000000000000000000000",
            INIT_6B => X"00000000000000000000004c0000000000000075000000000000000000000000",
            INIT_6C => X"0000001f00000000000000000000000000000000000000000000007a00000000",
            INIT_6D => X"0000000c00000000000000080000000000000000000000000000001a00000000",
            INIT_6E => X"00000000000000000000000d000000000000000c000000000000001000000000",
            INIT_6F => X"0000000000000000000000840000000000000071000000000000000000000000",
            INIT_70 => X"0000000600000000000000000000000000000002000000000000000000000000",
            INIT_71 => X"00000008000000000000000d0000000000000009000000000000000200000000",
            INIT_72 => X"00000000000000000000000e000000000000000f000000000000000600000000",
            INIT_73 => X"00000000000000000000000000000000000000bd000000000000001100000000",
            INIT_74 => X"0000000e00000000000000010000000000000000000000000000000c00000000",
            INIT_75 => X"000000040000000000000010000000000000000b000000000000000b00000000",
            INIT_76 => X"0000000c00000000000000000000000000000000000000000000002000000000",
            INIT_77 => X"0000002500000000000000000000000000000007000000000000002300000000",
            INIT_78 => X"00000000000000000000000b0000000000000006000000000000001800000000",
            INIT_79 => X"00000000000000000000002d000000000000000f000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000002500000000000000160000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000004000000000000001c00000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000e00000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE3;


    MEM_GOLD_LAYER0_INSTANCE4 : if BRAM_NAME = "gold_layer0_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000000000000c000000000000004500000000",
            INIT_01 => X"0000002700000000000000000000000000000018000000000000001d00000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_03 => X"00000001000000000000002b0000000000000025000000000000004e00000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000006000000000000001e00000000",
            INIT_06 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"00000000000000000000000a0000000000000010000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_0B => X"0000000000000000000000070000000000000009000000000000000000000000",
            INIT_0C => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000002900000000000000000000000000000000000000000000000a00000000",
            INIT_0E => X"0000000000000000000000000000000000000022000000000000006400000000",
            INIT_0F => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_11 => X"000000280000000000000000000000000000001a000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000600000000000000050000000000000000000000000000000000000000",
            INIT_16 => X"000000050000000000000000000000000000002b000000000000002000000000",
            INIT_17 => X"00000007000000000000000b0000000000000000000000000000000100000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000600000000000000540000000000000000000000000000000000000000",
            INIT_1A => X"0000003100000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"000000000000000000000000000000000000001f000000000000003a00000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_1D => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_1E => X"0000001a0000000000000037000000000000003f000000000000000000000000",
            INIT_1F => X"0000001000000000000000050000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"00000008000000000000002f0000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"000000320000000000000065000000000000002b000000000000002700000000",
            INIT_24 => X"0000006800000000000000500000000000000000000000000000000000000000",
            INIT_25 => X"00000013000000000000001e0000000000000043000000000000004600000000",
            INIT_26 => X"0000000000000000000000000000000000000009000000000000000500000000",
            INIT_27 => X"0000001900000000000000490000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000056000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_2B => X"0000004100000000000000510000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_2D => X"0000001300000000000000060000000000000000000000000000000200000000",
            INIT_2E => X"0000000000000000000000260000000000000000000000000000000800000000",
            INIT_2F => X"0000001f000000000000004e000000000000000b000000000000000000000000",
            INIT_30 => X"0000000000000000000000010000000000000024000000000000002400000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"000000a600000000000000a80000000000000000000000000000000000000000",
            INIT_33 => X"000000a400000000000000ad00000000000000ad00000000000000af00000000",
            INIT_34 => X"0000009100000000000000aa00000000000000b700000000000000b800000000",
            INIT_35 => X"00000096000000000000008f0000000000000086000000000000007b00000000",
            INIT_36 => X"000000b500000000000000b300000000000000ab000000000000008a00000000",
            INIT_37 => X"000000b300000000000000c400000000000000b400000000000000b200000000",
            INIT_38 => X"0000004f0000000000000057000000000000006400000000000000a000000000",
            INIT_39 => X"000000920000000000000080000000000000005d000000000000005200000000",
            INIT_3A => X"000000b100000000000000b6000000000000008d000000000000007200000000",
            INIT_3B => X"000000350000000000000054000000000000008b00000000000000b600000000",
            INIT_3C => X"0000003b00000000000000460000000000000065000000000000004100000000",
            INIT_3D => X"0000002a00000000000000850000000000000051000000000000003500000000",
            INIT_3E => X"000000a200000000000000b700000000000000b9000000000000009400000000",
            INIT_3F => X"00000034000000000000003f0000000000000071000000000000007f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000014000000000000003d0000000000000043000000000000006900000000",
            INIT_41 => X"000000a3000000000000002f0000000000000076000000000000001e00000000",
            INIT_42 => X"000000ac00000000000000c600000000000000bf00000000000000ad00000000",
            INIT_43 => X"00000063000000000000001c0000000000000036000000000000005a00000000",
            INIT_44 => X"0000001f000000000000003b0000000000000040000000000000006900000000",
            INIT_45 => X"000000a400000000000000770000000000000039000000000000004f00000000",
            INIT_46 => X"0000006800000000000000670000000000000057000000000000008400000000",
            INIT_47 => X"0000006200000000000000ac0000000000000021000000000000004900000000",
            INIT_48 => X"0000002f000000000000002c000000000000003e000000000000001f00000000",
            INIT_49 => X"00000077000000000000007c000000000000005a000000000000004400000000",
            INIT_4A => X"0000005d000000000000007b0000000000000095000000000000006e00000000",
            INIT_4B => X"0000002e000000000000003d000000000000009e000000000000002400000000",
            INIT_4C => X"0000005c00000000000000420000000000000043000000000000003500000000",
            INIT_4D => X"00000080000000000000007c0000000000000069000000000000005400000000",
            INIT_4E => X"0000002a0000000000000041000000000000004700000000000000ae00000000",
            INIT_4F => X"000000380000000000000022000000000000003e000000000000008f00000000",
            INIT_50 => X"0000006d000000000000005a0000000000000058000000000000004b00000000",
            INIT_51 => X"0000003600000000000000740000000000000065000000000000002b00000000",
            INIT_52 => X"00000064000000000000005f0000000000000048000000000000003b00000000",
            INIT_53 => X"0000005e00000000000000220000000000000004000000000000004400000000",
            INIT_54 => X"000000220000000000000069000000000000005a00000000000000a300000000",
            INIT_55 => X"000000630000000000000053000000000000004b000000000000005e00000000",
            INIT_56 => X"0000000800000000000000400000000000000059000000000000006a00000000",
            INIT_57 => X"0000009400000000000000a7000000000000004c000000000000000800000000",
            INIT_58 => X"000000b3000000000000001f0000000000000074000000000000006d00000000",
            INIT_59 => X"0000004d00000000000000850000000000000077000000000000007c00000000",
            INIT_5A => X"0000002000000000000000110000000000000015000000000000001f00000000",
            INIT_5B => X"00000024000000000000002d000000000000003c000000000000002900000000",
            INIT_5C => X"0000002200000000000000de0000000000000059000000000000004f00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"000000000000000000000000000000000000008d000000000000006f00000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000005a00000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000c00000000000000000000000000000000000000000000000900000000",
            INIT_6B => X"0000000e0000000000000011000000000000000b000000000000001100000000",
            INIT_6C => X"0000000d0000000000000011000000000000000d000000000000000900000000",
            INIT_6D => X"000000090000000000000003000000000000000e000000000000000d00000000",
            INIT_6E => X"0000000900000000000000060000000000000013000000000000000f00000000",
            INIT_6F => X"0000000000000000000000070000000000000014000000000000000800000000",
            INIT_70 => X"0000000000000000000000270000000000000009000000000000002100000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_72 => X"0000000900000000000000000000000000000013000000000000000b00000000",
            INIT_73 => X"0000003a000000000000000e0000000000000007000000000000001200000000",
            INIT_74 => X"0000003100000000000000000000000000000000000000000000001000000000",
            INIT_75 => X"000000000000000000000000000000000000002e000000000000002600000000",
            INIT_76 => X"00000001000000000000000a0000000000000000000000000000005e00000000",
            INIT_77 => X"0000002700000000000000140000000000000000000000000000000f00000000",
            INIT_78 => X"0000001a00000000000000540000000000000000000000000000001500000000",
            INIT_79 => X"0000007d00000000000000000000000000000013000000000000003500000000",
            INIT_7A => X"0000001800000000000000000000000000000037000000000000000000000000",
            INIT_7B => X"0000002200000000000000390000000000000052000000000000002800000000",
            INIT_7C => X"0000000700000000000000490000000000000023000000000000000000000000",
            INIT_7D => X"00000009000000000000006c0000000000000000000000000000002d00000000",
            INIT_7E => X"0000004c0000000000000000000000000000001b000000000000004e00000000",
            INIT_7F => X"000000000000000000000040000000000000003b000000000000005100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE4;


    MEM_GOLD_LAYER0_INSTANCE5 : if BRAM_NAME = "gold_layer0_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000270000000000000000000000000000005f000000000000006b00000000",
            INIT_01 => X"00000013000000000000003f0000000000000068000000000000001400000000",
            INIT_02 => X"0000004100000000000000000000000000000000000000000000004700000000",
            INIT_03 => X"0000007900000000000000000000000000000059000000000000004a00000000",
            INIT_04 => X"0000002800000000000000000000000000000002000000000000003900000000",
            INIT_05 => X"000000210000000000000023000000000000004e000000000000005700000000",
            INIT_06 => X"0000003200000000000000900000000000000000000000000000000000000000",
            INIT_07 => X"00000045000000000000005a0000000000000000000000000000004200000000",
            INIT_08 => X"00000065000000000000002c0000000000000013000000000000000000000000",
            INIT_09 => X"0000001d0000000000000000000000000000007d000000000000002400000000",
            INIT_0A => X"00000000000000000000000f0000000000000031000000000000002600000000",
            INIT_0B => X"00000000000000000000005b0000000000000000000000000000002800000000",
            INIT_0C => X"0000003000000000000000460000000000000000000000000000000000000000",
            INIT_0D => X"0000001500000000000000440000000000000000000000000000008f00000000",
            INIT_0E => X"0000002d0000000000000015000000000000002f000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000007000000000000005400000000",
            INIT_10 => X"00000089000000000000002c0000000000000000000000000000001700000000",
            INIT_11 => X"000000000000000000000023000000000000008d000000000000000000000000",
            INIT_12 => X"0000000000000000000000280000000000000069000000000000004e00000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"000000000000000000000054000000000000000c000000000000000000000000",
            INIT_15 => X"000000110000000000000010000000000000006400000000000000c200000000",
            INIT_16 => X"0000000800000000000000080000000000000009000000000000001c00000000",
            INIT_17 => X"00000021000000000000001b000000000000000f000000000000000c00000000",
            INIT_18 => X"000000b600000000000000410000000000000000000000000000000000000000",
            INIT_19 => X"000000110000000000000011000000000000001a000000000000001400000000",
            INIT_1A => X"0000001500000000000000030000000000000004000000000000000800000000",
            INIT_1B => X"0000000600000000000000310000000000000003000000000000001700000000",
            INIT_1C => X"0000000b00000000000000410000000000000091000000000000000000000000",
            INIT_1D => X"0000000c000000000000000e0000000000000010000000000000002000000000",
            INIT_1E => X"00000000000000000000001f0000000000000014000000000000001200000000",
            INIT_1F => X"0000000700000000000000110000000000000040000000000000003700000000",
            INIT_20 => X"000000150000000000000000000000000000001f000000000000001d00000000",
            INIT_21 => X"000000220000000000000011000000000000000b000000000000001a00000000",
            INIT_22 => X"00000050000000000000002f0000000000000000000000000000001000000000",
            INIT_23 => X"00000053000000000000004b0000000000000053000000000000004d00000000",
            INIT_24 => X"000000550000000000000054000000000000004a000000000000004f00000000",
            INIT_25 => X"000000400000000000000047000000000000004a000000000000004e00000000",
            INIT_26 => X"0000004a0000000000000049000000000000004b000000000000004800000000",
            INIT_27 => X"000000490000000000000058000000000000004a000000000000004f00000000",
            INIT_28 => X"00000054000000000000004f0000000000000068000000000000004c00000000",
            INIT_29 => X"0000002600000000000000340000000000000041000000000000002c00000000",
            INIT_2A => X"00000032000000000000004f0000000000000048000000000000003a00000000",
            INIT_2B => X"00000049000000000000004b0000000000000057000000000000005200000000",
            INIT_2C => X"00000009000000000000001f0000000000000040000000000000007c00000000",
            INIT_2D => X"0000001700000000000000530000000000000050000000000000006200000000",
            INIT_2E => X"0000005b0000000000000000000000000000008e000000000000003600000000",
            INIT_2F => X"00000056000000000000002f0000000000000059000000000000004700000000",
            INIT_30 => X"0000008e0000000000000000000000000000003a000000000000004500000000",
            INIT_31 => X"000000000000000000000036000000000000005c000000000000004300000000",
            INIT_32 => X"000000040000000000000082000000000000002500000000000000b200000000",
            INIT_33 => X"00000065000000000000008f0000000000000053000000000000007a00000000",
            INIT_34 => X"00000075000000000000006a0000000000000000000000000000004500000000",
            INIT_35 => X"0000009400000000000000000000000000000050000000000000003200000000",
            INIT_36 => X"00000044000000000000003b00000000000000a1000000000000006800000000",
            INIT_37 => X"0000006c000000000000006d00000000000000aa000000000000008900000000",
            INIT_38 => X"00000029000000000000008b00000000000000a9000000000000000000000000",
            INIT_39 => X"0000009500000000000000950000000000000036000000000000004a00000000",
            INIT_3A => X"0000003800000000000000000000000000000086000000000000006f00000000",
            INIT_3B => X"00000000000000000000008a0000000000000089000000000000009700000000",
            INIT_3C => X"0000002f000000000000002b000000000000006b00000000000000be00000000",
            INIT_3D => X"0000005600000000000000a40000000000000095000000000000005600000000",
            INIT_3E => X"000000be000000000000002a0000000000000009000000000000007700000000",
            INIT_3F => X"000000990000000000000000000000000000007b000000000000006700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005a0000000000000041000000000000001c000000000000007700000000",
            INIT_41 => X"0000004200000000000000b2000000000000007900000000000000ad00000000",
            INIT_42 => X"0000004d00000000000000740000000000000050000000000000005600000000",
            INIT_43 => X"00000077000000000000003e000000000000005c000000000000002900000000",
            INIT_44 => X"00000097000000000000003b0000000000000032000000000000001600000000",
            INIT_45 => X"0000008d000000000000000e00000000000000d6000000000000007a00000000",
            INIT_46 => X"0000003f0000000000000080000000000000002b000000000000002c00000000",
            INIT_47 => X"000000030000000000000021000000000000006d000000000000005d00000000",
            INIT_48 => X"0000007f0000000000000042000000000000005f000000000000002600000000",
            INIT_49 => X"0000006000000000000000ec000000000000000000000000000000ce00000000",
            INIT_4A => X"0000004a000000000000009d0000000000000092000000000000002300000000",
            INIT_4B => X"00000028000000000000000f000000000000000d000000000000001500000000",
            INIT_4C => X"0000009d00000000000000600000000000000006000000000000004300000000",
            INIT_4D => X"0000003f000000000000009e0000000000000111000000000000001600000000",
            INIT_4E => X"00000029000000000000002a000000000000004a000000000000004300000000",
            INIT_4F => X"0000004000000000000000300000000000000030000000000000002700000000",
            INIT_50 => X"000000ac00000000000000270000000000000001000000000000004300000000",
            INIT_51 => X"0000002f0000000000000036000000000000003600000000000000e100000000",
            INIT_52 => X"0000002800000000000000230000000000000025000000000000002e00000000",
            INIT_53 => X"0000005400000000000000300000000000000036000000000000003700000000",
            INIT_54 => X"0000006600000000000000f30000000000000000000000000000002a00000000",
            INIT_55 => X"00000028000000000000002f0000000000000042000000000000002b00000000",
            INIT_56 => X"0000003e0000000000000037000000000000002d000000000000002900000000",
            INIT_57 => X"0000002f000000000000005e0000000000000057000000000000001800000000",
            INIT_58 => X"0000001e000000000000003a0000000000000055000000000000002b00000000",
            INIT_59 => X"0000003600000000000000290000000000000038000000000000003200000000",
            INIT_5A => X"000000570000000000000014000000000000002b000000000000004100000000",
            INIT_5B => X"0000003b0000000000000034000000000000003a000000000000006f00000000",
            INIT_5C => X"0000004200000000000000340000000000000039000000000000003800000000",
            INIT_5D => X"0000002f000000000000002f0000000000000039000000000000004600000000",
            INIT_5E => X"0000002c00000000000000320000000000000032000000000000003400000000",
            INIT_5F => X"0000003b000000000000003a000000000000003b000000000000004000000000",
            INIT_60 => X"000000370000000000000039000000000000001f000000000000003700000000",
            INIT_61 => X"000000080000000000000000000000000000000c000000000000002700000000",
            INIT_62 => X"0000002400000000000000300000000000000037000000000000002300000000",
            INIT_63 => X"0000003c00000000000000400000000000000041000000000000004f00000000",
            INIT_64 => X"0000000100000000000000130000000000000025000000000000001100000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000001c0000000000000000000000000000002e000000000000001a00000000",
            INIT_67 => X"0000001f000000000000002e000000000000003d000000000000004400000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000003800000000000000000000000000000000000000000000002500000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"00000002000000000000003d0000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"00000000000000000000001c0000000000000047000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000022000000000000000400000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000001a00000000000000030000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE5;


    MEM_GOLD_LAYER0_INSTANCE6 : if BRAM_NAME = "gold_layer0_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000031000000000000001b000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000002400000000000000240000000000000000000000000000000000000000",
            INIT_14 => X"0000001c000000000000001f000000000000001e000000000000002000000000",
            INIT_15 => X"0000002400000000000000200000000000000029000000000000002700000000",
            INIT_16 => X"00000021000000000000001e0000000000000029000000000000002d00000000",
            INIT_17 => X"00000021000000000000001d000000000000001f000000000000001e00000000",
            INIT_18 => X"0000001d00000000000000000000000000000017000000000000002100000000",
            INIT_19 => X"000000000000000000000000000000000000003d000000000000002800000000",
            INIT_1A => X"00000019000000000000001d0000000000000023000000000000000700000000",
            INIT_1B => X"00000023000000000000001f0000000000000031000000000000003b00000000",
            INIT_1C => X"0000002200000000000000330000000000000042000000000000002400000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"000000000000000000000014000000000000001e000000000000000000000000",
            INIT_1F => X"0000001b000000000000001a0000000000000019000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000d0000000000000015000000000000000a000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000014000000000000001100000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_24 => X"0000000000000000000000180000000000000006000000000000000900000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000001e00000000000000000000000000000008000000000000002200000000",
            INIT_27 => X"00000000000000000000001f000000000000002b000000000000004400000000",
            INIT_28 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_2A => X"00000020000000000000002b0000000000000002000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_2C => X"00000000000000000000000c0000000000000000000000000000000100000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000a00000000000000250000000000000032000000000000000000000000",
            INIT_30 => X"00000000000000000000000d000000000000000d000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000013000000000000001000000000",
            INIT_32 => X"0000003800000000000000080000000000000000000000000000000c00000000",
            INIT_33 => X"0000001e00000000000000000000000000000000000000000000000d00000000",
            INIT_34 => X"000000000000000000000018000000000000003d000000000000001500000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_36 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_37 => X"000000330000000000000028000000000000000e000000000000000000000000",
            INIT_38 => X"0000001e00000000000000000000000000000000000000000000000700000000",
            INIT_39 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_3A => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_3C => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000004700000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"00000000000000000000000d0000000000000012000000000000002e00000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000100000000000000120000000000000017000000000000000700000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"00000000000000000000001c000000000000000e000000000000000000000000",
            INIT_52 => X"0000000c000000000000000d0000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000290000000000000022000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"00000004000000000000000e0000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_5A => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_5F => X"0000000900000000000000150000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_62 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"000000060000000000000014000000000000001d000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_6A => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"00000000000000000000000c0000000000000005000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000001400000000000000040000000000000000000000000000000000000000",
            INIT_6F => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000070000000000000000000000000000001600000000",
            INIT_71 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_72 => X"0000002f00000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000023000000000000002e00000000",
            INIT_74 => X"0000001b00000000000000190000000000000005000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000021000000000000002d00000000",
            INIT_76 => X"000000000000000000000000000000000000000e000000000000001500000000",
            INIT_77 => X"0000000000000000000000010000000000000002000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"00000003000000000000000b000000000000000b000000000000001c00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"000000000000000000000003000000000000001f000000000000003100000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE6;


    MEM_GOLD_LAYER0_INSTANCE7 : if BRAM_NAME = "gold_layer0_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_01 => X"0000000a00000000000000030000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE7;


    MEM_GOLD_LAYER1_INSTANCE0 : if BRAM_NAME = "gold_layer1_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_01 => X"000000d500000000000000040000000000000000000000000000002000000000",
            INIT_02 => X"0000006100000000000000080000000000000000000000000000002c00000000",
            INIT_03 => X"0000002a0000000000000042000000000000002a000000000000000700000000",
            INIT_04 => X"0000001e00000000000001540000000000000000000000000000000000000000",
            INIT_05 => X"00000000000000000000004e0000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000042000000000000002800000000",
            INIT_07 => X"00000000000000000000001e0000000000000140000000000000000000000000",
            INIT_08 => X"000000000000000000000000000000000000004c000000000000000000000000",
            INIT_09 => X"0000004200000000000000000000000000000032000000000000000000000000",
            INIT_0A => X"0000000000000000000000180000000000000000000000000000000f00000000",
            INIT_0B => X"000000040000000000000004000000000000000c000000000000003c00000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"000000020000000000000000000000000000007a000000000000007b00000000",
            INIT_0E => X"0000002900000000000000000000000000000000000000000000003b00000000",
            INIT_0F => X"0000000000000000000000760000000000000010000000000000000000000000",
            INIT_10 => X"0000007400000000000000000000000000000000000000000000007a00000000",
            INIT_11 => X"0000003000000000000000000000000000000000000000000000008400000000",
            INIT_12 => X"000000c700000000000000000000000000000067000000000000000000000000",
            INIT_13 => X"0000000f00000000000000a20000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000af000000000000005f000000000000000000000000",
            INIT_15 => X"00000021000000000000016d0000000000000000000000000000000000000000",
            INIT_16 => X"0000008b00000000000000000000000000000000000000000000004900000000",
            INIT_17 => X"0000000000000000000000190000000000000078000000000000000000000000",
            INIT_18 => X"0000003e00000000000000470000000000000000000000000000000400000000",
            INIT_19 => X"0000005d0000000000000044000000000000003c000000000000004a00000000",
            INIT_1A => X"00000067000000000000005b0000000000000068000000000000007500000000",
            INIT_1B => X"000000700000000000000067000000000000002d000000000000005a00000000",
            INIT_1C => X"0000005d000000000000004d000000000000003c000000000000004200000000",
            INIT_1D => X"000000000000000000000056000000000000004c000000000000000000000000",
            INIT_1E => X"00000035000000000000005c0000000000000012000000000000002800000000",
            INIT_1F => X"0000001000000000000000000000000000000092000000000000007300000000",
            INIT_20 => X"0000002800000000000000260000000000000032000000000000003c00000000",
            INIT_21 => X"0000000000000000000000000000000000000002000000000000007000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"000000000000000000000000000000000000001b000000000000000000000000",
            INIT_24 => X"0000003600000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000045000000000000007100000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000002a0000000000000000000000000000001f000000000000001200000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000001b00000000000000000000000000000000000000000000000e00000000",
            INIT_2A => X"0000001a00000000000000010000000000000000000000000000000000000000",
            INIT_2B => X"00000000000000000000004d0000000000000036000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"00000103000000000000000000000000000000b0000000000000000000000000",
            INIT_33 => X"0000000e00000000000000420000000000000077000000000000000000000000",
            INIT_34 => X"0000015000000000000000b50000000000000135000000000000004700000000",
            INIT_35 => X"0000005d0000000000000064000000000000003c000000000000000000000000",
            INIT_36 => X"0000000000000000000000390000000000000029000000000000000000000000",
            INIT_37 => X"000000000000000000000027000000000000013a000000000000000000000000",
            INIT_38 => X"00000000000000000000010f0000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000180000000000000010000000000000005300000000",
            INIT_3A => X"0000000000000000000000000000000000000062000000000000014500000000",
            INIT_3B => X"0000000000000000000001d40000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_3D => X"000000460000000000000086000000000000003c000000000000001c00000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_3F => X"0000001d00000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000700000000000000000000000000000032000000000000000000000000",
            INIT_41 => X"000000000000000000000040000000000000000e000000000000000000000000",
            INIT_42 => X"00000000000000000000001b0000000000000000000000000000004e00000000",
            INIT_43 => X"0000003400000000000000000000000000000069000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000031000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_4D => X"0000005500000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000005500000000000000000000000000000044000000000000000000000000",
            INIT_4F => X"0000000000000000000000270000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000540000000000000000000000000000002e00000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000003600000000",
            INIT_52 => X"000000c000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000039000000000000000000000000",
            INIT_54 => X"0000003800000000000000620000000000000000000000000000005d00000000",
            INIT_55 => X"0000000000000000000000450000000000000003000000000000002b00000000",
            INIT_56 => X"0000004400000000000000010000000000000025000000000000000000000000",
            INIT_57 => X"0000007500000000000000030000000000000000000000000000004600000000",
            INIT_58 => X"0000001000000000000000000000000000000030000000000000007300000000",
            INIT_59 => X"0000004d00000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000004400000000000000040000000000000000000000000000008600000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000008400000000",
            INIT_5C => X"0000005800000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"000000000000000000000092000000000000000c000000000000007400000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000006900000000000000100000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000005300000000",
            INIT_61 => X"0000000000000000000000000000000000000015000000000000000900000000",
            INIT_62 => X"0000008d00000000000000000000000000000005000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000200000000000000029000000000000000000000000",
            INIT_65 => X"0000000000000000000000010000000000000000000000000000004900000000",
            INIT_66 => X"0000006900000000000000000000000000000061000000000000000000000000",
            INIT_67 => X"0000004f00000000000000000000000000000048000000000000000000000000",
            INIT_68 => X"0000000000000000000000140000000000000000000000000000006700000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000005c00000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000006a00000000",
            INIT_6B => X"0000000000000000000000000000000000000023000000000000000000000000",
            INIT_6C => X"0000008d00000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000200000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000230000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000048000000000000003900000000",
            INIT_74 => X"0000004100000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"00000000000000000000002e0000000000000014000000000000001700000000",
            INIT_77 => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"000000000000000000000000000000000000000000000000000000ca00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000003400000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"000000450000000000000000000000000000000300000000000000a600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE0;


    MEM_GOLD_LAYER1_INSTANCE1 : if BRAM_NAME = "gold_layer1_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"00000107000000000000000c0000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000004f00000000",
            INIT_03 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_04 => X"00000027000000000000002e0000000000000022000000000000000000000000",
            INIT_05 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"00000000000000000000001e000000000000004b000000000000002800000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000970000000000000000000000000000000000000000",
            INIT_0A => X"00000000000000000000004e0000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000106000000000000000000000000",
            INIT_0C => X"00000000000000000000002e0000000000000000000000000000000000000000",
            INIT_0D => X"000000000000000000000000000000000000000000000000000000d800000000",
            INIT_0E => X"0000000000000000000000000000000000000028000000000000006500000000",
            INIT_0F => X"0000007100000000000000b80000000000000000000000000000000000000000",
            INIT_10 => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"000000000000000000000000000000000000014a000000000000002a00000000",
            INIT_12 => X"0000000f000000000000007f000000000000000e000000000000001000000000",
            INIT_13 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_17 => X"0000000000000000000000000000000000000051000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000900000000000000120000000000000000000000000000000000000000",
            INIT_1A => X"0000005a00000000000000060000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000001200000000000000000000000000000000000000000000004f00000000",
            INIT_1D => X"0000000000000000000000000000000000000003000000000000002200000000",
            INIT_1E => X"0000000200000000000000290000000000000023000000000000003c00000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000004900000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"00000000000000000000005c0000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000006100000000",
            INIT_24 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000009500000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000009500000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000001c00000000000000000000000000000038000000000000008300000000",
            INIT_36 => X"0000004d00000000000000830000000000000063000000000000001b00000000",
            INIT_37 => X"0000000000000000000000150000000000000046000000000000004300000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"000000000000000000000000000000000000000a000000000000006b00000000",
            INIT_4F => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000890000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000310000000000000000000000000000000000000000",
            INIT_52 => X"0000007200000000000000340000000000000014000000000000000000000000",
            INIT_53 => X"00000000000000000000000000000000000000a1000000000000000000000000",
            INIT_54 => X"0000000000000000000000c80000000000000000000000000000000000000000",
            INIT_55 => X"000000000000000000000080000000000000005f000000000000009000000000",
            INIT_56 => X"000000000000000000000000000000000000003b000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"00000000000000000000000f0000000000000013000000000000005600000000",
            INIT_5B => X"000000650000000000000069000000000000002b000000000000000000000000",
            INIT_5C => X"0000000000000000000000200000000000000000000000000000001f00000000",
            INIT_5D => X"0000005d00000000000000200000000000000028000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000006c00000000",
            INIT_5F => X"0000007300000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_61 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_63 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_64 => X"00000036000000000000001e0000000000000000000000000000000000000000",
            INIT_65 => X"00000039000000000000000000000000000000d8000000000000009500000000",
            INIT_66 => X"000000a300000000000000910000000000000065000000000000008500000000",
            INIT_67 => X"00000060000000000000005a0000000000000070000000000000010e00000000",
            INIT_68 => X"00000000000000000000004b000000000000007b000000000000006a00000000",
            INIT_69 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000350000000000000000000000000000002300000000",
            INIT_6B => X"000000180000000000000000000000000000001a000000000000005d00000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000b00000000000000000000000000000000000000000000001700000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000001000000000000000000000000000000023000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000007500000000",
            INIT_72 => X"0000002e00000000000000360000000000000052000000000000002700000000",
            INIT_73 => X"0000000000000000000000000000000000000027000000000000002500000000",
            INIT_74 => X"0000002600000000000000000000000000000020000000000000000000000000",
            INIT_75 => X"0000005200000000000000a70000000000000059000000000000004e00000000",
            INIT_76 => X"000000f100000000000000450000000000000059000000000000004b00000000",
            INIT_77 => X"000000d800000000000000800000000000000077000000000000006d00000000",
            INIT_78 => X"0000009c00000000000000bc0000000000000055000000000000009100000000",
            INIT_79 => X"00000078000000000000019a000000000000009d000000000000003e00000000",
            INIT_7A => X"000000da000000000000004e0000000000000037000000000000002400000000",
            INIT_7B => X"0000006e00000000000000640000000000000133000000000000008200000000",
            INIT_7C => X"00000053000000000000007b0000000000000112000000000000004a00000000",
            INIT_7D => X"0000000000000000000000530000000000000000000000000000002e00000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000014000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE1;


    MEM_GOLD_LAYER1_INSTANCE2 : if BRAM_NAME = "gold_layer1_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"00000039000000000000002c0000000000000036000000000000000000000000",
            INIT_02 => X"000000080000000000000000000000000000001f000000000000002b00000000",
            INIT_03 => X"000000000000000000000000000000000000000b000000000000006a00000000",
            INIT_04 => X"0000009100000000000000270000000000000000000000000000002600000000",
            INIT_05 => X"0000005200000000000000000000000000000034000000000000001400000000",
            INIT_06 => X"000000000000000000000035000000000000000c000000000000001900000000",
            INIT_07 => X"00000034000000000000005a0000000000000027000000000000000000000000",
            INIT_08 => X"0000000000000000000000770000000000000018000000000000004d00000000",
            INIT_09 => X"000000080000000000000032000000000000002c000000000000001400000000",
            INIT_0A => X"0000002e000000000000007d0000000000000085000000000000000000000000",
            INIT_0B => X"00000031000000000000004d0000000000000050000000000000003500000000",
            INIT_0C => X"0000003e000000000000004c0000000000000017000000000000003f00000000",
            INIT_0D => X"0000009100000000000000840000000000000065000000000000004800000000",
            INIT_0E => X"000000430000000000000051000000000000002e000000000000009300000000",
            INIT_0F => X"0000007400000000000000ca0000000000000078000000000000005a00000000",
            INIT_10 => X"0000005e0000000000000059000000000000008a000000000000006000000000",
            INIT_11 => X"0000005d000000000000006f000000000000006c000000000000008900000000",
            INIT_12 => X"0000003700000000000000600000000000000055000000000000009c00000000",
            INIT_13 => X"0000006b00000000000000220000000000000020000000000000007800000000",
            INIT_14 => X"000000cf0000000000000022000000000000008b000000000000005900000000",
            INIT_15 => X"0000000000000000000000000000000000000075000000000000005d00000000",
            INIT_16 => X"0000000000000000000000090000000000000000000000000000006e00000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000005700000000000000000000000000000059000000000000000000000000",
            INIT_1B => X"0000004000000000000000900000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000e50000000000000000000000000000000700000000",
            INIT_1D => X"0000002f00000000000000080000000000000025000000000000000000000000",
            INIT_1E => X"00000000000000000000000000000000000001e8000000000000000000000000",
            INIT_1F => X"0000000000000000000000bd0000000000000000000000000000000000000000",
            INIT_20 => X"00000000000000000000002b0000000000000000000000000000010a00000000",
            INIT_21 => X"000000000000000000000000000000000000000000000000000000ec00000000",
            INIT_22 => X"0000018a0000000000000057000000000000009b000000000000000000000000",
            INIT_23 => X"0000006b00000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000e0000000000000000000000000000008a000000000000003300000000",
            INIT_25 => X"0000009300000000000000570000000000000050000000000000001700000000",
            INIT_26 => X"0000005300000000000000000000000000000019000000000000000000000000",
            INIT_27 => X"000000000000000000000000000000000000004d000000000000000000000000",
            INIT_28 => X"0000000000000000000000a5000000000000000d000000000000000000000000",
            INIT_29 => X"00000000000000000000009e000000000000003b00000000000000bd00000000",
            INIT_2A => X"000000f300000000000000000000000000000131000000000000000000000000",
            INIT_2B => X"00000000000000000000000d0000000000000124000000000000004800000000",
            INIT_2C => X"0000000000000000000000b60000000000000000000000000000008900000000",
            INIT_2D => X"00000033000000000000001b000000000000000000000000000000cb00000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000006700000000",
            INIT_2F => X"0000002f000000000000000000000000000000e5000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000031000000000000003500000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000b0000000000000000000000000000002a000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000002e00000000",
            INIT_3A => X"0000000000000000000000720000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000007400000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_3E => X"0000000000000000000000260000000000000000000000000000000000000000",
            INIT_3F => X"000000420000000000000075000000000000009d000000000000000e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002300000000000000000000000000000000000000000000005900000000",
            INIT_41 => X"0000001800000000000000000000000000000000000000000000001a00000000",
            INIT_42 => X"000000000000000000000079000000000000006b000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_44 => X"0000000000000000000000350000000000000053000000000000001e00000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_46 => X"00000062000000000000009a0000000000000021000000000000000c00000000",
            INIT_47 => X"000000e4000000000000002300000000000000c0000000000000003f00000000",
            INIT_48 => X"0000001000000000000000000000000000000018000000000000008400000000",
            INIT_49 => X"0000000000000000000000370000000000000102000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000001700000000000000180000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"000000400000000000000009000000000000003d000000000000001e00000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000007a00000000",
            INIT_51 => X"0000009d00000000000000000000000000000024000000000000000000000000",
            INIT_52 => X"00000010000000000000005a0000000000000016000000000000008900000000",
            INIT_53 => X"000000a700000000000000fe0000000000000000000000000000004800000000",
            INIT_54 => X"0000011600000000000000f500000000000000f800000000000000b900000000",
            INIT_55 => X"00000117000000000000013c0000000000000122000000000000013c00000000",
            INIT_56 => X"000001530000000000000127000000000000011e000000000000010e00000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000004300000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"000000000000000000000087000000000000003c000000000000003200000000",
            INIT_5B => X"0000001f00000000000000a1000000000000001b000000000000000000000000",
            INIT_5C => X"00000000000000000000000b0000000000000057000000000000004100000000",
            INIT_5D => X"0000002e000000000000000000000000000000be000000000000000000000000",
            INIT_5E => X"0000001a0000000000000000000000000000005f000000000000005900000000",
            INIT_5F => X"0000000000000000000000480000000000000000000000000000000000000000",
            INIT_60 => X"0000007c0000000000000000000000000000000000000000000000b900000000",
            INIT_61 => X"0000000000000000000000f2000000000000005400000000000000ac00000000",
            INIT_62 => X"000000b200000000000000c900000000000000ab000000000000005d00000000",
            INIT_63 => X"000000b900000000000000aa000000000000008300000000000000c000000000",
            INIT_64 => X"0000006200000000000000600000000000000062000000000000007300000000",
            INIT_65 => X"0000005800000000000000a300000000000000b800000000000000a900000000",
            INIT_66 => X"000000000000000000000061000000000000001e000000000000006100000000",
            INIT_67 => X"0000007e000000000000000e0000000000000000000000000000008800000000",
            INIT_68 => X"0000006c00000000000000000000000000000039000000000000000400000000",
            INIT_69 => X"0000000000000000000000620000000000000000000000000000006500000000",
            INIT_6A => X"0000002b00000000000000110000000000000000000000000000003d00000000",
            INIT_6B => X"0000006c000000000000001f000000000000000b000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"000000e300000000000000fc0000000000000000000000000000000000000000",
            INIT_70 => X"0000005c000000000000008d00000000000000f0000000000000006b00000000",
            INIT_71 => X"0000007600000000000000c9000000000000004b00000000000000c700000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_77 => X"0000002000000000000000380000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE2;


    MEM_GOLD_LAYER1_INSTANCE3 : if BRAM_NAME = "gold_layer1_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_04 => X"0000001e00000000000001170000000000000000000000000000000000000000",
            INIT_05 => X"0000008c000000000000006500000000000000bd000000000000007a00000000",
            INIT_06 => X"0000008d000000000000011200000000000000c7000000000000009900000000",
            INIT_07 => X"000000cd00000000000000ce000000000000009b000000000000008800000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE3;


    MEM_GOLD_LAYER2_INSTANCE0 : if BRAM_NAME = "gold_layer2_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0001645600000000fffddf45fffffffffff9da94fffffffffffebef8ffffffff",
            INIT_01 => X"fffd7458fffffffffffccb7afffffffffffeb2bffffffffffffde323ffffffff",
            INIT_02 => X"fff94239fffffffffffd5829ffffffff",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER2_INSTANCE0;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE0 : if BRAM_NAME = "sampleifmap_layersamples_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a600000000000000a5000000000000009f000000000000009e00000000",
            INIT_01 => X"0000009f00000000000000a2000000000000009c00000000000000a000000000",
            INIT_02 => X"000000a000000000000000a1000000000000009f000000000000009e00000000",
            INIT_03 => X"000000aa00000000000000a900000000000000a600000000000000a100000000",
            INIT_04 => X"000000a000000000000000a000000000000000a200000000000000a700000000",
            INIT_05 => X"0000009400000000000000960000000000000095000000000000009c00000000",
            INIT_06 => X"0000008d000000000000008c000000000000008f000000000000009500000000",
            INIT_07 => X"00000074000000000000007e0000000000000089000000000000008f00000000",
            INIT_08 => X"000000a6000000000000009f0000000000000097000000000000009800000000",
            INIT_09 => X"000000a200000000000000a400000000000000a000000000000000a200000000",
            INIT_0A => X"0000009f000000000000009b000000000000009c00000000000000a300000000",
            INIT_0B => X"000000ab00000000000000ab00000000000000aa00000000000000a300000000",
            INIT_0C => X"00000097000000000000009a00000000000000a000000000000000a900000000",
            INIT_0D => X"0000008d000000000000008c000000000000008b000000000000009100000000",
            INIT_0E => X"0000008e00000000000000910000000000000093000000000000009500000000",
            INIT_0F => X"00000077000000000000007d0000000000000088000000000000008f00000000",
            INIT_10 => X"000000a7000000000000009e0000000000000097000000000000009700000000",
            INIT_11 => X"000000a500000000000000a500000000000000a300000000000000a000000000",
            INIT_12 => X"0000009d000000000000009e00000000000000a200000000000000a300000000",
            INIT_13 => X"000000a900000000000000a700000000000000a600000000000000a100000000",
            INIT_14 => X"000000790000000000000091000000000000009f00000000000000aa00000000",
            INIT_15 => X"0000007200000000000000650000000000000062000000000000006e00000000",
            INIT_16 => X"0000008c000000000000008f0000000000000086000000000000007800000000",
            INIT_17 => X"000000780000000000000082000000000000008b000000000000008e00000000",
            INIT_18 => X"000000ae00000000000000a0000000000000009b000000000000009b00000000",
            INIT_19 => X"000000a900000000000000a900000000000000a700000000000000a700000000",
            INIT_1A => X"000000bf00000000000000a700000000000000a500000000000000a500000000",
            INIT_1B => X"000000a400000000000000a2000000000000009d00000000000000b100000000",
            INIT_1C => X"0000006700000000000000680000000000000095000000000000009e00000000",
            INIT_1D => X"0000004a0000000000000050000000000000005c000000000000006200000000",
            INIT_1E => X"0000008400000000000000710000000000000053000000000000005600000000",
            INIT_1F => X"0000007f0000000000000088000000000000008c000000000000008c00000000",
            INIT_20 => X"000000aa00000000000000a1000000000000009c000000000000009b00000000",
            INIT_21 => X"000000a600000000000000a900000000000000a300000000000000a900000000",
            INIT_22 => X"000000f600000000000000ad00000000000000a400000000000000a400000000",
            INIT_23 => X"0000008e0000000000000092000000000000009700000000000000c300000000",
            INIT_24 => X"000000710000000000000055000000000000004e000000000000006f00000000",
            INIT_25 => X"0000005d0000000000000061000000000000006a000000000000007000000000",
            INIT_26 => X"0000006900000000000000550000000000000054000000000000004a00000000",
            INIT_27 => X"000000810000000000000085000000000000008a000000000000008000000000",
            INIT_28 => X"0000009300000000000000820000000000000085000000000000009400000000",
            INIT_29 => X"000000a700000000000000a700000000000000a500000000000000a100000000",
            INIT_2A => X"000000b400000000000000a300000000000000a500000000000000a300000000",
            INIT_2B => X"0000004200000000000000610000000000000080000000000000009d00000000",
            INIT_2C => X"0000007600000000000000590000000000000042000000000000004500000000",
            INIT_2D => X"0000005e00000000000000720000000000000077000000000000007a00000000",
            INIT_2E => X"00000043000000000000003a000000000000005b000000000000006300000000",
            INIT_2F => X"00000086000000000000008a000000000000008c000000000000006c00000000",
            INIT_30 => X"00000058000000000000002f000000000000006d000000000000007f00000000",
            INIT_31 => X"000000aa00000000000000a800000000000000aa000000000000009900000000",
            INIT_32 => X"0000009300000000000000a400000000000000a600000000000000a900000000",
            INIT_33 => X"000000440000000000000064000000000000007f000000000000008100000000",
            INIT_34 => X"0000008400000000000000530000000000000048000000000000004e00000000",
            INIT_35 => X"0000006b0000000000000069000000000000007c000000000000009200000000",
            INIT_36 => X"0000002e000000000000003f0000000000000055000000000000007300000000",
            INIT_37 => X"00000086000000000000008d0000000000000084000000000000004f00000000",
            INIT_38 => X"00000046000000000000002a0000000000000063000000000000008300000000",
            INIT_39 => X"000000a800000000000000a500000000000000a7000000000000008f00000000",
            INIT_3A => X"00000078000000000000008c00000000000000a100000000000000ab00000000",
            INIT_3B => X"0000005800000000000000740000000000000090000000000000008200000000",
            INIT_3C => X"0000007c000000000000004d0000000000000055000000000000005b00000000",
            INIT_3D => X"0000006a0000000000000066000000000000008800000000000000a300000000",
            INIT_3E => X"0000003100000000000000360000000000000055000000000000006400000000",
            INIT_3F => X"00000088000000000000008a000000000000006b000000000000003900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007c0000000000000036000000000000006700000000000000aa00000000",
            INIT_41 => X"000000a600000000000000a300000000000000a1000000000000009900000000",
            INIT_42 => X"0000007d000000000000007100000000000000ae00000000000000a500000000",
            INIT_43 => X"000000560000000000000079000000000000009c000000000000009d00000000",
            INIT_44 => X"0000005100000000000000500000000000000054000000000000005200000000",
            INIT_45 => X"0000005700000000000000710000000000000092000000000000008a00000000",
            INIT_46 => X"0000003800000000000000470000000000000056000000000000005300000000",
            INIT_47 => X"000000890000000000000085000000000000004a000000000000002800000000",
            INIT_48 => X"0000009a000000000000005e000000000000008600000000000000b400000000",
            INIT_49 => X"00000099000000000000009c000000000000009e00000000000000ae00000000",
            INIT_4A => X"0000009c00000000000000cf00000000000000ed00000000000000cf00000000",
            INIT_4B => X"0000005d000000000000007d000000000000009400000000000000ae00000000",
            INIT_4C => X"0000004c000000000000003b000000000000004a000000000000005600000000",
            INIT_4D => X"0000006a0000000000000085000000000000008f000000000000008900000000",
            INIT_4E => X"0000004b00000000000000540000000000000057000000000000005600000000",
            INIT_4F => X"00000084000000000000005f0000000000000028000000000000003200000000",
            INIT_50 => X"000000a5000000000000008e000000000000006c00000000000000b700000000",
            INIT_51 => X"0000007a000000000000009f000000000000009b00000000000000b100000000",
            INIT_52 => X"000000a400000000000000dc00000000000000ed00000000000000d500000000",
            INIT_53 => X"00000078000000000000007d000000000000009c00000000000000b700000000",
            INIT_54 => X"0000005b000000000000002d0000000000000050000000000000004e00000000",
            INIT_55 => X"0000006b000000000000009b000000000000009d00000000000000af00000000",
            INIT_56 => X"0000004e00000000000000580000000000000067000000000000005700000000",
            INIT_57 => X"00000068000000000000003b0000000000000029000000000000003b00000000",
            INIT_58 => X"000000aa0000000000000087000000000000006400000000000000bc00000000",
            INIT_59 => X"0000008600000000000000ad00000000000000a600000000000000bb00000000",
            INIT_5A => X"000000aa00000000000000c700000000000000c2000000000000007500000000",
            INIT_5B => X"00000075000000000000008600000000000000bd00000000000000b900000000",
            INIT_5C => X"0000007d00000000000000260000000000000054000000000000006600000000",
            INIT_5D => X"0000005d000000000000009200000000000000a000000000000000d200000000",
            INIT_5E => X"000000550000000000000068000000000000005e000000000000005300000000",
            INIT_5F => X"0000004c000000000000003e0000000000000037000000000000004900000000",
            INIT_60 => X"000000af000000000000007f000000000000005a00000000000000bd00000000",
            INIT_61 => X"0000009f00000000000000b200000000000000a600000000000000ae00000000",
            INIT_62 => X"0000008900000000000000a800000000000000a8000000000000006100000000",
            INIT_63 => X"0000007b00000000000000a000000000000000d800000000000000ba00000000",
            INIT_64 => X"0000009600000000000000320000000000000073000000000000007800000000",
            INIT_65 => X"0000005b000000000000007b000000000000009b00000000000000c200000000",
            INIT_66 => X"00000056000000000000005f0000000000000054000000000000005400000000",
            INIT_67 => X"00000049000000000000004f0000000000000049000000000000005400000000",
            INIT_68 => X"000000b90000000000000098000000000000005d00000000000000bd00000000",
            INIT_69 => X"000000a700000000000000ad0000000000000088000000000000007700000000",
            INIT_6A => X"000000a700000000000000910000000000000093000000000000006700000000",
            INIT_6B => X"0000008d00000000000000b400000000000000e200000000000000bd00000000",
            INIT_6C => X"0000009a00000000000000470000000000000075000000000000007e00000000",
            INIT_6D => X"000000570000000000000072000000000000009500000000000000ba00000000",
            INIT_6E => X"0000006300000000000000500000000000000048000000000000005000000000",
            INIT_6F => X"0000005e0000000000000061000000000000005a000000000000006400000000",
            INIT_70 => X"000000ba00000000000000a8000000000000006c00000000000000c200000000",
            INIT_71 => X"000000a7000000000000009c0000000000000063000000000000006900000000",
            INIT_72 => X"000000c6000000000000008a0000000000000073000000000000006400000000",
            INIT_73 => X"0000009a000000000000009100000000000000ac00000000000000be00000000",
            INIT_74 => X"0000009800000000000000470000000000000067000000000000009200000000",
            INIT_75 => X"0000006e0000000000000082000000000000008900000000000000b300000000",
            INIT_76 => X"0000006d000000000000005f000000000000005b000000000000005500000000",
            INIT_77 => X"0000007500000000000000610000000000000064000000000000007300000000",
            INIT_78 => X"000000b800000000000000ac000000000000008400000000000000c500000000",
            INIT_79 => X"0000009b000000000000008c000000000000004e000000000000008200000000",
            INIT_7A => X"000000e6000000000000008f0000000000000082000000000000007300000000",
            INIT_7B => X"000000830000000000000087000000000000009100000000000000f200000000",
            INIT_7C => X"00000090000000000000005f000000000000006c000000000000007900000000",
            INIT_7D => X"000000570000000000000070000000000000009800000000000000a800000000",
            INIT_7E => X"0000007000000000000000690000000000000057000000000000004700000000",
            INIT_7F => X"0000008800000000000000790000000000000067000000000000007800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE0;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE1 : if BRAM_NAME = "sampleifmap_layersamples_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bf00000000000000a8000000000000009200000000000000cb00000000",
            INIT_01 => X"0000008a000000000000007e000000000000004e00000000000000a800000000",
            INIT_02 => X"000000ad000000000000009a0000000000000060000000000000008a00000000",
            INIT_03 => X"000000710000000000000071000000000000008c00000000000000a200000000",
            INIT_04 => X"000000ab00000000000000700000000000000069000000000000006500000000",
            INIT_05 => X"0000006d00000000000000870000000000000094000000000000009c00000000",
            INIT_06 => X"00000065000000000000005e000000000000004f000000000000004e00000000",
            INIT_07 => X"000000900000000000000097000000000000007d000000000000006b00000000",
            INIT_08 => X"000000b700000000000000a400000000000000a300000000000000d600000000",
            INIT_09 => X"0000009c0000000000000060000000000000005e00000000000000b000000000",
            INIT_0A => X"000000760000000000000081000000000000006a000000000000009400000000",
            INIT_0B => X"0000007300000000000000660000000000000074000000000000007200000000",
            INIT_0C => X"0000007600000000000000900000000000000065000000000000005600000000",
            INIT_0D => X"0000004b00000000000000850000000000000080000000000000004400000000",
            INIT_0E => X"000000660000000000000047000000000000003a000000000000003c00000000",
            INIT_0F => X"0000008c0000000000000096000000000000008f000000000000007400000000",
            INIT_10 => X"000000ad00000000000000a700000000000000b200000000000000d400000000",
            INIT_11 => X"0000008d0000000000000056000000000000007c00000000000000b000000000",
            INIT_12 => X"0000004d00000000000000680000000000000087000000000000009900000000",
            INIT_13 => X"000000930000000000000081000000000000007c000000000000008600000000",
            INIT_14 => X"000000840000000000000096000000000000005c000000000000005500000000",
            INIT_15 => X"00000040000000000000004b000000000000006b000000000000007500000000",
            INIT_16 => X"0000008500000000000000560000000000000041000000000000002c00000000",
            INIT_17 => X"00000097000000000000009a00000000000000a0000000000000009b00000000",
            INIT_18 => X"000000ae00000000000000ab00000000000000bb00000000000000c700000000",
            INIT_19 => X"000000770000000000000056000000000000009000000000000000b100000000",
            INIT_1A => X"0000004600000000000000900000000000000089000000000000007a00000000",
            INIT_1B => X"000000b80000000000000091000000000000006c000000000000008100000000",
            INIT_1C => X"0000008900000000000000830000000000000049000000000000007400000000",
            INIT_1D => X"0000003400000000000000330000000000000059000000000000008600000000",
            INIT_1E => X"000000a30000000000000079000000000000005a000000000000002f00000000",
            INIT_1F => X"00000095000000000000009e00000000000000a400000000000000ab00000000",
            INIT_20 => X"000000b100000000000000b300000000000000c300000000000000a500000000",
            INIT_21 => X"000000830000000000000063000000000000009800000000000000b500000000",
            INIT_22 => X"00000050000000000000005d000000000000006700000000000000ab00000000",
            INIT_23 => X"000000bf00000000000000b2000000000000007a000000000000005d00000000",
            INIT_24 => X"0000005700000000000000590000000000000064000000000000009600000000",
            INIT_25 => X"000000180000000000000026000000000000002e000000000000003c00000000",
            INIT_26 => X"00000090000000000000006c000000000000003c000000000000002e00000000",
            INIT_27 => X"00000078000000000000007f0000000000000080000000000000009000000000",
            INIT_28 => X"000000b200000000000000b100000000000000c3000000000000007500000000",
            INIT_29 => X"000000960000000000000053000000000000008a00000000000000b500000000",
            INIT_2A => X"00000086000000000000008500000000000000db00000000000000f500000000",
            INIT_2B => X"000000c200000000000000be00000000000000b0000000000000009500000000",
            INIT_2C => X"0000003d000000000000006e000000000000007d00000000000000a800000000",
            INIT_2D => X"0000003a00000000000000310000000000000022000000000000002300000000",
            INIT_2E => X"000000480000000000000045000000000000003a000000000000003d00000000",
            INIT_2F => X"00000037000000000000003b0000000000000045000000000000004e00000000",
            INIT_30 => X"000000b000000000000000ae00000000000000af000000000000004f00000000",
            INIT_31 => X"000000d3000000000000006d000000000000008c00000000000000b100000000",
            INIT_32 => X"0000007c00000000000000d000000000000000fc00000000000000fd00000000",
            INIT_33 => X"0000007a0000000000000074000000000000007c000000000000007200000000",
            INIT_34 => X"0000003c00000000000000440000000000000044000000000000006800000000",
            INIT_35 => X"0000003800000000000000330000000000000032000000000000003400000000",
            INIT_36 => X"00000033000000000000002b0000000000000033000000000000003800000000",
            INIT_37 => X"0000002a000000000000002b0000000000000030000000000000003b00000000",
            INIT_38 => X"000000a800000000000000900000000000000060000000000000002900000000",
            INIT_39 => X"000000f600000000000000a500000000000000a500000000000000b200000000",
            INIT_3A => X"0000003c000000000000006e00000000000000e300000000000000fd00000000",
            INIT_3B => X"0000003000000000000000310000000000000031000000000000003500000000",
            INIT_3C => X"0000002a000000000000002e000000000000002a000000000000002d00000000",
            INIT_3D => X"0000002b000000000000002e000000000000002e000000000000002600000000",
            INIT_3E => X"00000032000000000000002e000000000000002e000000000000002a00000000",
            INIT_3F => X"0000002d00000000000000330000000000000035000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000083000000000000003b000000000000001d000000000000001d00000000",
            INIT_41 => X"000000fe00000000000000c2000000000000008400000000000000a600000000",
            INIT_42 => X"00000032000000000000003d000000000000008d00000000000000f100000000",
            INIT_43 => X"0000003200000000000000310000000000000033000000000000003200000000",
            INIT_44 => X"000000220000000000000027000000000000002a000000000000002f00000000",
            INIT_45 => X"0000002a00000000000000260000000000000027000000000000002300000000",
            INIT_46 => X"0000003b000000000000003e0000000000000038000000000000002d00000000",
            INIT_47 => X"00000033000000000000002e0000000000000032000000000000003800000000",
            INIT_48 => X"000000490000000000000022000000000000001e000000000000003000000000",
            INIT_49 => X"0000010000000000000000d70000000000000080000000000000008000000000",
            INIT_4A => X"000000320000000000000036000000000000004200000000000000bb00000000",
            INIT_4B => X"0000002d000000000000002e0000000000000034000000000000003400000000",
            INIT_4C => X"0000002700000000000000240000000000000029000000000000002b00000000",
            INIT_4D => X"0000002e000000000000002b0000000000000028000000000000002800000000",
            INIT_4E => X"0000003b0000000000000040000000000000003e000000000000003b00000000",
            INIT_4F => X"0000005300000000000000460000000000000032000000000000003600000000",
            INIT_50 => X"00000029000000000000001f0000000000000023000000000000003400000000",
            INIT_51 => X"000000f000000000000000e00000000000000080000000000000004200000000",
            INIT_52 => X"000000380000000000000031000000000000003a000000000000007c00000000",
            INIT_53 => X"0000002f000000000000002c000000000000002c000000000000003600000000",
            INIT_54 => X"0000002c000000000000002b000000000000002b000000000000002e00000000",
            INIT_55 => X"0000003a0000000000000036000000000000002d000000000000002c00000000",
            INIT_56 => X"00000024000000000000002b000000000000002e000000000000003600000000",
            INIT_57 => X"0000004c00000000000000550000000000000049000000000000003300000000",
            INIT_58 => X"00000023000000000000001d0000000000000023000000000000003200000000",
            INIT_59 => X"000000d300000000000000ca000000000000004e000000000000002c00000000",
            INIT_5A => X"0000003000000000000000360000000000000041000000000000006100000000",
            INIT_5B => X"0000002d00000000000000280000000000000030000000000000003a00000000",
            INIT_5C => X"0000002e000000000000002f0000000000000030000000000000002f00000000",
            INIT_5D => X"0000003000000000000000270000000000000027000000000000003300000000",
            INIT_5E => X"00000028000000000000001c0000000000000027000000000000002f00000000",
            INIT_5F => X"00000033000000000000002e0000000000000043000000000000004300000000",
            INIT_60 => X"0000002100000000000000200000000000000023000000000000003200000000",
            INIT_61 => X"000000aa0000000000000068000000000000002e000000000000002900000000",
            INIT_62 => X"0000003500000000000000340000000000000036000000000000004000000000",
            INIT_63 => X"0000002d0000000000000036000000000000003a000000000000003d00000000",
            INIT_64 => X"00000031000000000000002e0000000000000029000000000000002a00000000",
            INIT_65 => X"000000270000000000000028000000000000002a000000000000002e00000000",
            INIT_66 => X"0000003f000000000000002c0000000000000028000000000000002500000000",
            INIT_67 => X"00000033000000000000000f000000000000001f000000000000002f00000000",
            INIT_68 => X"00000026000000000000001f000000000000002a000000000000004400000000",
            INIT_69 => X"00000047000000000000002a000000000000002b000000000000002500000000",
            INIT_6A => X"00000026000000000000001b000000000000001f000000000000003100000000",
            INIT_6B => X"00000035000000000000003a0000000000000038000000000000003100000000",
            INIT_6C => X"000000350000000000000039000000000000003c000000000000003800000000",
            INIT_6D => X"000000210000000000000027000000000000002d000000000000003200000000",
            INIT_6E => X"00000049000000000000004f000000000000003e000000000000002a00000000",
            INIT_6F => X"00000028000000000000000d0000000000000026000000000000003800000000",
            INIT_70 => X"0000002b00000000000000230000000000000031000000000000003d00000000",
            INIT_71 => X"00000028000000000000002c000000000000002a000000000000002700000000",
            INIT_72 => X"0000001e0000000000000017000000000000001b000000000000002a00000000",
            INIT_73 => X"0000002f0000000000000024000000000000001d000000000000001b00000000",
            INIT_74 => X"0000004b0000000000000042000000000000003e000000000000003800000000",
            INIT_75 => X"0000002b000000000000002b0000000000000031000000000000004500000000",
            INIT_76 => X"0000005d000000000000006d0000000000000055000000000000003c00000000",
            INIT_77 => X"00000014000000000000001d000000000000001a000000000000003c00000000",
            INIT_78 => X"0000002b000000000000002d0000000000000038000000000000003600000000",
            INIT_79 => X"0000002600000000000000280000000000000028000000000000002800000000",
            INIT_7A => X"0000001d0000000000000016000000000000001a000000000000002400000000",
            INIT_7B => X"000000120000000000000013000000000000001d000000000000001900000000",
            INIT_7C => X"0000004a000000000000003d000000000000002f000000000000002000000000",
            INIT_7D => X"0000002d00000000000000340000000000000035000000000000004200000000",
            INIT_7E => X"0000005900000000000000690000000000000059000000000000004300000000",
            INIT_7F => X"0000001500000000000000220000000000000018000000000000003000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE1;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE2 : if BRAM_NAME = "sampleifmap_layersamples_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000760000000000000074000000000000006f000000000000007000000000",
            INIT_01 => X"000000710000000000000073000000000000006d000000000000007000000000",
            INIT_02 => X"0000006f00000000000000740000000000000071000000000000006f00000000",
            INIT_03 => X"0000007700000000000000750000000000000075000000000000006f00000000",
            INIT_04 => X"00000070000000000000006f0000000000000071000000000000007500000000",
            INIT_05 => X"0000006a000000000000006b000000000000006b000000000000006d00000000",
            INIT_06 => X"0000006100000000000000620000000000000065000000000000006b00000000",
            INIT_07 => X"00000055000000000000005b000000000000005f000000000000006100000000",
            INIT_08 => X"000000740000000000000072000000000000006e000000000000007000000000",
            INIT_09 => X"0000007200000000000000750000000000000071000000000000007000000000",
            INIT_0A => X"0000006e000000000000006f000000000000006e000000000000007400000000",
            INIT_0B => X"0000007300000000000000750000000000000077000000000000007100000000",
            INIT_0C => X"000000730000000000000070000000000000006f000000000000007300000000",
            INIT_0D => X"0000006400000000000000660000000000000068000000000000006e00000000",
            INIT_0E => X"0000006100000000000000660000000000000066000000000000006900000000",
            INIT_0F => X"00000058000000000000005b000000000000005f000000000000006200000000",
            INIT_10 => X"0000006f000000000000006f000000000000006d000000000000006e00000000",
            INIT_11 => X"0000007500000000000000750000000000000073000000000000006a00000000",
            INIT_12 => X"0000006d00000000000000720000000000000073000000000000007300000000",
            INIT_13 => X"0000007100000000000000720000000000000073000000000000006f00000000",
            INIT_14 => X"00000060000000000000006f0000000000000072000000000000007400000000",
            INIT_15 => X"00000055000000000000004d000000000000004e000000000000005a00000000",
            INIT_16 => X"0000006300000000000000670000000000000060000000000000005600000000",
            INIT_17 => X"00000059000000000000005f0000000000000062000000000000006300000000",
            INIT_18 => X"00000070000000000000006d000000000000006e000000000000006b00000000",
            INIT_19 => X"0000007700000000000000780000000000000075000000000000006e00000000",
            INIT_1A => X"00000092000000000000007b0000000000000075000000000000007300000000",
            INIT_1B => X"000000720000000000000073000000000000006f000000000000008200000000",
            INIT_1C => X"000000570000000000000050000000000000006f000000000000007000000000",
            INIT_1D => X"0000003f000000000000004b000000000000005a000000000000005a00000000",
            INIT_1E => X"000000620000000000000055000000000000003e000000000000004600000000",
            INIT_1F => X"0000005e00000000000000630000000000000065000000000000006600000000",
            INIT_20 => X"0000007200000000000000730000000000000072000000000000006b00000000",
            INIT_21 => X"0000007400000000000000780000000000000071000000000000007200000000",
            INIT_22 => X"000000d600000000000000800000000000000074000000000000007100000000",
            INIT_23 => X"0000006c000000000000006f0000000000000072000000000000009c00000000",
            INIT_24 => X"0000006700000000000000450000000000000035000000000000005000000000",
            INIT_25 => X"0000005e00000000000000660000000000000072000000000000006e00000000",
            INIT_26 => X"000000530000000000000049000000000000004e000000000000004800000000",
            INIT_27 => X"0000005d000000000000005e0000000000000065000000000000006000000000",
            INIT_28 => X"0000007000000000000000640000000000000068000000000000006d00000000",
            INIT_29 => X"0000007300000000000000740000000000000071000000000000007300000000",
            INIT_2A => X"0000008a00000000000000760000000000000074000000000000006f00000000",
            INIT_2B => X"00000032000000000000004b0000000000000066000000000000007a00000000",
            INIT_2C => X"0000007100000000000000530000000000000038000000000000003a00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007900000000",
            INIT_2E => X"0000003a000000000000003a000000000000005b000000000000006400000000",
            INIT_2F => X"0000005f00000000000000620000000000000069000000000000005400000000",
            INIT_30 => X"0000004a0000000000000025000000000000005f000000000000006400000000",
            INIT_31 => X"0000007600000000000000730000000000000076000000000000007500000000",
            INIT_32 => X"0000006b00000000000000780000000000000074000000000000007500000000",
            INIT_33 => X"000000430000000000000057000000000000006c000000000000006200000000",
            INIT_34 => X"000000820000000000000054000000000000004b000000000000005300000000",
            INIT_35 => X"0000006600000000000000630000000000000076000000000000008e00000000",
            INIT_36 => X"0000002f00000000000000470000000000000053000000000000006f00000000",
            INIT_37 => X"0000005d00000000000000630000000000000062000000000000003d00000000",
            INIT_38 => X"00000040000000000000002b0000000000000060000000000000007300000000",
            INIT_39 => X"0000007400000000000000720000000000000075000000000000006f00000000",
            INIT_3A => X"0000005e000000000000006d0000000000000071000000000000007700000000",
            INIT_3B => X"00000057000000000000006a0000000000000083000000000000006e00000000",
            INIT_3C => X"00000076000000000000004d0000000000000058000000000000005f00000000",
            INIT_3D => X"00000062000000000000005d000000000000007c000000000000009900000000",
            INIT_3E => X"00000035000000000000003c0000000000000051000000000000005d00000000",
            INIT_3F => X"0000006100000000000000670000000000000053000000000000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000079000000000000003a000000000000006900000000000000a100000000",
            INIT_41 => X"0000007a00000000000000750000000000000071000000000000007c00000000",
            INIT_42 => X"0000006900000000000000590000000000000087000000000000007900000000",
            INIT_43 => X"00000050000000000000006f000000000000008f000000000000008d00000000",
            INIT_44 => X"00000047000000000000004e0000000000000055000000000000005100000000",
            INIT_45 => X"0000004f00000000000000670000000000000087000000000000007d00000000",
            INIT_46 => X"0000003900000000000000490000000000000052000000000000004d00000000",
            INIT_47 => X"00000067000000000000006a000000000000003b000000000000002300000000",
            INIT_48 => X"0000009a0000000000000064000000000000008b00000000000000b000000000",
            INIT_49 => X"0000007600000000000000740000000000000074000000000000009500000000",
            INIT_4A => X"0000008300000000000000b400000000000000d600000000000000b400000000",
            INIT_4B => X"00000055000000000000006e0000000000000083000000000000009900000000",
            INIT_4C => X"000000440000000000000039000000000000004a000000000000005400000000",
            INIT_4D => X"00000062000000000000007c0000000000000085000000000000007d00000000",
            INIT_4E => X"0000004c00000000000000550000000000000055000000000000005100000000",
            INIT_4F => X"00000067000000000000004b000000000000001e000000000000003100000000",
            INIT_50 => X"000000a90000000000000097000000000000007400000000000000b700000000",
            INIT_51 => X"0000005900000000000000760000000000000070000000000000009c00000000",
            INIT_52 => X"0000008700000000000000bf00000000000000e000000000000000c500000000",
            INIT_53 => X"0000006f000000000000006c0000000000000089000000000000009f00000000",
            INIT_54 => X"00000055000000000000002c0000000000000050000000000000004c00000000",
            INIT_55 => X"000000640000000000000093000000000000009300000000000000a500000000",
            INIT_56 => X"0000004f00000000000000580000000000000066000000000000005300000000",
            INIT_57 => X"00000051000000000000002e0000000000000024000000000000003b00000000",
            INIT_58 => X"000000af0000000000000090000000000000006c00000000000000bf00000000",
            INIT_59 => X"0000005d000000000000007b000000000000007800000000000000a700000000",
            INIT_5A => X"0000008e00000000000000ab00000000000000b6000000000000005f00000000",
            INIT_5B => X"0000006b000000000000007700000000000000ab00000000000000a100000000",
            INIT_5C => X"0000007900000000000000260000000000000054000000000000006200000000",
            INIT_5D => X"00000059000000000000008b000000000000009800000000000000c900000000",
            INIT_5E => X"000000570000000000000068000000000000005d000000000000005000000000",
            INIT_5F => X"0000003800000000000000370000000000000035000000000000004b00000000",
            INIT_60 => X"000000b40000000000000086000000000000006000000000000000c200000000",
            INIT_61 => X"0000006d000000000000007b000000000000007b000000000000009c00000000",
            INIT_62 => X"000000720000000000000090000000000000009a000000000000004400000000",
            INIT_63 => X"00000071000000000000009500000000000000ca00000000000000a600000000",
            INIT_64 => X"0000009300000000000000320000000000000072000000000000007200000000",
            INIT_65 => X"000000580000000000000076000000000000009500000000000000bb00000000",
            INIT_66 => X"00000057000000000000005f0000000000000054000000000000005300000000",
            INIT_67 => X"00000037000000000000004a0000000000000049000000000000005700000000",
            INIT_68 => X"000000bc000000000000009a000000000000005f00000000000000c000000000",
            INIT_69 => X"00000074000000000000007c000000000000006a000000000000006e00000000",
            INIT_6A => X"00000095000000000000007d0000000000000084000000000000004800000000",
            INIT_6B => X"0000008300000000000000ac00000000000000d800000000000000ae00000000",
            INIT_6C => X"0000009800000000000000470000000000000072000000000000007500000000",
            INIT_6D => X"00000055000000000000006e000000000000009000000000000000b500000000",
            INIT_6E => X"0000006400000000000000500000000000000049000000000000005000000000",
            INIT_6F => X"0000004900000000000000590000000000000058000000000000006500000000",
            INIT_70 => X"000000ba00000000000000a7000000000000006b00000000000000c400000000",
            INIT_71 => X"0000007a00000000000000770000000000000059000000000000006d00000000",
            INIT_72 => X"000000b9000000000000007b000000000000006a000000000000004a00000000",
            INIT_73 => X"0000008f000000000000008c00000000000000a500000000000000b400000000",
            INIT_74 => X"0000009800000000000000470000000000000064000000000000008800000000",
            INIT_75 => X"0000006d0000000000000080000000000000008500000000000000af00000000",
            INIT_76 => X"0000006e0000000000000060000000000000005d000000000000005600000000",
            INIT_77 => X"0000005f00000000000000550000000000000060000000000000007400000000",
            INIT_78 => X"000000b200000000000000a7000000000000008100000000000000c500000000",
            INIT_79 => X"0000007d00000000000000780000000000000053000000000000008900000000",
            INIT_7A => X"000000dd00000000000000830000000000000078000000000000005e00000000",
            INIT_7B => X"000000790000000000000082000000000000008a00000000000000ec00000000",
            INIT_7C => X"0000008600000000000000580000000000000068000000000000007000000000",
            INIT_7D => X"00000055000000000000006c0000000000000093000000000000009f00000000",
            INIT_7E => X"0000006d00000000000000680000000000000058000000000000004800000000",
            INIT_7F => X"0000006800000000000000600000000000000056000000000000006e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE2;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE3 : if BRAM_NAME = "sampleifmap_layersamples_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b600000000000000a4000000000000009200000000000000cb00000000",
            INIT_01 => X"0000007e000000000000007d000000000000005600000000000000aa00000000",
            INIT_02 => X"000000a3000000000000008f0000000000000050000000000000007900000000",
            INIT_03 => X"0000006a000000000000006a0000000000000084000000000000009800000000",
            INIT_04 => X"0000008f000000000000005a0000000000000065000000000000006500000000",
            INIT_05 => X"000000690000000000000082000000000000008d000000000000008a00000000",
            INIT_06 => X"0000005b000000000000005d000000000000004f000000000000004c00000000",
            INIT_07 => X"00000068000000000000006c0000000000000058000000000000005300000000",
            INIT_08 => X"000000b800000000000000a700000000000000a600000000000000d700000000",
            INIT_09 => X"000000950000000000000060000000000000006600000000000000b600000000",
            INIT_0A => X"000000690000000000000074000000000000005d000000000000008900000000",
            INIT_0B => X"0000006e000000000000005b0000000000000069000000000000006600000000",
            INIT_0C => X"0000006000000000000000800000000000000067000000000000005b00000000",
            INIT_0D => X"00000045000000000000007e0000000000000078000000000000003800000000",
            INIT_0E => X"0000005d00000000000000460000000000000038000000000000003800000000",
            INIT_0F => X"0000006e00000000000000740000000000000070000000000000005e00000000",
            INIT_10 => X"000000b500000000000000af00000000000000b800000000000000d300000000",
            INIT_11 => X"0000008b0000000000000058000000000000008300000000000000b800000000",
            INIT_12 => X"00000040000000000000005a0000000000000080000000000000009400000000",
            INIT_13 => X"0000008f0000000000000075000000000000006f000000000000007900000000",
            INIT_14 => X"00000075000000000000008b0000000000000060000000000000005c00000000",
            INIT_15 => X"0000003b00000000000000440000000000000063000000000000006d00000000",
            INIT_16 => X"000000690000000000000045000000000000003e000000000000002900000000",
            INIT_17 => X"0000006f00000000000000730000000000000078000000000000007700000000",
            INIT_18 => X"000000b300000000000000b000000000000000bd00000000000000c000000000",
            INIT_19 => X"00000079000000000000005a000000000000009500000000000000b600000000",
            INIT_1A => X"0000003b00000000000000860000000000000088000000000000007c00000000",
            INIT_1B => X"000000b000000000000000860000000000000061000000000000007600000000",
            INIT_1C => X"0000007c0000000000000077000000000000004b000000000000007600000000",
            INIT_1D => X"0000003300000000000000310000000000000056000000000000008100000000",
            INIT_1E => X"00000076000000000000005b000000000000005a000000000000003100000000",
            INIT_1F => X"0000006b000000000000006f0000000000000071000000000000007900000000",
            INIT_20 => X"000000ad00000000000000b200000000000000c1000000000000009c00000000",
            INIT_21 => X"000000870000000000000067000000000000009d00000000000000b500000000",
            INIT_22 => X"0000004d000000000000005a000000000000006900000000000000af00000000",
            INIT_23 => X"000000b600000000000000ad0000000000000076000000000000005a00000000",
            INIT_24 => X"0000004d000000000000004e0000000000000064000000000000009400000000",
            INIT_25 => X"00000021000000000000002e0000000000000034000000000000003d00000000",
            INIT_26 => X"0000007d00000000000000640000000000000047000000000000003900000000",
            INIT_27 => X"000000690000000000000071000000000000006d000000000000007b00000000",
            INIT_28 => X"000000a900000000000000b200000000000000c8000000000000007800000000",
            INIT_29 => X"000000990000000000000057000000000000009000000000000000b300000000",
            INIT_2A => X"0000008d000000000000008c00000000000000de00000000000000f700000000",
            INIT_2B => X"000000c000000000000000c400000000000000b6000000000000009c00000000",
            INIT_2C => X"0000003e000000000000006d000000000000008500000000000000ac00000000",
            INIT_2D => X"0000005100000000000000460000000000000036000000000000003100000000",
            INIT_2E => X"0000006500000000000000630000000000000054000000000000005500000000",
            INIT_2F => X"0000005a000000000000005c0000000000000060000000000000006800000000",
            INIT_30 => X"000000ac00000000000000b700000000000000c5000000000000006900000000",
            INIT_31 => X"000000d30000000000000070000000000000009200000000000000b100000000",
            INIT_32 => X"0000008f00000000000000e000000000000000fd00000000000000fc00000000",
            INIT_33 => X"000000850000000000000085000000000000008d000000000000008400000000",
            INIT_34 => X"000000520000000000000057000000000000005d000000000000007c00000000",
            INIT_35 => X"0000005d00000000000000550000000000000054000000000000005400000000",
            INIT_36 => X"000000680000000000000060000000000000005b000000000000005e00000000",
            INIT_37 => X"0000005f00000000000000610000000000000061000000000000006c00000000",
            INIT_38 => X"000000ae00000000000000a80000000000000089000000000000005900000000",
            INIT_39 => X"000000f500000000000000a600000000000000aa00000000000000b600000000",
            INIT_3A => X"00000058000000000000008800000000000000e700000000000000fb00000000",
            INIT_3B => X"00000048000000000000004b000000000000004c000000000000005000000000",
            INIT_3C => X"0000005200000000000000510000000000000051000000000000004f00000000",
            INIT_3D => X"000000570000000000000059000000000000005a000000000000005600000000",
            INIT_3E => X"00000060000000000000005e000000000000005d000000000000005900000000",
            INIT_3F => X"0000005a000000000000005f000000000000005e000000000000006000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009900000000000000660000000000000057000000000000005b00000000",
            INIT_41 => X"000000fa00000000000000bd000000000000008800000000000000b300000000",
            INIT_42 => X"00000054000000000000005e000000000000009f00000000000000f500000000",
            INIT_43 => X"0000005400000000000000530000000000000055000000000000005400000000",
            INIT_44 => X"0000004f00000000000000520000000000000054000000000000005600000000",
            INIT_45 => X"0000005900000000000000550000000000000056000000000000005300000000",
            INIT_46 => X"0000006500000000000000670000000000000067000000000000005c00000000",
            INIT_47 => X"00000067000000000000005e0000000000000063000000000000006600000000",
            INIT_48 => X"0000006a0000000000000055000000000000005e000000000000006f00000000",
            INIT_49 => X"000000fd00000000000000d50000000000000088000000000000009400000000",
            INIT_4A => X"00000058000000000000005b000000000000005d00000000000000c600000000",
            INIT_4B => X"000000520000000000000053000000000000005a000000000000005a00000000",
            INIT_4C => X"0000005300000000000000500000000000000051000000000000005200000000",
            INIT_4D => X"0000005f000000000000005c0000000000000059000000000000005600000000",
            INIT_4E => X"0000006c000000000000006d000000000000006e000000000000006c00000000",
            INIT_4F => X"00000089000000000000007b0000000000000069000000000000006c00000000",
            INIT_50 => X"0000005300000000000000560000000000000063000000000000007200000000",
            INIT_51 => X"000000f500000000000000e50000000000000091000000000000005f00000000",
            INIT_52 => X"0000005e0000000000000057000000000000005c000000000000008f00000000",
            INIT_53 => X"0000005300000000000000520000000000000052000000000000005c00000000",
            INIT_54 => X"0000005800000000000000560000000000000053000000000000005400000000",
            INIT_55 => X"0000006e000000000000006a0000000000000061000000000000005a00000000",
            INIT_56 => X"0000005b000000000000005f0000000000000061000000000000006900000000",
            INIT_57 => X"0000007d000000000000008a0000000000000082000000000000006c00000000",
            INIT_58 => X"0000005600000000000000590000000000000062000000000000006e00000000",
            INIT_59 => X"000000e400000000000000db000000000000006a000000000000005300000000",
            INIT_5A => X"00000057000000000000005e0000000000000068000000000000007e00000000",
            INIT_5B => X"0000005200000000000000500000000000000057000000000000006100000000",
            INIT_5C => X"0000005900000000000000590000000000000057000000000000005400000000",
            INIT_5D => X"00000066000000000000005d000000000000005c000000000000006100000000",
            INIT_5E => X"000000650000000000000055000000000000005d000000000000006500000000",
            INIT_5F => X"000000600000000000000062000000000000007e000000000000008100000000",
            INIT_60 => X"00000058000000000000005c0000000000000061000000000000006c00000000",
            INIT_61 => X"000000c500000000000000850000000000000054000000000000005800000000",
            INIT_62 => X"0000005f000000000000005e0000000000000061000000000000006400000000",
            INIT_63 => X"0000005300000000000000600000000000000064000000000000006700000000",
            INIT_64 => X"0000005c00000000000000580000000000000050000000000000004f00000000",
            INIT_65 => X"0000005c000000000000005d000000000000005f000000000000005c00000000",
            INIT_66 => X"0000007d0000000000000066000000000000005d000000000000005a00000000",
            INIT_67 => X"0000005d000000000000003c000000000000005a000000000000006e00000000",
            INIT_68 => X"0000005b00000000000000580000000000000064000000000000007c00000000",
            INIT_69 => X"0000006b000000000000004f0000000000000059000000000000005700000000",
            INIT_6A => X"000000520000000000000047000000000000004d000000000000005900000000",
            INIT_6B => X"0000005c00000000000000660000000000000064000000000000005d00000000",
            INIT_6C => X"0000006100000000000000630000000000000063000000000000005e00000000",
            INIT_6D => X"000000530000000000000058000000000000005e000000000000005f00000000",
            INIT_6E => X"0000008300000000000000840000000000000070000000000000005b00000000",
            INIT_6F => X"0000005500000000000000400000000000000061000000000000007400000000",
            INIT_70 => X"0000005b00000000000000550000000000000066000000000000007400000000",
            INIT_71 => X"000000510000000000000058000000000000005c000000000000005a00000000",
            INIT_72 => X"0000004a00000000000000430000000000000048000000000000005500000000",
            INIT_73 => X"0000005600000000000000500000000000000049000000000000004700000000",
            INIT_74 => X"00000077000000000000006d0000000000000065000000000000005f00000000",
            INIT_75 => X"000000580000000000000058000000000000005f000000000000007100000000",
            INIT_76 => X"00000091000000000000009c0000000000000082000000000000006900000000",
            INIT_77 => X"0000004000000000000000520000000000000052000000000000007300000000",
            INIT_78 => X"0000005600000000000000590000000000000069000000000000006b00000000",
            INIT_79 => X"000000510000000000000057000000000000005c000000000000005900000000",
            INIT_7A => X"0000004900000000000000420000000000000045000000000000004f00000000",
            INIT_7B => X"0000003a000000000000003f0000000000000049000000000000004500000000",
            INIT_7C => X"0000007700000000000000680000000000000057000000000000004600000000",
            INIT_7D => X"00000057000000000000005f0000000000000060000000000000006f00000000",
            INIT_7E => X"0000008700000000000000920000000000000083000000000000006d00000000",
            INIT_7F => X"000000430000000000000054000000000000004d000000000000006300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE3;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE4 : if BRAM_NAME = "sampleifmap_layersamples_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000350000000000000033000000000000002f000000000000003100000000",
            INIT_01 => X"0000002d000000000000002f0000000000000029000000000000002e00000000",
            INIT_02 => X"0000003400000000000000290000000000000029000000000000002c00000000",
            INIT_03 => X"0000002c000000000000002d0000000000000029000000000000003100000000",
            INIT_04 => X"0000002b00000000000000270000000000000026000000000000002800000000",
            INIT_05 => X"0000002b000000000000002d000000000000002d000000000000002c00000000",
            INIT_06 => X"00000029000000000000002b0000000000000027000000000000002c00000000",
            INIT_07 => X"0000002100000000000000240000000000000024000000000000002600000000",
            INIT_08 => X"00000038000000000000002d0000000000000028000000000000003300000000",
            INIT_09 => X"0000002d000000000000002f000000000000002b000000000000003100000000",
            INIT_0A => X"0000003600000000000000290000000000000026000000000000002e00000000",
            INIT_0B => X"0000002100000000000000280000000000000029000000000000003400000000",
            INIT_0C => X"0000003200000000000000290000000000000021000000000000001e00000000",
            INIT_0D => X"0000003000000000000000340000000000000037000000000000003500000000",
            INIT_0E => X"00000026000000000000002d000000000000002e000000000000003200000000",
            INIT_0F => X"000000220000000000000020000000000000001f000000000000002200000000",
            INIT_10 => X"0000003000000000000000240000000000000021000000000000002f00000000",
            INIT_11 => X"0000002d000000000000002d000000000000002c000000000000002a00000000",
            INIT_12 => X"000000390000000000000030000000000000002b000000000000002b00000000",
            INIT_13 => X"0000002300000000000000250000000000000026000000000000003300000000",
            INIT_14 => X"000000310000000000000036000000000000002f000000000000002700000000",
            INIT_15 => X"00000032000000000000002f0000000000000032000000000000003400000000",
            INIT_16 => X"0000002700000000000000330000000000000037000000000000003000000000",
            INIT_17 => X"0000002100000000000000220000000000000022000000000000002300000000",
            INIT_18 => X"0000002c000000000000001f0000000000000020000000000000002800000000",
            INIT_19 => X"000000300000000000000030000000000000002e000000000000002b00000000",
            INIT_1A => X"0000005f0000000000000039000000000000002d000000000000002c00000000",
            INIT_1B => X"00000036000000000000002f0000000000000029000000000000004b00000000",
            INIT_1C => X"00000041000000000000002f0000000000000043000000000000003a00000000",
            INIT_1D => X"0000003200000000000000420000000000000054000000000000004c00000000",
            INIT_1E => X"0000002e000000000000002d0000000000000027000000000000003400000000",
            INIT_1F => X"0000002400000000000000270000000000000027000000000000002b00000000",
            INIT_20 => X"0000002f00000000000000310000000000000030000000000000002900000000",
            INIT_21 => X"0000002c000000000000002f0000000000000028000000000000002b00000000",
            INIT_22 => X"000000a4000000000000003b000000000000002a000000000000002900000000",
            INIT_23 => X"00000047000000000000003c0000000000000038000000000000006b00000000",
            INIT_24 => X"000000620000000000000038000000000000001f000000000000003200000000",
            INIT_25 => X"0000005d00000000000000690000000000000076000000000000006f00000000",
            INIT_26 => X"0000002d000000000000002f0000000000000046000000000000004300000000",
            INIT_27 => X"000000240000000000000024000000000000002e000000000000003000000000",
            INIT_28 => X"0000003500000000000000390000000000000040000000000000003600000000",
            INIT_29 => X"0000002900000000000000290000000000000027000000000000002c00000000",
            INIT_2A => X"00000055000000000000002a0000000000000027000000000000002500000000",
            INIT_2B => X"0000001f000000000000002b000000000000003a000000000000004e00000000",
            INIT_2C => X"0000006e000000000000004c000000000000002d000000000000002b00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007800000000",
            INIT_2E => X"00000025000000000000002f0000000000000056000000000000006100000000",
            INIT_2F => X"00000028000000000000002c000000000000003a000000000000003100000000",
            INIT_30 => X"0000001c00000000000000110000000000000050000000000000003900000000",
            INIT_31 => X"0000002b0000000000000028000000000000002b000000000000003000000000",
            INIT_32 => X"0000003400000000000000270000000000000025000000000000002a00000000",
            INIT_33 => X"000000390000000000000046000000000000004b000000000000003b00000000",
            INIT_34 => X"00000079000000000000004a0000000000000040000000000000004800000000",
            INIT_35 => X"0000005e000000000000005a000000000000006c000000000000008400000000",
            INIT_36 => X"000000270000000000000045000000000000004d000000000000006700000000",
            INIT_37 => X"000000270000000000000030000000000000003a000000000000002400000000",
            INIT_38 => X"000000290000000000000026000000000000005c000000000000005a00000000",
            INIT_39 => X"000000270000000000000024000000000000002a000000000000003800000000",
            INIT_3A => X"0000003100000000000000330000000000000033000000000000003100000000",
            INIT_3B => X"0000004f000000000000005d000000000000006b000000000000004d00000000",
            INIT_3C => X"0000006b00000000000000450000000000000052000000000000005800000000",
            INIT_3D => X"0000005800000000000000510000000000000070000000000000008c00000000",
            INIT_3E => X"00000031000000000000003a000000000000004a000000000000005400000000",
            INIT_3F => X"0000002700000000000000330000000000000032000000000000002000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000071000000000000003b0000000000000069000000000000009000000000",
            INIT_41 => X"000000320000000000000029000000000000002b000000000000005200000000",
            INIT_42 => X"0000004e000000000000003b000000000000005f000000000000004200000000",
            INIT_43 => X"0000004a00000000000000650000000000000080000000000000007900000000",
            INIT_44 => X"0000003d00000000000000490000000000000052000000000000004d00000000",
            INIT_45 => X"00000046000000000000005d000000000000007b000000000000007000000000",
            INIT_46 => X"000000350000000000000043000000000000004c000000000000004500000000",
            INIT_47 => X"0000002d000000000000003b0000000000000023000000000000001b00000000",
            INIT_48 => X"000000950000000000000069000000000000008f00000000000000a300000000",
            INIT_49 => X"0000003c000000000000002f0000000000000033000000000000007000000000",
            INIT_4A => X"0000007700000000000000a600000000000000c6000000000000009200000000",
            INIT_4B => X"0000004f000000000000006b000000000000007d000000000000009100000000",
            INIT_4C => X"0000003a00000000000000350000000000000047000000000000004f00000000",
            INIT_4D => X"000000590000000000000072000000000000007a000000000000007000000000",
            INIT_4E => X"00000047000000000000004e000000000000004e000000000000004a00000000",
            INIT_4F => X"00000039000000000000002c000000000000000f000000000000002b00000000",
            INIT_50 => X"000000a8000000000000009e000000000000007a00000000000000af00000000",
            INIT_51 => X"0000002f00000000000000330000000000000032000000000000007a00000000",
            INIT_52 => X"0000008300000000000000bc00000000000000e200000000000000b300000000",
            INIT_53 => X"0000006800000000000000680000000000000084000000000000009b00000000",
            INIT_54 => X"0000004d0000000000000028000000000000004d000000000000004500000000",
            INIT_55 => X"0000005c000000000000008a0000000000000089000000000000009a00000000",
            INIT_56 => X"00000049000000000000004f0000000000000060000000000000004d00000000",
            INIT_57 => X"0000002e000000000000001f0000000000000021000000000000003b00000000",
            INIT_58 => X"000000b20000000000000099000000000000007400000000000000bd00000000",
            INIT_59 => X"0000002c0000000000000037000000000000003b000000000000008800000000",
            INIT_5A => X"0000008500000000000000a400000000000000bc000000000000005000000000",
            INIT_5B => X"0000005f000000000000006a000000000000009f000000000000009700000000",
            INIT_5C => X"000000710000000000000022000000000000004f000000000000005900000000",
            INIT_5D => X"000000520000000000000082000000000000008e00000000000000c000000000",
            INIT_5E => X"00000051000000000000005e0000000000000058000000000000004b00000000",
            INIT_5F => X"0000001a00000000000000300000000000000037000000000000004e00000000",
            INIT_60 => X"000000b90000000000000090000000000000006900000000000000c200000000",
            INIT_61 => X"0000002f00000000000000350000000000000044000000000000008500000000",
            INIT_62 => X"0000005e000000000000007e0000000000000098000000000000002c00000000",
            INIT_63 => X"00000062000000000000008100000000000000b7000000000000009400000000",
            INIT_64 => X"0000008c000000000000002f000000000000006d000000000000006900000000",
            INIT_65 => X"00000053000000000000006f000000000000008c00000000000000b200000000",
            INIT_66 => X"0000005100000000000000550000000000000050000000000000004f00000000",
            INIT_67 => X"0000001800000000000000400000000000000049000000000000005900000000",
            INIT_68 => X"000000c000000000000000a3000000000000006700000000000000c100000000",
            INIT_69 => X"00000032000000000000003a0000000000000042000000000000006200000000",
            INIT_6A => X"0000007f00000000000000670000000000000078000000000000002700000000",
            INIT_6B => X"00000075000000000000009d00000000000000c8000000000000009b00000000",
            INIT_6C => X"000000930000000000000044000000000000006d000000000000006b00000000",
            INIT_6D => X"000000500000000000000068000000000000008800000000000000ae00000000",
            INIT_6E => X"0000005e00000000000000480000000000000046000000000000004c00000000",
            INIT_6F => X"0000002200000000000000450000000000000051000000000000006300000000",
            INIT_70 => X"000000bc00000000000000ac000000000000007000000000000000c400000000",
            INIT_71 => X"00000037000000000000003e0000000000000043000000000000006d00000000",
            INIT_72 => X"000000a900000000000000670000000000000058000000000000002200000000",
            INIT_73 => X"00000086000000000000008c000000000000009f00000000000000a900000000",
            INIT_74 => X"000000950000000000000046000000000000005f000000000000007d00000000",
            INIT_75 => X"00000069000000000000007a000000000000007f00000000000000aa00000000",
            INIT_76 => X"00000068000000000000005a000000000000005b000000000000005300000000",
            INIT_77 => X"0000002f00000000000000350000000000000050000000000000006f00000000",
            INIT_78 => X"000000b500000000000000ae000000000000008800000000000000c500000000",
            INIT_79 => X"0000004d0000000000000058000000000000004d000000000000008e00000000",
            INIT_7A => X"000000d30000000000000074000000000000005d000000000000003400000000",
            INIT_7B => X"000000700000000000000082000000000000008900000000000000e600000000",
            INIT_7C => X"00000076000000000000004b000000000000005f000000000000006500000000",
            INIT_7D => X"000000500000000000000065000000000000008a000000000000009200000000",
            INIT_7E => X"0000006300000000000000630000000000000057000000000000004400000000",
            INIT_7F => X"0000003000000000000000300000000000000036000000000000005d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE4;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE5 : if BRAM_NAME = "sampleifmap_layersamples_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bc00000000000000b200000000000000a000000000000000cc00000000",
            INIT_01 => X"00000071000000000000007e000000000000005a00000000000000ac00000000",
            INIT_02 => X"0000009b00000000000000850000000000000025000000000000005200000000",
            INIT_03 => X"0000005a00000000000000580000000000000075000000000000008d00000000",
            INIT_04 => X"00000068000000000000003a0000000000000057000000000000005c00000000",
            INIT_05 => X"000000610000000000000076000000000000007e000000000000006d00000000",
            INIT_06 => X"00000052000000000000005e000000000000004d000000000000004800000000",
            INIT_07 => X"0000002e0000000000000037000000000000002d000000000000003700000000",
            INIT_08 => X"000000c200000000000000b800000000000000b400000000000000d700000000",
            INIT_09 => X"000000910000000000000066000000000000006900000000000000ba00000000",
            INIT_0A => X"0000005f0000000000000069000000000000003d000000000000006f00000000",
            INIT_0B => X"0000006200000000000000490000000000000059000000000000005900000000",
            INIT_0C => X"000000400000000000000066000000000000005f000000000000005800000000",
            INIT_0D => X"0000003d00000000000000730000000000000069000000000000002000000000",
            INIT_0E => X"0000004e00000000000000410000000000000035000000000000003300000000",
            INIT_0F => X"0000003600000000000000400000000000000044000000000000004000000000",
            INIT_10 => X"000000c100000000000000bd00000000000000c000000000000000cd00000000",
            INIT_11 => X"0000008f0000000000000060000000000000008500000000000000bc00000000",
            INIT_12 => X"000000370000000000000050000000000000006f000000000000008d00000000",
            INIT_13 => X"0000008500000000000000640000000000000060000000000000006c00000000",
            INIT_14 => X"0000005d0000000000000078000000000000005d000000000000005d00000000",
            INIT_15 => X"00000034000000000000003a0000000000000056000000000000005c00000000",
            INIT_16 => X"0000003b0000000000000028000000000000003c000000000000002700000000",
            INIT_17 => X"0000002e000000000000002d0000000000000036000000000000003e00000000",
            INIT_18 => X"000000b900000000000000b500000000000000bb00000000000000b400000000",
            INIT_19 => X"000000840000000000000063000000000000009800000000000000b800000000",
            INIT_1A => X"00000033000000000000007e0000000000000087000000000000008200000000",
            INIT_1B => X"000000a8000000000000007b0000000000000056000000000000006c00000000",
            INIT_1C => X"0000006900000000000000670000000000000049000000000000007600000000",
            INIT_1D => X"00000032000000000000002c000000000000004e000000000000007600000000",
            INIT_1E => X"00000044000000000000003c000000000000005d000000000000003400000000",
            INIT_1F => X"0000002e00000000000000320000000000000034000000000000004000000000",
            INIT_20 => X"000000ac00000000000000af00000000000000bb000000000000009200000000",
            INIT_21 => X"00000092000000000000006f00000000000000a000000000000000b400000000",
            INIT_22 => X"000000490000000000000057000000000000006f00000000000000b900000000",
            INIT_23 => X"000000b100000000000000ad0000000000000074000000000000005600000000",
            INIT_24 => X"0000003f00000000000000420000000000000065000000000000009400000000",
            INIT_25 => X"0000002900000000000000330000000000000036000000000000003900000000",
            INIT_26 => X"00000052000000000000004b0000000000000053000000000000004500000000",
            INIT_27 => X"0000003f0000000000000045000000000000003d000000000000004c00000000",
            INIT_28 => X"000000a800000000000000b000000000000000c8000000000000007c00000000",
            INIT_29 => X"0000009f000000000000005b000000000000009300000000000000b300000000",
            INIT_2A => X"00000093000000000000009000000000000000e100000000000000fa00000000",
            INIT_2B => X"000000c500000000000000d000000000000000c000000000000000a400000000",
            INIT_2C => X"0000003e000000000000006d000000000000008f00000000000000b500000000",
            INIT_2D => X"0000006600000000000000570000000000000044000000000000003a00000000",
            INIT_2E => X"00000077000000000000007a000000000000006f000000000000006e00000000",
            INIT_2F => X"0000007300000000000000700000000000000070000000000000007800000000",
            INIT_30 => X"000000b100000000000000c000000000000000d5000000000000008500000000",
            INIT_31 => X"000000d10000000000000071000000000000009600000000000000b600000000",
            INIT_32 => X"0000009d00000000000000e800000000000000fc00000000000000f700000000",
            INIT_33 => X"00000098000000000000009c00000000000000a2000000000000009500000000",
            INIT_34 => X"0000006500000000000000680000000000000077000000000000009400000000",
            INIT_35 => X"0000007d0000000000000073000000000000006e000000000000006f00000000",
            INIT_36 => X"0000008d00000000000000870000000000000082000000000000008300000000",
            INIT_37 => X"0000008400000000000000890000000000000084000000000000008e00000000",
            INIT_38 => X"000000bc00000000000000bc00000000000000a8000000000000008700000000",
            INIT_39 => X"000000ed00000000000000a400000000000000ae00000000000000c000000000",
            INIT_3A => X"0000006f000000000000009900000000000000e400000000000000f100000000",
            INIT_3B => X"00000065000000000000006b0000000000000069000000000000006900000000",
            INIT_3C => X"0000007400000000000000710000000000000078000000000000007300000000",
            INIT_3D => X"00000080000000000000007e000000000000007d000000000000007d00000000",
            INIT_3E => X"000000890000000000000089000000000000008b000000000000008400000000",
            INIT_3F => X"00000085000000000000008b0000000000000086000000000000008700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b000000000000000860000000000000082000000000000008d00000000",
            INIT_41 => X"000000f200000000000000b5000000000000008900000000000000bf00000000",
            INIT_42 => X"00000076000000000000007f00000000000000af00000000000000f500000000",
            INIT_43 => X"0000007400000000000000780000000000000079000000000000007700000000",
            INIT_44 => X"0000007100000000000000730000000000000075000000000000007500000000",
            INIT_45 => X"00000082000000000000007d000000000000007d000000000000007800000000",
            INIT_46 => X"0000008e000000000000008e0000000000000091000000000000008600000000",
            INIT_47 => X"00000095000000000000008c0000000000000090000000000000009200000000",
            INIT_48 => X"00000088000000000000007c000000000000008c00000000000000a200000000",
            INIT_49 => X"000000f900000000000000d1000000000000008f00000000000000a700000000",
            INIT_4A => X"0000007d0000000000000080000000000000007600000000000000cd00000000",
            INIT_4B => X"000000730000000000000079000000000000007f000000000000007f00000000",
            INIT_4C => X"0000007500000000000000710000000000000070000000000000007100000000",
            INIT_4D => X"0000008a00000000000000860000000000000083000000000000007b00000000",
            INIT_4E => X"0000009500000000000000930000000000000098000000000000009600000000",
            INIT_4F => X"000000b600000000000000a70000000000000098000000000000009a00000000",
            INIT_50 => X"0000007a0000000000000082000000000000009300000000000000a500000000",
            INIT_51 => X"000000f700000000000000ea00000000000000a4000000000000007e00000000",
            INIT_52 => X"00000083000000000000007b0000000000000072000000000000009900000000",
            INIT_53 => X"0000007700000000000000770000000000000077000000000000008100000000",
            INIT_54 => X"0000007f000000000000007b0000000000000077000000000000007700000000",
            INIT_55 => X"0000009a0000000000000096000000000000008d000000000000008300000000",
            INIT_56 => X"0000008a000000000000008c000000000000008d000000000000009600000000",
            INIT_57 => X"000000a900000000000000b600000000000000b2000000000000009e00000000",
            INIT_58 => X"00000085000000000000008a000000000000009500000000000000a200000000",
            INIT_59 => X"000000ea00000000000000e9000000000000008a000000000000007e00000000",
            INIT_5A => X"0000007c0000000000000081000000000000007e000000000000008c00000000",
            INIT_5B => X"000000770000000000000074000000000000007b000000000000008500000000",
            INIT_5C => X"000000840000000000000082000000000000007e000000000000007a00000000",
            INIT_5D => X"00000094000000000000008b000000000000008a000000000000008c00000000",
            INIT_5E => X"000000990000000000000085000000000000008b000000000000009300000000",
            INIT_5F => X"0000008b000000000000008e00000000000000b000000000000000b600000000",
            INIT_60 => X"0000008d000000000000008f000000000000009300000000000000a100000000",
            INIT_61 => X"000000d3000000000000009f000000000000007d000000000000008a00000000",
            INIT_62 => X"0000008200000000000000800000000000000079000000000000007700000000",
            INIT_63 => X"0000007800000000000000830000000000000087000000000000008b00000000",
            INIT_64 => X"0000008700000000000000820000000000000078000000000000007600000000",
            INIT_65 => X"00000088000000000000008a000000000000008b000000000000008800000000",
            INIT_66 => X"000000b20000000000000097000000000000008a000000000000008700000000",
            INIT_67 => X"000000880000000000000067000000000000008c00000000000000a400000000",
            INIT_68 => X"000000920000000000000089000000000000009400000000000000b100000000",
            INIT_69 => X"0000008500000000000000710000000000000084000000000000008b00000000",
            INIT_6A => X"0000007500000000000000690000000000000069000000000000007200000000",
            INIT_6B => X"0000008000000000000000890000000000000087000000000000008000000000",
            INIT_6C => X"0000008a000000000000008b0000000000000089000000000000008300000000",
            INIT_6D => X"0000007d00000000000000830000000000000088000000000000008900000000",
            INIT_6E => X"000000b500000000000000b3000000000000009a000000000000008500000000",
            INIT_6F => X"0000007f000000000000006c000000000000009200000000000000a800000000",
            INIT_70 => X"0000008f0000000000000084000000000000009400000000000000a800000000",
            INIT_71 => X"00000070000000000000007d0000000000000086000000000000008b00000000",
            INIT_72 => X"0000006d00000000000000660000000000000068000000000000007300000000",
            INIT_73 => X"000000780000000000000073000000000000006c000000000000006a00000000",
            INIT_74 => X"0000009c00000000000000900000000000000087000000000000008000000000",
            INIT_75 => X"0000007f000000000000007f0000000000000086000000000000009800000000",
            INIT_76 => X"000000be00000000000000c500000000000000aa000000000000009000000000",
            INIT_77 => X"0000006b000000000000007e000000000000008200000000000000a400000000",
            INIT_78 => X"000000860000000000000084000000000000009500000000000000a000000000",
            INIT_79 => X"00000073000000000000007b0000000000000084000000000000008600000000",
            INIT_7A => X"0000006c00000000000000650000000000000069000000000000007200000000",
            INIT_7B => X"000000590000000000000062000000000000006c000000000000006800000000",
            INIT_7C => X"0000009800000000000000890000000000000076000000000000006400000000",
            INIT_7D => X"0000007b00000000000000820000000000000083000000000000009100000000",
            INIT_7E => X"000000af00000000000000b600000000000000a7000000000000009100000000",
            INIT_7F => X"0000006e0000000000000081000000000000007c000000000000009100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE5;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE6 : if BRAM_NAME = "sampleifmap_layersamples_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e800000000000000e800000000000000e700000000000000eb00000000",
            INIT_01 => X"000000e800000000000000e800000000000000e800000000000000e800000000",
            INIT_02 => X"000000e900000000000000e900000000000000e800000000000000e800000000",
            INIT_03 => X"000000e900000000000000e900000000000000e900000000000000e900000000",
            INIT_04 => X"000000e600000000000000e700000000000000e800000000000000e900000000",
            INIT_05 => X"000000e900000000000000e800000000000000e800000000000000e800000000",
            INIT_06 => X"000000e800000000000000e800000000000000e900000000000000e800000000",
            INIT_07 => X"000000e800000000000000e900000000000000e900000000000000e800000000",
            INIT_08 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_09 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_0A => X"000000ec00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_0B => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_0C => X"000000ea00000000000000ec00000000000000ec00000000000000ed00000000",
            INIT_0D => X"000000ec00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_0E => X"000000eb00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_0F => X"000000eb00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_10 => X"000000ea00000000000000ea00000000000000ea00000000000000ed00000000",
            INIT_11 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_12 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_13 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_14 => X"000000ea00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_15 => X"000000ea00000000000000e700000000000000e700000000000000e300000000",
            INIT_16 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_17 => X"000000ea00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_18 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_19 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_1A => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_1B => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_1C => X"000000df00000000000000e400000000000000e800000000000000e900000000",
            INIT_1D => X"000000e400000000000000cf00000000000000d100000000000000ba00000000",
            INIT_1E => X"000000ea00000000000000ea00000000000000ea00000000000000ec00000000",
            INIT_1F => X"000000eb00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_20 => X"000000eb00000000000000eb00000000000000ea00000000000000ed00000000",
            INIT_21 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_22 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_23 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_24 => X"000000cb00000000000000db00000000000000e900000000000000ec00000000",
            INIT_25 => X"000000e600000000000000d600000000000000c300000000000000a300000000",
            INIT_26 => X"000000eb00000000000000eb00000000000000eb00000000000000ed00000000",
            INIT_27 => X"000000ec00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_28 => X"000000ec00000000000000ec00000000000000ec00000000000000ef00000000",
            INIT_29 => X"000000eb00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_2A => X"000000ed00000000000000ed00000000000000eb00000000000000ea00000000",
            INIT_2B => X"000000e500000000000000eb00000000000000e800000000000000ea00000000",
            INIT_2C => X"000000ae00000000000000b900000000000000c200000000000000d000000000",
            INIT_2D => X"000000e200000000000000cf00000000000000b800000000000000a500000000",
            INIT_2E => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_2F => X"000000ed00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_30 => X"000000e700000000000000e800000000000000e400000000000000e400000000",
            INIT_31 => X"000000ec00000000000000ed00000000000000ed00000000000000ea00000000",
            INIT_32 => X"000000ef00000000000000ef00000000000000ed00000000000000ed00000000",
            INIT_33 => X"000000dd00000000000000e900000000000000e000000000000000e100000000",
            INIT_34 => X"0000009a000000000000009f00000000000000a100000000000000b700000000",
            INIT_35 => X"000000c6000000000000009c000000000000008f000000000000009000000000",
            INIT_36 => X"000000eb00000000000000eb00000000000000ec00000000000000e900000000",
            INIT_37 => X"000000ef00000000000000ed00000000000000ec00000000000000eb00000000",
            INIT_38 => X"000000e300000000000000e600000000000000e000000000000000d400000000",
            INIT_39 => X"000000ee00000000000000ed00000000000000ea00000000000000e500000000",
            INIT_3A => X"000000f000000000000000ef00000000000000ef00000000000000ef00000000",
            INIT_3B => X"000000d600000000000000e900000000000000db00000000000000c900000000",
            INIT_3C => X"000000ad00000000000000b800000000000000b900000000000000c100000000",
            INIT_3D => X"000000ba00000000000000a2000000000000009f00000000000000a500000000",
            INIT_3E => X"000000e900000000000000e900000000000000ea00000000000000e500000000",
            INIT_3F => X"000000ee00000000000000ed00000000000000ec00000000000000ea00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000e100000000000000e100000000000000dd00000000000000d800000000",
            INIT_41 => X"000000ee00000000000000ec00000000000000e700000000000000e300000000",
            INIT_42 => X"000000ef00000000000000ed00000000000000ee00000000000000ee00000000",
            INIT_43 => X"000000e600000000000000e900000000000000dc00000000000000c500000000",
            INIT_44 => X"000000d000000000000000db00000000000000d100000000000000d100000000",
            INIT_45 => X"000000da00000000000000d900000000000000d200000000000000d100000000",
            INIT_46 => X"000000e600000000000000e400000000000000e400000000000000e100000000",
            INIT_47 => X"000000ee00000000000000ed00000000000000eb00000000000000e600000000",
            INIT_48 => X"00000088000000000000007c0000000000000077000000000000007600000000",
            INIT_49 => X"000000ed00000000000000eb00000000000000e100000000000000ac00000000",
            INIT_4A => X"000000e900000000000000eb00000000000000eb00000000000000ec00000000",
            INIT_4B => X"000000ec00000000000000e800000000000000e200000000000000d600000000",
            INIT_4C => X"000000e100000000000000e700000000000000e300000000000000e400000000",
            INIT_4D => X"000000b900000000000000c900000000000000d900000000000000e100000000",
            INIT_4E => X"000000ba00000000000000a700000000000000a700000000000000ac00000000",
            INIT_4F => X"000000ee00000000000000ec00000000000000eb00000000000000df00000000",
            INIT_50 => X"0000006f000000000000006c0000000000000067000000000000006d00000000",
            INIT_51 => X"000000e500000000000000e300000000000000de000000000000009200000000",
            INIT_52 => X"000000e600000000000000e700000000000000ea00000000000000ec00000000",
            INIT_53 => X"000000e600000000000000e800000000000000e700000000000000e500000000",
            INIT_54 => X"000000df00000000000000e500000000000000e700000000000000e700000000",
            INIT_55 => X"00000089000000000000009200000000000000a400000000000000bf00000000",
            INIT_56 => X"0000009500000000000000790000000000000080000000000000008600000000",
            INIT_57 => X"000000ed00000000000000eb00000000000000ea00000000000000d800000000",
            INIT_58 => X"000000c800000000000000c700000000000000bc00000000000000c300000000",
            INIT_59 => X"000000d300000000000000d500000000000000df00000000000000d100000000",
            INIT_5A => X"000000d200000000000000db00000000000000dc00000000000000d800000000",
            INIT_5B => X"000000dc00000000000000d800000000000000d300000000000000d100000000",
            INIT_5C => X"000000da00000000000000e100000000000000e200000000000000e100000000",
            INIT_5D => X"000000b200000000000000b500000000000000af00000000000000b700000000",
            INIT_5E => X"000000b9000000000000008e00000000000000aa00000000000000ba00000000",
            INIT_5F => X"000000ec00000000000000ea00000000000000e700000000000000db00000000",
            INIT_60 => X"000000d600000000000000ca00000000000000bf00000000000000c100000000",
            INIT_61 => X"000000ab00000000000000cb00000000000000d600000000000000df00000000",
            INIT_62 => X"0000006200000000000000ae00000000000000cf00000000000000b100000000",
            INIT_63 => X"0000007a000000000000006f0000000000000065000000000000005d00000000",
            INIT_64 => X"000000df00000000000000ca0000000000000099000000000000008900000000",
            INIT_65 => X"000000d900000000000000df00000000000000dc00000000000000da00000000",
            INIT_66 => X"000000de00000000000000c400000000000000d400000000000000dd00000000",
            INIT_67 => X"000000eb00000000000000e800000000000000dd00000000000000db00000000",
            INIT_68 => X"0000007d0000000000000071000000000000006f000000000000007100000000",
            INIT_69 => X"000000be00000000000000bf00000000000000aa000000000000008a00000000",
            INIT_6A => X"00000036000000000000009e00000000000000d800000000000000d000000000",
            INIT_6B => X"0000004200000000000000350000000000000031000000000000002d00000000",
            INIT_6C => X"000000ea00000000000000dd000000000000009f000000000000006600000000",
            INIT_6D => X"000000cf00000000000000df00000000000000e300000000000000e900000000",
            INIT_6E => X"000000c700000000000000d400000000000000d300000000000000ca00000000",
            INIT_6F => X"000000dd00000000000000d300000000000000bc00000000000000b300000000",
            INIT_70 => X"00000044000000000000003f0000000000000045000000000000003d00000000",
            INIT_71 => X"000000c30000000000000097000000000000008b000000000000007b00000000",
            INIT_72 => X"0000006700000000000000a300000000000000ce00000000000000d600000000",
            INIT_73 => X"000000b5000000000000008a0000000000000065000000000000005f00000000",
            INIT_74 => X"000000cd00000000000000db00000000000000dd00000000000000cf00000000",
            INIT_75 => X"000000830000000000000093000000000000009e00000000000000b700000000",
            INIT_76 => X"0000008500000000000000880000000000000082000000000000007d00000000",
            INIT_77 => X"000000c500000000000000b6000000000000008a000000000000008000000000",
            INIT_78 => X"0000007f0000000000000055000000000000003a000000000000002800000000",
            INIT_79 => X"000000a300000000000000770000000000000060000000000000008400000000",
            INIT_7A => X"000000b500000000000000b600000000000000b800000000000000ad00000000",
            INIT_7B => X"000000c800000000000000da00000000000000c600000000000000b700000000",
            INIT_7C => X"000000840000000000000091000000000000009f00000000000000ae00000000",
            INIT_7D => X"00000063000000000000005e0000000000000062000000000000007400000000",
            INIT_7E => X"0000008a000000000000007a000000000000006b000000000000006900000000",
            INIT_7F => X"000000b900000000000000bc000000000000009d000000000000009600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE6;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE7 : if BRAM_NAME = "sampleifmap_layersamples_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ce0000000000000086000000000000001a000000000000000d00000000",
            INIT_01 => X"000000ac000000000000008d0000000000000076000000000000008a00000000",
            INIT_02 => X"000000e400000000000000dc00000000000000cf00000000000000b500000000",
            INIT_03 => X"000000b000000000000000e200000000000000e600000000000000e000000000",
            INIT_04 => X"00000091000000000000008e000000000000008a000000000000009000000000",
            INIT_05 => X"0000009a00000000000000950000000000000095000000000000009a00000000",
            INIT_06 => X"000000bb00000000000000ad00000000000000a0000000000000009d00000000",
            INIT_07 => X"0000009d00000000000000a500000000000000b200000000000000be00000000",
            INIT_08 => X"000000e100000000000000c8000000000000003a000000000000000500000000",
            INIT_09 => X"000000e200000000000000d400000000000000c700000000000000c500000000",
            INIT_0A => X"000000e600000000000000e800000000000000e900000000000000e500000000",
            INIT_0B => X"000000d200000000000000dd00000000000000df00000000000000d100000000",
            INIT_0C => X"000000bc00000000000000c100000000000000b400000000000000c600000000",
            INIT_0D => X"000000b800000000000000c000000000000000c200000000000000bd00000000",
            INIT_0E => X"0000009000000000000000a100000000000000ab00000000000000ac00000000",
            INIT_0F => X"0000008a00000000000000800000000000000083000000000000008800000000",
            INIT_10 => X"000000ba00000000000000be0000000000000091000000000000002700000000",
            INIT_11 => X"000000c200000000000000c200000000000000c000000000000000b800000000",
            INIT_12 => X"000000be00000000000000c000000000000000bf00000000000000c200000000",
            INIT_13 => X"00000093000000000000009a00000000000000b400000000000000b100000000",
            INIT_14 => X"000000710000000000000092000000000000009c000000000000009100000000",
            INIT_15 => X"0000006f000000000000007e0000000000000084000000000000007200000000",
            INIT_16 => X"0000005e000000000000005d000000000000005b000000000000005c00000000",
            INIT_17 => X"0000008100000000000000810000000000000079000000000000006900000000",
            INIT_18 => X"00000089000000000000008f00000000000000a2000000000000007a00000000",
            INIT_19 => X"00000082000000000000007f0000000000000080000000000000008300000000",
            INIT_1A => X"00000081000000000000007f0000000000000080000000000000008300000000",
            INIT_1B => X"000000640000000000000068000000000000007c000000000000008100000000",
            INIT_1C => X"0000005e00000000000000700000000000000076000000000000006600000000",
            INIT_1D => X"000000530000000000000057000000000000005e000000000000005e00000000",
            INIT_1E => X"00000065000000000000005d0000000000000053000000000000005000000000",
            INIT_1F => X"0000008200000000000000790000000000000073000000000000006c00000000",
            INIT_20 => X"00000050000000000000004d000000000000004c000000000000004900000000",
            INIT_21 => X"0000005a00000000000000570000000000000057000000000000005400000000",
            INIT_22 => X"00000071000000000000006b0000000000000066000000000000005e00000000",
            INIT_23 => X"0000007800000000000000760000000000000076000000000000007300000000",
            INIT_24 => X"00000064000000000000006a000000000000006e000000000000007300000000",
            INIT_25 => X"00000050000000000000004f0000000000000055000000000000005f00000000",
            INIT_26 => X"000000520000000000000050000000000000004d000000000000005000000000",
            INIT_27 => X"00000088000000000000007d0000000000000071000000000000005c00000000",
            INIT_28 => X"0000001200000000000000090000000000000003000000000000000d00000000",
            INIT_29 => X"0000001600000000000000140000000000000015000000000000001200000000",
            INIT_2A => X"00000030000000000000002a0000000000000022000000000000001a00000000",
            INIT_2B => X"000000460000000000000042000000000000003c000000000000003400000000",
            INIT_2C => X"0000003c00000000000000430000000000000048000000000000004700000000",
            INIT_2D => X"0000003900000000000000350000000000000035000000000000003700000000",
            INIT_2E => X"0000005700000000000000480000000000000039000000000000003900000000",
            INIT_2F => X"0000008900000000000000820000000000000078000000000000006800000000",
            INIT_30 => X"000000200000000000000008000000000000000b000000000000002400000000",
            INIT_31 => X"0000000300000000000000080000000000000016000000000000002400000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_33 => X"0000000300000000000000010000000000000005000000000000000600000000",
            INIT_34 => X"0000001500000000000000150000000000000018000000000000000d00000000",
            INIT_35 => X"00000027000000000000001e0000000000000016000000000000001500000000",
            INIT_36 => X"0000007b00000000000000710000000000000055000000000000003900000000",
            INIT_37 => X"000000990000000000000086000000000000007a000000000000007400000000",
            INIT_38 => X"0000001b000000000000000d000000000000001a000000000000002300000000",
            INIT_39 => X"0000001b00000000000000310000000000000046000000000000004700000000",
            INIT_3A => X"0000000000000000000000020000000000000005000000000000000f00000000",
            INIT_3B => X"0000000a000000000000001f0000000000000039000000000000001100000000",
            INIT_3C => X"0000000e00000000000000070000000000000004000000000000000400000000",
            INIT_3D => X"00000056000000000000003e0000000000000029000000000000001900000000",
            INIT_3E => X"0000007200000000000000840000000000000090000000000000007a00000000",
            INIT_3F => X"000000ac00000000000000920000000000000084000000000000007500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000030000000000000004000000000000000d000000000000001000000000",
            INIT_41 => X"0000002400000000000000360000000000000041000000000000002d00000000",
            INIT_42 => X"0000000000000000000000020000000000000004000000000000001200000000",
            INIT_43 => X"0000008300000000000000a10000000000000076000000000000000700000000",
            INIT_44 => X"0000006d00000000000000690000000000000069000000000000007000000000",
            INIT_45 => X"00000097000000000000009a000000000000008a000000000000007600000000",
            INIT_46 => X"00000078000000000000006a0000000000000069000000000000007f00000000",
            INIT_47 => X"000000b800000000000000a4000000000000008e000000000000008100000000",
            INIT_48 => X"000000000000000000000000000000000000000c000000000000002800000000",
            INIT_49 => X"000000150000000000000020000000000000001e000000000000000c00000000",
            INIT_4A => X"0000000300000000000000020000000000000002000000000000000700000000",
            INIT_4B => X"000000cd00000000000000b60000000000000044000000000000000000000000",
            INIT_4C => X"000000bb00000000000000c300000000000000c200000000000000c400000000",
            INIT_4D => X"00000067000000000000007b000000000000009600000000000000ac00000000",
            INIT_4E => X"00000081000000000000007a0000000000000068000000000000005f00000000",
            INIT_4F => X"000000b900000000000000ab0000000000000098000000000000008400000000",
            INIT_50 => X"000000010000000000000001000000000000001a000000000000004500000000",
            INIT_51 => X"0000000c0000000000000012000000000000000c000000000000000400000000",
            INIT_52 => X"0000000400000000000000020000000000000002000000000000000400000000",
            INIT_53 => X"000000cb00000000000000990000000000000020000000000000000100000000",
            INIT_54 => X"0000009b00000000000000b300000000000000bf00000000000000c300000000",
            INIT_55 => X"0000005e0000000000000051000000000000005b000000000000007700000000",
            INIT_56 => X"00000081000000000000007d000000000000007d000000000000007500000000",
            INIT_57 => X"000000b800000000000000ad00000000000000a2000000000000009000000000",
            INIT_58 => X"000000020000000000000001000000000000002f000000000000005300000000",
            INIT_59 => X"0000000400000000000000070000000000000005000000000000000200000000",
            INIT_5A => X"0000000300000000000000010000000000000001000000000000000100000000",
            INIT_5B => X"000000cd000000000000008e000000000000001b000000000000000100000000",
            INIT_5C => X"00000055000000000000007900000000000000a900000000000000c600000000",
            INIT_5D => X"0000007900000000000000660000000000000055000000000000004a00000000",
            INIT_5E => X"000000840000000000000079000000000000007a000000000000008000000000",
            INIT_5F => X"000000ba00000000000000b000000000000000a5000000000000009300000000",
            INIT_60 => X"0000000300000000000000060000000000000036000000000000005c00000000",
            INIT_61 => X"0000000100000000000000010000000000000001000000000000000200000000",
            INIT_62 => X"0000000100000000000000010000000000000001000000000000000100000000",
            INIT_63 => X"0000009d0000000000000066000000000000000f000000000000000000000000",
            INIT_64 => X"0000004a0000000000000038000000000000004a000000000000007500000000",
            INIT_65 => X"0000007c000000000000007a0000000000000073000000000000006300000000",
            INIT_66 => X"000000880000000000000080000000000000007d000000000000007b00000000",
            INIT_67 => X"000000bc00000000000000b100000000000000a2000000000000009400000000",
            INIT_68 => X"0000000b0000000000000013000000000000002b000000000000005700000000",
            INIT_69 => X"0000000200000000000000020000000000000005000000000000000800000000",
            INIT_6A => X"0000000200000000000000030000000000000003000000000000000300000000",
            INIT_6B => X"00000047000000000000002a0000000000000004000000000000000000000000",
            INIT_6C => X"0000007100000000000000500000000000000039000000000000003500000000",
            INIT_6D => X"00000074000000000000007b0000000000000086000000000000008400000000",
            INIT_6E => X"0000008f000000000000008b0000000000000083000000000000007800000000",
            INIT_6F => X"000000bc00000000000000b600000000000000a9000000000000009c00000000",
            INIT_70 => X"0000001f0000000000000024000000000000002e000000000000005200000000",
            INIT_71 => X"0000001000000000000000110000000000000016000000000000001b00000000",
            INIT_72 => X"0000001300000000000000140000000000000013000000000000001200000000",
            INIT_73 => X"0000004000000000000000250000000000000017000000000000001300000000",
            INIT_74 => X"0000008000000000000000740000000000000068000000000000005700000000",
            INIT_75 => X"0000007300000000000000750000000000000083000000000000008b00000000",
            INIT_76 => X"00000094000000000000008b0000000000000083000000000000007b00000000",
            INIT_77 => X"000000bb00000000000000b900000000000000ae000000000000009f00000000",
            INIT_78 => X"00000037000000000000003a000000000000003e000000000000005500000000",
            INIT_79 => X"00000030000000000000002e000000000000002f000000000000003300000000",
            INIT_7A => X"0000003700000000000000350000000000000033000000000000003100000000",
            INIT_7B => X"0000006800000000000000510000000000000044000000000000003b00000000",
            INIT_7C => X"0000007f0000000000000085000000000000007f000000000000007400000000",
            INIT_7D => X"0000007a00000000000000720000000000000076000000000000007f00000000",
            INIT_7E => X"00000095000000000000008d0000000000000088000000000000008100000000",
            INIT_7F => X"000000ba00000000000000b400000000000000a8000000000000009e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE7;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE8 : if BRAM_NAME = "sampleifmap_layersamples_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e800000000000000e800000000000000e700000000000000eb00000000",
            INIT_01 => X"000000e800000000000000e800000000000000e800000000000000e800000000",
            INIT_02 => X"000000e900000000000000e900000000000000e800000000000000e800000000",
            INIT_03 => X"000000e800000000000000e900000000000000e900000000000000e900000000",
            INIT_04 => X"000000e900000000000000e900000000000000e700000000000000e700000000",
            INIT_05 => X"000000e900000000000000e800000000000000e700000000000000e800000000",
            INIT_06 => X"000000e800000000000000e800000000000000e900000000000000e900000000",
            INIT_07 => X"000000e800000000000000e900000000000000e900000000000000e800000000",
            INIT_08 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_09 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_0A => X"000000ec00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_0B => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_0C => X"000000ec00000000000000ec00000000000000ea00000000000000ea00000000",
            INIT_0D => X"000000ec00000000000000ec00000000000000ea00000000000000eb00000000",
            INIT_0E => X"000000eb00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_0F => X"000000eb00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_10 => X"000000ea00000000000000ea00000000000000ea00000000000000ed00000000",
            INIT_11 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_12 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_13 => X"000000ea00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_14 => X"000000eb00000000000000eb00000000000000ea00000000000000e900000000",
            INIT_15 => X"000000ea00000000000000e900000000000000eb00000000000000e600000000",
            INIT_16 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_17 => X"000000ea00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_18 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_19 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_1A => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_1B => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_1C => X"000000e200000000000000e600000000000000e800000000000000e900000000",
            INIT_1D => X"000000e400000000000000d200000000000000d800000000000000c000000000",
            INIT_1E => X"000000ea00000000000000ea00000000000000ea00000000000000eb00000000",
            INIT_1F => X"000000eb00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_20 => X"000000eb00000000000000eb00000000000000ea00000000000000ed00000000",
            INIT_21 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_22 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_23 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_24 => X"000000d200000000000000e100000000000000ed00000000000000ee00000000",
            INIT_25 => X"000000e500000000000000da00000000000000cd00000000000000ac00000000",
            INIT_26 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_27 => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_28 => X"000000eb00000000000000eb00000000000000eb00000000000000ef00000000",
            INIT_29 => X"000000eb00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_2A => X"000000ec00000000000000ec00000000000000eb00000000000000ea00000000",
            INIT_2B => X"000000e700000000000000ed00000000000000e900000000000000eb00000000",
            INIT_2C => X"000000bc00000000000000c600000000000000cd00000000000000d800000000",
            INIT_2D => X"000000e400000000000000d700000000000000c400000000000000b300000000",
            INIT_2E => X"000000ec00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_2F => X"000000ed00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_30 => X"000000e400000000000000e600000000000000e300000000000000e500000000",
            INIT_31 => X"000000ed00000000000000ed00000000000000ec00000000000000e800000000",
            INIT_32 => X"000000ed00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_33 => X"000000e200000000000000ed00000000000000e400000000000000e500000000",
            INIT_34 => X"000000b000000000000000b400000000000000b400000000000000c500000000",
            INIT_35 => X"000000ce00000000000000a9000000000000009f00000000000000a300000000",
            INIT_36 => X"000000eb00000000000000ec00000000000000ed00000000000000ee00000000",
            INIT_37 => X"000000ed00000000000000ed00000000000000ee00000000000000ec00000000",
            INIT_38 => X"000000e800000000000000ea00000000000000e600000000000000dc00000000",
            INIT_39 => X"000000ed00000000000000ee00000000000000ed00000000000000ea00000000",
            INIT_3A => X"000000ee00000000000000ec00000000000000ed00000000000000ed00000000",
            INIT_3B => X"000000da00000000000000ec00000000000000de00000000000000cc00000000",
            INIT_3C => X"000000bf00000000000000c900000000000000c900000000000000cc00000000",
            INIT_3D => X"000000c700000000000000b000000000000000ae00000000000000b600000000",
            INIT_3E => X"000000ee00000000000000ee00000000000000ef00000000000000ef00000000",
            INIT_3F => X"000000ee00000000000000ef00000000000000ef00000000000000ef00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ef00000000000000ee00000000000000ec00000000000000ea00000000",
            INIT_41 => X"000000ec00000000000000ed00000000000000ee00000000000000f000000000",
            INIT_42 => X"000000ef00000000000000ed00000000000000ec00000000000000ec00000000",
            INIT_43 => X"000000e700000000000000ea00000000000000dd00000000000000c600000000",
            INIT_44 => X"000000da00000000000000e400000000000000d800000000000000d500000000",
            INIT_45 => X"000000eb00000000000000e900000000000000e000000000000000dd00000000",
            INIT_46 => X"000000f000000000000000ef00000000000000ee00000000000000f000000000",
            INIT_47 => X"000000ee00000000000000f000000000000000f000000000000000f000000000",
            INIT_48 => X"0000009b000000000000008e000000000000008a000000000000008c00000000",
            INIT_49 => X"000000ea00000000000000ec00000000000000ea00000000000000bc00000000",
            INIT_4A => X"000000ed00000000000000ed00000000000000eb00000000000000e900000000",
            INIT_4B => X"000000ed00000000000000ea00000000000000e400000000000000d800000000",
            INIT_4C => X"000000e800000000000000ec00000000000000e600000000000000e600000000",
            INIT_4D => X"000000cc00000000000000db00000000000000e900000000000000ed00000000",
            INIT_4E => X"000000c700000000000000b400000000000000b300000000000000bd00000000",
            INIT_4F => X"000000f000000000000000f000000000000000f100000000000000eb00000000",
            INIT_50 => X"0000007f000000000000007d0000000000000079000000000000008200000000",
            INIT_51 => X"000000e200000000000000e400000000000000e5000000000000009f00000000",
            INIT_52 => X"000000ed00000000000000ec00000000000000ea00000000000000e800000000",
            INIT_53 => X"000000eb00000000000000ed00000000000000eb00000000000000ea00000000",
            INIT_54 => X"000000e800000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_55 => X"0000009c00000000000000a500000000000000b800000000000000ce00000000",
            INIT_56 => X"000000a20000000000000085000000000000008c000000000000009500000000",
            INIT_57 => X"000000f000000000000000f000000000000000f100000000000000e400000000",
            INIT_58 => X"000000d300000000000000d300000000000000ca00000000000000d400000000",
            INIT_59 => X"000000d100000000000000d500000000000000e300000000000000d900000000",
            INIT_5A => X"000000dd00000000000000e200000000000000de00000000000000d500000000",
            INIT_5B => X"000000e500000000000000e100000000000000dd00000000000000db00000000",
            INIT_5C => X"000000e700000000000000ed00000000000000ec00000000000000ea00000000",
            INIT_5D => X"000000c200000000000000c800000000000000c600000000000000cc00000000",
            INIT_5E => X"000000c3000000000000009700000000000000b200000000000000c500000000",
            INIT_5F => X"000000f000000000000000f100000000000000f000000000000000e600000000",
            INIT_60 => X"000000d900000000000000d300000000000000ca00000000000000cf00000000",
            INIT_61 => X"000000ae00000000000000d000000000000000db00000000000000e100000000",
            INIT_62 => X"0000007000000000000000b800000000000000d500000000000000b400000000",
            INIT_63 => X"0000008a00000000000000810000000000000079000000000000007200000000",
            INIT_64 => X"000000ec00000000000000d800000000000000a7000000000000009800000000",
            INIT_65 => X"000000e200000000000000ea00000000000000e900000000000000e800000000",
            INIT_66 => X"000000e600000000000000cb00000000000000db00000000000000e400000000",
            INIT_67 => X"000000f100000000000000ef00000000000000e600000000000000e300000000",
            INIT_68 => X"00000083000000000000007d000000000000007d000000000000008200000000",
            INIT_69 => X"000000c700000000000000c900000000000000b6000000000000009100000000",
            INIT_6A => X"0000004700000000000000ac00000000000000e600000000000000db00000000",
            INIT_6B => X"0000005400000000000000490000000000000049000000000000004600000000",
            INIT_6C => X"000000ef00000000000000e300000000000000a8000000000000007200000000",
            INIT_6D => X"000000d300000000000000e400000000000000e700000000000000ed00000000",
            INIT_6E => X"000000ce00000000000000db00000000000000da00000000000000d000000000",
            INIT_6F => X"000000e700000000000000dd00000000000000c500000000000000ba00000000",
            INIT_70 => X"00000055000000000000004f0000000000000056000000000000005100000000",
            INIT_71 => X"000000c8000000000000009d000000000000009b000000000000008d00000000",
            INIT_72 => X"0000007900000000000000b400000000000000df00000000000000e400000000",
            INIT_73 => X"000000c000000000000000970000000000000075000000000000007000000000",
            INIT_74 => X"000000cb00000000000000db00000000000000de00000000000000d400000000",
            INIT_75 => X"0000008a000000000000009a00000000000000a600000000000000ba00000000",
            INIT_76 => X"0000008e0000000000000092000000000000008b000000000000008500000000",
            INIT_77 => X"000000d400000000000000c50000000000000099000000000000008900000000",
            INIT_78 => X"0000009000000000000000620000000000000046000000000000003500000000",
            INIT_79 => X"0000009e0000000000000073000000000000006b000000000000009700000000",
            INIT_7A => X"000000c100000000000000c200000000000000c200000000000000b400000000",
            INIT_7B => X"000000d200000000000000e400000000000000d100000000000000c200000000",
            INIT_7C => X"00000088000000000000009600000000000000a500000000000000b500000000",
            INIT_7D => X"0000006f000000000000006a000000000000006f000000000000007d00000000",
            INIT_7E => X"0000009700000000000000870000000000000079000000000000007600000000",
            INIT_7F => X"000000cb00000000000000ce00000000000000ae00000000000000a400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE8;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE9 : if BRAM_NAME = "sampleifmap_layersamples_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d8000000000000008c000000000000001d000000000000000f00000000",
            INIT_01 => X"000000a20000000000000085000000000000007b000000000000009600000000",
            INIT_02 => X"000000ea00000000000000e000000000000000d100000000000000b500000000",
            INIT_03 => X"000000bd00000000000000ee00000000000000f100000000000000ea00000000",
            INIT_04 => X"000000a3000000000000009e000000000000009a000000000000009f00000000",
            INIT_05 => X"000000ab00000000000000a500000000000000a500000000000000ab00000000",
            INIT_06 => X"000000cc00000000000000be00000000000000b100000000000000ae00000000",
            INIT_07 => X"000000af00000000000000b700000000000000c400000000000000cf00000000",
            INIT_08 => X"000000e800000000000000cf000000000000003e000000000000000500000000",
            INIT_09 => X"000000e000000000000000d400000000000000cf00000000000000cd00000000",
            INIT_0A => X"000000ee00000000000000ee00000000000000ec00000000000000e600000000",
            INIT_0B => X"000000e400000000000000ee00000000000000ee00000000000000dd00000000",
            INIT_0C => X"000000d500000000000000d800000000000000c800000000000000d900000000",
            INIT_0D => X"000000cc00000000000000d400000000000000d600000000000000d400000000",
            INIT_0E => X"000000a500000000000000b500000000000000bf00000000000000c100000000",
            INIT_0F => X"0000009a000000000000008f0000000000000092000000000000009c00000000",
            INIT_10 => X"000000c400000000000000cc000000000000009b000000000000002d00000000",
            INIT_11 => X"000000d000000000000000d300000000000000d300000000000000c500000000",
            INIT_12 => X"000000cf00000000000000cf00000000000000cb00000000000000ce00000000",
            INIT_13 => X"000000a900000000000000b000000000000000c600000000000000c100000000",
            INIT_14 => X"0000008500000000000000a300000000000000ab00000000000000a100000000",
            INIT_15 => X"000000870000000000000096000000000000009d000000000000008900000000",
            INIT_16 => X"0000007400000000000000720000000000000070000000000000007300000000",
            INIT_17 => X"0000008e000000000000008d0000000000000085000000000000007d00000000",
            INIT_18 => X"0000009a00000000000000a000000000000000b3000000000000008700000000",
            INIT_19 => X"0000009600000000000000960000000000000098000000000000009800000000",
            INIT_1A => X"0000009500000000000000930000000000000093000000000000009600000000",
            INIT_1B => X"0000007a000000000000007e0000000000000091000000000000009500000000",
            INIT_1C => X"0000006d00000000000000800000000000000086000000000000007800000000",
            INIT_1D => X"0000006700000000000000700000000000000075000000000000007000000000",
            INIT_1E => X"00000075000000000000006f0000000000000067000000000000006100000000",
            INIT_1F => X"000000900000000000000085000000000000007d000000000000007900000000",
            INIT_20 => X"0000005d000000000000005a000000000000005a000000000000005700000000",
            INIT_21 => X"0000006900000000000000660000000000000066000000000000006200000000",
            INIT_22 => X"00000083000000000000007c0000000000000077000000000000006f00000000",
            INIT_23 => X"0000008500000000000000840000000000000088000000000000008900000000",
            INIT_24 => X"00000077000000000000007f0000000000000085000000000000008800000000",
            INIT_25 => X"0000005c00000000000000610000000000000065000000000000006d00000000",
            INIT_26 => X"0000006200000000000000640000000000000064000000000000005e00000000",
            INIT_27 => X"0000009500000000000000870000000000000077000000000000006800000000",
            INIT_28 => X"0000001a0000000000000010000000000000000b000000000000001900000000",
            INIT_29 => X"0000001e00000000000000190000000000000019000000000000001a00000000",
            INIT_2A => X"0000003b0000000000000033000000000000002b000000000000002400000000",
            INIT_2B => X"0000004f000000000000004d000000000000004b000000000000004500000000",
            INIT_2C => X"0000004800000000000000510000000000000058000000000000005700000000",
            INIT_2D => X"0000004500000000000000450000000000000044000000000000004300000000",
            INIT_2E => X"000000640000000000000059000000000000004e000000000000004700000000",
            INIT_2F => X"000000920000000000000088000000000000007c000000000000007100000000",
            INIT_30 => X"0000002c000000000000000d0000000000000010000000000000002e00000000",
            INIT_31 => X"00000008000000000000000b0000000000000019000000000000002d00000000",
            INIT_32 => X"0000000400000000000000020000000000000002000000000000000400000000",
            INIT_33 => X"0000001700000000000000130000000000000012000000000000000d00000000",
            INIT_34 => X"0000001f00000000000000210000000000000026000000000000001d00000000",
            INIT_35 => X"0000003a0000000000000032000000000000002c000000000000002600000000",
            INIT_36 => X"0000007b0000000000000073000000000000005a000000000000004600000000",
            INIT_37 => X"000000a0000000000000008b000000000000007b000000000000007300000000",
            INIT_38 => X"000000290000000000000013000000000000001b000000000000002900000000",
            INIT_39 => X"0000001f00000000000000320000000000000046000000000000005100000000",
            INIT_3A => X"0000000000000000000000020000000000000005000000000000000f00000000",
            INIT_3B => X"0000002400000000000000320000000000000040000000000000001100000000",
            INIT_3C => X"00000023000000000000001e000000000000001e000000000000001e00000000",
            INIT_3D => X"0000006100000000000000470000000000000037000000000000002b00000000",
            INIT_3E => X"0000006900000000000000780000000000000083000000000000007c00000000",
            INIT_3F => X"000000b300000000000000980000000000000086000000000000006f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000c000000000000000a000000000000000a000000000000000f00000000",
            INIT_41 => X"00000021000000000000002b0000000000000034000000000000002c00000000",
            INIT_42 => X"0000000100000000000000020000000000000004000000000000001200000000",
            INIT_43 => X"00000080000000000000009e0000000000000075000000000000000800000000",
            INIT_44 => X"0000006900000000000000670000000000000069000000000000007000000000",
            INIT_45 => X"0000007e000000000000007e0000000000000073000000000000006b00000000",
            INIT_46 => X"00000074000000000000005e0000000000000056000000000000006a00000000",
            INIT_47 => X"000000c200000000000000ac0000000000000093000000000000008200000000",
            INIT_48 => X"000000040000000000000003000000000000000a000000000000002800000000",
            INIT_49 => X"0000000a000000000000000c000000000000000c000000000000000600000000",
            INIT_4A => X"0000000200000000000000010000000000000001000000000000000600000000",
            INIT_4B => X"000000820000000000000080000000000000003a000000000000000000000000",
            INIT_4C => X"000000710000000000000077000000000000007b000000000000007f00000000",
            INIT_4D => X"00000042000000000000004b0000000000000060000000000000006e00000000",
            INIT_4E => X"000000840000000000000076000000000000005d000000000000004700000000",
            INIT_4F => X"000000c500000000000000b600000000000000a2000000000000008d00000000",
            INIT_50 => X"000000010000000000000001000000000000001d000000000000004d00000000",
            INIT_51 => X"0000000200000000000000030000000000000002000000000000000100000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_53 => X"0000002f000000000000002d000000000000000c000000000000000100000000",
            INIT_54 => X"0000003100000000000000320000000000000030000000000000002e00000000",
            INIT_55 => X"0000004d00000000000000300000000000000026000000000000002a00000000",
            INIT_56 => X"000000870000000000000080000000000000007e000000000000006e00000000",
            INIT_57 => X"000000c600000000000000bb00000000000000b0000000000000009900000000",
            INIT_58 => X"0000000100000000000000010000000000000034000000000000005e00000000",
            INIT_59 => X"0000000000000000000000010000000000000001000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000002000000000000000190000000000000003000000000000000200000000",
            INIT_5C => X"0000001d00000000000000190000000000000019000000000000001900000000",
            INIT_5D => X"00000071000000000000005c0000000000000042000000000000002900000000",
            INIT_5E => X"0000008b000000000000007f000000000000007e000000000000007c00000000",
            INIT_5F => X"000000c900000000000000bf00000000000000b3000000000000009d00000000",
            INIT_60 => X"000000020000000000000007000000000000003c000000000000006600000000",
            INIT_61 => X"0000000200000000000000030000000000000003000000000000000200000000",
            INIT_62 => X"0000000100000000000000000000000000000000000000000000000100000000",
            INIT_63 => X"0000001f00000000000000130000000000000001000000000000000300000000",
            INIT_64 => X"0000003a000000000000001b000000000000000d000000000000001100000000",
            INIT_65 => X"0000007c000000000000007e0000000000000073000000000000005a00000000",
            INIT_66 => X"0000009100000000000000870000000000000082000000000000007b00000000",
            INIT_67 => X"000000ca00000000000000c000000000000000b0000000000000009f00000000",
            INIT_68 => X"0000000c00000000000000170000000000000033000000000000006300000000",
            INIT_69 => X"00000007000000000000000a000000000000000b000000000000000a00000000",
            INIT_6A => X"0000000300000000000000040000000000000004000000000000000400000000",
            INIT_6B => X"00000015000000000000000d0000000000000005000000000000000600000000",
            INIT_6C => X"00000062000000000000004d0000000000000032000000000000001b00000000",
            INIT_6D => X"0000007d000000000000007e000000000000007e000000000000007100000000",
            INIT_6E => X"0000009a0000000000000094000000000000008a000000000000008000000000",
            INIT_6F => X"000000ca00000000000000c500000000000000b800000000000000a800000000",
            INIT_70 => X"00000023000000000000002c0000000000000039000000000000006000000000",
            INIT_71 => X"00000017000000000000001a000000000000001c000000000000001e00000000",
            INIT_72 => X"0000001700000000000000160000000000000015000000000000001500000000",
            INIT_73 => X"000000370000000000000028000000000000001f000000000000001b00000000",
            INIT_74 => X"0000007000000000000000660000000000000058000000000000004600000000",
            INIT_75 => X"0000007f000000000000007a000000000000007a000000000000007900000000",
            INIT_76 => X"000000a00000000000000095000000000000008b000000000000008500000000",
            INIT_77 => X"000000ca00000000000000c800000000000000bd00000000000000ac00000000",
            INIT_78 => X"0000003d0000000000000043000000000000004b000000000000006500000000",
            INIT_79 => X"0000003700000000000000350000000000000035000000000000003800000000",
            INIT_7A => X"0000003e000000000000003a0000000000000038000000000000003700000000",
            INIT_7B => X"0000006000000000000000540000000000000047000000000000004300000000",
            INIT_7C => X"000000790000000000000074000000000000006d000000000000006700000000",
            INIT_7D => X"00000083000000000000007d000000000000007c000000000000007f00000000",
            INIT_7E => X"000000a200000000000000980000000000000091000000000000008800000000",
            INIT_7F => X"000000c800000000000000c300000000000000b700000000000000ab00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE9;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE10 : if BRAM_NAME = "sampleifmap_layersamples_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e800000000000000e800000000000000e700000000000000eb00000000",
            INIT_01 => X"000000e800000000000000e800000000000000e800000000000000e800000000",
            INIT_02 => X"000000e900000000000000e900000000000000e800000000000000e800000000",
            INIT_03 => X"000000e900000000000000e900000000000000e900000000000000e900000000",
            INIT_04 => X"000000e800000000000000e900000000000000e900000000000000e900000000",
            INIT_05 => X"000000e600000000000000e800000000000000ea00000000000000ea00000000",
            INIT_06 => X"000000e800000000000000e800000000000000e900000000000000e700000000",
            INIT_07 => X"000000e800000000000000e900000000000000e900000000000000e800000000",
            INIT_08 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_09 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_0A => X"000000ec00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_0B => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_0C => X"000000ea00000000000000ea00000000000000e900000000000000e900000000",
            INIT_0D => X"000000eb00000000000000ed00000000000000ee00000000000000ed00000000",
            INIT_0E => X"000000eb00000000000000eb00000000000000ec00000000000000ea00000000",
            INIT_0F => X"000000eb00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_10 => X"000000ea00000000000000ea00000000000000ea00000000000000ed00000000",
            INIT_11 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_12 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_13 => X"000000ea00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_14 => X"000000ec00000000000000ea00000000000000e700000000000000e700000000",
            INIT_15 => X"000000ea00000000000000eb00000000000000ee00000000000000e900000000",
            INIT_16 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_17 => X"000000ea00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_18 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_19 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_1A => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_1B => X"000000ea00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_1C => X"000000e700000000000000e800000000000000e700000000000000e600000000",
            INIT_1D => X"000000e600000000000000d500000000000000db00000000000000c500000000",
            INIT_1E => X"000000ea00000000000000ea00000000000000ea00000000000000eb00000000",
            INIT_1F => X"000000eb00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_20 => X"000000eb00000000000000eb00000000000000ea00000000000000ed00000000",
            INIT_21 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_22 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_23 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_24 => X"000000db00000000000000e600000000000000ed00000000000000ec00000000",
            INIT_25 => X"000000e800000000000000dd00000000000000d000000000000000b300000000",
            INIT_26 => X"000000eb00000000000000eb00000000000000eb00000000000000ed00000000",
            INIT_27 => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_28 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_29 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_2A => X"000000ec00000000000000ec00000000000000eb00000000000000ea00000000",
            INIT_2B => X"000000e800000000000000ed00000000000000ea00000000000000ec00000000",
            INIT_2C => X"000000c800000000000000cf00000000000000d200000000000000da00000000",
            INIT_2D => X"000000e800000000000000dc00000000000000ca00000000000000bd00000000",
            INIT_2E => X"000000eb00000000000000eb00000000000000eb00000000000000ed00000000",
            INIT_2F => X"000000ed00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_30 => X"000000e600000000000000e700000000000000e400000000000000e500000000",
            INIT_31 => X"000000eb00000000000000eb00000000000000ec00000000000000e900000000",
            INIT_32 => X"000000ee00000000000000ed00000000000000ec00000000000000ec00000000",
            INIT_33 => X"000000e400000000000000ee00000000000000e500000000000000e600000000",
            INIT_34 => X"000000be00000000000000bf00000000000000be00000000000000cc00000000",
            INIT_35 => X"000000d300000000000000b100000000000000ab00000000000000b100000000",
            INIT_36 => X"000000eb00000000000000e900000000000000ea00000000000000ef00000000",
            INIT_37 => X"000000ee00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_38 => X"000000ea00000000000000ee00000000000000e900000000000000de00000000",
            INIT_39 => X"000000ec00000000000000eb00000000000000ec00000000000000ea00000000",
            INIT_3A => X"000000ef00000000000000ed00000000000000ee00000000000000ee00000000",
            INIT_3B => X"000000da00000000000000eb00000000000000dd00000000000000cb00000000",
            INIT_3C => X"000000cb00000000000000d300000000000000d200000000000000d200000000",
            INIT_3D => X"000000cc00000000000000b900000000000000bb00000000000000c400000000",
            INIT_3E => X"000000ee00000000000000ed00000000000000ee00000000000000f000000000",
            INIT_3F => X"000000ee00000000000000ee00000000000000ee00000000000000ee00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f300000000000000f600000000000000f300000000000000f100000000",
            INIT_41 => X"000000eb00000000000000eb00000000000000ed00000000000000f000000000",
            INIT_42 => X"000000ef00000000000000ed00000000000000ed00000000000000ed00000000",
            INIT_43 => X"000000e500000000000000e700000000000000da00000000000000c400000000",
            INIT_44 => X"000000e300000000000000eb00000000000000de00000000000000d900000000",
            INIT_45 => X"000000f100000000000000f000000000000000eb00000000000000ea00000000",
            INIT_46 => X"000000f000000000000000f000000000000000f000000000000000f300000000",
            INIT_47 => X"000000ee00000000000000ef00000000000000ef00000000000000ef00000000",
            INIT_48 => X"000000a100000000000000990000000000000094000000000000009500000000",
            INIT_49 => X"000000e800000000000000e900000000000000e900000000000000bf00000000",
            INIT_4A => X"000000eb00000000000000ec00000000000000eb00000000000000ea00000000",
            INIT_4B => X"000000ec00000000000000e800000000000000e200000000000000d600000000",
            INIT_4C => X"000000ef00000000000000f100000000000000eb00000000000000e800000000",
            INIT_4D => X"000000d300000000000000e200000000000000f300000000000000f700000000",
            INIT_4E => X"000000c900000000000000b900000000000000ba00000000000000c300000000",
            INIT_4F => X"000000ef00000000000000ef00000000000000ef00000000000000eb00000000",
            INIT_50 => X"0000008900000000000000890000000000000085000000000000008d00000000",
            INIT_51 => X"000000e000000000000000e100000000000000e700000000000000a500000000",
            INIT_52 => X"000000eb00000000000000ea00000000000000ea00000000000000e900000000",
            INIT_53 => X"000000ec00000000000000ee00000000000000ec00000000000000eb00000000",
            INIT_54 => X"000000ee00000000000000f100000000000000f000000000000000ee00000000",
            INIT_55 => X"000000a300000000000000ac00000000000000bf00000000000000d500000000",
            INIT_56 => X"000000a6000000000000008f0000000000000099000000000000009f00000000",
            INIT_57 => X"000000ef00000000000000ee00000000000000ef00000000000000e500000000",
            INIT_58 => X"000000df00000000000000e000000000000000d700000000000000e000000000",
            INIT_59 => X"000000ce00000000000000d300000000000000e700000000000000e300000000",
            INIT_5A => X"000000db00000000000000e100000000000000de00000000000000d600000000",
            INIT_5B => X"000000e900000000000000e600000000000000e100000000000000df00000000",
            INIT_5C => X"000000ed00000000000000f100000000000000ef00000000000000ed00000000",
            INIT_5D => X"000000ca00000000000000cf00000000000000cb00000000000000d000000000",
            INIT_5E => X"000000ca00000000000000a400000000000000c400000000000000d300000000",
            INIT_5F => X"000000ef00000000000000ef00000000000000ee00000000000000e900000000",
            INIT_60 => X"000000ea00000000000000e000000000000000d900000000000000de00000000",
            INIT_61 => X"000000ae00000000000000d000000000000000e300000000000000f100000000",
            INIT_62 => X"0000007900000000000000bc00000000000000d600000000000000b700000000",
            INIT_63 => X"00000093000000000000008b0000000000000084000000000000007e00000000",
            INIT_64 => X"000000ed00000000000000dc00000000000000ae00000000000000a100000000",
            INIT_65 => X"000000e900000000000000f000000000000000ee00000000000000eb00000000",
            INIT_66 => X"000000ed00000000000000d400000000000000e500000000000000ed00000000",
            INIT_67 => X"000000f200000000000000f200000000000000e900000000000000ea00000000",
            INIT_68 => X"00000097000000000000008d0000000000000093000000000000009800000000",
            INIT_69 => X"000000cc00000000000000cd00000000000000c100000000000000a500000000",
            INIT_6A => X"0000005c00000000000000b700000000000000ea00000000000000e200000000",
            INIT_6B => X"00000062000000000000005a000000000000005b000000000000005b00000000",
            INIT_6C => X"000000f100000000000000e900000000000000b3000000000000008100000000",
            INIT_6D => X"000000d900000000000000e900000000000000ed00000000000000f100000000",
            INIT_6E => X"000000d600000000000000df00000000000000dc00000000000000d400000000",
            INIT_6F => X"000000ea00000000000000e300000000000000cd00000000000000c400000000",
            INIT_70 => X"0000006600000000000000640000000000000072000000000000006c00000000",
            INIT_71 => X"000000cf00000000000000a400000000000000a4000000000000009b00000000",
            INIT_72 => X"0000008a00000000000000be00000000000000e400000000000000ea00000000",
            INIT_73 => X"000000cf00000000000000a80000000000000087000000000000008300000000",
            INIT_74 => X"000000d400000000000000e300000000000000e800000000000000df00000000",
            INIT_75 => X"0000009300000000000000a300000000000000ae00000000000000c300000000",
            INIT_76 => X"0000009700000000000000980000000000000090000000000000008c00000000",
            INIT_77 => X"000000d800000000000000cb00000000000000a0000000000000009300000000",
            INIT_78 => X"000000990000000000000074000000000000005e000000000000004d00000000",
            INIT_79 => X"000000a10000000000000076000000000000006e000000000000009c00000000",
            INIT_7A => X"000000c800000000000000c600000000000000c500000000000000b600000000",
            INIT_7B => X"000000d900000000000000ec00000000000000d900000000000000ca00000000",
            INIT_7C => X"00000095000000000000009f00000000000000ac00000000000000ba00000000",
            INIT_7D => X"0000007b0000000000000076000000000000007b000000000000008a00000000",
            INIT_7E => X"000000a100000000000000910000000000000082000000000000008000000000",
            INIT_7F => X"000000d000000000000000d500000000000000b800000000000000ae00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE10;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE11 : if BRAM_NAME = "sampleifmap_layersamples_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000dc0000000000000097000000000000002f000000000000002300000000",
            INIT_01 => X"000000a20000000000000086000000000000007b000000000000009600000000",
            INIT_02 => X"000000e900000000000000e100000000000000d300000000000000b400000000",
            INIT_03 => X"000000be00000000000000ee00000000000000f000000000000000e800000000",
            INIT_04 => X"000000b100000000000000aa00000000000000a200000000000000a300000000",
            INIT_05 => X"000000bb00000000000000b600000000000000b600000000000000bb00000000",
            INIT_06 => X"000000d900000000000000cc00000000000000bf00000000000000bd00000000",
            INIT_07 => X"000000b700000000000000c100000000000000d000000000000000da00000000",
            INIT_08 => X"000000ef00000000000000d9000000000000004f000000000000001800000000",
            INIT_09 => X"000000e500000000000000da00000000000000d300000000000000d400000000",
            INIT_0A => X"000000ef00000000000000f500000000000000f600000000000000ed00000000",
            INIT_0B => X"000000ea00000000000000f100000000000000ef00000000000000dc00000000",
            INIT_0C => X"000000e500000000000000e600000000000000d600000000000000e400000000",
            INIT_0D => X"000000e000000000000000e800000000000000ea00000000000000e700000000",
            INIT_0E => X"000000b300000000000000c500000000000000d100000000000000d400000000",
            INIT_0F => X"000000a5000000000000009e00000000000000a100000000000000a900000000",
            INIT_10 => X"000000d800000000000000de00000000000000b3000000000000004700000000",
            INIT_11 => X"000000e300000000000000e600000000000000e500000000000000d900000000",
            INIT_12 => X"000000dd00000000000000e400000000000000e400000000000000e300000000",
            INIT_13 => X"000000bc00000000000000c100000000000000d700000000000000cf00000000",
            INIT_14 => X"0000009c00000000000000ba00000000000000c300000000000000b800000000",
            INIT_15 => X"0000009e00000000000000ad00000000000000b400000000000000a100000000",
            INIT_16 => X"0000008300000000000000850000000000000087000000000000008a00000000",
            INIT_17 => X"0000009c000000000000009e0000000000000097000000000000008c00000000",
            INIT_18 => X"000000bd00000000000000c200000000000000cf00000000000000a100000000",
            INIT_19 => X"000000c100000000000000c000000000000000be00000000000000bb00000000",
            INIT_1A => X"000000bd00000000000000bd00000000000000be00000000000000c000000000",
            INIT_1B => X"0000009a00000000000000a300000000000000ba00000000000000bc00000000",
            INIT_1C => X"0000009100000000000000a300000000000000aa000000000000009a00000000",
            INIT_1D => X"0000008800000000000000900000000000000099000000000000009400000000",
            INIT_1E => X"0000008d000000000000008b0000000000000086000000000000008200000000",
            INIT_1F => X"0000009c00000000000000940000000000000092000000000000009000000000",
            INIT_20 => X"0000007f000000000000007a0000000000000071000000000000006d00000000",
            INIT_21 => X"000000960000000000000093000000000000008e000000000000008600000000",
            INIT_22 => X"000000ac00000000000000a500000000000000a0000000000000009800000000",
            INIT_23 => X"000000af00000000000000b400000000000000ba00000000000000b500000000",
            INIT_24 => X"0000009b00000000000000a300000000000000a800000000000000ac00000000",
            INIT_25 => X"0000007f0000000000000084000000000000008b000000000000009400000000",
            INIT_26 => X"0000007a00000000000000810000000000000085000000000000008100000000",
            INIT_27 => X"0000009c0000000000000092000000000000008a000000000000007e00000000",
            INIT_28 => X"0000003000000000000000230000000000000019000000000000002900000000",
            INIT_29 => X"0000003d000000000000003a0000000000000038000000000000003400000000",
            INIT_2A => X"00000057000000000000004d0000000000000046000000000000003e00000000",
            INIT_2B => X"0000007e000000000000007e0000000000000079000000000000006a00000000",
            INIT_2C => X"000000700000000000000078000000000000007e000000000000007f00000000",
            INIT_2D => X"0000006600000000000000670000000000000068000000000000006a00000000",
            INIT_2E => X"000000770000000000000073000000000000006e000000000000006900000000",
            INIT_2F => X"00000095000000000000008d0000000000000088000000000000008000000000",
            INIT_30 => X"0000003500000000000000130000000000000014000000000000003700000000",
            INIT_31 => X"00000018000000000000001e0000000000000029000000000000003a00000000",
            INIT_32 => X"00000014000000000000000f000000000000000f000000000000001100000000",
            INIT_33 => X"0000003e000000000000003c0000000000000038000000000000002a00000000",
            INIT_34 => X"0000004c000000000000004d0000000000000051000000000000004700000000",
            INIT_35 => X"0000005a0000000000000053000000000000004f000000000000004e00000000",
            INIT_36 => X"0000008a000000000000008a0000000000000076000000000000006500000000",
            INIT_37 => X"0000009e00000000000000890000000000000080000000000000007d00000000",
            INIT_38 => X"000000290000000000000012000000000000001a000000000000002d00000000",
            INIT_39 => X"000000250000000000000039000000000000004c000000000000005400000000",
            INIT_3A => X"000000070000000000000007000000000000000b000000000000001500000000",
            INIT_3B => X"0000003e000000000000004e000000000000005b000000000000002300000000",
            INIT_3C => X"00000045000000000000003f000000000000003e000000000000003c00000000",
            INIT_3D => X"0000007b00000000000000630000000000000053000000000000004a00000000",
            INIT_3E => X"0000007200000000000000870000000000000095000000000000009200000000",
            INIT_3F => X"000000af00000000000000920000000000000085000000000000007400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000b00000000000000080000000000000009000000000000001100000000",
            INIT_41 => X"00000023000000000000002f0000000000000039000000000000002e00000000",
            INIT_42 => X"0000000300000000000000040000000000000007000000000000001400000000",
            INIT_43 => X"0000009400000000000000b30000000000000086000000000000000f00000000",
            INIT_44 => X"0000007f000000000000007c000000000000007d000000000000008300000000",
            INIT_45 => X"0000008d00000000000000900000000000000085000000000000007e00000000",
            INIT_46 => X"000000740000000000000061000000000000005b000000000000007400000000",
            INIT_47 => X"000000be00000000000000a50000000000000090000000000000008100000000",
            INIT_48 => X"0000000400000000000000030000000000000007000000000000002300000000",
            INIT_49 => X"0000000c00000000000000110000000000000011000000000000000700000000",
            INIT_4A => X"0000000300000000000000020000000000000003000000000000000700000000",
            INIT_4B => X"0000009400000000000000920000000000000040000000000000000200000000",
            INIT_4C => X"000000810000000000000089000000000000008d000000000000009000000000",
            INIT_4D => X"000000450000000000000053000000000000006a000000000000007a00000000",
            INIT_4E => X"0000007e00000000000000710000000000000058000000000000004600000000",
            INIT_4F => X"000000c200000000000000b0000000000000009e000000000000008700000000",
            INIT_50 => X"0000000200000000000000010000000000000015000000000000004000000000",
            INIT_51 => X"0000000500000000000000090000000000000005000000000000000000000000",
            INIT_52 => X"0000000100000000000000000000000000000000000000000000000200000000",
            INIT_53 => X"00000044000000000000003b000000000000000b000000000000000100000000",
            INIT_54 => X"0000003b00000000000000430000000000000045000000000000004300000000",
            INIT_55 => X"00000047000000000000002e000000000000002a000000000000003100000000",
            INIT_56 => X"0000008000000000000000780000000000000074000000000000006600000000",
            INIT_57 => X"000000c400000000000000b700000000000000ab000000000000009300000000",
            INIT_58 => X"000000020000000000000001000000000000002b000000000000005200000000",
            INIT_59 => X"0000000200000000000000050000000000000002000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000003600000000000000260000000000000002000000000000000000000000",
            INIT_5C => X"000000220000000000000024000000000000002b000000000000002e00000000",
            INIT_5D => X"0000006900000000000000520000000000000038000000000000002700000000",
            INIT_5E => X"0000008300000000000000760000000000000073000000000000007300000000",
            INIT_5F => X"000000c700000000000000bb00000000000000ae000000000000009600000000",
            INIT_60 => X"0000000100000000000000030000000000000032000000000000005d00000000",
            INIT_61 => X"0000000200000000000000030000000000000001000000000000000000000000",
            INIT_62 => X"0000000100000000000000000000000000000000000000000000000100000000",
            INIT_63 => X"0000002f000000000000001c0000000000000000000000000000000200000000",
            INIT_64 => X"000000370000000000000016000000000000000c000000000000001700000000",
            INIT_65 => X"00000070000000000000006f0000000000000063000000000000005100000000",
            INIT_66 => X"00000089000000000000007e0000000000000077000000000000007100000000",
            INIT_67 => X"000000c900000000000000bc00000000000000ab000000000000009700000000",
            INIT_68 => X"00000004000000000000000b0000000000000025000000000000005900000000",
            INIT_69 => X"0000000200000000000000040000000000000004000000000000000200000000",
            INIT_6A => X"0000000200000000000000010000000000000001000000000000000100000000",
            INIT_6B => X"00000018000000000000000d0000000000000002000000000000000600000000",
            INIT_6C => X"00000052000000000000003e0000000000000029000000000000001900000000",
            INIT_6D => X"0000006f00000000000000700000000000000071000000000000006500000000",
            INIT_6E => X"000000910000000000000089000000000000007e000000000000007300000000",
            INIT_6F => X"000000c900000000000000c100000000000000b300000000000000a100000000",
            INIT_70 => X"0000001100000000000000160000000000000024000000000000005200000000",
            INIT_71 => X"0000000c000000000000000d000000000000000f000000000000000f00000000",
            INIT_72 => X"0000000f000000000000000e000000000000000d000000000000000c00000000",
            INIT_73 => X"0000002d000000000000001b0000000000000015000000000000001400000000",
            INIT_74 => X"0000005800000000000000550000000000000051000000000000004300000000",
            INIT_75 => X"00000070000000000000006b000000000000006e000000000000006900000000",
            INIT_76 => X"00000097000000000000008a000000000000007f000000000000007700000000",
            INIT_77 => X"000000c800000000000000c400000000000000b700000000000000a400000000",
            INIT_78 => X"0000002500000000000000260000000000000030000000000000005300000000",
            INIT_79 => X"0000002600000000000000220000000000000021000000000000002300000000",
            INIT_7A => X"0000002e000000000000002c0000000000000029000000000000002800000000",
            INIT_7B => X"0000004a000000000000003b0000000000000030000000000000002d00000000",
            INIT_7C => X"000000610000000000000061000000000000005c000000000000005300000000",
            INIT_7D => X"00000075000000000000006c000000000000006a000000000000006b00000000",
            INIT_7E => X"00000099000000000000008d0000000000000085000000000000007b00000000",
            INIT_7F => X"000000c700000000000000bf00000000000000b200000000000000a300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE11;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE12 : if BRAM_NAME = "sampleifmap_layersamples_instance12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000084000000000000008b000000000000009e000000000000009e00000000",
            INIT_01 => X"000000c100000000000000bb00000000000000b600000000000000a600000000",
            INIT_02 => X"000000ce00000000000000d100000000000000cd00000000000000c700000000",
            INIT_03 => X"000000e600000000000000e300000000000000df00000000000000da00000000",
            INIT_04 => X"000000eb00000000000000e700000000000000e200000000000000d500000000",
            INIT_05 => X"000000ea00000000000000ea00000000000000e800000000000000ec00000000",
            INIT_06 => X"000000ee00000000000000e600000000000000e200000000000000ec00000000",
            INIT_07 => X"000000ee00000000000000ed00000000000000e400000000000000e800000000",
            INIT_08 => X"00000089000000000000009700000000000000ac00000000000000aa00000000",
            INIT_09 => X"000000c700000000000000c500000000000000c100000000000000ae00000000",
            INIT_0A => X"000000d200000000000000d900000000000000d700000000000000ce00000000",
            INIT_0B => X"000000ed00000000000000e900000000000000e700000000000000e100000000",
            INIT_0C => X"000000f200000000000000e800000000000000e400000000000000db00000000",
            INIT_0D => X"000000f200000000000000ec00000000000000ea00000000000000f500000000",
            INIT_0E => X"000000f300000000000000eb00000000000000e400000000000000f100000000",
            INIT_0F => X"000000f600000000000000f600000000000000e800000000000000e900000000",
            INIT_10 => X"0000008e000000000000009d00000000000000b000000000000000ae00000000",
            INIT_11 => X"000000c700000000000000ce00000000000000c900000000000000b500000000",
            INIT_12 => X"000000d400000000000000da00000000000000df00000000000000d100000000",
            INIT_13 => X"000000ef00000000000000e600000000000000e600000000000000e000000000",
            INIT_14 => X"000000ef00000000000000e900000000000000e400000000000000dd00000000",
            INIT_15 => X"000000f300000000000000ec00000000000000d500000000000000e800000000",
            INIT_16 => X"000000f800000000000000ee00000000000000e700000000000000f500000000",
            INIT_17 => X"000000f500000000000000fa00000000000000e600000000000000ed00000000",
            INIT_18 => X"0000009300000000000000a000000000000000b200000000000000b400000000",
            INIT_19 => X"000000cf00000000000000d400000000000000cb00000000000000ba00000000",
            INIT_1A => X"000000d600000000000000dd00000000000000e400000000000000d600000000",
            INIT_1B => X"000000f000000000000000df00000000000000e700000000000000dc00000000",
            INIT_1C => X"000000e400000000000000e900000000000000e400000000000000e000000000",
            INIT_1D => X"000000f300000000000000e600000000000000ac00000000000000b100000000",
            INIT_1E => X"000000fa00000000000000ee00000000000000e800000000000000f800000000",
            INIT_1F => X"000000f400000000000000f900000000000000e400000000000000ee00000000",
            INIT_20 => X"0000009300000000000000a500000000000000b900000000000000ba00000000",
            INIT_21 => X"000000cf00000000000000d900000000000000cc00000000000000bd00000000",
            INIT_22 => X"000000d600000000000000de00000000000000e700000000000000d300000000",
            INIT_23 => X"000000eb00000000000000d300000000000000e700000000000000da00000000",
            INIT_24 => X"000000d400000000000000e800000000000000e000000000000000e200000000",
            INIT_25 => X"000000ed00000000000000e000000000000000a8000000000000009f00000000",
            INIT_26 => X"000000f600000000000000eb00000000000000e700000000000000f700000000",
            INIT_27 => X"000000f200000000000000f800000000000000ea00000000000000e800000000",
            INIT_28 => X"0000008e00000000000000aa00000000000000be00000000000000c100000000",
            INIT_29 => X"000000d300000000000000db00000000000000cb00000000000000bf00000000",
            INIT_2A => X"000000d600000000000000dd00000000000000ea00000000000000d700000000",
            INIT_2B => X"000000cd00000000000000c700000000000000e400000000000000d600000000",
            INIT_2C => X"000000c100000000000000eb00000000000000ce00000000000000cf00000000",
            INIT_2D => X"000000e600000000000000de000000000000009e000000000000007000000000",
            INIT_2E => X"000000f100000000000000e200000000000000e500000000000000f500000000",
            INIT_2F => X"000000eb00000000000000f300000000000000e700000000000000e400000000",
            INIT_30 => X"0000008500000000000000ac00000000000000bf00000000000000c400000000",
            INIT_31 => X"000000d900000000000000de00000000000000ca00000000000000bf00000000",
            INIT_32 => X"000000d600000000000000da00000000000000eb00000000000000df00000000",
            INIT_33 => X"000000b000000000000000bc00000000000000e300000000000000d700000000",
            INIT_34 => X"000000bb00000000000000cd00000000000000ba00000000000000bb00000000",
            INIT_35 => X"000000b700000000000000ac0000000000000089000000000000007800000000",
            INIT_36 => X"000000eb00000000000000d800000000000000df00000000000000db00000000",
            INIT_37 => X"000000eb00000000000000f000000000000000e100000000000000e200000000",
            INIT_38 => X"0000008c00000000000000ae00000000000000c500000000000000cc00000000",
            INIT_39 => X"000000e000000000000000e000000000000000da00000000000000cb00000000",
            INIT_3A => X"000000dc00000000000000dc00000000000000ed00000000000000e800000000",
            INIT_3B => X"000000cd00000000000000c900000000000000dd00000000000000dc00000000",
            INIT_3C => X"000000530000000000000064000000000000008a00000000000000ac00000000",
            INIT_3D => X"0000003c0000000000000041000000000000003e000000000000004700000000",
            INIT_3E => X"000000e400000000000000d100000000000000b6000000000000006800000000",
            INIT_3F => X"000000ec00000000000000ef00000000000000d400000000000000da00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000089000000000000009d00000000000000aa00000000000000af00000000",
            INIT_41 => X"000000c500000000000000af00000000000000ba00000000000000b000000000",
            INIT_42 => X"000000d200000000000000ce00000000000000d400000000000000d100000000",
            INIT_43 => X"000000c100000000000000c100000000000000c900000000000000d400000000",
            INIT_44 => X"0000005b00000000000000590000000000000069000000000000008e00000000",
            INIT_45 => X"00000045000000000000005e0000000000000053000000000000005400000000",
            INIT_46 => X"000000b700000000000000a20000000000000079000000000000004e00000000",
            INIT_47 => X"000000c300000000000000cf00000000000000a300000000000000ae00000000",
            INIT_48 => X"0000006800000000000000710000000000000073000000000000007200000000",
            INIT_49 => X"00000080000000000000006f000000000000006b000000000000006900000000",
            INIT_4A => X"0000009b00000000000000970000000000000092000000000000008b00000000",
            INIT_4B => X"0000009600000000000000970000000000000093000000000000009d00000000",
            INIT_4C => X"0000006300000000000000630000000000000064000000000000007600000000",
            INIT_4D => X"0000005300000000000000560000000000000056000000000000005500000000",
            INIT_4E => X"00000099000000000000009a0000000000000080000000000000008b00000000",
            INIT_4F => X"0000007b0000000000000084000000000000006d000000000000007600000000",
            INIT_50 => X"00000044000000000000004b000000000000004c000000000000004200000000",
            INIT_51 => X"0000005a0000000000000054000000000000005a000000000000005300000000",
            INIT_52 => X"000000670000000000000066000000000000006a000000000000005d00000000",
            INIT_53 => X"0000006c0000000000000072000000000000006b000000000000006a00000000",
            INIT_54 => X"00000055000000000000005b000000000000005a000000000000005a00000000",
            INIT_55 => X"00000072000000000000005f0000000000000042000000000000004800000000",
            INIT_56 => X"000000c70000000000000093000000000000006e000000000000008000000000",
            INIT_57 => X"0000005e000000000000005c0000000000000067000000000000007d00000000",
            INIT_58 => X"0000004d000000000000004b0000000000000041000000000000003500000000",
            INIT_59 => X"000000460000000000000055000000000000006a000000000000006f00000000",
            INIT_5A => X"0000005d000000000000005f0000000000000071000000000000005d00000000",
            INIT_5B => X"00000061000000000000006b0000000000000073000000000000006c00000000",
            INIT_5C => X"000000610000000000000062000000000000005f000000000000006200000000",
            INIT_5D => X"000000bb00000000000000950000000000000055000000000000005a00000000",
            INIT_5E => X"000000cc0000000000000070000000000000009200000000000000b300000000",
            INIT_5F => X"000000550000000000000057000000000000005f000000000000009a00000000",
            INIT_60 => X"0000004a000000000000005e0000000000000056000000000000003a00000000",
            INIT_61 => X"00000055000000000000004d0000000000000064000000000000006400000000",
            INIT_62 => X"0000006c000000000000007f0000000000000085000000000000007800000000",
            INIT_63 => X"000000570000000000000062000000000000006e000000000000006900000000",
            INIT_64 => X"0000005f00000000000000570000000000000051000000000000005100000000",
            INIT_65 => X"000000c300000000000000aa0000000000000070000000000000005f00000000",
            INIT_66 => X"000000ad000000000000007f00000000000000c100000000000000d000000000",
            INIT_67 => X"0000004f0000000000000055000000000000005000000000000000b200000000",
            INIT_68 => X"0000004b00000000000000570000000000000059000000000000004a00000000",
            INIT_69 => X"0000005000000000000000470000000000000044000000000000005200000000",
            INIT_6A => X"0000006f00000000000000760000000000000067000000000000005900000000",
            INIT_6B => X"000000620000000000000069000000000000006a000000000000006500000000",
            INIT_6C => X"0000006d00000000000000620000000000000062000000000000006000000000",
            INIT_6D => X"000000b800000000000000b4000000000000008e000000000000007200000000",
            INIT_6E => X"0000008400000000000000a000000000000000c000000000000000bf00000000",
            INIT_6F => X"00000043000000000000003c000000000000005000000000000000aa00000000",
            INIT_70 => X"0000004e0000000000000052000000000000004f000000000000004d00000000",
            INIT_71 => X"0000005600000000000000460000000000000048000000000000004f00000000",
            INIT_72 => X"0000008500000000000000810000000000000079000000000000006d00000000",
            INIT_73 => X"0000008300000000000000870000000000000088000000000000008900000000",
            INIT_74 => X"0000009600000000000000920000000000000094000000000000009200000000",
            INIT_75 => X"000000b500000000000000b300000000000000a3000000000000009400000000",
            INIT_76 => X"0000006500000000000000aa00000000000000b000000000000000b900000000",
            INIT_77 => X"0000003b00000000000000370000000000000049000000000000005a00000000",
            INIT_78 => X"00000068000000000000006a000000000000005e000000000000006000000000",
            INIT_79 => X"0000008a00000000000000840000000000000083000000000000006d00000000",
            INIT_7A => X"0000009a000000000000009b0000000000000098000000000000009000000000",
            INIT_7B => X"00000094000000000000009e000000000000009b000000000000009b00000000",
            INIT_7C => X"00000092000000000000009c000000000000009d000000000000009600000000",
            INIT_7D => X"000000a900000000000000920000000000000082000000000000007700000000",
            INIT_7E => X"0000006900000000000000a700000000000000a800000000000000b100000000",
            INIT_7F => X"0000004800000000000000560000000000000062000000000000004500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE12;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE13 : if BRAM_NAME = "sampleifmap_layersamples_instance13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000008300000000000000730000000000000065000000000000006a00000000",
            INIT_01 => X"0000008f00000000000000900000000000000087000000000000008100000000",
            INIT_02 => X"0000009a000000000000009a0000000000000096000000000000009200000000",
            INIT_03 => X"0000009000000000000000970000000000000099000000000000009a00000000",
            INIT_04 => X"0000007f000000000000008b0000000000000086000000000000008200000000",
            INIT_05 => X"0000009f00000000000000920000000000000075000000000000005e00000000",
            INIT_06 => X"0000008400000000000000a200000000000000a300000000000000a700000000",
            INIT_07 => X"00000069000000000000009a00000000000000c0000000000000009000000000",
            INIT_08 => X"0000006d0000000000000076000000000000006c000000000000005f00000000",
            INIT_09 => X"000000910000000000000081000000000000005d000000000000005f00000000",
            INIT_0A => X"0000009000000000000000960000000000000097000000000000009500000000",
            INIT_0B => X"0000007b000000000000007a000000000000007e000000000000008600000000",
            INIT_0C => X"00000094000000000000009b0000000000000085000000000000007a00000000",
            INIT_0D => X"0000009c00000000000000a20000000000000093000000000000008300000000",
            INIT_0E => X"0000009500000000000000990000000000000097000000000000009d00000000",
            INIT_0F => X"00000094000000000000009d00000000000000a4000000000000009f00000000",
            INIT_10 => X"0000004600000000000000490000000000000059000000000000006600000000",
            INIT_11 => X"0000008c000000000000007b000000000000006f000000000000005600000000",
            INIT_12 => X"0000007500000000000000780000000000000081000000000000008f00000000",
            INIT_13 => X"0000008d0000000000000085000000000000007e000000000000007800000000",
            INIT_14 => X"0000009f0000000000000099000000000000008e000000000000009600000000",
            INIT_15 => X"000000a100000000000000a5000000000000009d000000000000009700000000",
            INIT_16 => X"00000090000000000000009a0000000000000098000000000000009900000000",
            INIT_17 => X"00000095000000000000007d0000000000000079000000000000008300000000",
            INIT_18 => X"0000006e0000000000000047000000000000003d000000000000005600000000",
            INIT_19 => X"0000007b0000000000000082000000000000008a000000000000008000000000",
            INIT_1A => X"000000840000000000000076000000000000006c000000000000007600000000",
            INIT_1B => X"00000099000000000000009c0000000000000098000000000000008f00000000",
            INIT_1C => X"0000009a00000000000000910000000000000089000000000000009500000000",
            INIT_1D => X"000000a400000000000000a0000000000000009a000000000000009900000000",
            INIT_1E => X"00000069000000000000007d0000000000000090000000000000009800000000",
            INIT_1F => X"000000840000000000000056000000000000004b000000000000005c00000000",
            INIT_20 => X"00000072000000000000006b0000000000000067000000000000006800000000",
            INIT_21 => X"00000076000000000000007b0000000000000074000000000000007300000000",
            INIT_22 => X"00000090000000000000008d0000000000000086000000000000007400000000",
            INIT_23 => X"000000750000000000000085000000000000008d000000000000008f00000000",
            INIT_24 => X"0000009600000000000000820000000000000059000000000000006200000000",
            INIT_25 => X"000000910000000000000098000000000000009a000000000000009700000000",
            INIT_26 => X"00000050000000000000005a0000000000000060000000000000007500000000",
            INIT_27 => X"0000004100000000000000490000000000000047000000000000004100000000",
            INIT_28 => X"0000006f000000000000006f000000000000006b000000000000006300000000",
            INIT_29 => X"0000007e000000000000007d0000000000000077000000000000007200000000",
            INIT_2A => X"00000081000000000000007d000000000000007d000000000000007500000000",
            INIT_2B => X"0000003d000000000000005b0000000000000082000000000000008300000000",
            INIT_2C => X"0000009400000000000000730000000000000038000000000000003900000000",
            INIT_2D => X"0000005f00000000000000720000000000000082000000000000008b00000000",
            INIT_2E => X"0000003a00000000000000490000000000000053000000000000005600000000",
            INIT_2F => X"0000001b0000000000000033000000000000004b000000000000003c00000000",
            INIT_30 => X"0000007200000000000000740000000000000068000000000000003e00000000",
            INIT_31 => X"0000005b00000000000000660000000000000075000000000000007400000000",
            INIT_32 => X"00000070000000000000004e0000000000000051000000000000005400000000",
            INIT_33 => X"0000004c00000000000000600000000000000082000000000000008500000000",
            INIT_34 => X"0000006c000000000000006b0000000000000056000000000000005300000000",
            INIT_35 => X"0000005100000000000000530000000000000058000000000000006000000000",
            INIT_36 => X"0000002d0000000000000033000000000000003d000000000000004600000000",
            INIT_37 => X"00000018000000000000001e000000000000002e000000000000003400000000",
            INIT_38 => X"00000069000000000000006a0000000000000060000000000000003900000000",
            INIT_39 => X"0000003500000000000000410000000000000068000000000000006b00000000",
            INIT_3A => X"0000006e00000000000000440000000000000040000000000000003b00000000",
            INIT_3B => X"0000006200000000000000730000000000000085000000000000008700000000",
            INIT_3C => X"00000050000000000000004e000000000000004f000000000000005800000000",
            INIT_3D => X"0000003700000000000000460000000000000050000000000000005100000000",
            INIT_3E => X"00000029000000000000002d0000000000000031000000000000002c00000000",
            INIT_3F => X"00000018000000000000001b000000000000001e000000000000002200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000690000000000000068000000000000005a000000000000004100000000",
            INIT_41 => X"00000049000000000000004f000000000000006d000000000000006d00000000",
            INIT_42 => X"0000006a00000000000000620000000000000058000000000000005500000000",
            INIT_43 => X"0000004100000000000000440000000000000053000000000000006200000000",
            INIT_44 => X"000000520000000000000051000000000000004a000000000000004600000000",
            INIT_45 => X"0000002c00000000000000290000000000000033000000000000004800000000",
            INIT_46 => X"0000002300000000000000270000000000000037000000000000003d00000000",
            INIT_47 => X"00000019000000000000001b000000000000001e000000000000002000000000",
            INIT_48 => X"0000006700000000000000690000000000000057000000000000004300000000",
            INIT_49 => X"0000005100000000000000580000000000000063000000000000006600000000",
            INIT_4A => X"00000039000000000000003b0000000000000045000000000000004c00000000",
            INIT_4B => X"000000460000000000000042000000000000003f000000000000003a00000000",
            INIT_4C => X"00000036000000000000003e0000000000000044000000000000004800000000",
            INIT_4D => X"0000002c0000000000000031000000000000002f000000000000002e00000000",
            INIT_4E => X"0000001c000000000000001e000000000000002e000000000000003800000000",
            INIT_4F => X"0000001e00000000000000180000000000000019000000000000001d00000000",
            INIT_50 => X"0000003a0000000000000041000000000000003a000000000000003600000000",
            INIT_51 => X"0000002c000000000000002d0000000000000032000000000000003700000000",
            INIT_52 => X"0000003a00000000000000370000000000000033000000000000002e00000000",
            INIT_53 => X"0000003a000000000000003e0000000000000040000000000000003e00000000",
            INIT_54 => X"0000003000000000000000250000000000000026000000000000003300000000",
            INIT_55 => X"00000026000000000000002a0000000000000030000000000000003100000000",
            INIT_56 => X"0000001c000000000000001b0000000000000020000000000000002900000000",
            INIT_57 => X"0000001f000000000000001c0000000000000019000000000000001b00000000",
            INIT_58 => X"0000001b000000000000001a000000000000001d000000000000001e00000000",
            INIT_59 => X"0000002700000000000000210000000000000020000000000000001f00000000",
            INIT_5A => X"0000003300000000000000350000000000000034000000000000003100000000",
            INIT_5B => X"0000002800000000000000260000000000000028000000000000002e00000000",
            INIT_5C => X"000000370000000000000042000000000000002c000000000000002600000000",
            INIT_5D => X"0000002500000000000000240000000000000025000000000000002900000000",
            INIT_5E => X"0000001b000000000000001a000000000000001b000000000000001f00000000",
            INIT_5F => X"000000170000000000000021000000000000001e000000000000001c00000000",
            INIT_60 => X"0000001c000000000000001b000000000000001f000000000000002100000000",
            INIT_61 => X"00000020000000000000001f000000000000001e000000000000001c00000000",
            INIT_62 => X"0000001e000000000000001e0000000000000021000000000000002300000000",
            INIT_63 => X"0000002d00000000000000290000000000000027000000000000002200000000",
            INIT_64 => X"0000003100000000000000490000000000000034000000000000002a00000000",
            INIT_65 => X"0000002000000000000000260000000000000023000000000000001e00000000",
            INIT_66 => X"0000001d000000000000001b000000000000001a000000000000001b00000000",
            INIT_67 => X"0000000d000000000000001a0000000000000026000000000000001e00000000",
            INIT_68 => X"0000001a000000000000001a000000000000001e000000000000001f00000000",
            INIT_69 => X"0000001b000000000000001a0000000000000019000000000000001900000000",
            INIT_6A => X"0000002800000000000000250000000000000020000000000000001d00000000",
            INIT_6B => X"0000002a00000000000000280000000000000029000000000000002a00000000",
            INIT_6C => X"000000260000000000000040000000000000002e000000000000002700000000",
            INIT_6D => X"0000001d000000000000001e0000000000000024000000000000001c00000000",
            INIT_6E => X"0000001c000000000000001b0000000000000019000000000000001a00000000",
            INIT_6F => X"0000000400000000000000090000000000000025000000000000002100000000",
            INIT_70 => X"0000001c0000000000000019000000000000001b000000000000001700000000",
            INIT_71 => X"0000002500000000000000220000000000000020000000000000001e00000000",
            INIT_72 => X"0000002700000000000000280000000000000027000000000000002700000000",
            INIT_73 => X"00000021000000000000001e0000000000000023000000000000002600000000",
            INIT_74 => X"0000002400000000000000390000000000000024000000000000001c00000000",
            INIT_75 => X"0000001d000000000000001d000000000000001d000000000000001e00000000",
            INIT_76 => X"0000001b00000000000000170000000000000018000000000000001800000000",
            INIT_77 => X"0000000500000000000000040000000000000013000000000000002400000000",
            INIT_78 => X"000000220000000000000020000000000000001e000000000000001c00000000",
            INIT_79 => X"0000002500000000000000230000000000000022000000000000002100000000",
            INIT_7A => X"0000002200000000000000240000000000000026000000000000002600000000",
            INIT_7B => X"0000000c000000000000000f0000000000000018000000000000001e00000000",
            INIT_7C => X"00000020000000000000002d0000000000000013000000000000000800000000",
            INIT_7D => X"0000001c000000000000001b000000000000001b000000000000001900000000",
            INIT_7E => X"0000002200000000000000140000000000000015000000000000001800000000",
            INIT_7F => X"0000000700000000000000040000000000000005000000000000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE13;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE14 : if BRAM_NAME = "sampleifmap_layersamples_instance14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009e00000000000000a600000000000000bb00000000000000be00000000",
            INIT_01 => X"000000d800000000000000d300000000000000d000000000000000c100000000",
            INIT_02 => X"000000da00000000000000de00000000000000dd00000000000000db00000000",
            INIT_03 => X"000000ed00000000000000eb00000000000000e800000000000000e500000000",
            INIT_04 => X"000000ef00000000000000ee00000000000000e900000000000000dc00000000",
            INIT_05 => X"000000f100000000000000f100000000000000ef00000000000000f100000000",
            INIT_06 => X"000000f300000000000000eb00000000000000e700000000000000f200000000",
            INIT_07 => X"000000f100000000000000ef00000000000000e700000000000000ed00000000",
            INIT_08 => X"000000a000000000000000b000000000000000c700000000000000c800000000",
            INIT_09 => X"000000da00000000000000da00000000000000d900000000000000c700000000",
            INIT_0A => X"000000db00000000000000e500000000000000e500000000000000df00000000",
            INIT_0B => X"000000f300000000000000ef00000000000000ee00000000000000e900000000",
            INIT_0C => X"000000f500000000000000ee00000000000000ea00000000000000e100000000",
            INIT_0D => X"000000f500000000000000ef00000000000000ed00000000000000f700000000",
            INIT_0E => X"000000f800000000000000ef00000000000000e900000000000000f500000000",
            INIT_0F => X"000000f700000000000000f600000000000000e800000000000000ec00000000",
            INIT_10 => X"000000a200000000000000b300000000000000c800000000000000c900000000",
            INIT_11 => X"000000d600000000000000df00000000000000dc00000000000000c900000000",
            INIT_12 => X"000000db00000000000000e200000000000000e900000000000000dd00000000",
            INIT_13 => X"000000f400000000000000ea00000000000000ea00000000000000e500000000",
            INIT_14 => X"000000f300000000000000ee00000000000000e900000000000000e200000000",
            INIT_15 => X"000000f100000000000000ea00000000000000d600000000000000eb00000000",
            INIT_16 => X"000000fa00000000000000f000000000000000e900000000000000f700000000",
            INIT_17 => X"000000f400000000000000f900000000000000e500000000000000ee00000000",
            INIT_18 => X"000000a400000000000000b300000000000000c700000000000000cb00000000",
            INIT_19 => X"000000d900000000000000e100000000000000d900000000000000c900000000",
            INIT_1A => X"000000d900000000000000e300000000000000eb00000000000000df00000000",
            INIT_1B => X"000000f400000000000000e200000000000000e800000000000000dd00000000",
            INIT_1C => X"000000eb00000000000000ed00000000000000e700000000000000e400000000",
            INIT_1D => X"000000f100000000000000e400000000000000af00000000000000b800000000",
            INIT_1E => X"000000fa00000000000000ee00000000000000e800000000000000f800000000",
            INIT_1F => X"000000f200000000000000f700000000000000e300000000000000ed00000000",
            INIT_20 => X"000000a100000000000000b500000000000000cc00000000000000cf00000000",
            INIT_21 => X"000000d500000000000000e100000000000000d600000000000000c900000000",
            INIT_22 => X"000000d700000000000000e200000000000000ed00000000000000d700000000",
            INIT_23 => X"000000ec00000000000000d400000000000000e500000000000000d900000000",
            INIT_24 => X"000000e100000000000000ec00000000000000e100000000000000e300000000",
            INIT_25 => X"000000ec00000000000000e000000000000000ae00000000000000aa00000000",
            INIT_26 => X"000000f600000000000000eb00000000000000e700000000000000f700000000",
            INIT_27 => X"000000ef00000000000000f500000000000000e700000000000000e700000000",
            INIT_28 => X"0000009a00000000000000b700000000000000cd00000000000000d000000000",
            INIT_29 => X"000000d700000000000000e200000000000000d400000000000000c900000000",
            INIT_2A => X"000000d700000000000000df00000000000000ee00000000000000da00000000",
            INIT_2B => X"000000cd00000000000000c700000000000000e500000000000000d700000000",
            INIT_2C => X"000000cc00000000000000ef00000000000000d000000000000000d100000000",
            INIT_2D => X"000000e900000000000000e300000000000000a7000000000000007c00000000",
            INIT_2E => X"000000ef00000000000000e100000000000000e500000000000000f600000000",
            INIT_2F => X"000000e800000000000000f100000000000000e600000000000000e200000000",
            INIT_30 => X"0000008b00000000000000b300000000000000c700000000000000cc00000000",
            INIT_31 => X"000000d500000000000000dd00000000000000cb00000000000000c200000000",
            INIT_32 => X"000000d400000000000000d800000000000000e900000000000000db00000000",
            INIT_33 => X"000000b000000000000000bc00000000000000e600000000000000d800000000",
            INIT_34 => X"000000c000000000000000d400000000000000c000000000000000be00000000",
            INIT_35 => X"000000be00000000000000b70000000000000097000000000000008100000000",
            INIT_36 => X"000000e500000000000000d600000000000000e000000000000000e000000000",
            INIT_37 => X"000000e000000000000000eb00000000000000de00000000000000db00000000",
            INIT_38 => X"0000008a00000000000000af00000000000000c600000000000000cd00000000",
            INIT_39 => X"000000cc00000000000000ce00000000000000cb00000000000000c000000000",
            INIT_3A => X"000000d200000000000000d000000000000000df00000000000000d400000000",
            INIT_3B => X"000000ce00000000000000c700000000000000d800000000000000d500000000",
            INIT_3C => X"0000005d0000000000000071000000000000009500000000000000b200000000",
            INIT_3D => X"0000004500000000000000500000000000000050000000000000005500000000",
            INIT_3E => X"000000de00000000000000ce00000000000000b7000000000000006c00000000",
            INIT_3F => X"000000d400000000000000dd00000000000000c500000000000000d000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000085000000000000009a00000000000000a800000000000000ad00000000",
            INIT_41 => X"000000b300000000000000a000000000000000ac00000000000000a500000000",
            INIT_42 => X"000000c300000000000000bd00000000000000c200000000000000be00000000",
            INIT_43 => X"000000c600000000000000c100000000000000bf00000000000000c700000000",
            INIT_44 => X"0000006c000000000000006b0000000000000079000000000000009800000000",
            INIT_45 => X"0000004f000000000000006e0000000000000068000000000000006800000000",
            INIT_46 => X"000000af000000000000009f000000000000007a000000000000005200000000",
            INIT_47 => X"000000af00000000000000be000000000000009500000000000000a300000000",
            INIT_48 => X"0000006900000000000000720000000000000074000000000000007300000000",
            INIT_49 => X"0000007f0000000000000070000000000000006e000000000000006d00000000",
            INIT_4A => X"00000093000000000000008c0000000000000088000000000000008700000000",
            INIT_4B => X"000000a1000000000000009e000000000000008f000000000000009700000000",
            INIT_4C => X"0000007800000000000000780000000000000077000000000000008600000000",
            INIT_4D => X"0000005c0000000000000066000000000000006c000000000000006c00000000",
            INIT_4E => X"0000009100000000000000970000000000000080000000000000008f00000000",
            INIT_4F => X"000000780000000000000082000000000000006a000000000000006e00000000",
            INIT_50 => X"0000005200000000000000560000000000000057000000000000004e00000000",
            INIT_51 => X"0000006400000000000000610000000000000069000000000000006300000000",
            INIT_52 => X"0000006f000000000000006a000000000000006d000000000000006500000000",
            INIT_53 => X"0000007f00000000000000840000000000000076000000000000007200000000",
            INIT_54 => X"0000006b000000000000006e000000000000006d000000000000006d00000000",
            INIT_55 => X"00000077000000000000006c0000000000000057000000000000006000000000",
            INIT_56 => X"000000bf0000000000000090000000000000006f000000000000008400000000",
            INIT_57 => X"000000680000000000000066000000000000006f000000000000007800000000",
            INIT_58 => X"00000062000000000000005f0000000000000055000000000000004a00000000",
            INIT_59 => X"000000510000000000000062000000000000007a000000000000008000000000",
            INIT_5A => X"0000007300000000000000710000000000000081000000000000006800000000",
            INIT_5B => X"0000007b0000000000000086000000000000008b000000000000008400000000",
            INIT_5C => X"0000007700000000000000740000000000000073000000000000007800000000",
            INIT_5D => X"000000bd000000000000009e0000000000000068000000000000007100000000",
            INIT_5E => X"000000c5000000000000006d000000000000009400000000000000b700000000",
            INIT_5F => X"0000006300000000000000630000000000000067000000000000009500000000",
            INIT_60 => X"0000005d0000000000000071000000000000006b000000000000005100000000",
            INIT_61 => X"00000066000000000000005d0000000000000073000000000000007500000000",
            INIT_62 => X"0000008300000000000000950000000000000098000000000000008900000000",
            INIT_63 => X"00000071000000000000007d0000000000000088000000000000008200000000",
            INIT_64 => X"0000007b0000000000000072000000000000006c000000000000006c00000000",
            INIT_65 => X"000000c200000000000000af000000000000007f000000000000007600000000",
            INIT_66 => X"000000a2000000000000007600000000000000bd00000000000000ce00000000",
            INIT_67 => X"000000650000000000000062000000000000005000000000000000a700000000",
            INIT_68 => X"0000005d000000000000006a000000000000006e000000000000006100000000",
            INIT_69 => X"0000006400000000000000590000000000000054000000000000006200000000",
            INIT_6A => X"00000086000000000000008a000000000000007b000000000000006e00000000",
            INIT_6B => X"0000007c00000000000000820000000000000083000000000000007e00000000",
            INIT_6C => X"00000087000000000000007e000000000000007f000000000000007b00000000",
            INIT_6D => X"000000b400000000000000b50000000000000099000000000000008600000000",
            INIT_6E => X"0000007a000000000000009700000000000000b700000000000000b800000000",
            INIT_6F => X"000000590000000000000048000000000000004d00000000000000a000000000",
            INIT_70 => X"0000006100000000000000660000000000000065000000000000006600000000",
            INIT_71 => X"0000006b00000000000000580000000000000058000000000000005f00000000",
            INIT_72 => X"0000009e0000000000000097000000000000008e000000000000008200000000",
            INIT_73 => X"0000009d00000000000000a100000000000000a400000000000000a300000000",
            INIT_74 => X"000000a900000000000000aa00000000000000ad00000000000000ab00000000",
            INIT_75 => X"000000ae00000000000000b100000000000000a900000000000000a200000000",
            INIT_76 => X"0000006200000000000000a400000000000000a800000000000000b000000000",
            INIT_77 => X"0000004b000000000000003f0000000000000046000000000000005700000000",
            INIT_78 => X"0000007c000000000000007f0000000000000076000000000000007b00000000",
            INIT_79 => X"000000a000000000000000980000000000000094000000000000007e00000000",
            INIT_7A => X"000000b400000000000000b300000000000000af00000000000000a700000000",
            INIT_7B => X"000000ae00000000000000b900000000000000b800000000000000b700000000",
            INIT_7C => X"000000a000000000000000af00000000000000b200000000000000ad00000000",
            INIT_7D => X"000000a1000000000000008e0000000000000085000000000000008000000000",
            INIT_7E => X"0000006c00000000000000a600000000000000a200000000000000a900000000",
            INIT_7F => X"000000520000000000000059000000000000005f000000000000004600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE14;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE15 : if BRAM_NAME = "sampleifmap_layersamples_instance15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000098000000000000008a000000000000007d000000000000008500000000",
            INIT_01 => X"000000a700000000000000a6000000000000009a000000000000009400000000",
            INIT_02 => X"000000b600000000000000b300000000000000ae00000000000000aa00000000",
            INIT_03 => X"000000ab00000000000000b500000000000000b900000000000000b900000000",
            INIT_04 => X"0000008b000000000000009a0000000000000098000000000000009800000000",
            INIT_05 => X"0000009b00000000000000900000000000000078000000000000006600000000",
            INIT_06 => X"0000008800000000000000a300000000000000a200000000000000a500000000",
            INIT_07 => X"0000006c000000000000009900000000000000bb000000000000009100000000",
            INIT_08 => X"00000083000000000000008d0000000000000085000000000000007c00000000",
            INIT_09 => X"000000aa00000000000000980000000000000072000000000000007400000000",
            INIT_0A => X"000000ad00000000000000b000000000000000af00000000000000af00000000",
            INIT_0B => X"00000097000000000000009a00000000000000a000000000000000a700000000",
            INIT_0C => X"000000a000000000000000a80000000000000096000000000000009000000000",
            INIT_0D => X"0000009e00000000000000a50000000000000098000000000000008c00000000",
            INIT_0E => X"00000097000000000000009c000000000000009b00000000000000a300000000",
            INIT_0F => X"000000930000000000000098000000000000009e000000000000009e00000000",
            INIT_10 => X"0000005d00000000000000600000000000000071000000000000008100000000",
            INIT_11 => X"000000a400000000000000940000000000000087000000000000006e00000000",
            INIT_12 => X"000000920000000000000096000000000000009f00000000000000a900000000",
            INIT_13 => X"000000a5000000000000009f0000000000000099000000000000009400000000",
            INIT_14 => X"000000ac00000000000000a800000000000000a000000000000000aa00000000",
            INIT_15 => X"000000a400000000000000a800000000000000a400000000000000a100000000",
            INIT_16 => X"00000092000000000000009e000000000000009e00000000000000a000000000",
            INIT_17 => X"00000096000000000000007d0000000000000079000000000000008400000000",
            INIT_18 => X"0000008700000000000000600000000000000055000000000000007000000000",
            INIT_19 => X"00000093000000000000009c00000000000000a5000000000000009b00000000",
            INIT_1A => X"000000a00000000000000097000000000000008d000000000000008e00000000",
            INIT_1B => X"000000ab00000000000000ae00000000000000ad00000000000000a700000000",
            INIT_1C => X"000000a800000000000000a2000000000000009b00000000000000a700000000",
            INIT_1D => X"000000a600000000000000a300000000000000a100000000000000a300000000",
            INIT_1E => X"0000006f00000000000000820000000000000097000000000000009e00000000",
            INIT_1F => X"0000008a000000000000005c0000000000000052000000000000006200000000",
            INIT_20 => X"0000008f00000000000000870000000000000084000000000000008500000000",
            INIT_21 => X"0000008e0000000000000096000000000000008f000000000000008f00000000",
            INIT_22 => X"000000ab00000000000000a900000000000000a1000000000000008a00000000",
            INIT_23 => X"00000086000000000000009700000000000000a500000000000000a900000000",
            INIT_24 => X"000000a40000000000000094000000000000006b000000000000007400000000",
            INIT_25 => X"00000098000000000000009f00000000000000a300000000000000a300000000",
            INIT_26 => X"0000005b0000000000000066000000000000006c000000000000008000000000",
            INIT_27 => X"000000480000000000000050000000000000004e000000000000004b00000000",
            INIT_28 => X"0000008f0000000000000090000000000000008c000000000000008400000000",
            INIT_29 => X"0000009600000000000000970000000000000093000000000000009000000000",
            INIT_2A => X"0000009a00000000000000940000000000000092000000000000008b00000000",
            INIT_2B => X"0000004e000000000000006e000000000000009c000000000000009f00000000",
            INIT_2C => X"000000a30000000000000084000000000000004a000000000000004b00000000",
            INIT_2D => X"0000006d000000000000007e000000000000008f000000000000009900000000",
            INIT_2E => X"0000004c000000000000005a0000000000000064000000000000006700000000",
            INIT_2F => X"0000002100000000000000390000000000000052000000000000004b00000000",
            INIT_30 => X"0000009200000000000000940000000000000089000000000000005e00000000",
            INIT_31 => X"0000007300000000000000810000000000000091000000000000009200000000",
            INIT_32 => X"0000008700000000000000630000000000000066000000000000006a00000000",
            INIT_33 => X"0000005d0000000000000072000000000000009a000000000000009d00000000",
            INIT_34 => X"0000007c000000000000007d0000000000000068000000000000006500000000",
            INIT_35 => X"000000650000000000000066000000000000006a000000000000007100000000",
            INIT_36 => X"0000003f0000000000000045000000000000004f000000000000005800000000",
            INIT_37 => X"0000001f00000000000000250000000000000035000000000000004300000000",
            INIT_38 => X"000000860000000000000086000000000000007d000000000000005600000000",
            INIT_39 => X"0000004d000000000000005c0000000000000085000000000000008900000000",
            INIT_3A => X"00000083000000000000005c0000000000000059000000000000005200000000",
            INIT_3B => X"0000007300000000000000840000000000000096000000000000009900000000",
            INIT_3C => X"0000006100000000000000600000000000000061000000000000006a00000000",
            INIT_3D => X"0000004f000000000000005f0000000000000065000000000000006300000000",
            INIT_3E => X"00000039000000000000003c0000000000000040000000000000003c00000000",
            INIT_3F => X"0000001f00000000000000220000000000000026000000000000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008300000000000000810000000000000074000000000000005a00000000",
            INIT_41 => X"00000061000000000000006a000000000000008a000000000000008900000000",
            INIT_42 => X"0000007e000000000000007c0000000000000074000000000000006c00000000",
            INIT_43 => X"000000530000000000000054000000000000005f000000000000007100000000",
            INIT_44 => X"000000640000000000000062000000000000005c000000000000005900000000",
            INIT_45 => X"000000450000000000000043000000000000004a000000000000005c00000000",
            INIT_46 => X"0000002e00000000000000330000000000000042000000000000004a00000000",
            INIT_47 => X"0000002000000000000000230000000000000026000000000000002b00000000",
            INIT_48 => X"0000007f00000000000000820000000000000070000000000000005c00000000",
            INIT_49 => X"00000066000000000000006e0000000000000078000000000000007c00000000",
            INIT_4A => X"0000004c0000000000000050000000000000005a000000000000006100000000",
            INIT_4B => X"0000005b00000000000000540000000000000050000000000000004b00000000",
            INIT_4C => X"0000004900000000000000510000000000000059000000000000005f00000000",
            INIT_4D => X"0000003d00000000000000430000000000000041000000000000004100000000",
            INIT_4E => X"00000028000000000000002a000000000000003a000000000000004500000000",
            INIT_4F => X"0000002500000000000000230000000000000028000000000000002a00000000",
            INIT_50 => X"0000004e0000000000000056000000000000004f000000000000004c00000000",
            INIT_51 => X"0000003f00000000000000400000000000000045000000000000004a00000000",
            INIT_52 => X"0000004d000000000000004a0000000000000046000000000000004100000000",
            INIT_53 => X"0000005000000000000000510000000000000052000000000000005100000000",
            INIT_54 => X"000000440000000000000037000000000000003b000000000000004900000000",
            INIT_55 => X"000000320000000000000036000000000000003f000000000000004300000000",
            INIT_56 => X"000000280000000000000028000000000000002d000000000000003600000000",
            INIT_57 => X"0000002500000000000000270000000000000028000000000000002900000000",
            INIT_58 => X"0000002a0000000000000028000000000000002b000000000000002d00000000",
            INIT_59 => X"0000003a00000000000000350000000000000034000000000000003100000000",
            INIT_5A => X"0000004600000000000000480000000000000047000000000000004400000000",
            INIT_5B => X"0000003b000000000000003a000000000000003b000000000000004100000000",
            INIT_5C => X"000000490000000000000055000000000000003f000000000000003800000000",
            INIT_5D => X"0000002f000000000000002f0000000000000033000000000000003900000000",
            INIT_5E => X"0000002800000000000000270000000000000028000000000000002c00000000",
            INIT_5F => X"0000001d000000000000002a000000000000002a000000000000002900000000",
            INIT_60 => X"0000002600000000000000240000000000000028000000000000002b00000000",
            INIT_61 => X"0000003200000000000000310000000000000030000000000000002c00000000",
            INIT_62 => X"0000003100000000000000310000000000000034000000000000003500000000",
            INIT_63 => X"0000003d000000000000003e000000000000003b000000000000003500000000",
            INIT_64 => X"00000042000000000000005e0000000000000045000000000000003700000000",
            INIT_65 => X"00000028000000000000002f000000000000002e000000000000002c00000000",
            INIT_66 => X"0000002a00000000000000280000000000000027000000000000002700000000",
            INIT_67 => X"000000120000000000000020000000000000002e000000000000002900000000",
            INIT_68 => X"0000002400000000000000230000000000000027000000000000002800000000",
            INIT_69 => X"0000002b00000000000000290000000000000029000000000000002700000000",
            INIT_6A => X"0000003a00000000000000380000000000000033000000000000002e00000000",
            INIT_6B => X"00000037000000000000003c000000000000003d000000000000003d00000000",
            INIT_6C => X"000000360000000000000055000000000000003c000000000000002e00000000",
            INIT_6D => X"000000240000000000000025000000000000002e000000000000002800000000",
            INIT_6E => X"0000002a00000000000000280000000000000026000000000000002600000000",
            INIT_6F => X"00000007000000000000000d0000000000000028000000000000002b00000000",
            INIT_70 => X"0000002800000000000000240000000000000026000000000000002200000000",
            INIT_71 => X"000000330000000000000031000000000000002f000000000000002c00000000",
            INIT_72 => X"00000039000000000000003b0000000000000039000000000000003600000000",
            INIT_73 => X"0000002b00000000000000330000000000000037000000000000003900000000",
            INIT_74 => X"00000032000000000000004e0000000000000030000000000000001f00000000",
            INIT_75 => X"0000002300000000000000230000000000000025000000000000002900000000",
            INIT_76 => X"0000002900000000000000240000000000000025000000000000002500000000",
            INIT_77 => X"0000000700000000000000060000000000000014000000000000002d00000000",
            INIT_78 => X"0000002f000000000000002d000000000000002b000000000000002900000000",
            INIT_79 => X"0000003100000000000000300000000000000030000000000000003000000000",
            INIT_7A => X"0000002d00000000000000310000000000000033000000000000003200000000",
            INIT_7B => X"00000011000000000000001a0000000000000022000000000000002800000000",
            INIT_7C => X"0000002c000000000000003f000000000000001b000000000000000800000000",
            INIT_7D => X"0000002300000000000000220000000000000022000000000000002100000000",
            INIT_7E => X"0000002c00000000000000220000000000000022000000000000002300000000",
            INIT_7F => X"0000000800000000000000050000000000000006000000000000001f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE15;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE16 : if BRAM_NAME = "sampleifmap_layersamples_instance16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ba00000000000000c200000000000000da00000000000000de00000000",
            INIT_01 => X"000000f100000000000000ee00000000000000ec00000000000000de00000000",
            INIT_02 => X"000000eb00000000000000f400000000000000f500000000000000f300000000",
            INIT_03 => X"000000f500000000000000f200000000000000f100000000000000f000000000",
            INIT_04 => X"000000f800000000000000f500000000000000f000000000000000e300000000",
            INIT_05 => X"000000f300000000000000f300000000000000f300000000000000f900000000",
            INIT_06 => X"000000f700000000000000ef00000000000000eb00000000000000f500000000",
            INIT_07 => X"000000f600000000000000f300000000000000ea00000000000000f100000000",
            INIT_08 => X"000000b800000000000000c900000000000000e200000000000000e500000000",
            INIT_09 => X"000000ee00000000000000f000000000000000f000000000000000df00000000",
            INIT_0A => X"000000e800000000000000f500000000000000f700000000000000f300000000",
            INIT_0B => X"000000f800000000000000f500000000000000f500000000000000f300000000",
            INIT_0C => X"000000fb00000000000000f300000000000000ef00000000000000e600000000",
            INIT_0D => X"000000f400000000000000ee00000000000000ee00000000000000fb00000000",
            INIT_0E => X"000000fc00000000000000f300000000000000ec00000000000000f800000000",
            INIT_0F => X"000000fb00000000000000fa00000000000000ec00000000000000f000000000",
            INIT_10 => X"000000b500000000000000c700000000000000de00000000000000e100000000",
            INIT_11 => X"000000e400000000000000ef00000000000000ee00000000000000db00000000",
            INIT_12 => X"000000e400000000000000ec00000000000000f400000000000000eb00000000",
            INIT_13 => X"000000f700000000000000ee00000000000000ef00000000000000eb00000000",
            INIT_14 => X"000000f600000000000000f100000000000000ec00000000000000e500000000",
            INIT_15 => X"000000ef00000000000000e800000000000000d700000000000000ec00000000",
            INIT_16 => X"000000fc00000000000000f200000000000000eb00000000000000f800000000",
            INIT_17 => X"000000f700000000000000fb00000000000000e800000000000000f100000000",
            INIT_18 => X"000000b300000000000000c200000000000000d800000000000000de00000000",
            INIT_19 => X"000000e100000000000000eb00000000000000e400000000000000d600000000",
            INIT_1A => X"000000dd00000000000000e600000000000000ef00000000000000e500000000",
            INIT_1B => X"000000f700000000000000e600000000000000ec00000000000000e100000000",
            INIT_1C => X"000000ee00000000000000f000000000000000ea00000000000000e600000000",
            INIT_1D => X"000000f100000000000000e500000000000000b000000000000000ba00000000",
            INIT_1E => X"000000fb00000000000000ef00000000000000e900000000000000f800000000",
            INIT_1F => X"000000f300000000000000f800000000000000e400000000000000ee00000000",
            INIT_20 => X"000000ac00000000000000c100000000000000d900000000000000df00000000",
            INIT_21 => X"000000d900000000000000e700000000000000dd00000000000000d200000000",
            INIT_22 => X"000000d700000000000000e100000000000000eb00000000000000da00000000",
            INIT_23 => X"000000ee00000000000000d600000000000000e800000000000000db00000000",
            INIT_24 => X"000000e400000000000000ee00000000000000e300000000000000e500000000",
            INIT_25 => X"000000ef00000000000000e500000000000000b200000000000000b000000000",
            INIT_26 => X"000000f500000000000000ea00000000000000e700000000000000f700000000",
            INIT_27 => X"000000f000000000000000f600000000000000e800000000000000e700000000",
            INIT_28 => X"000000a400000000000000bf00000000000000d500000000000000dc00000000",
            INIT_29 => X"000000d500000000000000e100000000000000d500000000000000ce00000000",
            INIT_2A => X"000000d600000000000000da00000000000000e600000000000000d600000000",
            INIT_2B => X"000000ce00000000000000c800000000000000e300000000000000d600000000",
            INIT_2C => X"000000cf00000000000000ed00000000000000ce00000000000000d000000000",
            INIT_2D => X"000000e900000000000000e600000000000000ad000000000000008200000000",
            INIT_2E => X"000000e800000000000000db00000000000000e100000000000000f400000000",
            INIT_2F => X"000000e600000000000000f200000000000000e700000000000000dd00000000",
            INIT_30 => X"0000009600000000000000b900000000000000ca00000000000000d400000000",
            INIT_31 => X"000000d000000000000000d900000000000000c900000000000000c400000000",
            INIT_32 => X"000000d300000000000000d000000000000000db00000000000000d300000000",
            INIT_33 => X"000000af00000000000000b900000000000000dd00000000000000d400000000",
            INIT_34 => X"000000c500000000000000d200000000000000bd00000000000000bb00000000",
            INIT_35 => X"000000bb00000000000000b8000000000000009d000000000000008900000000",
            INIT_36 => X"000000da00000000000000ce00000000000000dc00000000000000dd00000000",
            INIT_37 => X"000000d800000000000000e700000000000000db00000000000000d100000000",
            INIT_38 => X"0000009300000000000000b300000000000000c900000000000000d300000000",
            INIT_39 => X"000000cb00000000000000ce00000000000000cc00000000000000c500000000",
            INIT_3A => X"000000cd00000000000000c600000000000000d200000000000000d000000000",
            INIT_3B => X"000000cb00000000000000c000000000000000ce00000000000000ce00000000",
            INIT_3C => X"0000006a000000000000007a000000000000009b00000000000000b300000000",
            INIT_3D => X"000000490000000000000058000000000000005e000000000000006400000000",
            INIT_3E => X"000000d700000000000000ca00000000000000b7000000000000006f00000000",
            INIT_3F => X"000000c100000000000000ce00000000000000b900000000000000c600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008c00000000000000a000000000000000ad00000000000000b300000000",
            INIT_41 => X"000000b300000000000000a100000000000000af00000000000000aa00000000",
            INIT_42 => X"000000bd00000000000000b400000000000000b800000000000000bb00000000",
            INIT_43 => X"000000c400000000000000ba00000000000000b900000000000000c300000000",
            INIT_44 => X"0000008000000000000000800000000000000089000000000000009f00000000",
            INIT_45 => X"0000005a0000000000000080000000000000007e000000000000007e00000000",
            INIT_46 => X"000000ac000000000000009e000000000000007c000000000000005800000000",
            INIT_47 => X"0000009f00000000000000b00000000000000089000000000000009c00000000",
            INIT_48 => X"00000070000000000000007b000000000000007e000000000000007b00000000",
            INIT_49 => X"0000008000000000000000720000000000000072000000000000007200000000",
            INIT_4A => X"0000009000000000000000890000000000000086000000000000008600000000",
            INIT_4B => X"000000a700000000000000a00000000000000092000000000000009800000000",
            INIT_4C => X"0000008c0000000000000090000000000000008b000000000000009300000000",
            INIT_4D => X"0000006800000000000000780000000000000083000000000000008200000000",
            INIT_4E => X"0000008d00000000000000960000000000000083000000000000009500000000",
            INIT_4F => X"0000007500000000000000800000000000000069000000000000006a00000000",
            INIT_50 => X"0000005800000000000000620000000000000066000000000000005900000000",
            INIT_51 => X"0000006a00000000000000680000000000000073000000000000006b00000000",
            INIT_52 => X"0000007300000000000000710000000000000076000000000000006b00000000",
            INIT_53 => X"0000009200000000000000970000000000000086000000000000007b00000000",
            INIT_54 => X"00000078000000000000007f000000000000007f000000000000008000000000",
            INIT_55 => X"00000080000000000000007a0000000000000068000000000000006f00000000",
            INIT_56 => X"000000b6000000000000008b000000000000006e000000000000008600000000",
            INIT_57 => X"00000070000000000000006d0000000000000075000000000000007200000000",
            INIT_58 => X"0000006a000000000000006e0000000000000068000000000000005800000000",
            INIT_59 => X"0000005e00000000000000710000000000000089000000000000008e00000000",
            INIT_5A => X"0000007d000000000000007f0000000000000092000000000000007400000000",
            INIT_5B => X"0000009700000000000000a500000000000000a5000000000000009400000000",
            INIT_5C => X"0000007f000000000000007f0000000000000082000000000000008e00000000",
            INIT_5D => X"000000bf00000000000000a50000000000000072000000000000007b00000000",
            INIT_5E => X"000000b80000000000000064000000000000008e00000000000000b400000000",
            INIT_5F => X"0000006c000000000000006c000000000000006d000000000000008c00000000",
            INIT_60 => X"0000006800000000000000840000000000000082000000000000006400000000",
            INIT_61 => X"00000076000000000000006d0000000000000082000000000000008100000000",
            INIT_62 => X"0000009700000000000000a800000000000000ab000000000000009a00000000",
            INIT_63 => X"0000008b000000000000009a00000000000000a5000000000000009b00000000",
            INIT_64 => X"0000008c0000000000000081000000000000007d000000000000008200000000",
            INIT_65 => X"000000c100000000000000b30000000000000089000000000000008600000000",
            INIT_66 => X"00000098000000000000007000000000000000b900000000000000cb00000000",
            INIT_67 => X"0000006d0000000000000069000000000000005400000000000000a000000000",
            INIT_68 => X"0000006a000000000000007e0000000000000086000000000000007800000000",
            INIT_69 => X"00000079000000000000006c0000000000000065000000000000007100000000",
            INIT_6A => X"0000009f00000000000000a10000000000000091000000000000008300000000",
            INIT_6B => X"00000095000000000000009e00000000000000a1000000000000009900000000",
            INIT_6C => X"0000009b00000000000000910000000000000093000000000000009200000000",
            INIT_6D => X"000000b100000000000000b600000000000000a1000000000000009600000000",
            INIT_6E => X"00000076000000000000009400000000000000b500000000000000b500000000",
            INIT_6F => X"00000060000000000000004e0000000000000050000000000000009d00000000",
            INIT_70 => X"00000072000000000000007d0000000000000080000000000000007f00000000",
            INIT_71 => X"0000008600000000000000730000000000000071000000000000007400000000",
            INIT_72 => X"000000b800000000000000b000000000000000a8000000000000009f00000000",
            INIT_73 => X"000000b900000000000000be00000000000000bf00000000000000be00000000",
            INIT_74 => X"000000b800000000000000be00000000000000c400000000000000c500000000",
            INIT_75 => X"000000a800000000000000af00000000000000ad00000000000000ac00000000",
            INIT_76 => X"0000006300000000000000a300000000000000a500000000000000ab00000000",
            INIT_77 => X"0000005100000000000000430000000000000047000000000000005700000000",
            INIT_78 => X"00000091000000000000009a0000000000000095000000000000009700000000",
            INIT_79 => X"000000c100000000000000b800000000000000b3000000000000009900000000",
            INIT_7A => X"000000d000000000000000cf00000000000000cd00000000000000c900000000",
            INIT_7B => X"000000c800000000000000d400000000000000d200000000000000d100000000",
            INIT_7C => X"000000ab00000000000000c300000000000000c900000000000000c600000000",
            INIT_7D => X"0000009b000000000000008b0000000000000087000000000000008600000000",
            INIT_7E => X"0000007100000000000000a800000000000000a100000000000000a500000000",
            INIT_7F => X"00000056000000000000005a000000000000005c000000000000004900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE16;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE17 : if BRAM_NAME = "sampleifmap_layersamples_instance17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b000000000000000a7000000000000009f00000000000000a500000000",
            INIT_01 => X"000000c900000000000000c600000000000000b900000000000000af00000000",
            INIT_02 => X"000000d200000000000000d200000000000000d000000000000000cd00000000",
            INIT_03 => X"000000be00000000000000c900000000000000d000000000000000d200000000",
            INIT_04 => X"0000009400000000000000a900000000000000aa00000000000000aa00000000",
            INIT_05 => X"00000099000000000000008e000000000000007a000000000000006c00000000",
            INIT_06 => X"0000008e00000000000000a700000000000000a500000000000000a700000000",
            INIT_07 => X"0000006f000000000000009800000000000000b5000000000000009300000000",
            INIT_08 => X"0000009d00000000000000ae00000000000000aa000000000000009d00000000",
            INIT_09 => X"000000ca00000000000000b6000000000000008f000000000000008d00000000",
            INIT_0A => X"000000ca00000000000000d100000000000000d300000000000000d000000000",
            INIT_0B => X"000000a200000000000000a700000000000000b500000000000000bf00000000",
            INIT_0C => X"000000a900000000000000b200000000000000a0000000000000009b00000000",
            INIT_0D => X"000000a000000000000000a7000000000000009d000000000000009300000000",
            INIT_0E => X"0000009c00000000000000a100000000000000a200000000000000a900000000",
            INIT_0F => X"0000009400000000000000960000000000000096000000000000009e00000000",
            INIT_10 => X"000000790000000000000080000000000000009400000000000000a200000000",
            INIT_11 => X"000000c200000000000000b100000000000000a4000000000000008a00000000",
            INIT_12 => X"000000ab00000000000000b200000000000000bc00000000000000c700000000",
            INIT_13 => X"000000b000000000000000ac00000000000000ac00000000000000aa00000000",
            INIT_14 => X"000000b500000000000000b000000000000000a800000000000000b400000000",
            INIT_15 => X"000000ac00000000000000af00000000000000ad00000000000000aa00000000",
            INIT_16 => X"0000009600000000000000a300000000000000a500000000000000a800000000",
            INIT_17 => X"00000099000000000000007d0000000000000076000000000000008500000000",
            INIT_18 => X"000000a6000000000000007f0000000000000075000000000000008f00000000",
            INIT_19 => X"000000b000000000000000ba00000000000000c500000000000000bc00000000",
            INIT_1A => X"000000b200000000000000ab00000000000000a300000000000000a900000000",
            INIT_1B => X"000000ba00000000000000bf00000000000000be00000000000000b900000000",
            INIT_1C => X"000000b100000000000000ac00000000000000a500000000000000b400000000",
            INIT_1D => X"000000b200000000000000af00000000000000ac00000000000000ad00000000",
            INIT_1E => X"000000740000000000000088000000000000009c00000000000000a400000000",
            INIT_1F => X"0000009000000000000000620000000000000057000000000000006700000000",
            INIT_20 => X"000000b000000000000000a800000000000000a500000000000000a600000000",
            INIT_21 => X"000000aa00000000000000b300000000000000ae00000000000000b000000000",
            INIT_22 => X"000000bd00000000000000be00000000000000b800000000000000a400000000",
            INIT_23 => X"0000009600000000000000a800000000000000b500000000000000b900000000",
            INIT_24 => X"000000ad000000000000009d0000000000000076000000000000008100000000",
            INIT_25 => X"000000a200000000000000ab00000000000000ad00000000000000ad00000000",
            INIT_26 => X"0000005f000000000000006a0000000000000070000000000000008500000000",
            INIT_27 => X"0000004e00000000000000560000000000000054000000000000005000000000",
            INIT_28 => X"000000af00000000000000b100000000000000ac00000000000000a500000000",
            INIT_29 => X"000000b000000000000000b300000000000000b000000000000000ae00000000",
            INIT_2A => X"000000ad00000000000000ab00000000000000ab00000000000000a400000000",
            INIT_2B => X"0000005e000000000000007e00000000000000ab00000000000000af00000000",
            INIT_2C => X"000000ac000000000000008e0000000000000055000000000000005800000000",
            INIT_2D => X"000000750000000000000088000000000000009800000000000000a200000000",
            INIT_2E => X"00000050000000000000005e0000000000000068000000000000006c00000000",
            INIT_2F => X"00000027000000000000003f0000000000000058000000000000004f00000000",
            INIT_30 => X"000000af00000000000000b200000000000000a6000000000000007c00000000",
            INIT_31 => X"0000008b000000000000009a00000000000000ad00000000000000af00000000",
            INIT_32 => X"0000009a000000000000007a000000000000007e000000000000008200000000",
            INIT_33 => X"0000006c000000000000008300000000000000a900000000000000ae00000000",
            INIT_34 => X"0000008500000000000000860000000000000072000000000000007200000000",
            INIT_35 => X"0000006c000000000000006d0000000000000071000000000000007900000000",
            INIT_36 => X"00000045000000000000004b0000000000000056000000000000005f00000000",
            INIT_37 => X"00000026000000000000002b000000000000003b000000000000004900000000",
            INIT_38 => X"0000009f00000000000000a00000000000000096000000000000006f00000000",
            INIT_39 => X"000000640000000000000074000000000000009e00000000000000a300000000",
            INIT_3A => X"0000009700000000000000730000000000000070000000000000006800000000",
            INIT_3B => X"00000083000000000000009500000000000000a800000000000000ac00000000",
            INIT_3C => X"0000006a000000000000006a000000000000006b000000000000007700000000",
            INIT_3D => X"000000540000000000000064000000000000006c000000000000006a00000000",
            INIT_3E => X"0000004100000000000000440000000000000049000000000000004500000000",
            INIT_3F => X"000000250000000000000028000000000000002c000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009a0000000000000097000000000000008a000000000000007100000000",
            INIT_41 => X"00000077000000000000008000000000000000a200000000000000a100000000",
            INIT_42 => X"0000009200000000000000900000000000000088000000000000008100000000",
            INIT_43 => X"0000006200000000000000650000000000000072000000000000008400000000",
            INIT_44 => X"0000006c000000000000006d0000000000000067000000000000006500000000",
            INIT_45 => X"0000004b00000000000000480000000000000050000000000000006300000000",
            INIT_46 => X"0000003a000000000000003d000000000000004d000000000000005500000000",
            INIT_47 => X"000000270000000000000029000000000000002d000000000000003400000000",
            INIT_48 => X"00000097000000000000009a0000000000000088000000000000007400000000",
            INIT_49 => X"0000007c0000000000000084000000000000008f000000000000009400000000",
            INIT_4A => X"00000057000000000000005b0000000000000067000000000000007600000000",
            INIT_4B => X"000000650000000000000063000000000000005b000000000000005600000000",
            INIT_4C => X"00000052000000000000005e0000000000000063000000000000006500000000",
            INIT_4D => X"00000045000000000000004a0000000000000048000000000000004800000000",
            INIT_4E => X"0000003200000000000000340000000000000044000000000000004e00000000",
            INIT_4F => X"00000030000000000000002f0000000000000030000000000000003300000000",
            INIT_50 => X"00000063000000000000006a0000000000000064000000000000006000000000",
            INIT_51 => X"0000005100000000000000520000000000000056000000000000005c00000000",
            INIT_52 => X"000000540000000000000051000000000000004f000000000000005200000000",
            INIT_53 => X"00000058000000000000005e000000000000005b000000000000005700000000",
            INIT_54 => X"0000004c00000000000000440000000000000044000000000000004d00000000",
            INIT_55 => X"0000003b00000000000000400000000000000048000000000000004a00000000",
            INIT_56 => X"0000003200000000000000310000000000000036000000000000003f00000000",
            INIT_57 => X"0000003000000000000000340000000000000030000000000000003100000000",
            INIT_58 => X"0000003700000000000000360000000000000039000000000000003b00000000",
            INIT_59 => X"00000044000000000000003e000000000000003d000000000000003c00000000",
            INIT_5A => X"0000004d000000000000004f000000000000004f000000000000004e00000000",
            INIT_5B => X"0000004200000000000000450000000000000044000000000000004800000000",
            INIT_5C => X"0000005200000000000000610000000000000047000000000000003d00000000",
            INIT_5D => X"000000390000000000000038000000000000003c000000000000004100000000",
            INIT_5E => X"0000003100000000000000300000000000000031000000000000003500000000",
            INIT_5F => X"0000002300000000000000320000000000000032000000000000003200000000",
            INIT_60 => X"0000002d000000000000002c0000000000000030000000000000003200000000",
            INIT_61 => X"0000003700000000000000350000000000000035000000000000003100000000",
            INIT_62 => X"000000380000000000000038000000000000003b000000000000003a00000000",
            INIT_63 => X"0000004400000000000000470000000000000042000000000000003c00000000",
            INIT_64 => X"0000004b0000000000000068000000000000004b000000000000003b00000000",
            INIT_65 => X"00000033000000000000003a0000000000000038000000000000003500000000",
            INIT_66 => X"0000003300000000000000310000000000000030000000000000003100000000",
            INIT_67 => X"0000001400000000000000250000000000000035000000000000003200000000",
            INIT_68 => X"000000290000000000000028000000000000002c000000000000002d00000000",
            INIT_69 => X"00000030000000000000002e000000000000002e000000000000002c00000000",
            INIT_6A => X"00000041000000000000003f0000000000000039000000000000003300000000",
            INIT_6B => X"0000003d00000000000000440000000000000044000000000000004400000000",
            INIT_6C => X"0000003f000000000000005d0000000000000042000000000000003200000000",
            INIT_6D => X"0000002f00000000000000300000000000000038000000000000003100000000",
            INIT_6E => X"000000330000000000000031000000000000002f000000000000002f00000000",
            INIT_6F => X"00000005000000000000000e000000000000002e000000000000003400000000",
            INIT_70 => X"0000002d0000000000000029000000000000002b000000000000002700000000",
            INIT_71 => X"0000003b00000000000000380000000000000036000000000000003200000000",
            INIT_72 => X"0000004000000000000000420000000000000040000000000000003e00000000",
            INIT_73 => X"00000031000000000000003a000000000000003d000000000000004000000000",
            INIT_74 => X"0000003b00000000000000550000000000000035000000000000002400000000",
            INIT_75 => X"0000002f000000000000002f0000000000000030000000000000003200000000",
            INIT_76 => X"00000032000000000000002d000000000000002e000000000000002e00000000",
            INIT_77 => X"0000000300000000000000030000000000000018000000000000003600000000",
            INIT_78 => X"0000003600000000000000340000000000000032000000000000002f00000000",
            INIT_79 => X"0000003a00000000000000380000000000000038000000000000003800000000",
            INIT_7A => X"0000003200000000000000350000000000000037000000000000003a00000000",
            INIT_7B => X"00000014000000000000001e0000000000000027000000000000002d00000000",
            INIT_7C => X"0000003600000000000000480000000000000021000000000000000b00000000",
            INIT_7D => X"0000002e000000000000002d000000000000002d000000000000002c00000000",
            INIT_7E => X"00000034000000000000002b000000000000002c000000000000002c00000000",
            INIT_7F => X"0000000700000000000000030000000000000008000000000000002500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE17;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE18 : if BRAM_NAME = "sampleifmap_layersamples_instance18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000be00000000000000b000000000000000a7000000000000009b00000000",
            INIT_01 => X"000000a600000000000000a800000000000000a600000000000000b100000000",
            INIT_02 => X"000000bb00000000000000bb00000000000000b300000000000000aa00000000",
            INIT_03 => X"000000b800000000000000b800000000000000bb00000000000000bb00000000",
            INIT_04 => X"000000ba00000000000000b800000000000000b400000000000000b600000000",
            INIT_05 => X"000000bd00000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_06 => X"000000c300000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_07 => X"000000c000000000000000ca00000000000000c900000000000000c900000000",
            INIT_08 => X"000000bb00000000000000ab00000000000000a3000000000000009900000000",
            INIT_09 => X"0000009f000000000000009a000000000000009b00000000000000b300000000",
            INIT_0A => X"000000af00000000000000ab00000000000000a5000000000000009f00000000",
            INIT_0B => X"000000a500000000000000a200000000000000ab00000000000000a900000000",
            INIT_0C => X"000000a500000000000000a600000000000000a400000000000000aa00000000",
            INIT_0D => X"000000a800000000000000a900000000000000ad00000000000000a700000000",
            INIT_0E => X"000000ca00000000000000be00000000000000ad00000000000000a900000000",
            INIT_0F => X"000000bd00000000000000cb00000000000000ca00000000000000cc00000000",
            INIT_10 => X"000000b800000000000000a800000000000000a0000000000000009b00000000",
            INIT_11 => X"000000bc00000000000000b000000000000000ae00000000000000bb00000000",
            INIT_12 => X"000000be00000000000000b100000000000000b300000000000000b600000000",
            INIT_13 => X"000000b900000000000000bc00000000000000c200000000000000c000000000",
            INIT_14 => X"000000c200000000000000c100000000000000c200000000000000c100000000",
            INIT_15 => X"000000bf00000000000000c100000000000000c500000000000000c300000000",
            INIT_16 => X"000000cf00000000000000ce00000000000000c500000000000000bf00000000",
            INIT_17 => X"000000bd00000000000000cc00000000000000ce00000000000000d000000000",
            INIT_18 => X"000000b100000000000000a6000000000000009d000000000000009700000000",
            INIT_19 => X"000000c500000000000000c700000000000000b900000000000000b400000000",
            INIT_1A => X"000000c600000000000000cd00000000000000cc00000000000000b600000000",
            INIT_1B => X"000000cb00000000000000c400000000000000c500000000000000d200000000",
            INIT_1C => X"000000cb00000000000000d200000000000000cf00000000000000cd00000000",
            INIT_1D => X"000000cc00000000000000c500000000000000d200000000000000cf00000000",
            INIT_1E => X"000000c900000000000000cc00000000000000c600000000000000d000000000",
            INIT_1F => X"000000c000000000000000ce00000000000000cf00000000000000d100000000",
            INIT_20 => X"000000ae00000000000000a8000000000000009e000000000000009700000000",
            INIT_21 => X"000000c400000000000000bf00000000000000b500000000000000b100000000",
            INIT_22 => X"000000b900000000000000bd00000000000000c200000000000000b700000000",
            INIT_23 => X"000000ca00000000000000b900000000000000b900000000000000c400000000",
            INIT_24 => X"000000c000000000000000c800000000000000c700000000000000c700000000",
            INIT_25 => X"000000bc00000000000000be00000000000000c700000000000000c300000000",
            INIT_26 => X"000000c400000000000000c900000000000000c700000000000000c900000000",
            INIT_27 => X"000000c400000000000000cf00000000000000cc00000000000000ce00000000",
            INIT_28 => X"000000ae00000000000000a7000000000000009c000000000000009400000000",
            INIT_29 => X"000000c300000000000000c400000000000000ae00000000000000ab00000000",
            INIT_2A => X"000000b800000000000000bd00000000000000be00000000000000c000000000",
            INIT_2B => X"000000bf00000000000000bd00000000000000bd00000000000000bb00000000",
            INIT_2C => X"000000c600000000000000bb00000000000000c300000000000000be00000000",
            INIT_2D => X"000000c100000000000000c000000000000000bc00000000000000c000000000",
            INIT_2E => X"000000d100000000000000cb00000000000000ce00000000000000cd00000000",
            INIT_2F => X"000000c400000000000000d100000000000000d000000000000000d400000000",
            INIT_30 => X"000000ae00000000000000a50000000000000099000000000000009400000000",
            INIT_31 => X"000000c300000000000000cb00000000000000b000000000000000a800000000",
            INIT_32 => X"000000be00000000000000bb00000000000000bc00000000000000bc00000000",
            INIT_33 => X"000000c300000000000000c500000000000000c200000000000000b600000000",
            INIT_34 => X"000000cd00000000000000c800000000000000c100000000000000c400000000",
            INIT_35 => X"000000c900000000000000c500000000000000c500000000000000c600000000",
            INIT_36 => X"000000c300000000000000c600000000000000c800000000000000c500000000",
            INIT_37 => X"000000c300000000000000cf00000000000000cb00000000000000c500000000",
            INIT_38 => X"000000ac00000000000000a3000000000000009b000000000000009900000000",
            INIT_39 => X"000000d100000000000000c700000000000000bc00000000000000ac00000000",
            INIT_3A => X"000000bf00000000000000bd00000000000000be00000000000000c400000000",
            INIT_3B => X"000000c400000000000000bb00000000000000bc00000000000000c100000000",
            INIT_3C => X"000000ce00000000000000c400000000000000c200000000000000ca00000000",
            INIT_3D => X"000000c800000000000000c400000000000000c900000000000000c200000000",
            INIT_3E => X"000000c900000000000000c800000000000000bb00000000000000b500000000",
            INIT_3F => X"000000bd00000000000000c700000000000000c400000000000000c800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ac00000000000000a3000000000000009f00000000000000a000000000",
            INIT_41 => X"000000be00000000000000b000000000000000b000000000000000ae00000000",
            INIT_42 => X"000000b000000000000000b000000000000000af00000000000000b400000000",
            INIT_43 => X"000000b600000000000000ac00000000000000aa00000000000000b500000000",
            INIT_44 => X"000000bb00000000000000b500000000000000b200000000000000bb00000000",
            INIT_45 => X"000000bb00000000000000b400000000000000bc00000000000000b100000000",
            INIT_46 => X"000000bc00000000000000bc00000000000000c400000000000000c700000000",
            INIT_47 => X"000000b800000000000000c200000000000000c000000000000000c500000000",
            INIT_48 => X"000000ac00000000000000a200000000000000a700000000000000ab00000000",
            INIT_49 => X"000000b000000000000000b400000000000000ab00000000000000aa00000000",
            INIT_4A => X"0000009c0000000000000096000000000000009c000000000000009b00000000",
            INIT_4B => X"0000009e00000000000000990000000000000092000000000000009600000000",
            INIT_4C => X"0000009d00000000000000a400000000000000a600000000000000a600000000",
            INIT_4D => X"000000a6000000000000009c00000000000000a2000000000000009d00000000",
            INIT_4E => X"000000bd00000000000000bc00000000000000c700000000000000c800000000",
            INIT_4F => X"000000b600000000000000c200000000000000c100000000000000c500000000",
            INIT_50 => X"000000b000000000000000a800000000000000b400000000000000af00000000",
            INIT_51 => X"000000ae00000000000000b600000000000000b100000000000000ad00000000",
            INIT_52 => X"0000009a000000000000009f00000000000000a0000000000000009c00000000",
            INIT_53 => X"000000ad00000000000000a800000000000000a3000000000000009f00000000",
            INIT_54 => X"000000a200000000000000a000000000000000a400000000000000aa00000000",
            INIT_55 => X"000000ac00000000000000a700000000000000a800000000000000a000000000",
            INIT_56 => X"000000c400000000000000c400000000000000c300000000000000c200000000",
            INIT_57 => X"000000b700000000000000c100000000000000bf00000000000000c500000000",
            INIT_58 => X"000000bb00000000000000b200000000000000bb00000000000000b500000000",
            INIT_59 => X"000000b600000000000000ae00000000000000aa00000000000000b700000000",
            INIT_5A => X"000000b500000000000000b400000000000000b300000000000000b300000000",
            INIT_5B => X"000000c100000000000000c100000000000000bb00000000000000b800000000",
            INIT_5C => X"000000b900000000000000bc00000000000000c000000000000000c100000000",
            INIT_5D => X"000000c000000000000000c000000000000000ba00000000000000b800000000",
            INIT_5E => X"000000bd00000000000000c000000000000000bc00000000000000bb00000000",
            INIT_5F => X"000000ba00000000000000c400000000000000bf00000000000000be00000000",
            INIT_60 => X"000000ab00000000000000ba00000000000000be00000000000000b900000000",
            INIT_61 => X"000000c100000000000000950000000000000084000000000000009900000000",
            INIT_62 => X"000000bc00000000000000ba00000000000000bf00000000000000c600000000",
            INIT_63 => X"000000c400000000000000c300000000000000c100000000000000bf00000000",
            INIT_64 => X"000000bc00000000000000be00000000000000c000000000000000c300000000",
            INIT_65 => X"000000bf00000000000000c000000000000000be00000000000000bc00000000",
            INIT_66 => X"000000c500000000000000c300000000000000c100000000000000bf00000000",
            INIT_67 => X"000000c100000000000000cc00000000000000ca00000000000000ca00000000",
            INIT_68 => X"0000009e00000000000000bc00000000000000c200000000000000ba00000000",
            INIT_69 => X"0000006d000000000000005e0000000000000074000000000000008400000000",
            INIT_6A => X"000000c200000000000000c200000000000000b1000000000000009100000000",
            INIT_6B => X"000000c700000000000000c400000000000000c100000000000000bf00000000",
            INIT_6C => X"000000c600000000000000c800000000000000c700000000000000c700000000",
            INIT_6D => X"000000c600000000000000c700000000000000c400000000000000c400000000",
            INIT_6E => X"000000c400000000000000c400000000000000c400000000000000c500000000",
            INIT_6F => X"000000b900000000000000c600000000000000c500000000000000c600000000",
            INIT_70 => X"000000c600000000000000c400000000000000c500000000000000ba00000000",
            INIT_71 => X"0000005c000000000000008d00000000000000b800000000000000c200000000",
            INIT_72 => X"000000b3000000000000008e0000000000000068000000000000005400000000",
            INIT_73 => X"000000cc00000000000000cc00000000000000c900000000000000c300000000",
            INIT_74 => X"000000c700000000000000cc00000000000000cc00000000000000cc00000000",
            INIT_75 => X"000000bf00000000000000c200000000000000c200000000000000c200000000",
            INIT_76 => X"000000be00000000000000be00000000000000be00000000000000bd00000000",
            INIT_77 => X"000000b500000000000000c000000000000000be00000000000000bf00000000",
            INIT_78 => X"000000c800000000000000c600000000000000c700000000000000b800000000",
            INIT_79 => X"000000b100000000000000c900000000000000c800000000000000c500000000",
            INIT_7A => X"00000080000000000000005d0000000000000054000000000000007500000000",
            INIT_7B => X"000000cd00000000000000d000000000000000ca00000000000000ad00000000",
            INIT_7C => X"000000c700000000000000c700000000000000c800000000000000ca00000000",
            INIT_7D => X"000000c300000000000000c500000000000000c400000000000000c300000000",
            INIT_7E => X"000000bf00000000000000c200000000000000c300000000000000c100000000",
            INIT_7F => X"000000b200000000000000be00000000000000bd00000000000000bf00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE18;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE19 : if BRAM_NAME = "sampleifmap_layersamples_instance19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d000000000000000cb00000000000000c900000000000000b900000000",
            INIT_01 => X"000000d600000000000000d000000000000000ce00000000000000cd00000000",
            INIT_02 => X"0000005b000000000000004c000000000000005c00000000000000af00000000",
            INIT_03 => X"000000cb00000000000000b5000000000000008c000000000000006900000000",
            INIT_04 => X"000000c200000000000000c500000000000000ca00000000000000ce00000000",
            INIT_05 => X"000000c200000000000000c200000000000000c200000000000000c100000000",
            INIT_06 => X"000000bf00000000000000c100000000000000c300000000000000c200000000",
            INIT_07 => X"000000b400000000000000be00000000000000be00000000000000c100000000",
            INIT_08 => X"000000d600000000000000cf00000000000000cc00000000000000bb00000000",
            INIT_09 => X"000000d000000000000000d300000000000000d400000000000000d400000000",
            INIT_0A => X"000000570000000000000047000000000000007c00000000000000cb00000000",
            INIT_0B => X"0000008400000000000000630000000000000054000000000000005400000000",
            INIT_0C => X"000000cb00000000000000cb00000000000000be00000000000000a700000000",
            INIT_0D => X"000000c400000000000000c500000000000000c000000000000000c300000000",
            INIT_0E => X"000000bf00000000000000c000000000000000c200000000000000c200000000",
            INIT_0F => X"000000b700000000000000c000000000000000bf00000000000000c100000000",
            INIT_10 => X"000000d600000000000000cf00000000000000cf00000000000000be00000000",
            INIT_11 => X"000000d000000000000000d300000000000000d300000000000000d400000000",
            INIT_12 => X"000000570000000000000048000000000000008900000000000000d300000000",
            INIT_13 => X"0000005300000000000000560000000000000054000000000000005300000000",
            INIT_14 => X"0000009b0000000000000083000000000000006b000000000000005900000000",
            INIT_15 => X"000000cc00000000000000cb00000000000000b600000000000000a300000000",
            INIT_16 => X"000000bf00000000000000c200000000000000c600000000000000ca00000000",
            INIT_17 => X"000000b600000000000000bf00000000000000c000000000000000c100000000",
            INIT_18 => X"000000d700000000000000d100000000000000d200000000000000bf00000000",
            INIT_19 => X"000000d500000000000000d400000000000000d400000000000000d500000000",
            INIT_1A => X"0000003a000000000000002f000000000000007100000000000000cc00000000",
            INIT_1B => X"0000005d0000000000000057000000000000004c000000000000003f00000000",
            INIT_1C => X"0000003e00000000000000460000000000000050000000000000005a00000000",
            INIT_1D => X"0000009f000000000000007a000000000000004d000000000000003a00000000",
            INIT_1E => X"000000c800000000000000c900000000000000c200000000000000b400000000",
            INIT_1F => X"000000b900000000000000c400000000000000c400000000000000c800000000",
            INIT_20 => X"000000d300000000000000cf00000000000000d000000000000000bf00000000",
            INIT_21 => X"000000d400000000000000d100000000000000d200000000000000d100000000",
            INIT_22 => X"0000002500000000000000410000000000000065000000000000009d00000000",
            INIT_23 => X"00000058000000000000004a0000000000000044000000000000003300000000",
            INIT_24 => X"0000004900000000000000550000000000000056000000000000005b00000000",
            INIT_25 => X"00000048000000000000003e000000000000002e000000000000003700000000",
            INIT_26 => X"0000009e0000000000000085000000000000006b000000000000004e00000000",
            INIT_27 => X"000000ba00000000000000c400000000000000c300000000000000b800000000",
            INIT_28 => X"000000d100000000000000cb00000000000000ca00000000000000ba00000000",
            INIT_29 => X"000000c800000000000000d100000000000000ce00000000000000cf00000000",
            INIT_2A => X"000000640000000000000097000000000000008c000000000000009500000000",
            INIT_2B => X"0000006000000000000000320000000000000035000000000000002d00000000",
            INIT_2C => X"00000048000000000000008000000000000000a0000000000000009c00000000",
            INIT_2D => X"0000004200000000000000590000000000000070000000000000006200000000",
            INIT_2E => X"000000a300000000000000a60000000000000083000000000000004300000000",
            INIT_2F => X"000000b200000000000000bc00000000000000b700000000000000ad00000000",
            INIT_30 => X"000000d200000000000000ca00000000000000c900000000000000b900000000",
            INIT_31 => X"000000d100000000000000d100000000000000d000000000000000d200000000",
            INIT_32 => X"000000bd00000000000000d700000000000000d300000000000000d200000000",
            INIT_33 => X"000000a800000000000000940000000000000092000000000000009000000000",
            INIT_34 => X"0000009a00000000000000c000000000000000ce00000000000000ca00000000",
            INIT_35 => X"0000009f00000000000000b100000000000000b200000000000000a300000000",
            INIT_36 => X"000000c200000000000000bf00000000000000b2000000000000009c00000000",
            INIT_37 => X"000000b000000000000000bc00000000000000c100000000000000c400000000",
            INIT_38 => X"000000c400000000000000c000000000000000bc00000000000000b000000000",
            INIT_39 => X"000000b700000000000000b900000000000000bc00000000000000c000000000",
            INIT_3A => X"000000ad00000000000000b300000000000000b200000000000000b600000000",
            INIT_3B => X"000000ad00000000000000ab00000000000000aa00000000000000aa00000000",
            INIT_3C => X"000000a700000000000000a100000000000000a000000000000000a900000000",
            INIT_3D => X"000000aa00000000000000a500000000000000a100000000000000a500000000",
            INIT_3E => X"00000096000000000000009800000000000000a000000000000000aa00000000",
            INIT_3F => X"0000009c00000000000000a400000000000000a3000000000000009d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006b000000000000006e0000000000000063000000000000007200000000",
            INIT_41 => X"0000005d000000000000005e0000000000000061000000000000006600000000",
            INIT_42 => X"0000005000000000000000580000000000000055000000000000005800000000",
            INIT_43 => X"000000650000000000000053000000000000004e000000000000004d00000000",
            INIT_44 => X"0000006b000000000000006a000000000000006c000000000000007100000000",
            INIT_45 => X"00000071000000000000006f000000000000006e000000000000006c00000000",
            INIT_46 => X"0000007700000000000000780000000000000077000000000000007500000000",
            INIT_47 => X"0000007c000000000000007a0000000000000079000000000000007800000000",
            INIT_48 => X"000000750000000000000071000000000000006d000000000000007a00000000",
            INIT_49 => X"0000007100000000000000720000000000000070000000000000007300000000",
            INIT_4A => X"0000006d000000000000006f0000000000000070000000000000006f00000000",
            INIT_4B => X"0000006c000000000000006e000000000000006d000000000000006e00000000",
            INIT_4C => X"0000006b00000000000000690000000000000070000000000000007300000000",
            INIT_4D => X"000000680000000000000065000000000000006a000000000000006c00000000",
            INIT_4E => X"0000006d000000000000006d000000000000006b000000000000006a00000000",
            INIT_4F => X"00000065000000000000005e0000000000000066000000000000006700000000",
            INIT_50 => X"00000070000000000000006b0000000000000061000000000000007800000000",
            INIT_51 => X"0000005e00000000000000620000000000000068000000000000006d00000000",
            INIT_52 => X"000000560000000000000058000000000000005d000000000000005e00000000",
            INIT_53 => X"0000004e0000000000000050000000000000004f000000000000005200000000",
            INIT_54 => X"000000450000000000000048000000000000004f000000000000005000000000",
            INIT_55 => X"0000004100000000000000410000000000000042000000000000004300000000",
            INIT_56 => X"0000004000000000000000420000000000000041000000000000004000000000",
            INIT_57 => X"0000004d0000000000000035000000000000003f000000000000004300000000",
            INIT_58 => X"0000004500000000000000410000000000000037000000000000005b00000000",
            INIT_59 => X"0000003d000000000000003f0000000000000042000000000000004200000000",
            INIT_5A => X"00000039000000000000003c0000000000000040000000000000004200000000",
            INIT_5B => X"0000003f000000000000003d000000000000003c000000000000003900000000",
            INIT_5C => X"0000003a00000000000000400000000000000042000000000000003f00000000",
            INIT_5D => X"0000003c000000000000003b0000000000000039000000000000003800000000",
            INIT_5E => X"0000003900000000000000380000000000000039000000000000003a00000000",
            INIT_5F => X"0000005c000000000000004b0000000000000031000000000000003400000000",
            INIT_60 => X"000000440000000000000042000000000000003c000000000000005d00000000",
            INIT_61 => X"0000004100000000000000400000000000000043000000000000004300000000",
            INIT_62 => X"0000003b000000000000003e0000000000000041000000000000004500000000",
            INIT_63 => X"0000003d000000000000003c000000000000003b000000000000003b00000000",
            INIT_64 => X"00000038000000000000003a000000000000003f000000000000004000000000",
            INIT_65 => X"0000003800000000000000380000000000000037000000000000003700000000",
            INIT_66 => X"000000350000000000000038000000000000003a000000000000003900000000",
            INIT_67 => X"000000510000000000000061000000000000005d000000000000004100000000",
            INIT_68 => X"00000039000000000000003d0000000000000039000000000000005900000000",
            INIT_69 => X"0000003b0000000000000039000000000000003b000000000000003900000000",
            INIT_6A => X"000000360000000000000038000000000000003a000000000000003c00000000",
            INIT_6B => X"0000003d000000000000003b000000000000003d000000000000003c00000000",
            INIT_6C => X"00000039000000000000003a000000000000003d000000000000004100000000",
            INIT_6D => X"0000003d000000000000003d000000000000003c000000000000003c00000000",
            INIT_6E => X"000000460000000000000039000000000000003e000000000000004200000000",
            INIT_6F => X"00000043000000000000003b0000000000000059000000000000006100000000",
            INIT_70 => X"0000003e000000000000003f000000000000003c000000000000005900000000",
            INIT_71 => X"0000003f000000000000003e000000000000003e000000000000003e00000000",
            INIT_72 => X"000000520000000000000041000000000000003d000000000000003e00000000",
            INIT_73 => X"00000051000000000000004e0000000000000051000000000000005400000000",
            INIT_74 => X"0000005300000000000000550000000000000054000000000000005800000000",
            INIT_75 => X"0000004000000000000000420000000000000043000000000000005000000000",
            INIT_76 => X"0000006700000000000000560000000000000038000000000000003400000000",
            INIT_77 => X"0000004b000000000000003d0000000000000039000000000000004c00000000",
            INIT_78 => X"0000003c000000000000003d000000000000003c000000000000005c00000000",
            INIT_79 => X"0000004100000000000000430000000000000042000000000000003f00000000",
            INIT_7A => X"0000004800000000000000410000000000000043000000000000004200000000",
            INIT_7B => X"0000004600000000000000480000000000000049000000000000004900000000",
            INIT_7C => X"0000004b000000000000004b000000000000004a000000000000004900000000",
            INIT_7D => X"0000003e00000000000000400000000000000040000000000000004b00000000",
            INIT_7E => X"0000004000000000000000580000000000000056000000000000004100000000",
            INIT_7F => X"000000490000000000000040000000000000003c000000000000003900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE19;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE20 : if BRAM_NAME = "sampleifmap_layersamples_instance20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000c000000000000000b300000000000000b0000000000000009c00000000",
            INIT_01 => X"000000ad00000000000000ad00000000000000ab00000000000000b900000000",
            INIT_02 => X"000000b800000000000000b600000000000000b300000000000000af00000000",
            INIT_03 => X"000000b500000000000000b600000000000000b800000000000000b900000000",
            INIT_04 => X"000000b900000000000000b700000000000000b300000000000000b300000000",
            INIT_05 => X"000000bd00000000000000bb00000000000000ba00000000000000ba00000000",
            INIT_06 => X"000000c300000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_07 => X"000000b700000000000000ca00000000000000c400000000000000c500000000",
            INIT_08 => X"000000c300000000000000b800000000000000b3000000000000009b00000000",
            INIT_09 => X"000000a4000000000000009f00000000000000a200000000000000be00000000",
            INIT_0A => X"000000b000000000000000a900000000000000a500000000000000a300000000",
            INIT_0B => X"000000a700000000000000a400000000000000ae00000000000000ab00000000",
            INIT_0C => X"000000a600000000000000a800000000000000a600000000000000ac00000000",
            INIT_0D => X"000000a900000000000000ab00000000000000af00000000000000a900000000",
            INIT_0E => X"000000cc00000000000000bf00000000000000ae00000000000000aa00000000",
            INIT_0F => X"000000be00000000000000d700000000000000d000000000000000ce00000000",
            INIT_10 => X"000000c400000000000000b900000000000000b2000000000000009a00000000",
            INIT_11 => X"000000a800000000000000b200000000000000c100000000000000cb00000000",
            INIT_12 => X"000000c400000000000000be00000000000000af00000000000000a000000000",
            INIT_13 => X"000000bc00000000000000be00000000000000c500000000000000c300000000",
            INIT_14 => X"000000c300000000000000c200000000000000c300000000000000c400000000",
            INIT_15 => X"000000bf00000000000000c100000000000000c600000000000000c400000000",
            INIT_16 => X"000000cd00000000000000cd00000000000000c400000000000000c000000000",
            INIT_17 => X"000000bf00000000000000d700000000000000d000000000000000ce00000000",
            INIT_18 => X"000000c300000000000000bc00000000000000b2000000000000009a00000000",
            INIT_19 => X"0000008000000000000000bc00000000000000c500000000000000ca00000000",
            INIT_1A => X"0000009b000000000000009a0000000000000098000000000000006c00000000",
            INIT_1B => X"0000009400000000000000950000000000000095000000000000009e00000000",
            INIT_1C => X"000000ad00000000000000a300000000000000a100000000000000a700000000",
            INIT_1D => X"0000009f00000000000000ae00000000000000a300000000000000a800000000",
            INIT_1E => X"000000ce00000000000000cc00000000000000d000000000000000bc00000000",
            INIT_1F => X"000000bc00000000000000d400000000000000cd00000000000000cc00000000",
            INIT_20 => X"000000bf00000000000000bb00000000000000b1000000000000009a00000000",
            INIT_21 => X"0000007e00000000000000bd00000000000000c400000000000000c600000000",
            INIT_22 => X"0000006b000000000000006a000000000000008b000000000000008000000000",
            INIT_23 => X"0000007100000000000000760000000000000078000000000000007300000000",
            INIT_24 => X"0000007e00000000000000720000000000000072000000000000007700000000",
            INIT_25 => X"0000007000000000000000880000000000000070000000000000007600000000",
            INIT_26 => X"000000ce00000000000000c900000000000000cb00000000000000a000000000",
            INIT_27 => X"000000be00000000000000d600000000000000cd00000000000000ce00000000",
            INIT_28 => X"000000bd00000000000000bb00000000000000ae000000000000009700000000",
            INIT_29 => X"0000009300000000000000b700000000000000c800000000000000c500000000",
            INIT_2A => X"000000a5000000000000009100000000000000a800000000000000a900000000",
            INIT_2B => X"0000009d0000000000000095000000000000009200000000000000aa00000000",
            INIT_2C => X"000000bd00000000000000b000000000000000b200000000000000b400000000",
            INIT_2D => X"000000b100000000000000bc00000000000000b300000000000000b000000000",
            INIT_2E => X"000000d000000000000000cf00000000000000d000000000000000c400000000",
            INIT_2F => X"000000be00000000000000d800000000000000d100000000000000d000000000",
            INIT_30 => X"000000bd00000000000000b900000000000000ac000000000000009800000000",
            INIT_31 => X"00000060000000000000009300000000000000c600000000000000c200000000",
            INIT_32 => X"0000009800000000000000900000000000000097000000000000009500000000",
            INIT_33 => X"0000008b00000000000000800000000000000079000000000000009800000000",
            INIT_34 => X"000000a200000000000000aa0000000000000097000000000000009c00000000",
            INIT_35 => X"000000a4000000000000009600000000000000ad000000000000009600000000",
            INIT_36 => X"000000d200000000000000cc00000000000000a6000000000000009c00000000",
            INIT_37 => X"000000bc00000000000000d400000000000000cf00000000000000d300000000",
            INIT_38 => X"000000bb00000000000000b600000000000000ac000000000000009b00000000",
            INIT_39 => X"00000065000000000000007700000000000000b500000000000000c200000000",
            INIT_3A => X"0000007800000000000000830000000000000083000000000000007b00000000",
            INIT_3B => X"0000007f00000000000000870000000000000087000000000000009200000000",
            INIT_3C => X"0000007b0000000000000083000000000000007b000000000000007b00000000",
            INIT_3D => X"0000009f000000000000007b0000000000000084000000000000006d00000000",
            INIT_3E => X"000000c700000000000000bf0000000000000084000000000000007b00000000",
            INIT_3F => X"000000ba00000000000000d000000000000000c900000000000000c900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b900000000000000b400000000000000af00000000000000a100000000",
            INIT_41 => X"000000af00000000000000ab00000000000000ba00000000000000c000000000",
            INIT_42 => X"000000a600000000000000ac00000000000000a500000000000000a200000000",
            INIT_43 => X"000000aa00000000000000ad00000000000000ac00000000000000af00000000",
            INIT_44 => X"000000af00000000000000b200000000000000b200000000000000ac00000000",
            INIT_45 => X"000000be00000000000000b200000000000000ac00000000000000a300000000",
            INIT_46 => X"000000cd00000000000000c800000000000000b000000000000000ac00000000",
            INIT_47 => X"000000b900000000000000d100000000000000c900000000000000c800000000",
            INIT_48 => X"000000ba00000000000000b400000000000000b700000000000000ac00000000",
            INIT_49 => X"000000b700000000000000c200000000000000c000000000000000be00000000",
            INIT_4A => X"000000a300000000000000a200000000000000a500000000000000a000000000",
            INIT_4B => X"000000a200000000000000a4000000000000009e000000000000009f00000000",
            INIT_4C => X"000000a200000000000000ac00000000000000ae00000000000000a700000000",
            INIT_4D => X"000000b600000000000000a500000000000000a300000000000000a000000000",
            INIT_4E => X"000000cd00000000000000ca00000000000000c600000000000000c800000000",
            INIT_4F => X"000000b800000000000000d000000000000000ca00000000000000ca00000000",
            INIT_50 => X"000000be00000000000000ba00000000000000c400000000000000b100000000",
            INIT_51 => X"000000b700000000000000c100000000000000c100000000000000c000000000",
            INIT_52 => X"0000009f00000000000000a500000000000000a700000000000000a300000000",
            INIT_53 => X"000000ac00000000000000aa00000000000000a600000000000000a400000000",
            INIT_54 => X"000000ab00000000000000a600000000000000a600000000000000a800000000",
            INIT_55 => X"000000b200000000000000ab00000000000000ad00000000000000a800000000",
            INIT_56 => X"000000c700000000000000c700000000000000c600000000000000c700000000",
            INIT_57 => X"000000b800000000000000d000000000000000c800000000000000c800000000",
            INIT_58 => X"000000c800000000000000c300000000000000cc00000000000000b700000000",
            INIT_59 => X"000000c600000000000000be00000000000000bb00000000000000c900000000",
            INIT_5A => X"000000c100000000000000c100000000000000c100000000000000c200000000",
            INIT_5B => X"000000c600000000000000c600000000000000c200000000000000c100000000",
            INIT_5C => X"000000c600000000000000c300000000000000c300000000000000c600000000",
            INIT_5D => X"000000c500000000000000c400000000000000c400000000000000c500000000",
            INIT_5E => X"000000c900000000000000c900000000000000cb00000000000000c900000000",
            INIT_5F => X"000000bb00000000000000d100000000000000c800000000000000ca00000000",
            INIT_60 => X"000000b200000000000000c600000000000000cd00000000000000b900000000",
            INIT_61 => X"000000c4000000000000009a000000000000008d00000000000000a600000000",
            INIT_62 => X"000000c500000000000000c700000000000000ca00000000000000ca00000000",
            INIT_63 => X"000000ca00000000000000c900000000000000c700000000000000c500000000",
            INIT_64 => X"000000c400000000000000c600000000000000c700000000000000c900000000",
            INIT_65 => X"000000c600000000000000c700000000000000c600000000000000c400000000",
            INIT_66 => X"000000ce00000000000000cb00000000000000ca00000000000000c700000000",
            INIT_67 => X"000000bd00000000000000d400000000000000ce00000000000000cf00000000",
            INIT_68 => X"000000a500000000000000c800000000000000d000000000000000ba00000000",
            INIT_69 => X"0000006b000000000000005f000000000000007c000000000000009000000000",
            INIT_6A => X"000000c700000000000000c700000000000000b3000000000000008f00000000",
            INIT_6B => X"000000cc00000000000000c900000000000000c600000000000000c500000000",
            INIT_6C => X"000000cc00000000000000ce00000000000000cd00000000000000cc00000000",
            INIT_6D => X"000000cd00000000000000cd00000000000000c900000000000000c900000000",
            INIT_6E => X"000000cb00000000000000cb00000000000000cb00000000000000cc00000000",
            INIT_6F => X"000000b700000000000000cf00000000000000ca00000000000000ca00000000",
            INIT_70 => X"000000cc00000000000000d000000000000000d400000000000000ba00000000",
            INIT_71 => X"0000005b000000000000008f00000000000000c100000000000000ce00000000",
            INIT_72 => X"000000b5000000000000008e0000000000000065000000000000005100000000",
            INIT_73 => X"000000cf00000000000000cf00000000000000cc00000000000000c600000000",
            INIT_74 => X"000000ca00000000000000cf00000000000000cf00000000000000cf00000000",
            INIT_75 => X"000000c500000000000000c600000000000000c500000000000000c500000000",
            INIT_76 => X"000000c500000000000000c500000000000000c500000000000000c500000000",
            INIT_77 => X"000000b500000000000000cc00000000000000c500000000000000c400000000",
            INIT_78 => X"000000ce00000000000000d200000000000000d600000000000000b800000000",
            INIT_79 => X"000000b300000000000000cf00000000000000d400000000000000d100000000",
            INIT_7A => X"00000080000000000000005d0000000000000053000000000000007400000000",
            INIT_7B => X"000000ce00000000000000d200000000000000cb00000000000000ae00000000",
            INIT_7C => X"000000c900000000000000ca00000000000000ca00000000000000cc00000000",
            INIT_7D => X"000000c900000000000000c900000000000000c700000000000000c600000000",
            INIT_7E => X"000000c700000000000000c900000000000000ca00000000000000c800000000",
            INIT_7F => X"000000b400000000000000cb00000000000000c600000000000000c600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE20;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE21 : if BRAM_NAME = "sampleifmap_layersamples_instance21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d500000000000000d600000000000000d700000000000000ba00000000",
            INIT_01 => X"000000d900000000000000d400000000000000d600000000000000d600000000",
            INIT_02 => X"000000560000000000000049000000000000005b00000000000000af00000000",
            INIT_03 => X"000000cc00000000000000b5000000000000008a000000000000006500000000",
            INIT_04 => X"000000c600000000000000c700000000000000cb00000000000000d000000000",
            INIT_05 => X"000000c800000000000000c900000000000000c900000000000000c700000000",
            INIT_06 => X"000000c900000000000000c900000000000000ca00000000000000c800000000",
            INIT_07 => X"000000b600000000000000cc00000000000000c800000000000000ca00000000",
            INIT_08 => X"000000d900000000000000d800000000000000d800000000000000bb00000000",
            INIT_09 => X"000000d300000000000000d600000000000000d900000000000000db00000000",
            INIT_0A => X"000000520000000000000044000000000000007b00000000000000cc00000000",
            INIT_0B => X"0000008200000000000000610000000000000051000000000000004f00000000",
            INIT_0C => X"000000ca00000000000000c900000000000000bc00000000000000a500000000",
            INIT_0D => X"000000c600000000000000c700000000000000c100000000000000c400000000",
            INIT_0E => X"000000c800000000000000c800000000000000c700000000000000c600000000",
            INIT_0F => X"000000b600000000000000cc00000000000000c700000000000000c900000000",
            INIT_10 => X"000000d600000000000000d500000000000000d900000000000000bc00000000",
            INIT_11 => X"000000d200000000000000d600000000000000d800000000000000d800000000",
            INIT_12 => X"000000530000000000000046000000000000008800000000000000d400000000",
            INIT_13 => X"0000004d00000000000000500000000000000050000000000000004e00000000",
            INIT_14 => X"00000097000000000000007e0000000000000066000000000000005300000000",
            INIT_15 => X"000000cc00000000000000c900000000000000b2000000000000009f00000000",
            INIT_16 => X"000000c600000000000000c800000000000000c900000000000000cb00000000",
            INIT_17 => X"000000b400000000000000c900000000000000c500000000000000c700000000",
            INIT_18 => X"000000d500000000000000d600000000000000da00000000000000bb00000000",
            INIT_19 => X"000000d800000000000000d700000000000000d800000000000000d700000000",
            INIT_1A => X"00000037000000000000002d000000000000007000000000000000cc00000000",
            INIT_1B => X"00000051000000000000004d0000000000000045000000000000003a00000000",
            INIT_1C => X"0000003e0000000000000046000000000000004d000000000000005000000000",
            INIT_1D => X"000000a0000000000000007c000000000000004f000000000000003b00000000",
            INIT_1E => X"000000cd00000000000000cd00000000000000c400000000000000b500000000",
            INIT_1F => X"000000b400000000000000ca00000000000000c800000000000000cb00000000",
            INIT_20 => X"000000d100000000000000d200000000000000d800000000000000bc00000000",
            INIT_21 => X"000000d400000000000000d400000000000000d600000000000000d300000000",
            INIT_22 => X"00000021000000000000003a000000000000005f000000000000009a00000000",
            INIT_23 => X"0000004d0000000000000041000000000000003e000000000000003000000000",
            INIT_24 => X"0000004800000000000000540000000000000054000000000000005200000000",
            INIT_25 => X"00000048000000000000003f000000000000002f000000000000003800000000",
            INIT_26 => X"0000009e0000000000000084000000000000006b000000000000004e00000000",
            INIT_27 => X"000000b600000000000000ca00000000000000c100000000000000b500000000",
            INIT_28 => X"000000cf00000000000000ce00000000000000d200000000000000b800000000",
            INIT_29 => X"000000c800000000000000d400000000000000d300000000000000d100000000",
            INIT_2A => X"00000061000000000000008f0000000000000085000000000000009100000000",
            INIT_2B => X"0000005a000000000000002e0000000000000032000000000000002d00000000",
            INIT_2C => X"00000047000000000000007f000000000000009e000000000000009600000000",
            INIT_2D => X"0000004100000000000000580000000000000070000000000000006100000000",
            INIT_2E => X"000000a200000000000000a50000000000000082000000000000004300000000",
            INIT_2F => X"000000b000000000000000c500000000000000b500000000000000a800000000",
            INIT_30 => X"000000d000000000000000cd00000000000000d200000000000000b700000000",
            INIT_31 => X"000000d200000000000000d500000000000000d400000000000000d300000000",
            INIT_32 => X"000000bf00000000000000d400000000000000d100000000000000d100000000",
            INIT_33 => X"000000a600000000000000930000000000000093000000000000009400000000",
            INIT_34 => X"0000009d00000000000000c300000000000000d000000000000000c800000000",
            INIT_35 => X"000000a200000000000000b400000000000000b500000000000000a600000000",
            INIT_36 => X"000000c500000000000000c100000000000000b4000000000000009f00000000",
            INIT_37 => X"000000b100000000000000c700000000000000c100000000000000c300000000",
            INIT_38 => X"000000c200000000000000c300000000000000c400000000000000ae00000000",
            INIT_39 => X"000000b900000000000000bb00000000000000be00000000000000c200000000",
            INIT_3A => X"000000b500000000000000b700000000000000b500000000000000b800000000",
            INIT_3B => X"000000ad00000000000000ae00000000000000b000000000000000b200000000",
            INIT_3C => X"000000ac00000000000000a600000000000000a400000000000000aa00000000",
            INIT_3D => X"000000b000000000000000aa00000000000000a600000000000000aa00000000",
            INIT_3E => X"0000009b000000000000009d00000000000000a500000000000000af00000000",
            INIT_3F => X"0000009e00000000000000af00000000000000a3000000000000009d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000690000000000000070000000000000006c000000000000007000000000",
            INIT_41 => X"0000006000000000000000610000000000000064000000000000006700000000",
            INIT_42 => X"00000057000000000000005e000000000000005a000000000000005c00000000",
            INIT_43 => X"0000006700000000000000570000000000000053000000000000005400000000",
            INIT_44 => X"00000070000000000000006f0000000000000070000000000000007300000000",
            INIT_45 => X"0000007600000000000000740000000000000073000000000000007100000000",
            INIT_46 => X"0000007b000000000000007c000000000000007b000000000000007a00000000",
            INIT_47 => X"0000007c0000000000000084000000000000007a000000000000007900000000",
            INIT_48 => X"0000007000000000000000710000000000000073000000000000007500000000",
            INIT_49 => X"000000710000000000000071000000000000006f000000000000007100000000",
            INIT_4A => X"0000006e000000000000006f0000000000000070000000000000006f00000000",
            INIT_4B => X"0000006b000000000000006e000000000000006d000000000000006e00000000",
            INIT_4C => X"0000006e000000000000006c0000000000000073000000000000007300000000",
            INIT_4D => X"0000006b0000000000000068000000000000006d000000000000006f00000000",
            INIT_4E => X"000000700000000000000070000000000000006e000000000000006d00000000",
            INIT_4F => X"000000650000000000000062000000000000005f000000000000006400000000",
            INIT_50 => X"0000006a00000000000000690000000000000066000000000000007100000000",
            INIT_51 => X"0000005d00000000000000610000000000000066000000000000006a00000000",
            INIT_52 => X"000000550000000000000059000000000000005e000000000000005f00000000",
            INIT_53 => X"0000004e000000000000004f000000000000004e000000000000005200000000",
            INIT_54 => X"000000440000000000000047000000000000004f000000000000005000000000",
            INIT_55 => X"0000004100000000000000410000000000000041000000000000004300000000",
            INIT_56 => X"0000004100000000000000420000000000000042000000000000004100000000",
            INIT_57 => X"0000006400000000000000470000000000000037000000000000003c00000000",
            INIT_58 => X"000000400000000000000041000000000000003c000000000000005400000000",
            INIT_59 => X"0000003c000000000000003e0000000000000040000000000000004000000000",
            INIT_5A => X"00000038000000000000003d0000000000000040000000000000004200000000",
            INIT_5B => X"0000003f000000000000003d000000000000003c000000000000003900000000",
            INIT_5C => X"0000003b00000000000000410000000000000043000000000000004000000000",
            INIT_5D => X"0000003c000000000000003b000000000000003a000000000000003800000000",
            INIT_5E => X"0000003800000000000000380000000000000039000000000000003a00000000",
            INIT_5F => X"0000008000000000000000750000000000000048000000000000003800000000",
            INIT_60 => X"0000003e000000000000003f000000000000003b000000000000005300000000",
            INIT_61 => X"0000003f000000000000003d0000000000000041000000000000003f00000000",
            INIT_62 => X"00000039000000000000003c000000000000003e000000000000004300000000",
            INIT_63 => X"0000003d000000000000003c000000000000003a000000000000003a00000000",
            INIT_64 => X"0000003e00000000000000400000000000000044000000000000004100000000",
            INIT_65 => X"0000003d000000000000003e000000000000003c000000000000003d00000000",
            INIT_66 => X"00000041000000000000003d000000000000003a000000000000003a00000000",
            INIT_67 => X"0000006300000000000000890000000000000088000000000000005b00000000",
            INIT_68 => X"00000039000000000000003d0000000000000035000000000000004f00000000",
            INIT_69 => X"0000003c000000000000003a000000000000003b000000000000003700000000",
            INIT_6A => X"000000370000000000000039000000000000003c000000000000003d00000000",
            INIT_6B => X"0000003f000000000000003d000000000000003e000000000000003c00000000",
            INIT_6C => X"0000003b000000000000003c000000000000003f000000000000004300000000",
            INIT_6D => X"0000003f0000000000000040000000000000003e000000000000003e00000000",
            INIT_6E => X"0000006e0000000000000047000000000000003c000000000000003e00000000",
            INIT_6F => X"0000004a000000000000004f0000000000000077000000000000008e00000000",
            INIT_70 => X"000000410000000000000042000000000000003a000000000000005200000000",
            INIT_71 => X"0000003e000000000000003e000000000000003e000000000000003f00000000",
            INIT_72 => X"0000004f0000000000000041000000000000003e000000000000003f00000000",
            INIT_73 => X"0000004d000000000000004a000000000000004c000000000000004f00000000",
            INIT_74 => X"0000004e00000000000000500000000000000050000000000000005400000000",
            INIT_75 => X"00000041000000000000003e000000000000003f000000000000004c00000000",
            INIT_76 => X"0000008d000000000000007c0000000000000056000000000000004200000000",
            INIT_77 => X"0000004500000000000000400000000000000042000000000000006600000000",
            INIT_78 => X"0000003a000000000000003a0000000000000034000000000000004e00000000",
            INIT_79 => X"00000039000000000000003b000000000000003a000000000000003a00000000",
            INIT_7A => X"00000045000000000000003a000000000000003b000000000000003a00000000",
            INIT_7B => X"0000004500000000000000460000000000000047000000000000004700000000",
            INIT_7C => X"0000004a00000000000000490000000000000048000000000000004800000000",
            INIT_7D => X"00000044000000000000003f000000000000003f000000000000004900000000",
            INIT_7E => X"0000005800000000000000800000000000000080000000000000005a00000000",
            INIT_7F => X"000000440000000000000041000000000000003f000000000000004200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE21;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE22 : if BRAM_NAME = "sampleifmap_layersamples_instance22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000cd00000000000000c100000000000000bb000000000000009500000000",
            INIT_01 => X"000000b400000000000000b500000000000000b700000000000000ca00000000",
            INIT_02 => X"000000c000000000000000c100000000000000bd00000000000000b600000000",
            INIT_03 => X"000000bd00000000000000bd00000000000000c000000000000000c000000000",
            INIT_04 => X"000000c000000000000000bd00000000000000b900000000000000ba00000000",
            INIT_05 => X"000000be00000000000000c000000000000000c100000000000000c100000000",
            INIT_06 => X"000000c300000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_07 => X"000000ab00000000000000d400000000000000d100000000000000ca00000000",
            INIT_08 => X"000000e300000000000000d700000000000000cc000000000000009d00000000",
            INIT_09 => X"000000b300000000000000b300000000000000be00000000000000e000000000",
            INIT_0A => X"000000c300000000000000c300000000000000bb00000000000000b300000000",
            INIT_0B => X"000000b700000000000000b400000000000000be00000000000000bb00000000",
            INIT_0C => X"000000b700000000000000b800000000000000b700000000000000bc00000000",
            INIT_0D => X"000000bc00000000000000bc00000000000000bf00000000000000b900000000",
            INIT_0E => X"000000e000000000000000d300000000000000c200000000000000be00000000",
            INIT_0F => X"000000b700000000000000e300000000000000de00000000000000df00000000",
            INIT_10 => X"000000db00000000000000d500000000000000c9000000000000009900000000",
            INIT_11 => X"000000b800000000000000c400000000000000d500000000000000df00000000",
            INIT_12 => X"000000d400000000000000d300000000000000c300000000000000b100000000",
            INIT_13 => X"000000ca00000000000000cc00000000000000d200000000000000d000000000",
            INIT_14 => X"000000d100000000000000d000000000000000d100000000000000d100000000",
            INIT_15 => X"000000d000000000000000d000000000000000d400000000000000d200000000",
            INIT_16 => X"000000df00000000000000de00000000000000d500000000000000d000000000",
            INIT_17 => X"000000b800000000000000e000000000000000d700000000000000da00000000",
            INIT_18 => X"000000de00000000000000d300000000000000cf00000000000000a600000000",
            INIT_19 => X"0000008300000000000000c900000000000000dc00000000000000e200000000",
            INIT_1A => X"000000b100000000000000a6000000000000009e000000000000007700000000",
            INIT_1B => X"000000ab00000000000000a600000000000000a700000000000000b200000000",
            INIT_1C => X"000000ba00000000000000b200000000000000b200000000000000b700000000",
            INIT_1D => X"000000a500000000000000b400000000000000ba00000000000000b900000000",
            INIT_1E => X"000000dd00000000000000dc00000000000000e400000000000000cf00000000",
            INIT_1F => X"000000ba00000000000000e600000000000000df00000000000000e000000000",
            INIT_20 => X"000000da00000000000000ca00000000000000cb00000000000000a700000000",
            INIT_21 => X"0000008e00000000000000d600000000000000e100000000000000e000000000",
            INIT_22 => X"0000008100000000000000780000000000000098000000000000009900000000",
            INIT_23 => X"00000083000000000000007c000000000000007e000000000000008100000000",
            INIT_24 => X"0000008a00000000000000820000000000000084000000000000008600000000",
            INIT_25 => X"0000007b000000000000008d0000000000000088000000000000008800000000",
            INIT_26 => X"000000d900000000000000da00000000000000e300000000000000ba00000000",
            INIT_27 => X"000000b900000000000000e300000000000000dc00000000000000de00000000",
            INIT_28 => X"000000d900000000000000cb00000000000000c900000000000000a400000000",
            INIT_29 => X"000000a500000000000000d100000000000000da00000000000000dc00000000",
            INIT_2A => X"000000b4000000000000009c00000000000000b500000000000000c400000000",
            INIT_2B => X"000000ac00000000000000a300000000000000a000000000000000b300000000",
            INIT_2C => X"000000c900000000000000be00000000000000c100000000000000bf00000000",
            INIT_2D => X"000000be00000000000000c600000000000000c000000000000000bf00000000",
            INIT_2E => X"000000e100000000000000e100000000000000e100000000000000d400000000",
            INIT_2F => X"000000bc00000000000000e800000000000000e100000000000000df00000000",
            INIT_30 => X"000000d900000000000000c800000000000000c600000000000000a400000000",
            INIT_31 => X"0000006800000000000000ac00000000000000d600000000000000d900000000",
            INIT_32 => X"000000af00000000000000a600000000000000a5000000000000009e00000000",
            INIT_33 => X"000000a00000000000000097000000000000009000000000000000a500000000",
            INIT_34 => X"000000b600000000000000bd00000000000000ad00000000000000b200000000",
            INIT_35 => X"000000b900000000000000ad00000000000000b700000000000000aa00000000",
            INIT_36 => X"000000e200000000000000dc00000000000000b200000000000000a600000000",
            INIT_37 => X"000000bc00000000000000e700000000000000e000000000000000dd00000000",
            INIT_38 => X"000000d800000000000000c700000000000000c900000000000000a900000000",
            INIT_39 => X"0000006f000000000000009200000000000000cb00000000000000da00000000",
            INIT_3A => X"00000090000000000000009d0000000000000095000000000000008600000000",
            INIT_3B => X"00000090000000000000008f000000000000008f000000000000009b00000000",
            INIT_3C => X"0000008e0000000000000094000000000000008e000000000000009300000000",
            INIT_3D => X"000000b0000000000000008e000000000000008d000000000000007f00000000",
            INIT_3E => X"000000dc00000000000000d10000000000000095000000000000008900000000",
            INIT_3F => X"000000ba00000000000000e400000000000000dc00000000000000d900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d900000000000000c700000000000000ce00000000000000b100000000",
            INIT_41 => X"000000c500000000000000c100000000000000cd00000000000000db00000000",
            INIT_42 => X"000000b800000000000000bb00000000000000b700000000000000b800000000",
            INIT_43 => X"000000bd00000000000000bb00000000000000ba00000000000000c000000000",
            INIT_44 => X"000000bf00000000000000c200000000000000c200000000000000c000000000",
            INIT_45 => X"000000c800000000000000bc00000000000000ba00000000000000b200000000",
            INIT_46 => X"000000db00000000000000d600000000000000c600000000000000c100000000",
            INIT_47 => X"000000b900000000000000e400000000000000dd00000000000000db00000000",
            INIT_48 => X"000000d600000000000000c500000000000000d400000000000000ba00000000",
            INIT_49 => X"000000d200000000000000dc00000000000000d600000000000000d700000000",
            INIT_4A => X"000000ba00000000000000b600000000000000bb00000000000000b900000000",
            INIT_4B => X"000000ba00000000000000b900000000000000b400000000000000b600000000",
            INIT_4C => X"000000b800000000000000c300000000000000c600000000000000c100000000",
            INIT_4D => X"000000c600000000000000b600000000000000b600000000000000b500000000",
            INIT_4E => X"000000df00000000000000dd00000000000000de00000000000000de00000000",
            INIT_4F => X"000000b700000000000000e300000000000000de00000000000000df00000000",
            INIT_50 => X"000000d800000000000000c800000000000000de00000000000000bc00000000",
            INIT_51 => X"000000cc00000000000000d600000000000000d400000000000000d700000000",
            INIT_52 => X"000000b000000000000000b600000000000000b800000000000000b500000000",
            INIT_53 => X"000000bf00000000000000bc00000000000000b800000000000000b500000000",
            INIT_54 => X"000000b900000000000000b800000000000000ba00000000000000bd00000000",
            INIT_55 => X"000000c900000000000000ba00000000000000b800000000000000b600000000",
            INIT_56 => X"000000db00000000000000dc00000000000000dd00000000000000df00000000",
            INIT_57 => X"000000b800000000000000e300000000000000dc00000000000000db00000000",
            INIT_58 => X"000000e000000000000000cf00000000000000e200000000000000bf00000000",
            INIT_59 => X"000000de00000000000000d700000000000000d100000000000000dc00000000",
            INIT_5A => X"000000d700000000000000d600000000000000d700000000000000d900000000",
            INIT_5B => X"000000df00000000000000df00000000000000db00000000000000d900000000",
            INIT_5C => X"000000da00000000000000db00000000000000dd00000000000000df00000000",
            INIT_5D => X"000000db00000000000000d900000000000000d600000000000000d800000000",
            INIT_5E => X"000000d600000000000000d900000000000000db00000000000000db00000000",
            INIT_5F => X"000000ba00000000000000e300000000000000db00000000000000d700000000",
            INIT_60 => X"000000ce00000000000000d400000000000000dc00000000000000bc00000000",
            INIT_61 => X"000000d900000000000000ac000000000000009900000000000000b500000000",
            INIT_62 => X"000000dc00000000000000dd00000000000000e100000000000000e200000000",
            INIT_63 => X"000000e200000000000000e100000000000000df00000000000000de00000000",
            INIT_64 => X"000000da00000000000000dc00000000000000dd00000000000000e100000000",
            INIT_65 => X"000000da00000000000000dc00000000000000db00000000000000d900000000",
            INIT_66 => X"000000e000000000000000de00000000000000dc00000000000000d900000000",
            INIT_67 => X"000000bb00000000000000e600000000000000e000000000000000e000000000",
            INIT_68 => X"000000c100000000000000d600000000000000df00000000000000bd00000000",
            INIT_69 => X"000000730000000000000063000000000000007e000000000000009d00000000",
            INIT_6A => X"000000dd00000000000000dd00000000000000c6000000000000009d00000000",
            INIT_6B => X"000000e200000000000000df00000000000000dc00000000000000da00000000",
            INIT_6C => X"000000df00000000000000e100000000000000e000000000000000e200000000",
            INIT_6D => X"000000e000000000000000e000000000000000dd00000000000000dc00000000",
            INIT_6E => X"000000de00000000000000de00000000000000de00000000000000df00000000",
            INIT_6F => X"000000b700000000000000e200000000000000dd00000000000000dd00000000",
            INIT_70 => X"000000e900000000000000de00000000000000e200000000000000bd00000000",
            INIT_71 => X"0000005a000000000000009200000000000000c400000000000000dc00000000",
            INIT_72 => X"000000ca00000000000000a10000000000000071000000000000005400000000",
            INIT_73 => X"000000e400000000000000e300000000000000e000000000000000da00000000",
            INIT_74 => X"000000dc00000000000000e000000000000000e100000000000000e200000000",
            INIT_75 => X"000000d900000000000000d800000000000000d700000000000000d700000000",
            INIT_76 => X"000000d800000000000000d800000000000000d800000000000000d800000000",
            INIT_77 => X"000000b600000000000000e100000000000000da00000000000000d700000000",
            INIT_78 => X"000000ea00000000000000e000000000000000e500000000000000bb00000000",
            INIT_79 => X"000000b300000000000000da00000000000000e100000000000000e100000000",
            INIT_7A => X"00000091000000000000006a0000000000000058000000000000007300000000",
            INIT_7B => X"000000e100000000000000e400000000000000dd00000000000000c000000000",
            INIT_7C => X"000000d900000000000000da00000000000000db00000000000000df00000000",
            INIT_7D => X"000000db00000000000000d900000000000000d600000000000000d600000000",
            INIT_7E => X"000000da00000000000000dc00000000000000dd00000000000000db00000000",
            INIT_7F => X"000000b700000000000000e200000000000000dc00000000000000d900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE22;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE23 : if BRAM_NAME = "sampleifmap_layersamples_instance23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e900000000000000de00000000000000e900000000000000be00000000",
            INIT_01 => X"000000e100000000000000e000000000000000e200000000000000e400000000",
            INIT_02 => X"0000005b0000000000000050000000000000006200000000000000b500000000",
            INIT_03 => X"000000d900000000000000c00000000000000092000000000000006a00000000",
            INIT_04 => X"000000da00000000000000dd00000000000000e100000000000000e000000000",
            INIT_05 => X"000000d900000000000000da00000000000000da00000000000000d900000000",
            INIT_06 => X"000000dd00000000000000dd00000000000000dd00000000000000da00000000",
            INIT_07 => X"000000bc00000000000000e300000000000000dc00000000000000dd00000000",
            INIT_08 => X"000000e900000000000000dd00000000000000ea00000000000000bf00000000",
            INIT_09 => X"000000dd00000000000000e200000000000000e300000000000000e700000000",
            INIT_0A => X"0000004f0000000000000049000000000000008200000000000000d500000000",
            INIT_0B => X"0000008800000000000000640000000000000050000000000000004b00000000",
            INIT_0C => X"000000dc00000000000000d700000000000000c800000000000000ad00000000",
            INIT_0D => X"000000de00000000000000df00000000000000d900000000000000d900000000",
            INIT_0E => X"000000db00000000000000db00000000000000dd00000000000000dd00000000",
            INIT_0F => X"000000bd00000000000000e300000000000000db00000000000000da00000000",
            INIT_10 => X"000000e400000000000000d900000000000000e800000000000000bd00000000",
            INIT_11 => X"000000dc00000000000000e200000000000000e100000000000000e300000000",
            INIT_12 => X"00000050000000000000004a000000000000009000000000000000dd00000000",
            INIT_13 => X"0000004c000000000000004e000000000000004c000000000000004a00000000",
            INIT_14 => X"000000a100000000000000810000000000000064000000000000005300000000",
            INIT_15 => X"000000e200000000000000e100000000000000c900000000000000b000000000",
            INIT_16 => X"000000d700000000000000d900000000000000dc00000000000000df00000000",
            INIT_17 => X"000000bb00000000000000e100000000000000d900000000000000d700000000",
            INIT_18 => X"000000e100000000000000d700000000000000e800000000000000bb00000000",
            INIT_19 => X"000000e200000000000000e300000000000000e100000000000000e000000000",
            INIT_1A => X"000000380000000000000032000000000000007700000000000000d500000000",
            INIT_1B => X"00000052000000000000004d0000000000000045000000000000003b00000000",
            INIT_1C => X"0000003f00000000000000420000000000000048000000000000005000000000",
            INIT_1D => X"000000a20000000000000085000000000000005b000000000000004100000000",
            INIT_1E => X"000000df00000000000000da00000000000000cc00000000000000b800000000",
            INIT_1F => X"000000bc00000000000000e300000000000000dd00000000000000dd00000000",
            INIT_20 => X"000000df00000000000000de00000000000000e700000000000000b700000000",
            INIT_21 => X"000000e100000000000000e400000000000000e600000000000000df00000000",
            INIT_22 => X"00000027000000000000003c000000000000006200000000000000a200000000",
            INIT_23 => X"0000004e00000000000000440000000000000043000000000000003500000000",
            INIT_24 => X"0000004800000000000000530000000000000052000000000000005100000000",
            INIT_25 => X"00000043000000000000003f0000000000000031000000000000003900000000",
            INIT_26 => X"000000a8000000000000008b000000000000006d000000000000004b00000000",
            INIT_27 => X"000000c300000000000000df00000000000000d700000000000000c600000000",
            INIT_28 => X"000000de00000000000000e200000000000000e200000000000000b000000000",
            INIT_29 => X"000000d400000000000000e200000000000000e200000000000000de00000000",
            INIT_2A => X"0000006a0000000000000096000000000000008b000000000000009b00000000",
            INIT_2B => X"0000005e00000000000000330000000000000039000000000000003500000000",
            INIT_2C => X"00000049000000000000008200000000000000a1000000000000009a00000000",
            INIT_2D => X"00000043000000000000005a0000000000000072000000000000006300000000",
            INIT_2E => X"000000a900000000000000ab0000000000000086000000000000004500000000",
            INIT_2F => X"000000be00000000000000d000000000000000c500000000000000b700000000",
            INIT_30 => X"000000df00000000000000e100000000000000e100000000000000af00000000",
            INIT_31 => X"000000de00000000000000de00000000000000de00000000000000df00000000",
            INIT_32 => X"000000cc00000000000000e400000000000000e000000000000000de00000000",
            INIT_33 => X"000000b300000000000000a0000000000000009f000000000000009f00000000",
            INIT_34 => X"000000a900000000000000cf00000000000000dc00000000000000d600000000",
            INIT_35 => X"000000ad00000000000000c000000000000000c100000000000000b200000000",
            INIT_36 => X"000000d600000000000000d200000000000000c300000000000000ab00000000",
            INIT_37 => X"000000bd00000000000000d200000000000000d100000000000000d800000000",
            INIT_38 => X"000000d100000000000000d700000000000000d400000000000000a600000000",
            INIT_39 => X"000000c700000000000000c900000000000000cc00000000000000ce00000000",
            INIT_3A => X"000000c200000000000000c500000000000000c300000000000000c700000000",
            INIT_3B => X"000000c400000000000000c200000000000000c100000000000000c000000000",
            INIT_3C => X"000000ca00000000000000c400000000000000c200000000000000c400000000",
            INIT_3D => X"000000cd00000000000000c800000000000000c400000000000000c800000000",
            INIT_3E => X"000000bf00000000000000c000000000000000c500000000000000ce00000000",
            INIT_3F => X"000000b500000000000000c900000000000000c500000000000000c500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007800000000000000820000000000000078000000000000006500000000",
            INIT_41 => X"0000006a000000000000006b0000000000000070000000000000007600000000",
            INIT_42 => X"0000006300000000000000660000000000000062000000000000006500000000",
            INIT_43 => X"00000080000000000000006c0000000000000065000000000000006200000000",
            INIT_44 => X"0000009300000000000000920000000000000092000000000000009000000000",
            INIT_45 => X"0000009e00000000000000980000000000000096000000000000009400000000",
            INIT_46 => X"000000a800000000000000a800000000000000a600000000000000a400000000",
            INIT_47 => X"0000009200000000000000a700000000000000a500000000000000a800000000",
            INIT_48 => X"0000008600000000000000860000000000000082000000000000006f00000000",
            INIT_49 => X"0000008800000000000000890000000000000088000000000000008a00000000",
            INIT_4A => X"0000007e00000000000000830000000000000086000000000000008400000000",
            INIT_4B => X"0000008300000000000000830000000000000080000000000000007f00000000",
            INIT_4C => X"00000081000000000000007f0000000000000086000000000000008a00000000",
            INIT_4D => X"0000007e000000000000007c0000000000000080000000000000008100000000",
            INIT_4E => X"0000008400000000000000840000000000000082000000000000008100000000",
            INIT_4F => X"0000006000000000000000730000000000000073000000000000007700000000",
            INIT_50 => X"0000007800000000000000780000000000000071000000000000006800000000",
            INIT_51 => X"00000064000000000000006c0000000000000076000000000000007a00000000",
            INIT_52 => X"000000590000000000000055000000000000005b000000000000006000000000",
            INIT_53 => X"0000005600000000000000570000000000000055000000000000005800000000",
            INIT_54 => X"000000430000000000000046000000000000004f000000000000005600000000",
            INIT_55 => X"0000003c000000000000003f0000000000000041000000000000004200000000",
            INIT_56 => X"0000003b000000000000003c000000000000003c000000000000003b00000000",
            INIT_57 => X"0000004b000000000000003f0000000000000032000000000000003600000000",
            INIT_58 => X"00000039000000000000003d0000000000000037000000000000003d00000000",
            INIT_59 => X"00000036000000000000003b000000000000003f000000000000003a00000000",
            INIT_5A => X"0000002f000000000000002f0000000000000033000000000000003800000000",
            INIT_5B => X"0000003200000000000000310000000000000032000000000000003000000000",
            INIT_5C => X"0000002f00000000000000350000000000000037000000000000003300000000",
            INIT_5D => X"000000370000000000000032000000000000002e000000000000002d00000000",
            INIT_5E => X"0000003400000000000000340000000000000034000000000000003600000000",
            INIT_5F => X"000000680000000000000068000000000000003a000000000000003000000000",
            INIT_60 => X"0000003c0000000000000041000000000000003d000000000000004400000000",
            INIT_61 => X"000000390000000000000037000000000000003d000000000000003e00000000",
            INIT_62 => X"0000003a00000000000000370000000000000038000000000000003d00000000",
            INIT_63 => X"0000003600000000000000380000000000000038000000000000003b00000000",
            INIT_64 => X"000000340000000000000037000000000000003b000000000000003900000000",
            INIT_65 => X"0000003400000000000000340000000000000033000000000000003300000000",
            INIT_66 => X"0000003900000000000000370000000000000035000000000000003300000000",
            INIT_67 => X"0000004b00000000000000780000000000000071000000000000004b00000000",
            INIT_68 => X"00000035000000000000003b0000000000000034000000000000003e00000000",
            INIT_69 => X"0000003600000000000000340000000000000039000000000000003900000000",
            INIT_6A => X"0000003200000000000000300000000000000032000000000000003600000000",
            INIT_6B => X"0000003500000000000000340000000000000038000000000000003900000000",
            INIT_6C => X"0000003300000000000000340000000000000036000000000000003900000000",
            INIT_6D => X"0000003000000000000000350000000000000037000000000000003600000000",
            INIT_6E => X"0000005f000000000000003d0000000000000034000000000000003200000000",
            INIT_6F => X"00000032000000000000003e0000000000000065000000000000007c00000000",
            INIT_70 => X"00000037000000000000003a0000000000000035000000000000003e00000000",
            INIT_71 => X"0000003c000000000000003c000000000000003d000000000000003b00000000",
            INIT_72 => X"0000004b000000000000003a0000000000000037000000000000003900000000",
            INIT_73 => X"0000004500000000000000440000000000000048000000000000004c00000000",
            INIT_74 => X"00000049000000000000004b000000000000004a000000000000004b00000000",
            INIT_75 => X"000000350000000000000037000000000000003a000000000000004600000000",
            INIT_76 => X"0000007f000000000000006b0000000000000045000000000000003300000000",
            INIT_77 => X"000000330000000000000036000000000000003a000000000000005b00000000",
            INIT_78 => X"0000002e00000000000000330000000000000033000000000000004000000000",
            INIT_79 => X"0000003500000000000000390000000000000038000000000000003300000000",
            INIT_7A => X"0000003e00000000000000320000000000000033000000000000003400000000",
            INIT_7B => X"00000039000000000000003c000000000000003e000000000000004000000000",
            INIT_7C => X"000000400000000000000040000000000000003e000000000000003c00000000",
            INIT_7D => X"0000003700000000000000340000000000000035000000000000004000000000",
            INIT_7E => X"0000004800000000000000690000000000000067000000000000004600000000",
            INIT_7F => X"0000003200000000000000340000000000000032000000000000003500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE23;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE24 : if BRAM_NAME = "sampleifmap_layersamples_instance24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001e00000000000000300000000000000046000000000000004100000000",
            INIT_01 => X"0000002d000000000000002c0000000000000028000000000000001700000000",
            INIT_02 => X"0000000f000000000000000a0000000000000028000000000000002d00000000",
            INIT_03 => X"0000003000000000000000330000000000000035000000000000002c00000000",
            INIT_04 => X"0000005b000000000000005d000000000000005a000000000000004100000000",
            INIT_05 => X"00000037000000000000003c0000000000000051000000000000005f00000000",
            INIT_06 => X"000000440000000000000029000000000000006f000000000000007000000000",
            INIT_07 => X"0000004300000000000000360000000000000033000000000000004d00000000",
            INIT_08 => X"0000001e000000000000003c000000000000004f000000000000004500000000",
            INIT_09 => X"0000003100000000000000310000000000000041000000000000002900000000",
            INIT_0A => X"0000001900000000000000070000000000000023000000000000003100000000",
            INIT_0B => X"0000003100000000000000370000000000000045000000000000004100000000",
            INIT_0C => X"0000005000000000000000530000000000000055000000000000004d00000000",
            INIT_0D => X"0000003b00000000000000370000000000000051000000000000005700000000",
            INIT_0E => X"0000002f000000000000001f0000000000000079000000000000008300000000",
            INIT_0F => X"0000003d00000000000000410000000000000036000000000000003800000000",
            INIT_10 => X"0000002900000000000000480000000000000054000000000000004900000000",
            INIT_11 => X"000000360000000000000032000000000000004a000000000000004000000000",
            INIT_12 => X"00000024000000000000000b0000000000000020000000000000003600000000",
            INIT_13 => X"00000027000000000000002f0000000000000043000000000000003c00000000",
            INIT_14 => X"0000003e000000000000003b000000000000004d000000000000004b00000000",
            INIT_15 => X"0000003f00000000000000300000000000000055000000000000005300000000",
            INIT_16 => X"0000002900000000000000170000000000000080000000000000008b00000000",
            INIT_17 => X"000000300000000000000049000000000000004e000000000000004600000000",
            INIT_18 => X"000000360000000000000050000000000000004b000000000000005800000000",
            INIT_19 => X"0000003f00000000000000370000000000000044000000000000005000000000",
            INIT_1A => X"000000250000000000000011000000000000001c000000000000003a00000000",
            INIT_1B => X"0000002700000000000000280000000000000033000000000000002b00000000",
            INIT_1C => X"00000046000000000000004b0000000000000062000000000000005500000000",
            INIT_1D => X"0000004400000000000000320000000000000054000000000000005600000000",
            INIT_1E => X"0000004b000000000000002f0000000000000089000000000000008e00000000",
            INIT_1F => X"000000260000000000000041000000000000005d000000000000006400000000",
            INIT_20 => X"00000042000000000000006f0000000000000059000000000000005f00000000",
            INIT_21 => X"00000044000000000000003d000000000000003d000000000000005100000000",
            INIT_22 => X"00000016000000000000000f0000000000000016000000000000003e00000000",
            INIT_23 => X"0000003f00000000000000330000000000000023000000000000001f00000000",
            INIT_24 => X"000000470000000000000048000000000000004b000000000000004800000000",
            INIT_25 => X"0000004e00000000000000330000000000000053000000000000004d00000000",
            INIT_26 => X"000000570000000000000057000000000000009c000000000000009500000000",
            INIT_27 => X"00000058000000000000004b000000000000005f000000000000006300000000",
            INIT_28 => X"0000004d00000000000000520000000000000053000000000000005200000000",
            INIT_29 => X"000000390000000000000040000000000000003a000000000000004700000000",
            INIT_2A => X"0000001c00000000000000110000000000000014000000000000003b00000000",
            INIT_2B => X"000000470000000000000047000000000000003d000000000000003200000000",
            INIT_2C => X"0000003800000000000000440000000000000043000000000000004500000000",
            INIT_2D => X"0000004e00000000000000460000000000000053000000000000002900000000",
            INIT_2E => X"00000059000000000000006200000000000000ac000000000000009c00000000",
            INIT_2F => X"000000630000000000000070000000000000006f000000000000005e00000000",
            INIT_30 => X"0000003b00000000000000200000000000000040000000000000004500000000",
            INIT_31 => X"000000310000000000000049000000000000004a000000000000004800000000",
            INIT_32 => X"0000003e000000000000001d0000000000000012000000000000003100000000",
            INIT_33 => X"0000003f00000000000000560000000000000055000000000000005200000000",
            INIT_34 => X"0000002b000000000000005f0000000000000034000000000000002200000000",
            INIT_35 => X"0000004e0000000000000055000000000000005e000000000000001900000000",
            INIT_36 => X"0000006b000000000000006d00000000000000b400000000000000a600000000",
            INIT_37 => X"0000002f00000000000000560000000000000083000000000000006c00000000",
            INIT_38 => X"0000004600000000000000190000000000000035000000000000003b00000000",
            INIT_39 => X"0000003d0000000000000050000000000000004e000000000000005100000000",
            INIT_3A => X"0000005e0000000000000035000000000000000a000000000000002800000000",
            INIT_3B => X"00000019000000000000004b0000000000000058000000000000005700000000",
            INIT_3C => X"00000039000000000000005c000000000000002d000000000000000d00000000",
            INIT_3D => X"0000006200000000000000590000000000000065000000000000003200000000",
            INIT_3E => X"0000007c000000000000007800000000000000b3000000000000009000000000",
            INIT_3F => X"0000001800000000000000340000000000000080000000000000007c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000660000000000000031000000000000002f000000000000004400000000",
            INIT_41 => X"0000004f000000000000003f0000000000000059000000000000007700000000",
            INIT_42 => X"0000006000000000000000510000000000000022000000000000004200000000",
            INIT_43 => X"0000000e0000000000000029000000000000005a000000000000005900000000",
            INIT_44 => X"000000470000000000000043000000000000005c000000000000003400000000",
            INIT_45 => X"00000073000000000000006e0000000000000071000000000000006f00000000",
            INIT_46 => X"0000007f0000000000000079000000000000009c000000000000008800000000",
            INIT_47 => X"00000016000000000000001f0000000000000073000000000000007c00000000",
            INIT_48 => X"0000007200000000000000370000000000000035000000000000004d00000000",
            INIT_49 => X"000000370000000000000041000000000000007b000000000000008000000000",
            INIT_4A => X"0000006e000000000000006f0000000000000052000000000000004f00000000",
            INIT_4B => X"0000002500000000000000140000000000000045000000000000006a00000000",
            INIT_4C => X"0000006100000000000000530000000000000069000000000000005c00000000",
            INIT_4D => X"0000005c00000000000000730000000000000078000000000000007600000000",
            INIT_4E => X"0000007f000000000000007d0000000000000093000000000000009000000000",
            INIT_4F => X"00000017000000000000000e000000000000005f000000000000007700000000",
            INIT_50 => X"000000700000000000000036000000000000003a000000000000005500000000",
            INIT_51 => X"0000003100000000000000640000000000000084000000000000008100000000",
            INIT_52 => X"0000006d00000000000000680000000000000054000000000000002700000000",
            INIT_53 => X"00000053000000000000003f000000000000005d000000000000007d00000000",
            INIT_54 => X"0000006e0000000000000068000000000000005e000000000000006100000000",
            INIT_55 => X"000000390000000000000055000000000000007f000000000000006d00000000",
            INIT_56 => X"0000007c000000000000007b0000000000000096000000000000009800000000",
            INIT_57 => X"00000015000000000000000c000000000000005d000000000000007200000000",
            INIT_58 => X"0000006b00000000000000320000000000000035000000000000006c00000000",
            INIT_59 => X"0000004b00000000000000800000000000000083000000000000007e00000000",
            INIT_5A => X"0000006b0000000000000055000000000000005b000000000000003300000000",
            INIT_5B => X"000000930000000000000081000000000000006e000000000000008a00000000",
            INIT_5C => X"0000007700000000000000710000000000000078000000000000008400000000",
            INIT_5D => X"0000005d000000000000005a0000000000000073000000000000007500000000",
            INIT_5E => X"0000007d0000000000000071000000000000008d00000000000000a000000000",
            INIT_5F => X"00000009000000000000000e0000000000000065000000000000007900000000",
            INIT_60 => X"0000005c000000000000002b000000000000002a000000000000006000000000",
            INIT_61 => X"0000007700000000000000820000000000000080000000000000006a00000000",
            INIT_62 => X"000000890000000000000072000000000000007b000000000000007800000000",
            INIT_63 => X"000000840000000000000069000000000000006e000000000000009400000000",
            INIT_64 => X"0000008600000000000000800000000000000087000000000000009200000000",
            INIT_65 => X"00000077000000000000007e0000000000000078000000000000008c00000000",
            INIT_66 => X"0000006a00000000000000630000000000000091000000000000009800000000",
            INIT_67 => X"0000002800000000000000120000000000000063000000000000008200000000",
            INIT_68 => X"00000059000000000000003b0000000000000042000000000000006100000000",
            INIT_69 => X"000000880000000000000085000000000000006f000000000000006400000000",
            INIT_6A => X"000000910000000000000096000000000000008c000000000000009300000000",
            INIT_6B => X"0000007f00000000000000830000000000000088000000000000008e00000000",
            INIT_6C => X"000000930000000000000088000000000000007b000000000000007d00000000",
            INIT_6D => X"00000088000000000000009c000000000000008e000000000000009700000000",
            INIT_6E => X"00000070000000000000006d0000000000000090000000000000009200000000",
            INIT_6F => X"000000530000000000000032000000000000005c000000000000008200000000",
            INIT_70 => X"0000005f000000000000004b0000000000000048000000000000006900000000",
            INIT_71 => X"000000850000000000000085000000000000005e000000000000006800000000",
            INIT_72 => X"0000008500000000000000800000000000000087000000000000008f00000000",
            INIT_73 => X"0000009800000000000000a00000000000000096000000000000009300000000",
            INIT_74 => X"0000008700000000000000840000000000000090000000000000009100000000",
            INIT_75 => X"000000a500000000000000a2000000000000008a000000000000008a00000000",
            INIT_76 => X"00000077000000000000007e000000000000007f00000000000000a300000000",
            INIT_77 => X"0000004d000000000000003b000000000000005f000000000000007600000000",
            INIT_78 => X"0000005b00000000000000440000000000000044000000000000005e00000000",
            INIT_79 => X"00000083000000000000007b0000000000000062000000000000006500000000",
            INIT_7A => X"0000004f000000000000008a00000000000000c1000000000000009300000000",
            INIT_7B => X"000000a200000000000000930000000000000093000000000000007c00000000",
            INIT_7C => X"00000090000000000000009800000000000000ab00000000000000b400000000",
            INIT_7D => X"000000b300000000000000940000000000000079000000000000009000000000",
            INIT_7E => X"0000007b000000000000008000000000000000a000000000000000b400000000",
            INIT_7F => X"00000054000000000000001a000000000000003f000000000000007000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE24;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE25 : if BRAM_NAME = "sampleifmap_layersamples_instance25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000059000000000000004a000000000000004f000000000000005800000000",
            INIT_01 => X"0000008100000000000000780000000000000078000000000000006e00000000",
            INIT_02 => X"0000005700000000000000c000000000000000b8000000000000007800000000",
            INIT_03 => X"000000a600000000000000a4000000000000009c000000000000007200000000",
            INIT_04 => X"000000b600000000000000b700000000000000a1000000000000009a00000000",
            INIT_05 => X"0000008f000000000000009400000000000000ad00000000000000bb00000000",
            INIT_06 => X"0000007c000000000000008e00000000000000c300000000000000b500000000",
            INIT_07 => X"000000760000000000000029000000000000002c000000000000006b00000000",
            INIT_08 => X"0000006000000000000000670000000000000059000000000000005b00000000",
            INIT_09 => X"0000006a000000000000006f0000000000000064000000000000007400000000",
            INIT_0A => X"000000a800000000000000bb0000000000000080000000000000007200000000",
            INIT_0B => X"000000ac00000000000000ac0000000000000099000000000000008c00000000",
            INIT_0C => X"000000a3000000000000009d00000000000000a400000000000000a700000000",
            INIT_0D => X"0000009c00000000000000ab00000000000000a500000000000000a100000000",
            INIT_0E => X"0000007200000000000000a7000000000000009100000000000000a100000000",
            INIT_0F => X"0000005e000000000000002a000000000000004a000000000000006a00000000",
            INIT_10 => X"0000007a00000000000000780000000000000061000000000000006500000000",
            INIT_11 => X"0000005b000000000000005f000000000000004e000000000000007200000000",
            INIT_12 => X"000000cc0000000000000081000000000000006e000000000000007300000000",
            INIT_13 => X"0000009900000000000000a0000000000000008900000000000000a700000000",
            INIT_14 => X"000000b200000000000000aa00000000000000ba00000000000000b300000000",
            INIT_15 => X"000000a500000000000000a2000000000000009c00000000000000b300000000",
            INIT_16 => X"000000480000000000000068000000000000008c000000000000009c00000000",
            INIT_17 => X"0000007200000000000000460000000000000059000000000000005400000000",
            INIT_18 => X"00000060000000000000007a000000000000006b000000000000006e00000000",
            INIT_19 => X"000000640000000000000048000000000000004c000000000000005a00000000",
            INIT_1A => X"0000008c0000000000000057000000000000007f000000000000006d00000000",
            INIT_1B => X"000000b400000000000000a6000000000000009f00000000000000bd00000000",
            INIT_1C => X"000000bc00000000000000be00000000000000ad00000000000000ae00000000",
            INIT_1D => X"000000a100000000000000a2000000000000009900000000000000a200000000",
            INIT_1E => X"0000004a000000000000004b0000000000000095000000000000009900000000",
            INIT_1F => X"0000008a0000000000000070000000000000003e000000000000004200000000",
            INIT_20 => X"0000004e0000000000000059000000000000006a000000000000007700000000",
            INIT_21 => X"00000067000000000000003c0000000000000047000000000000005900000000",
            INIT_22 => X"000000420000000000000072000000000000005f000000000000004b00000000",
            INIT_23 => X"000000be00000000000000ae00000000000000b5000000000000007f00000000",
            INIT_24 => X"000000c100000000000000b800000000000000ab00000000000000ba00000000",
            INIT_25 => X"000000a500000000000000ab00000000000000a000000000000000a400000000",
            INIT_26 => X"0000005c0000000000000068000000000000008b000000000000009200000000",
            INIT_27 => X"000000730000000000000070000000000000005e000000000000004d00000000",
            INIT_28 => X"00000067000000000000003a000000000000005e000000000000007e00000000",
            INIT_29 => X"0000005f0000000000000048000000000000004c000000000000006a00000000",
            INIT_2A => X"0000006300000000000000780000000000000041000000000000005e00000000",
            INIT_2B => X"000000bc00000000000000c400000000000000a1000000000000005b00000000",
            INIT_2C => X"000000a700000000000000a700000000000000c100000000000000b600000000",
            INIT_2D => X"000000a1000000000000009a00000000000000a000000000000000aa00000000",
            INIT_2E => X"00000051000000000000006e000000000000008a000000000000009100000000",
            INIT_2F => X"00000064000000000000006d0000000000000088000000000000006900000000",
            INIT_30 => X"0000006800000000000000460000000000000052000000000000006f00000000",
            INIT_31 => X"000000540000000000000045000000000000005e000000000000007100000000",
            INIT_32 => X"0000007d0000000000000055000000000000006d000000000000007400000000",
            INIT_33 => X"000000c800000000000000ba000000000000009b000000000000007f00000000",
            INIT_34 => X"0000009d00000000000000b100000000000000bb00000000000000bb00000000",
            INIT_35 => X"000000a600000000000000a400000000000000a2000000000000009400000000",
            INIT_36 => X"000000610000000000000079000000000000009500000000000000a200000000",
            INIT_37 => X"0000006100000000000000610000000000000073000000000000007800000000",
            INIT_38 => X"000000b4000000000000008c000000000000005c000000000000006500000000",
            INIT_39 => X"0000004c0000000000000055000000000000007b000000000000009700000000",
            INIT_3A => X"00000054000000000000005a000000000000007c000000000000006700000000",
            INIT_3B => X"000000c800000000000000ad00000000000000af000000000000009200000000",
            INIT_3C => X"0000009f00000000000000ad00000000000000ad00000000000000bc00000000",
            INIT_3D => X"000000ad00000000000000a300000000000000ac000000000000009f00000000",
            INIT_3E => X"000000830000000000000083000000000000008b00000000000000a400000000",
            INIT_3F => X"000000600000000000000064000000000000005f000000000000007000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d100000000000000c00000000000000090000000000000007700000000",
            INIT_41 => X"0000006c000000000000007f000000000000009d00000000000000c200000000",
            INIT_42 => X"0000006f000000000000006a000000000000005e000000000000006a00000000",
            INIT_43 => X"000000c500000000000000b000000000000000af000000000000007c00000000",
            INIT_44 => X"000000a500000000000000b000000000000000aa00000000000000b800000000",
            INIT_45 => X"000000a300000000000000af00000000000000c5000000000000009c00000000",
            INIT_46 => X"00000065000000000000007a0000000000000083000000000000009300000000",
            INIT_47 => X"00000066000000000000006b0000000000000060000000000000006400000000",
            INIT_48 => X"000000a9000000000000008a0000000000000074000000000000006e00000000",
            INIT_49 => X"0000008800000000000000a000000000000000c400000000000000c500000000",
            INIT_4A => X"0000008a000000000000005c0000000000000063000000000000008100000000",
            INIT_4B => X"000000a900000000000000b4000000000000009f000000000000009200000000",
            INIT_4C => X"000000b200000000000000af000000000000008d000000000000008e00000000",
            INIT_4D => X"0000009700000000000000b300000000000000bc00000000000000a600000000",
            INIT_4E => X"0000003a0000000000000070000000000000009a000000000000008f00000000",
            INIT_4F => X"0000004900000000000000660000000000000065000000000000005b00000000",
            INIT_50 => X"0000006b000000000000004a0000000000000057000000000000005b00000000",
            INIT_51 => X"000000a300000000000000bf00000000000000b900000000000000a500000000",
            INIT_52 => X"00000066000000000000006a0000000000000080000000000000008600000000",
            INIT_53 => X"0000007400000000000000920000000000000084000000000000007600000000",
            INIT_54 => X"000000b600000000000000a10000000000000063000000000000004d00000000",
            INIT_55 => X"000000a700000000000000ad000000000000009f00000000000000b700000000",
            INIT_56 => X"0000002b000000000000005e0000000000000087000000000000009c00000000",
            INIT_57 => X"0000004d0000000000000044000000000000005c000000000000005b00000000",
            INIT_58 => X"0000002c0000000000000032000000000000005f000000000000005100000000",
            INIT_59 => X"000000bb00000000000000a60000000000000094000000000000005f00000000",
            INIT_5A => X"00000072000000000000007e000000000000009000000000000000ae00000000",
            INIT_5B => X"0000006b00000000000000770000000000000072000000000000006800000000",
            INIT_5C => X"000000b6000000000000009d0000000000000052000000000000005100000000",
            INIT_5D => X"0000009600000000000000a900000000000000b200000000000000a900000000",
            INIT_5E => X"0000003f000000000000002c000000000000006c000000000000009800000000",
            INIT_5F => X"0000005600000000000000500000000000000045000000000000006100000000",
            INIT_60 => X"000000150000000000000034000000000000005f000000000000005a00000000",
            INIT_61 => X"000000b00000000000000092000000000000006d000000000000001c00000000",
            INIT_62 => X"0000007f000000000000008e00000000000000b500000000000000ca00000000",
            INIT_63 => X"0000008200000000000000720000000000000077000000000000007800000000",
            INIT_64 => X"000000a900000000000000900000000000000076000000000000008100000000",
            INIT_65 => X"0000009800000000000000b400000000000000ad000000000000009f00000000",
            INIT_66 => X"00000055000000000000002c0000000000000044000000000000007700000000",
            INIT_67 => X"0000006a00000000000000a70000000000000072000000000000003300000000",
            INIT_68 => X"000000340000000000000039000000000000005b000000000000005f00000000",
            INIT_69 => X"0000009c00000000000000770000000000000031000000000000001800000000",
            INIT_6A => X"0000009b00000000000000ba00000000000000cb00000000000000bb00000000",
            INIT_6B => X"0000007500000000000000740000000000000085000000000000008d00000000",
            INIT_6C => X"00000099000000000000008b0000000000000077000000000000006d00000000",
            INIT_6D => X"0000007d000000000000009c00000000000000a7000000000000009f00000000",
            INIT_6E => X"0000004000000000000000440000000000000041000000000000006500000000",
            INIT_6F => X"0000007a00000000000000aa0000000000000090000000000000003700000000",
            INIT_70 => X"000000490000000000000020000000000000004b000000000000005e00000000",
            INIT_71 => X"0000007300000000000000360000000000000021000000000000002e00000000",
            INIT_72 => X"000000c200000000000000c300000000000000b0000000000000009600000000",
            INIT_73 => X"000000920000000000000088000000000000009b00000000000000b100000000",
            INIT_74 => X"00000077000000000000005e0000000000000065000000000000008b00000000",
            INIT_75 => X"000000690000000000000060000000000000005f000000000000006500000000",
            INIT_76 => X"0000006d000000000000006b0000000000000076000000000000008300000000",
            INIT_77 => X"0000006a000000000000009a000000000000008f000000000000008000000000",
            INIT_78 => X"0000004c00000000000000180000000000000023000000000000004e00000000",
            INIT_79 => X"0000003b000000000000001b0000000000000028000000000000004100000000",
            INIT_7A => X"000000b000000000000000960000000000000088000000000000007800000000",
            INIT_7B => X"000000ba00000000000000a500000000000000b700000000000000c000000000",
            INIT_7C => X"00000056000000000000006b00000000000000aa00000000000000cf00000000",
            INIT_7D => X"0000008c00000000000000700000000000000055000000000000004200000000",
            INIT_7E => X"000000890000000000000089000000000000009500000000000000a900000000",
            INIT_7F => X"00000080000000000000009a000000000000008f000000000000009600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE25;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE26 : if BRAM_NAME = "sampleifmap_layersamples_instance26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002e00000000000000400000000000000051000000000000004400000000",
            INIT_01 => X"00000050000000000000004b0000000000000039000000000000002100000000",
            INIT_02 => X"0000002200000000000000140000000000000046000000000000005300000000",
            INIT_03 => X"000000420000000000000046000000000000004b000000000000004700000000",
            INIT_04 => X"00000079000000000000007c0000000000000078000000000000005700000000",
            INIT_05 => X"000000520000000000000054000000000000006c000000000000007e00000000",
            INIT_06 => X"0000005b000000000000003b0000000000000081000000000000008800000000",
            INIT_07 => X"00000057000000000000004c0000000000000043000000000000006000000000",
            INIT_08 => X"0000002f000000000000004a0000000000000066000000000000005000000000",
            INIT_09 => X"000000540000000000000054000000000000005c000000000000003800000000",
            INIT_0A => X"000000300000000000000012000000000000003e000000000000005800000000",
            INIT_0B => X"00000049000000000000004d000000000000005c000000000000005d00000000",
            INIT_0C => X"0000006a000000000000006f0000000000000075000000000000006b00000000",
            INIT_0D => X"00000053000000000000004d000000000000006c000000000000007500000000",
            INIT_0E => X"00000041000000000000002d000000000000008b000000000000009700000000",
            INIT_0F => X"00000051000000000000005a0000000000000042000000000000004700000000",
            INIT_10 => X"000000380000000000000058000000000000006d000000000000005f00000000",
            INIT_11 => X"0000005a00000000000000560000000000000069000000000000005400000000",
            INIT_12 => X"0000003c00000000000000140000000000000035000000000000005c00000000",
            INIT_13 => X"0000003c00000000000000420000000000000058000000000000005900000000",
            INIT_14 => X"00000054000000000000004e0000000000000066000000000000006700000000",
            INIT_15 => X"0000005600000000000000420000000000000072000000000000007200000000",
            INIT_16 => X"000000370000000000000023000000000000008f000000000000009e00000000",
            INIT_17 => X"0000003b00000000000000620000000000000062000000000000005400000000",
            INIT_18 => X"0000004900000000000000640000000000000064000000000000007400000000",
            INIT_19 => X"0000006000000000000000580000000000000066000000000000006d00000000",
            INIT_1A => X"00000038000000000000001a000000000000002d000000000000005e00000000",
            INIT_1B => X"0000003700000000000000360000000000000043000000000000004100000000",
            INIT_1C => X"0000006200000000000000610000000000000075000000000000006a00000000",
            INIT_1D => X"0000005b00000000000000450000000000000072000000000000007600000000",
            INIT_1E => X"0000005d0000000000000040000000000000009600000000000000a000000000",
            INIT_1F => X"00000032000000000000005e000000000000007e000000000000007800000000",
            INIT_20 => X"0000005d00000000000000800000000000000068000000000000007800000000",
            INIT_21 => X"0000005e000000000000005a000000000000005e000000000000007200000000",
            INIT_22 => X"00000024000000000000001a0000000000000027000000000000005d00000000",
            INIT_23 => X"0000005600000000000000490000000000000037000000000000002f00000000",
            INIT_24 => X"00000065000000000000006b0000000000000071000000000000006900000000",
            INIT_25 => X"00000067000000000000004a000000000000006d000000000000006700000000",
            INIT_26 => X"00000074000000000000007000000000000000ac00000000000000a200000000",
            INIT_27 => X"0000006c00000000000000670000000000000084000000000000008100000000",
            INIT_28 => X"0000006200000000000000620000000000000066000000000000006900000000",
            INIT_29 => X"0000004e000000000000005b0000000000000059000000000000005f00000000",
            INIT_2A => X"0000002b000000000000001b0000000000000023000000000000005800000000",
            INIT_2B => X"0000006c000000000000006a000000000000005d000000000000004d00000000",
            INIT_2C => X"0000004e00000000000000640000000000000065000000000000006700000000",
            INIT_2D => X"000000660000000000000062000000000000006e000000000000003900000000",
            INIT_2E => X"0000007f000000000000008200000000000000ba00000000000000a700000000",
            INIT_2F => X"0000007800000000000000840000000000000090000000000000008100000000",
            INIT_30 => X"0000004f00000000000000300000000000000060000000000000005e00000000",
            INIT_31 => X"0000003f000000000000005d0000000000000064000000000000005a00000000",
            INIT_32 => X"0000005a0000000000000026000000000000001d000000000000004a00000000",
            INIT_33 => X"0000006300000000000000820000000000000081000000000000007e00000000",
            INIT_34 => X"0000003900000000000000730000000000000047000000000000003a00000000",
            INIT_35 => X"0000006a0000000000000071000000000000007b000000000000002500000000",
            INIT_36 => X"0000008c000000000000008d00000000000000c100000000000000b700000000",
            INIT_37 => X"0000003b000000000000006500000000000000a0000000000000008900000000",
            INIT_38 => X"00000069000000000000002f0000000000000054000000000000005600000000",
            INIT_39 => X"00000047000000000000005e0000000000000061000000000000006700000000",
            INIT_3A => X"0000008b00000000000000490000000000000014000000000000003800000000",
            INIT_3B => X"000000290000000000000072000000000000008c000000000000008a00000000",
            INIT_3C => X"0000004f00000000000000730000000000000041000000000000001a00000000",
            INIT_3D => X"0000008c0000000000000078000000000000007d000000000000003b00000000",
            INIT_3E => X"00000094000000000000009600000000000000c300000000000000b000000000",
            INIT_3F => X"00000018000000000000003f000000000000009b000000000000009000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008c000000000000004a000000000000004e000000000000006200000000",
            INIT_41 => X"0000005c00000000000000500000000000000072000000000000009500000000",
            INIT_42 => X"000000900000000000000071000000000000002c000000000000004700000000",
            INIT_43 => X"00000017000000000000003f0000000000000086000000000000008800000000",
            INIT_44 => X"00000056000000000000005e000000000000007c000000000000004500000000",
            INIT_45 => X"000000a5000000000000009b000000000000008b000000000000007000000000",
            INIT_46 => X"00000096000000000000009600000000000000b100000000000000aa00000000",
            INIT_47 => X"000000160000000000000029000000000000008e000000000000009200000000",
            INIT_48 => X"00000094000000000000004e0000000000000051000000000000007400000000",
            INIT_49 => X"000000450000000000000054000000000000009b00000000000000a300000000",
            INIT_4A => X"0000008e0000000000000089000000000000005a000000000000005100000000",
            INIT_4B => X"000000380000000000000021000000000000005d000000000000008a00000000",
            INIT_4C => X"000000800000000000000073000000000000008f000000000000007c00000000",
            INIT_4D => X"00000081000000000000009c000000000000009c000000000000009700000000",
            INIT_4E => X"0000009a000000000000009800000000000000ad00000000000000a700000000",
            INIT_4F => X"0000001800000000000000160000000000000079000000000000009400000000",
            INIT_50 => X"000000910000000000000049000000000000004f000000000000007800000000",
            INIT_51 => X"00000041000000000000007f00000000000000a600000000000000a500000000",
            INIT_52 => X"0000007f000000000000008e0000000000000072000000000000003600000000",
            INIT_53 => X"0000006c0000000000000047000000000000005d000000000000007e00000000",
            INIT_54 => X"000000a100000000000000920000000000000085000000000000008700000000",
            INIT_55 => X"00000057000000000000007500000000000000a5000000000000009c00000000",
            INIT_56 => X"0000009c000000000000009700000000000000af00000000000000a900000000",
            INIT_57 => X"0000001700000000000000130000000000000074000000000000009100000000",
            INIT_58 => X"0000008a00000000000000420000000000000045000000000000007b00000000",
            INIT_59 => X"0000005f00000000000000a500000000000000a800000000000000a100000000",
            INIT_5A => X"00000070000000000000008a000000000000008c000000000000004b00000000",
            INIT_5B => X"000000a200000000000000880000000000000066000000000000006d00000000",
            INIT_5C => X"000000870000000000000097000000000000009a000000000000009900000000",
            INIT_5D => X"0000008800000000000000760000000000000085000000000000007c00000000",
            INIT_5E => X"0000009d000000000000009200000000000000aa00000000000000bd00000000",
            INIT_5F => X"0000000b00000000000000140000000000000077000000000000009400000000",
            INIT_60 => X"00000079000000000000003c0000000000000039000000000000006a00000000",
            INIT_61 => X"0000009800000000000000ad00000000000000a4000000000000008700000000",
            INIT_62 => X"00000076000000000000007f0000000000000093000000000000009000000000",
            INIT_63 => X"0000008b0000000000000066000000000000005c000000000000007300000000",
            INIT_64 => X"000000740000000000000085000000000000008a000000000000008d00000000",
            INIT_65 => X"000000880000000000000077000000000000006b000000000000007800000000",
            INIT_66 => X"00000091000000000000008700000000000000ae00000000000000b000000000",
            INIT_67 => X"0000002b000000000000001a000000000000007200000000000000a100000000",
            INIT_68 => X"00000074000000000000004e0000000000000055000000000000007400000000",
            INIT_69 => X"000000ab00000000000000ac000000000000008c000000000000007f00000000",
            INIT_6A => X"000000780000000000000082000000000000007c000000000000009900000000",
            INIT_6B => X"0000006e00000000000000710000000000000076000000000000007700000000",
            INIT_6C => X"0000007d0000000000000077000000000000006c000000000000006900000000",
            INIT_6D => X"000000750000000000000081000000000000007a000000000000008300000000",
            INIT_6E => X"0000009a000000000000008d00000000000000a2000000000000009000000000",
            INIT_6F => X"0000005f0000000000000041000000000000007000000000000000a600000000",
            INIT_70 => X"0000007800000000000000630000000000000060000000000000008400000000",
            INIT_71 => X"000000a800000000000000a50000000000000072000000000000008200000000",
            INIT_72 => X"000000700000000000000068000000000000006b000000000000008b00000000",
            INIT_73 => X"00000084000000000000008e0000000000000081000000000000007c00000000",
            INIT_74 => X"0000006f000000000000006b0000000000000077000000000000007a00000000",
            INIT_75 => X"00000090000000000000008d0000000000000076000000000000007300000000",
            INIT_76 => X"0000009f0000000000000092000000000000007b000000000000008e00000000",
            INIT_77 => X"0000005e00000000000000480000000000000070000000000000009d00000000",
            INIT_78 => X"00000076000000000000005d000000000000005a000000000000007900000000",
            INIT_79 => X"000000a60000000000000097000000000000007c000000000000007f00000000",
            INIT_7A => X"00000045000000000000007900000000000000ab000000000000009900000000",
            INIT_7B => X"0000008b000000000000007b000000000000007c000000000000006b00000000",
            INIT_7C => X"0000007700000000000000800000000000000090000000000000009b00000000",
            INIT_7D => X"000000a700000000000000830000000000000067000000000000007a00000000",
            INIT_7E => X"000000a00000000000000080000000000000008c000000000000009f00000000",
            INIT_7F => X"000000680000000000000022000000000000004b000000000000009500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE26;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE27 : if BRAM_NAME = "sampleifmap_layersamples_instance27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007e00000000000000640000000000000064000000000000007000000000",
            INIT_01 => X"000000a300000000000000950000000000000098000000000000008d00000000",
            INIT_02 => X"0000004700000000000000a600000000000000a3000000000000008a00000000",
            INIT_03 => X"0000008d000000000000008b0000000000000085000000000000006400000000",
            INIT_04 => X"0000009e00000000000000a00000000000000088000000000000008100000000",
            INIT_05 => X"0000007e000000000000007d000000000000009700000000000000a300000000",
            INIT_06 => X"0000008f000000000000007a00000000000000b100000000000000a900000000",
            INIT_07 => X"0000008b0000000000000033000000000000003d000000000000008f00000000",
            INIT_08 => X"0000008100000000000000830000000000000070000000000000007000000000",
            INIT_09 => X"000000890000000000000090000000000000007c000000000000009300000000",
            INIT_0A => X"0000009900000000000000a80000000000000079000000000000008f00000000",
            INIT_0B => X"000000930000000000000092000000000000007f000000000000007a00000000",
            INIT_0C => X"0000008a0000000000000084000000000000008b000000000000008d00000000",
            INIT_0D => X"000000860000000000000099000000000000008f000000000000008600000000",
            INIT_0E => X"0000007a00000000000000920000000000000082000000000000009100000000",
            INIT_0F => X"0000006f000000000000003a0000000000000064000000000000008600000000",
            INIT_10 => X"0000008e00000000000000950000000000000076000000000000007900000000",
            INIT_11 => X"00000076000000000000007b0000000000000061000000000000008d00000000",
            INIT_12 => X"000000bb0000000000000079000000000000007e000000000000008f00000000",
            INIT_13 => X"000000820000000000000088000000000000006e000000000000009100000000",
            INIT_14 => X"0000009a000000000000009400000000000000a1000000000000009a00000000",
            INIT_15 => X"0000009100000000000000960000000000000086000000000000009700000000",
            INIT_16 => X"000000570000000000000061000000000000007b000000000000008600000000",
            INIT_17 => X"0000008600000000000000610000000000000077000000000000006700000000",
            INIT_18 => X"0000006f00000000000000970000000000000087000000000000008800000000",
            INIT_19 => X"0000007d000000000000005d0000000000000065000000000000007a00000000",
            INIT_1A => X"0000007d00000000000000600000000000000099000000000000008600000000",
            INIT_1B => X"000000a00000000000000092000000000000008800000000000000a900000000",
            INIT_1C => X"000000a700000000000000a60000000000000094000000000000009600000000",
            INIT_1D => X"0000009100000000000000900000000000000080000000000000008d00000000",
            INIT_1E => X"0000005e000000000000004b0000000000000082000000000000008400000000",
            INIT_1F => X"000000a900000000000000950000000000000057000000000000005300000000",
            INIT_20 => X"0000005e0000000000000070000000000000008c000000000000009400000000",
            INIT_21 => X"0000008200000000000000540000000000000068000000000000007900000000",
            INIT_22 => X"0000004a000000000000008d0000000000000074000000000000006600000000",
            INIT_23 => X"000000aa000000000000009b00000000000000a3000000000000007600000000",
            INIT_24 => X"000000a7000000000000009d000000000000009500000000000000a500000000",
            INIT_25 => X"0000009100000000000000930000000000000089000000000000009200000000",
            INIT_26 => X"00000071000000000000006d000000000000007c000000000000007f00000000",
            INIT_27 => X"000000a1000000000000009c0000000000000077000000000000006000000000",
            INIT_28 => X"0000007d00000000000000480000000000000077000000000000009800000000",
            INIT_29 => X"0000007900000000000000630000000000000065000000000000008100000000",
            INIT_2A => X"0000007d000000000000009a000000000000005b000000000000007800000000",
            INIT_2B => X"000000a900000000000000b50000000000000096000000000000005d00000000",
            INIT_2C => X"0000008f000000000000009100000000000000ad00000000000000a200000000",
            INIT_2D => X"0000008b00000000000000810000000000000087000000000000008f00000000",
            INIT_2E => X"0000006600000000000000750000000000000078000000000000007d00000000",
            INIT_2F => X"00000099000000000000009a00000000000000ab000000000000008100000000",
            INIT_30 => X"0000007b00000000000000520000000000000068000000000000008800000000",
            INIT_31 => X"0000007300000000000000620000000000000076000000000000008800000000",
            INIT_32 => X"000000940000000000000075000000000000008d000000000000009600000000",
            INIT_33 => X"000000b300000000000000ad0000000000000095000000000000008100000000",
            INIT_34 => X"0000008f000000000000009f00000000000000a800000000000000a500000000",
            INIT_35 => X"0000008d000000000000008c000000000000008b000000000000007e00000000",
            INIT_36 => X"0000006d000000000000007a0000000000000085000000000000008800000000",
            INIT_37 => X"00000095000000000000009600000000000000a4000000000000009800000000",
            INIT_38 => X"000000bf0000000000000096000000000000006f000000000000007d00000000",
            INIT_39 => X"0000006f0000000000000079000000000000009e00000000000000ac00000000",
            INIT_3A => X"0000006900000000000000730000000000000099000000000000009100000000",
            INIT_3B => X"000000ac000000000000009a00000000000000a1000000000000009400000000",
            INIT_3C => X"0000008d000000000000009c000000000000009b00000000000000a100000000",
            INIT_3D => X"0000008f00000000000000880000000000000093000000000000008900000000",
            INIT_3E => X"00000086000000000000007b000000000000008c000000000000008900000000",
            INIT_3F => X"00000095000000000000009e0000000000000095000000000000009c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000dc00000000000000c800000000000000a2000000000000009500000000",
            INIT_41 => X"0000009300000000000000aa00000000000000bd00000000000000d100000000",
            INIT_42 => X"00000088000000000000007d000000000000007a000000000000009100000000",
            INIT_43 => X"000000a40000000000000096000000000000009f000000000000008b00000000",
            INIT_44 => X"0000008e000000000000009f000000000000009b000000000000009b00000000",
            INIT_45 => X"00000088000000000000009300000000000000a9000000000000008500000000",
            INIT_46 => X"00000072000000000000006b000000000000007e000000000000007f00000000",
            INIT_47 => X"0000009c00000000000000a0000000000000008f000000000000009a00000000",
            INIT_48 => X"000000be000000000000009d0000000000000089000000000000008b00000000",
            INIT_49 => X"000000b000000000000000bf00000000000000d700000000000000d500000000",
            INIT_4A => X"000000a30000000000000075000000000000008400000000000000a900000000",
            INIT_4B => X"0000008f000000000000009a000000000000009700000000000000ad00000000",
            INIT_4C => X"0000009800000000000000990000000000000081000000000000007c00000000",
            INIT_4D => X"0000007c000000000000009500000000000000a3000000000000009100000000",
            INIT_4E => X"0000004a00000000000000600000000000000083000000000000007700000000",
            INIT_4F => X"0000007800000000000000970000000000000095000000000000009100000000",
            INIT_50 => X"000000860000000000000061000000000000006f000000000000007300000000",
            INIT_51 => X"000000c100000000000000d300000000000000cf00000000000000bf00000000",
            INIT_52 => X"0000007f000000000000009100000000000000ad00000000000000b100000000",
            INIT_53 => X"000000680000000000000086000000000000008f000000000000009000000000",
            INIT_54 => X"0000009b000000000000008b000000000000005c000000000000004900000000",
            INIT_55 => X"0000008e0000000000000094000000000000008a00000000000000a100000000",
            INIT_56 => X"0000003c00000000000000550000000000000075000000000000008300000000",
            INIT_57 => X"0000006d000000000000006f0000000000000091000000000000009200000000",
            INIT_58 => X"0000004000000000000000410000000000000072000000000000006a00000000",
            INIT_59 => X"000000d500000000000000c300000000000000b2000000000000007800000000",
            INIT_5A => X"0000009900000000000000ad00000000000000b900000000000000ca00000000",
            INIT_5B => X"0000007d000000000000008d0000000000000096000000000000008e00000000",
            INIT_5C => X"0000009a000000000000008e0000000000000060000000000000006c00000000",
            INIT_5D => X"0000007f000000000000009500000000000000a1000000000000009000000000",
            INIT_5E => X"0000006100000000000000310000000000000062000000000000008300000000",
            INIT_5F => X"000000750000000000000076000000000000006c000000000000009300000000",
            INIT_60 => X"00000026000000000000003e0000000000000070000000000000007400000000",
            INIT_61 => X"000000c700000000000000b40000000000000087000000000000002900000000",
            INIT_62 => X"000000b200000000000000b700000000000000cc00000000000000d400000000",
            INIT_63 => X"000000a1000000000000009e00000000000000a400000000000000ab00000000",
            INIT_64 => X"0000008d0000000000000087000000000000008b000000000000009d00000000",
            INIT_65 => X"0000007e000000000000009c0000000000000099000000000000008700000000",
            INIT_66 => X"0000007c000000000000003b0000000000000042000000000000006700000000",
            INIT_67 => X"0000008300000000000000c50000000000000088000000000000005400000000",
            INIT_68 => X"0000004e000000000000004f000000000000007b000000000000007f00000000",
            INIT_69 => X"000000bf00000000000000950000000000000042000000000000002500000000",
            INIT_6A => X"000000c200000000000000d600000000000000db00000000000000d000000000",
            INIT_6B => X"0000009f00000000000000a500000000000000b400000000000000b800000000",
            INIT_6C => X"00000083000000000000007b000000000000007d000000000000008700000000",
            INIT_6D => X"0000007200000000000000870000000000000093000000000000008a00000000",
            INIT_6E => X"0000005b0000000000000055000000000000004f000000000000006c00000000",
            INIT_6F => X"0000008f00000000000000c900000000000000ac000000000000004e00000000",
            INIT_70 => X"0000006b00000000000000340000000000000068000000000000007d00000000",
            INIT_71 => X"00000097000000000000004e0000000000000030000000000000004300000000",
            INIT_72 => X"000000da00000000000000d900000000000000cb00000000000000bd00000000",
            INIT_73 => X"000000b600000000000000b400000000000000c300000000000000cd00000000",
            INIT_74 => X"0000007a000000000000005e000000000000007400000000000000a500000000",
            INIT_75 => X"0000006f00000000000000590000000000000059000000000000006100000000",
            INIT_76 => X"000000860000000000000082000000000000008a000000000000009600000000",
            INIT_77 => X"0000008100000000000000bc00000000000000b5000000000000009f00000000",
            INIT_78 => X"0000007300000000000000280000000000000033000000000000006600000000",
            INIT_79 => X"0000004e0000000000000029000000000000003a000000000000006000000000",
            INIT_7A => X"000000cf00000000000000b900000000000000b500000000000000a000000000",
            INIT_7B => X"000000ce00000000000000c400000000000000d200000000000000da00000000",
            INIT_7C => X"00000071000000000000007c00000000000000b400000000000000d600000000",
            INIT_7D => X"000000a000000000000000840000000000000066000000000000005600000000",
            INIT_7E => X"000000a700000000000000a700000000000000a700000000000000ba00000000",
            INIT_7F => X"0000009c00000000000000b900000000000000b300000000000000b400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE27;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE28 : if BRAM_NAME = "sampleifmap_layersamples_instance28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001e000000000000002e0000000000000040000000000000003200000000",
            INIT_01 => X"0000003900000000000000370000000000000024000000000000001600000000",
            INIT_02 => X"00000012000000000000000c0000000000000036000000000000003b00000000",
            INIT_03 => X"000000320000000000000031000000000000002c000000000000002b00000000",
            INIT_04 => X"0000004d0000000000000051000000000000004d000000000000003a00000000",
            INIT_05 => X"000000390000000000000038000000000000004e000000000000005300000000",
            INIT_06 => X"0000003a000000000000001f000000000000005d000000000000006100000000",
            INIT_07 => X"0000004200000000000000350000000000000029000000000000004100000000",
            INIT_08 => X"0000001d00000000000000390000000000000051000000000000003a00000000",
            INIT_09 => X"0000003c000000000000003b000000000000003d000000000000002300000000",
            INIT_0A => X"0000001b0000000000000007000000000000002f000000000000004000000000",
            INIT_0B => X"0000002f000000000000003b000000000000003e000000000000003800000000",
            INIT_0C => X"00000044000000000000004a000000000000004a000000000000004400000000",
            INIT_0D => X"0000003c00000000000000330000000000000051000000000000004e00000000",
            INIT_0E => X"0000002700000000000000150000000000000060000000000000006f00000000",
            INIT_0F => X"000000420000000000000045000000000000002c000000000000002d00000000",
            INIT_10 => X"0000002300000000000000460000000000000057000000000000004800000000",
            INIT_11 => X"00000041000000000000003c0000000000000048000000000000003500000000",
            INIT_12 => X"0000002300000000000000070000000000000026000000000000004500000000",
            INIT_13 => X"0000002100000000000000300000000000000041000000000000003400000000",
            INIT_14 => X"0000003700000000000000320000000000000042000000000000004300000000",
            INIT_15 => X"0000003e000000000000002d0000000000000052000000000000004d00000000",
            INIT_16 => X"0000002600000000000000100000000000000063000000000000007400000000",
            INIT_17 => X"00000033000000000000004d000000000000004b000000000000003f00000000",
            INIT_18 => X"0000002f0000000000000050000000000000004c000000000000005e00000000",
            INIT_19 => X"0000004a00000000000000410000000000000048000000000000004700000000",
            INIT_1A => X"00000022000000000000000c000000000000001e000000000000004800000000",
            INIT_1B => X"0000001e00000000000000230000000000000034000000000000002800000000",
            INIT_1C => X"0000004500000000000000440000000000000057000000000000004b00000000",
            INIT_1D => X"00000043000000000000002e000000000000004d000000000000005100000000",
            INIT_1E => X"00000049000000000000002a000000000000006b000000000000007700000000",
            INIT_1F => X"0000002200000000000000440000000000000060000000000000005f00000000",
            INIT_20 => X"0000003c000000000000006a000000000000004f000000000000006100000000",
            INIT_21 => X"0000004c00000000000000480000000000000044000000000000004b00000000",
            INIT_22 => X"00000011000000000000000c0000000000000018000000000000004900000000",
            INIT_23 => X"0000003b00000000000000330000000000000025000000000000001c00000000",
            INIT_24 => X"00000047000000000000004b000000000000004f000000000000004800000000",
            INIT_25 => X"0000004d000000000000002d0000000000000049000000000000004700000000",
            INIT_26 => X"0000005500000000000000520000000000000081000000000000008000000000",
            INIT_27 => X"0000005000000000000000490000000000000061000000000000005e00000000",
            INIT_28 => X"00000043000000000000004b000000000000004d000000000000005200000000",
            INIT_29 => X"0000003d000000000000004d0000000000000045000000000000003d00000000",
            INIT_2A => X"00000016000000000000000d0000000000000013000000000000004300000000",
            INIT_2B => X"000000490000000000000047000000000000003b000000000000002c00000000",
            INIT_2C => X"0000003500000000000000490000000000000048000000000000004800000000",
            INIT_2D => X"0000004d000000000000003e0000000000000049000000000000002200000000",
            INIT_2E => X"0000005b00000000000000600000000000000093000000000000008800000000",
            INIT_2F => X"0000005c0000000000000068000000000000006e000000000000005c00000000",
            INIT_30 => X"0000003300000000000000190000000000000046000000000000004800000000",
            INIT_31 => X"00000032000000000000004f000000000000004f000000000000003e00000000",
            INIT_32 => X"000000360000000000000018000000000000000f000000000000003800000000",
            INIT_33 => X"0000003e000000000000004d000000000000004b000000000000004900000000",
            INIT_34 => X"0000002a00000000000000600000000000000033000000000000002200000000",
            INIT_35 => X"0000004a00000000000000480000000000000058000000000000001600000000",
            INIT_36 => X"0000006c000000000000006800000000000000a1000000000000009500000000",
            INIT_37 => X"0000002b00000000000000510000000000000083000000000000006b00000000",
            INIT_38 => X"000000460000000000000015000000000000003b000000000000003f00000000",
            INIT_39 => X"0000003a000000000000004b0000000000000048000000000000004d00000000",
            INIT_3A => X"00000051000000000000002f0000000000000008000000000000002900000000",
            INIT_3B => X"00000012000000000000003e000000000000004b000000000000004b00000000",
            INIT_3C => X"0000004000000000000000590000000000000027000000000000000600000000",
            INIT_3D => X"000000530000000000000048000000000000005e000000000000002a00000000",
            INIT_3E => X"00000078000000000000007200000000000000a2000000000000008300000000",
            INIT_3F => X"0000001500000000000000340000000000000085000000000000007600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006800000000000000310000000000000035000000000000004900000000",
            INIT_41 => X"0000004600000000000000390000000000000058000000000000007900000000",
            INIT_42 => X"0000005300000000000000470000000000000017000000000000003300000000",
            INIT_43 => X"000000070000000000000022000000000000004f000000000000004e00000000",
            INIT_44 => X"0000003e000000000000003c0000000000000051000000000000002800000000",
            INIT_45 => X"0000005d000000000000005b0000000000000063000000000000005000000000",
            INIT_46 => X"000000790000000000000078000000000000008d000000000000007300000000",
            INIT_47 => X"000000140000000000000021000000000000007c000000000000007900000000",
            INIT_48 => X"000000760000000000000038000000000000003a000000000000005600000000",
            INIT_49 => X"000000330000000000000040000000000000007f000000000000008300000000",
            INIT_4A => X"0000006300000000000000610000000000000040000000000000003b00000000",
            INIT_4B => X"0000001c000000000000000d000000000000003a000000000000005e00000000",
            INIT_4C => X"000000500000000000000049000000000000005d000000000000005300000000",
            INIT_4D => X"0000004a000000000000005f0000000000000069000000000000006200000000",
            INIT_4E => X"0000007e00000000000000770000000000000084000000000000007400000000",
            INIT_4F => X"00000017000000000000000d0000000000000065000000000000007f00000000",
            INIT_50 => X"000000740000000000000035000000000000003b000000000000005b00000000",
            INIT_51 => X"0000003000000000000000670000000000000087000000000000008400000000",
            INIT_52 => X"000000610000000000000060000000000000004b000000000000002000000000",
            INIT_53 => X"000000490000000000000032000000000000004a000000000000006600000000",
            INIT_54 => X"0000006100000000000000590000000000000052000000000000005a00000000",
            INIT_55 => X"000000310000000000000047000000000000006c000000000000006200000000",
            INIT_56 => X"0000008a0000000000000077000000000000007c000000000000007700000000",
            INIT_57 => X"00000014000000000000000a000000000000005b000000000000007b00000000",
            INIT_58 => X"0000006e000000000000002f0000000000000033000000000000006500000000",
            INIT_59 => X"0000004800000000000000870000000000000087000000000000008100000000",
            INIT_5A => X"0000004f00000000000000520000000000000054000000000000002e00000000",
            INIT_5B => X"0000008700000000000000750000000000000056000000000000005e00000000",
            INIT_5C => X"0000005e000000000000005d0000000000000066000000000000007800000000",
            INIT_5D => X"00000058000000000000004a0000000000000058000000000000005c00000000",
            INIT_5E => X"0000008d00000000000000760000000000000073000000000000008400000000",
            INIT_5F => X"00000007000000000000000b000000000000005b000000000000007700000000",
            INIT_60 => X"0000006000000000000000280000000000000028000000000000005800000000",
            INIT_61 => X"00000077000000000000008b0000000000000083000000000000006b00000000",
            INIT_62 => X"0000005900000000000000570000000000000066000000000000006b00000000",
            INIT_63 => X"0000006c0000000000000051000000000000004a000000000000005f00000000",
            INIT_64 => X"0000005d0000000000000064000000000000006e000000000000007600000000",
            INIT_65 => X"0000005f00000000000000570000000000000055000000000000006600000000",
            INIT_66 => X"0000007100000000000000650000000000000078000000000000007c00000000",
            INIT_67 => X"00000020000000000000000f0000000000000059000000000000007b00000000",
            INIT_68 => X"0000005c0000000000000037000000000000003f000000000000005f00000000",
            INIT_69 => X"00000089000000000000008b000000000000006e000000000000006400000000",
            INIT_6A => X"0000005c00000000000000650000000000000061000000000000007b00000000",
            INIT_6B => X"0000005600000000000000560000000000000058000000000000005a00000000",
            INIT_6C => X"0000006c00000000000000640000000000000058000000000000005500000000",
            INIT_6D => X"0000005f000000000000006e000000000000006c000000000000007200000000",
            INIT_6E => X"00000073000000000000006b0000000000000075000000000000006d00000000",
            INIT_6F => X"0000004c00000000000000310000000000000058000000000000008000000000",
            INIT_70 => X"0000006000000000000000470000000000000045000000000000006a00000000",
            INIT_71 => X"0000008700000000000000860000000000000056000000000000006800000000",
            INIT_72 => X"0000005800000000000000510000000000000057000000000000007400000000",
            INIT_73 => X"0000006a000000000000006e0000000000000060000000000000006000000000",
            INIT_74 => X"0000005c0000000000000057000000000000005f000000000000006200000000",
            INIT_75 => X"00000080000000000000007f000000000000006b000000000000006100000000",
            INIT_76 => X"000000770000000000000074000000000000005e000000000000007a00000000",
            INIT_77 => X"000000460000000000000035000000000000005c000000000000007a00000000",
            INIT_78 => X"0000005c00000000000000400000000000000040000000000000006000000000",
            INIT_79 => X"000000850000000000000079000000000000005f000000000000006700000000",
            INIT_7A => X"0000003300000000000000640000000000000096000000000000008100000000",
            INIT_7B => X"0000007100000000000000620000000000000065000000000000005800000000",
            INIT_7C => X"0000005f00000000000000650000000000000077000000000000008300000000",
            INIT_7D => X"0000009800000000000000710000000000000053000000000000006000000000",
            INIT_7E => X"0000007c00000000000000620000000000000078000000000000009400000000",
            INIT_7F => X"00000048000000000000000d0000000000000039000000000000007600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE28;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE29 : if BRAM_NAME = "sampleifmap_layersamples_instance29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005a0000000000000047000000000000004c000000000000005700000000",
            INIT_01 => X"000000820000000000000078000000000000007c000000000000007300000000",
            INIT_02 => X"0000003a0000000000000096000000000000008e000000000000006e00000000",
            INIT_03 => X"0000007800000000000000770000000000000074000000000000005400000000",
            INIT_04 => X"0000008600000000000000850000000000000071000000000000006c00000000",
            INIT_05 => X"0000006e0000000000000067000000000000007e000000000000008900000000",
            INIT_06 => X"00000072000000000000006300000000000000a3000000000000009f00000000",
            INIT_07 => X"0000006b0000000000000021000000000000002a000000000000007500000000",
            INIT_08 => X"0000005d00000000000000640000000000000058000000000000005600000000",
            INIT_09 => X"0000006900000000000000750000000000000063000000000000007500000000",
            INIT_0A => X"0000008b000000000000009b0000000000000066000000000000006e00000000",
            INIT_0B => X"000000810000000000000081000000000000006f000000000000006b00000000",
            INIT_0C => X"00000076000000000000006d0000000000000077000000000000007c00000000",
            INIT_0D => X"00000071000000000000007c0000000000000076000000000000007100000000",
            INIT_0E => X"0000006300000000000000830000000000000075000000000000008300000000",
            INIT_0F => X"0000005700000000000000270000000000000048000000000000006900000000",
            INIT_10 => X"0000007300000000000000780000000000000060000000000000005f00000000",
            INIT_11 => X"0000005600000000000000630000000000000047000000000000006d00000000",
            INIT_12 => X"000000b0000000000000006a0000000000000063000000000000006c00000000",
            INIT_13 => X"00000075000000000000007b000000000000005e000000000000008200000000",
            INIT_14 => X"000000880000000000000081000000000000008d000000000000008900000000",
            INIT_15 => X"000000790000000000000078000000000000006f000000000000008300000000",
            INIT_16 => X"000000430000000000000050000000000000006b000000000000007500000000",
            INIT_17 => X"0000006e00000000000000430000000000000051000000000000004800000000",
            INIT_18 => X"00000057000000000000007d0000000000000070000000000000006d00000000",
            INIT_19 => X"0000005e00000000000000470000000000000048000000000000005800000000",
            INIT_1A => X"0000007300000000000000490000000000000079000000000000006400000000",
            INIT_1B => X"0000009400000000000000870000000000000076000000000000009800000000",
            INIT_1C => X"0000009500000000000000940000000000000082000000000000008500000000",
            INIT_1D => X"0000007a00000000000000790000000000000071000000000000007d00000000",
            INIT_1E => X"0000004e000000000000003a0000000000000071000000000000007200000000",
            INIT_1F => X"0000008a00000000000000730000000000000038000000000000003d00000000",
            INIT_20 => X"0000004300000000000000590000000000000074000000000000007700000000",
            INIT_21 => X"00000066000000000000003c0000000000000048000000000000005800000000",
            INIT_22 => X"00000037000000000000006d0000000000000057000000000000004800000000",
            INIT_23 => X"0000009c000000000000008d0000000000000092000000000000006500000000",
            INIT_24 => X"00000098000000000000008c0000000000000088000000000000009800000000",
            INIT_25 => X"0000007c000000000000007f000000000000007b000000000000008600000000",
            INIT_26 => X"00000062000000000000005d0000000000000069000000000000006d00000000",
            INIT_27 => X"00000077000000000000007a0000000000000062000000000000004d00000000",
            INIT_28 => X"0000005d00000000000000320000000000000061000000000000007e00000000",
            INIT_29 => X"00000060000000000000004b0000000000000046000000000000006000000000",
            INIT_2A => X"000000610000000000000076000000000000003b000000000000005a00000000",
            INIT_2B => X"0000009700000000000000a20000000000000083000000000000004900000000",
            INIT_2C => X"0000007f000000000000008400000000000000a3000000000000009600000000",
            INIT_2D => X"00000075000000000000006e0000000000000076000000000000007d00000000",
            INIT_2E => X"0000004f000000000000005e0000000000000066000000000000006900000000",
            INIT_2F => X"0000006a0000000000000070000000000000008e000000000000006b00000000",
            INIT_30 => X"0000005900000000000000370000000000000051000000000000007000000000",
            INIT_31 => X"000000590000000000000045000000000000004e000000000000005c00000000",
            INIT_32 => X"000000760000000000000053000000000000006b000000000000007700000000",
            INIT_33 => X"0000009c0000000000000097000000000000007d000000000000006b00000000",
            INIT_34 => X"0000007e0000000000000094000000000000009b000000000000009400000000",
            INIT_35 => X"000000750000000000000078000000000000007b000000000000006c00000000",
            INIT_36 => X"0000005600000000000000540000000000000066000000000000007200000000",
            INIT_37 => X"0000006900000000000000630000000000000079000000000000008100000000",
            INIT_38 => X"0000009a00000000000000780000000000000056000000000000006200000000",
            INIT_39 => X"0000004e0000000000000045000000000000005f000000000000007700000000",
            INIT_3A => X"0000004e0000000000000057000000000000007e000000000000007300000000",
            INIT_3B => X"000000960000000000000084000000000000008b000000000000007d00000000",
            INIT_3C => X"0000007e0000000000000092000000000000008e000000000000008d00000000",
            INIT_3D => X"0000007b00000000000000760000000000000084000000000000007900000000",
            INIT_3E => X"0000006f00000000000000520000000000000058000000000000007300000000",
            INIT_3F => X"00000067000000000000006a0000000000000065000000000000007900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b600000000000000a70000000000000088000000000000007400000000",
            INIT_41 => X"0000005c00000000000000600000000000000077000000000000009f00000000",
            INIT_42 => X"0000006f0000000000000066000000000000005a000000000000006600000000",
            INIT_43 => X"0000008f00000000000000830000000000000088000000000000007000000000",
            INIT_44 => X"000000800000000000000096000000000000008e000000000000008600000000",
            INIT_45 => X"000000770000000000000084000000000000009c000000000000007500000000",
            INIT_46 => X"00000053000000000000004e0000000000000059000000000000006600000000",
            INIT_47 => X"0000006c00000000000000710000000000000060000000000000006a00000000",
            INIT_48 => X"000000920000000000000071000000000000006d000000000000006c00000000",
            INIT_49 => X"00000069000000000000007b000000000000009e00000000000000a600000000",
            INIT_4A => X"0000008c00000000000000550000000000000052000000000000006600000000",
            INIT_4B => X"0000007b0000000000000086000000000000007e000000000000009100000000",
            INIT_4C => X"00000089000000000000008a0000000000000073000000000000006800000000",
            INIT_4D => X"0000006a000000000000008a0000000000000096000000000000008300000000",
            INIT_4E => X"0000002d000000000000004a000000000000006f000000000000006100000000",
            INIT_4F => X"0000004b00000000000000690000000000000065000000000000006000000000",
            INIT_50 => X"0000005600000000000000370000000000000055000000000000005800000000",
            INIT_51 => X"0000007e00000000000000970000000000000097000000000000008b00000000",
            INIT_52 => X"0000005700000000000000570000000000000068000000000000006800000000",
            INIT_53 => X"00000052000000000000006e000000000000006e000000000000006f00000000",
            INIT_54 => X"0000008c0000000000000079000000000000004b000000000000003500000000",
            INIT_55 => X"0000007a00000000000000810000000000000078000000000000009100000000",
            INIT_56 => X"00000020000000000000003e0000000000000062000000000000007400000000",
            INIT_57 => X"0000004000000000000000410000000000000062000000000000006100000000",
            INIT_58 => X"000000200000000000000022000000000000005c000000000000005200000000",
            INIT_59 => X"0000009c00000000000000860000000000000075000000000000004b00000000",
            INIT_5A => X"000000570000000000000062000000000000006d000000000000008d00000000",
            INIT_5B => X"0000005f000000000000005b000000000000005a000000000000005200000000",
            INIT_5C => X"0000008b00000000000000790000000000000046000000000000005200000000",
            INIT_5D => X"0000006b0000000000000080000000000000008f000000000000008100000000",
            INIT_5E => X"0000003f000000000000001d000000000000004e000000000000007100000000",
            INIT_5F => X"0000004200000000000000470000000000000047000000000000006300000000",
            INIT_60 => X"0000000d00000000000000230000000000000056000000000000005a00000000",
            INIT_61 => X"000000940000000000000072000000000000004e000000000000000f00000000",
            INIT_62 => X"00000062000000000000006f000000000000008b00000000000000a200000000",
            INIT_63 => X"000000710000000000000056000000000000005b000000000000006100000000",
            INIT_64 => X"0000007e0000000000000073000000000000006a000000000000007800000000",
            INIT_65 => X"0000006a00000000000000870000000000000087000000000000007600000000",
            INIT_66 => X"0000005b0000000000000026000000000000002a000000000000004f00000000",
            INIT_67 => X"0000005300000000000000990000000000000060000000000000002c00000000",
            INIT_68 => X"00000025000000000000002d0000000000000056000000000000005c00000000",
            INIT_69 => X"0000007a0000000000000057000000000000001f000000000000000d00000000",
            INIT_6A => X"0000007a000000000000009e00000000000000ad000000000000009600000000",
            INIT_6B => X"0000005c000000000000005d0000000000000072000000000000007500000000",
            INIT_6C => X"0000007100000000000000670000000000000055000000000000004d00000000",
            INIT_6D => X"0000005b00000000000000730000000000000085000000000000007e00000000",
            INIT_6E => X"0000003c000000000000003b0000000000000032000000000000004e00000000",
            INIT_6F => X"000000620000000000000086000000000000006c000000000000002a00000000",
            INIT_70 => X"0000003800000000000000180000000000000047000000000000005200000000",
            INIT_71 => X"0000005400000000000000230000000000000017000000000000002400000000",
            INIT_72 => X"000000a500000000000000a50000000000000092000000000000007600000000",
            INIT_73 => X"00000079000000000000006f0000000000000082000000000000009600000000",
            INIT_74 => X"00000062000000000000003f0000000000000042000000000000006c00000000",
            INIT_75 => X"0000005600000000000000460000000000000045000000000000004e00000000",
            INIT_76 => X"000000620000000000000060000000000000006c000000000000007500000000",
            INIT_77 => X"00000059000000000000007b0000000000000074000000000000007800000000",
            INIT_78 => X"000000400000000000000011000000000000001b000000000000004100000000",
            INIT_79 => X"00000025000000000000000f000000000000001d000000000000003400000000",
            INIT_7A => X"0000009600000000000000740000000000000064000000000000005900000000",
            INIT_7B => X"0000009c0000000000000088000000000000009800000000000000aa00000000",
            INIT_7C => X"0000004a0000000000000045000000000000007900000000000000a600000000",
            INIT_7D => X"0000007f00000000000000660000000000000047000000000000002f00000000",
            INIT_7E => X"000000820000000000000083000000000000008b000000000000009c00000000",
            INIT_7F => X"0000007500000000000000920000000000000088000000000000009300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE29;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE30 : if BRAM_NAME = "sampleifmap_layersamples_instance30" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000058000000000000004d000000000000008b00000000000000b300000000",
            INIT_01 => X"00000097000000000000009c000000000000009d000000000000008d00000000",
            INIT_02 => X"000000970000000000000090000000000000009e000000000000009c00000000",
            INIT_03 => X"0000007600000000000000790000000000000088000000000000009700000000",
            INIT_04 => X"000000540000000000000054000000000000006c000000000000007e00000000",
            INIT_05 => X"00000053000000000000005e0000000000000062000000000000006200000000",
            INIT_06 => X"0000006000000000000000540000000000000056000000000000005a00000000",
            INIT_07 => X"0000004d000000000000004c0000000000000057000000000000007500000000",
            INIT_08 => X"000000920000000000000080000000000000008500000000000000b800000000",
            INIT_09 => X"000000a7000000000000009e000000000000009f000000000000009f00000000",
            INIT_0A => X"0000009a000000000000009900000000000000a200000000000000a500000000",
            INIT_0B => X"0000007d00000000000000880000000000000096000000000000009600000000",
            INIT_0C => X"00000052000000000000005a000000000000006d000000000000008100000000",
            INIT_0D => X"00000058000000000000005e0000000000000062000000000000005d00000000",
            INIT_0E => X"0000006a000000000000005b000000000000004c000000000000004e00000000",
            INIT_0F => X"0000005a000000000000005b0000000000000062000000000000007600000000",
            INIT_10 => X"000000aa00000000000000b0000000000000009800000000000000b400000000",
            INIT_11 => X"000000a4000000000000009b000000000000009800000000000000a400000000",
            INIT_12 => X"0000009f00000000000000a200000000000000aa00000000000000a200000000",
            INIT_13 => X"0000008c00000000000000920000000000000097000000000000009c00000000",
            INIT_14 => X"000000470000000000000058000000000000007c000000000000009200000000",
            INIT_15 => X"0000006b00000000000000670000000000000062000000000000005500000000",
            INIT_16 => X"0000006f000000000000006f000000000000006d000000000000006500000000",
            INIT_17 => X"0000005f000000000000005d0000000000000065000000000000006f00000000",
            INIT_18 => X"000000b500000000000000b800000000000000ae00000000000000af00000000",
            INIT_19 => X"000000a300000000000000a4000000000000009800000000000000a800000000",
            INIT_1A => X"000000a800000000000000a700000000000000b300000000000000a600000000",
            INIT_1B => X"000000a4000000000000009f00000000000000a200000000000000ae00000000",
            INIT_1C => X"0000003a00000000000000590000000000000089000000000000009700000000",
            INIT_1D => X"0000006b0000000000000063000000000000005a000000000000004800000000",
            INIT_1E => X"00000079000000000000007d0000000000000080000000000000007500000000",
            INIT_1F => X"0000006f000000000000006d0000000000000061000000000000006900000000",
            INIT_20 => X"000000ac00000000000000a700000000000000ae00000000000000af00000000",
            INIT_21 => X"000000af00000000000000b000000000000000a100000000000000a200000000",
            INIT_22 => X"000000b400000000000000b300000000000000b200000000000000b200000000",
            INIT_23 => X"000000a400000000000000a000000000000000a800000000000000b000000000",
            INIT_24 => X"000000450000000000000078000000000000009c00000000000000ad00000000",
            INIT_25 => X"0000005e0000000000000063000000000000005a000000000000004200000000",
            INIT_26 => X"0000007b000000000000007f000000000000007c000000000000006900000000",
            INIT_27 => X"0000007400000000000000710000000000000068000000000000007000000000",
            INIT_28 => X"000000aa000000000000009000000000000000ae00000000000000b500000000",
            INIT_29 => X"000000b300000000000000b000000000000000a600000000000000a900000000",
            INIT_2A => X"000000b500000000000000b400000000000000b400000000000000b400000000",
            INIT_2B => X"00000096000000000000009f00000000000000ae00000000000000b000000000",
            INIT_2C => X"00000074000000000000009b00000000000000af00000000000000b500000000",
            INIT_2D => X"000000700000000000000083000000000000007d000000000000006000000000",
            INIT_2E => X"00000079000000000000007a0000000000000078000000000000007500000000",
            INIT_2F => X"0000007c00000000000000760000000000000078000000000000007900000000",
            INIT_30 => X"000000b2000000000000008a000000000000009c00000000000000c000000000",
            INIT_31 => X"000000af00000000000000b000000000000000ae00000000000000af00000000",
            INIT_32 => X"000000b800000000000000ba00000000000000b400000000000000b800000000",
            INIT_33 => X"0000009900000000000000ad00000000000000bb00000000000000bb00000000",
            INIT_34 => X"000000a700000000000000ad00000000000000ad00000000000000a600000000",
            INIT_35 => X"0000007900000000000000940000000000000095000000000000009600000000",
            INIT_36 => X"0000006f000000000000006d0000000000000075000000000000007300000000",
            INIT_37 => X"00000080000000000000007b000000000000007a000000000000007800000000",
            INIT_38 => X"000000ab000000000000009c000000000000007d00000000000000b900000000",
            INIT_39 => X"000000b800000000000000af00000000000000af00000000000000ad00000000",
            INIT_3A => X"000000c200000000000000c100000000000000b700000000000000bc00000000",
            INIT_3B => X"000000a600000000000000b800000000000000b900000000000000bd00000000",
            INIT_3C => X"000000b000000000000000b100000000000000ac00000000000000a400000000",
            INIT_3D => X"0000007a000000000000008f000000000000008900000000000000aa00000000",
            INIT_3E => X"000000670000000000000060000000000000006e000000000000006b00000000",
            INIT_3F => X"0000007d000000000000007b0000000000000076000000000000007500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a0000000000000009f0000000000000095000000000000009b00000000",
            INIT_41 => X"000000b400000000000000b200000000000000ad00000000000000ac00000000",
            INIT_42 => X"000000bf00000000000000ba00000000000000ba00000000000000bb00000000",
            INIT_43 => X"000000a000000000000000ac00000000000000af00000000000000bb00000000",
            INIT_44 => X"000000b000000000000000a60000000000000097000000000000009a00000000",
            INIT_45 => X"0000008500000000000000a6000000000000009b00000000000000b700000000",
            INIT_46 => X"0000007700000000000000700000000000000068000000000000006800000000",
            INIT_47 => X"0000007d000000000000007a000000000000007a000000000000007600000000",
            INIT_48 => X"000000a900000000000000930000000000000098000000000000009a00000000",
            INIT_49 => X"000000aa00000000000000b700000000000000b200000000000000b200000000",
            INIT_4A => X"000000c100000000000000c600000000000000bc00000000000000b000000000",
            INIT_4B => X"000000a900000000000000a500000000000000a700000000000000ae00000000",
            INIT_4C => X"000000a90000000000000092000000000000008c000000000000009d00000000",
            INIT_4D => X"0000008d00000000000000ab00000000000000a000000000000000b300000000",
            INIT_4E => X"0000007700000000000000750000000000000068000000000000005f00000000",
            INIT_4F => X"0000007d0000000000000076000000000000007b000000000000007400000000",
            INIT_50 => X"000000b1000000000000009f0000000000000070000000000000008600000000",
            INIT_51 => X"000000ba00000000000000b800000000000000b800000000000000ae00000000",
            INIT_52 => X"000000b000000000000000bf00000000000000c200000000000000ba00000000",
            INIT_53 => X"000000bb00000000000000a7000000000000009e000000000000009b00000000",
            INIT_54 => X"000000970000000000000086000000000000009300000000000000ae00000000",
            INIT_55 => X"0000007c000000000000009b000000000000009c00000000000000a000000000",
            INIT_56 => X"0000006600000000000000690000000000000066000000000000004a00000000",
            INIT_57 => X"0000007f000000000000007b0000000000000075000000000000006b00000000",
            INIT_58 => X"0000009d00000000000000ae000000000000005b000000000000004100000000",
            INIT_59 => X"000000be00000000000000bf00000000000000b1000000000000009300000000",
            INIT_5A => X"000000b000000000000000ac00000000000000b000000000000000bc00000000",
            INIT_5B => X"000000a3000000000000009400000000000000ae00000000000000b800000000",
            INIT_5C => X"000000950000000000000085000000000000009a00000000000000b000000000",
            INIT_5D => X"0000005000000000000000830000000000000095000000000000009800000000",
            INIT_5E => X"0000006600000000000000670000000000000061000000000000004200000000",
            INIT_5F => X"0000007d00000000000000780000000000000071000000000000006700000000",
            INIT_60 => X"000000b100000000000000bf000000000000005c000000000000001500000000",
            INIT_61 => X"000000b600000000000000bd00000000000000ca00000000000000bc00000000",
            INIT_62 => X"000000bc00000000000000a5000000000000009c00000000000000b300000000",
            INIT_63 => X"00000072000000000000009800000000000000ae00000000000000c800000000",
            INIT_64 => X"000000890000000000000078000000000000007f000000000000005f00000000",
            INIT_65 => X"0000004e00000000000000720000000000000088000000000000009700000000",
            INIT_66 => X"0000006200000000000000590000000000000049000000000000004000000000",
            INIT_67 => X"0000007600000000000000750000000000000071000000000000006200000000",
            INIT_68 => X"000000ad00000000000000a80000000000000063000000000000002c00000000",
            INIT_69 => X"000000bb00000000000000bc00000000000000c300000000000000c800000000",
            INIT_6A => X"000000c200000000000000b4000000000000009500000000000000a500000000",
            INIT_6B => X"0000009a00000000000000a800000000000000a800000000000000b900000000",
            INIT_6C => X"0000008a00000000000000910000000000000092000000000000006b00000000",
            INIT_6D => X"000000480000000000000064000000000000007f000000000000009c00000000",
            INIT_6E => X"0000006000000000000000530000000000000040000000000000003900000000",
            INIT_6F => X"0000006f000000000000006c000000000000006a000000000000006200000000",
            INIT_70 => X"0000009f00000000000000750000000000000076000000000000006900000000",
            INIT_71 => X"000000bb00000000000000b400000000000000be00000000000000c400000000",
            INIT_72 => X"000000c100000000000000c600000000000000ad00000000000000ad00000000",
            INIT_73 => X"000000bc00000000000000b400000000000000a500000000000000ab00000000",
            INIT_74 => X"000000b300000000000000ad00000000000000bb00000000000000ae00000000",
            INIT_75 => X"000000480000000000000069000000000000008000000000000000a000000000",
            INIT_76 => X"0000006c00000000000000570000000000000045000000000000004300000000",
            INIT_77 => X"0000006600000000000000610000000000000064000000000000006300000000",
            INIT_78 => X"0000009d00000000000000680000000000000071000000000000008a00000000",
            INIT_79 => X"000000a800000000000000b400000000000000c400000000000000c600000000",
            INIT_7A => X"000000cd00000000000000cb00000000000000bf00000000000000b400000000",
            INIT_7B => X"000000c800000000000000c400000000000000bf00000000000000d200000000",
            INIT_7C => X"000000be00000000000000bc00000000000000bb00000000000000c000000000",
            INIT_7D => X"000000500000000000000071000000000000009900000000000000a800000000",
            INIT_7E => X"0000008700000000000000600000000000000040000000000000004600000000",
            INIT_7F => X"00000062000000000000005a000000000000005a000000000000007800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE30;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE31 : if BRAM_NAME = "sampleifmap_layersamples_instance31" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000930000000000000073000000000000008a000000000000009600000000",
            INIT_01 => X"0000009600000000000000b000000000000000bb00000000000000be00000000",
            INIT_02 => X"000000c600000000000000d300000000000000c700000000000000ab00000000",
            INIT_03 => X"000000cb00000000000000be00000000000000c200000000000000d300000000",
            INIT_04 => X"000000bd00000000000000b800000000000000ba00000000000000bf00000000",
            INIT_05 => X"00000046000000000000006400000000000000a600000000000000be00000000",
            INIT_06 => X"0000008f000000000000006a0000000000000038000000000000002f00000000",
            INIT_07 => X"0000005e000000000000004a000000000000005c000000000000009500000000",
            INIT_08 => X"000000a50000000000000092000000000000009b000000000000009b00000000",
            INIT_09 => X"0000009100000000000000bf00000000000000c000000000000000bd00000000",
            INIT_0A => X"0000009500000000000000a900000000000000d2000000000000009c00000000",
            INIT_0B => X"000000a800000000000000b200000000000000c200000000000000c000000000",
            INIT_0C => X"000000a700000000000000aa00000000000000b500000000000000a900000000",
            INIT_0D => X"0000002b00000000000000430000000000000075000000000000009a00000000",
            INIT_0E => X"0000008f00000000000000680000000000000031000000000000002200000000",
            INIT_0F => X"00000050000000000000003f000000000000006a000000000000009c00000000",
            INIT_10 => X"000000a6000000000000008a00000000000000a200000000000000a500000000",
            INIT_11 => X"0000008900000000000000ba00000000000000be00000000000000c400000000",
            INIT_12 => X"000000a9000000000000009d00000000000000c9000000000000007400000000",
            INIT_13 => X"0000008f000000000000008000000000000000b600000000000000d200000000",
            INIT_14 => X"00000061000000000000007f0000000000000093000000000000007c00000000",
            INIT_15 => X"00000033000000000000002f0000000000000038000000000000005200000000",
            INIT_16 => X"0000009d00000000000000690000000000000040000000000000002b00000000",
            INIT_17 => X"000000410000000000000039000000000000007b000000000000009d00000000",
            INIT_18 => X"0000009e0000000000000078000000000000009600000000000000a900000000",
            INIT_19 => X"0000009800000000000000be00000000000000be00000000000000be00000000",
            INIT_1A => X"000000b900000000000000bc0000000000000099000000000000003c00000000",
            INIT_1B => X"000000ce000000000000009000000000000000a500000000000000c300000000",
            INIT_1C => X"0000003d0000000000000065000000000000008900000000000000b100000000",
            INIT_1D => X"0000005000000000000000470000000000000033000000000000003700000000",
            INIT_1E => X"000000a0000000000000006e000000000000004a000000000000003700000000",
            INIT_1F => X"000000320000000000000036000000000000008e00000000000000b000000000",
            INIT_20 => X"000000a6000000000000009600000000000000a000000000000000aa00000000",
            INIT_21 => X"0000009a00000000000000ba00000000000000bc00000000000000ba00000000",
            INIT_22 => X"00000092000000000000007e0000000000000031000000000000002000000000",
            INIT_23 => X"000000c0000000000000008c000000000000008c000000000000009b00000000",
            INIT_24 => X"0000003e0000000000000061000000000000009c00000000000000cc00000000",
            INIT_25 => X"0000005700000000000000520000000000000049000000000000004900000000",
            INIT_26 => X"000000a6000000000000006b000000000000003e000000000000003a00000000",
            INIT_27 => X"00000033000000000000004800000000000000a700000000000000bc00000000",
            INIT_28 => X"0000009c000000000000009700000000000000ab00000000000000b200000000",
            INIT_29 => X"0000007c00000000000000a300000000000000b200000000000000b500000000",
            INIT_2A => X"000000370000000000000028000000000000001d000000000000002400000000",
            INIT_2B => X"0000008200000000000000650000000000000063000000000000004e00000000",
            INIT_2C => X"00000037000000000000005f000000000000007b000000000000009000000000",
            INIT_2D => X"00000055000000000000003c0000000000000033000000000000003400000000",
            INIT_2E => X"000000990000000000000066000000000000004d000000000000004e00000000",
            INIT_2F => X"00000037000000000000005900000000000000b100000000000000bb00000000",
            INIT_30 => X"00000098000000000000009200000000000000ab00000000000000b500000000",
            INIT_31 => X"00000069000000000000009500000000000000a700000000000000a900000000",
            INIT_32 => X"0000002e0000000000000042000000000000005e000000000000004f00000000",
            INIT_33 => X"00000078000000000000005c0000000000000047000000000000002f00000000",
            INIT_34 => X"0000002900000000000000380000000000000037000000000000005a00000000",
            INIT_35 => X"00000037000000000000001e0000000000000022000000000000002300000000",
            INIT_36 => X"0000007700000000000000610000000000000056000000000000005200000000",
            INIT_37 => X"0000003c000000000000006a00000000000000ae00000000000000ad00000000",
            INIT_38 => X"000000a3000000000000009e000000000000009c00000000000000b100000000",
            INIT_39 => X"00000089000000000000009400000000000000a0000000000000009c00000000",
            INIT_3A => X"0000006b00000000000000660000000000000076000000000000008f00000000",
            INIT_3B => X"00000067000000000000007d000000000000006d000000000000006e00000000",
            INIT_3C => X"0000001300000000000000100000000000000011000000000000002f00000000",
            INIT_3D => X"00000013000000000000000e000000000000001c000000000000001800000000",
            INIT_3E => X"0000006300000000000000600000000000000041000000000000002b00000000",
            INIT_3F => X"00000043000000000000008500000000000000ad000000000000008c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b600000000000000a7000000000000008b000000000000009e00000000",
            INIT_41 => X"000000c000000000000000ab000000000000008c000000000000009700000000",
            INIT_42 => X"000000880000000000000085000000000000007400000000000000ac00000000",
            INIT_43 => X"00000065000000000000007f000000000000008d000000000000009200000000",
            INIT_44 => X"0000001900000000000000200000000000000025000000000000004100000000",
            INIT_45 => X"0000000f000000000000000a0000000000000011000000000000001800000000",
            INIT_46 => X"0000004e00000000000000610000000000000042000000000000001400000000",
            INIT_47 => X"00000069000000000000009c0000000000000094000000000000006200000000",
            INIT_48 => X"000000ab00000000000000ae00000000000000a400000000000000a000000000",
            INIT_49 => X"000000b100000000000000940000000000000088000000000000009e00000000",
            INIT_4A => X"0000009700000000000000a9000000000000009300000000000000b800000000",
            INIT_4B => X"0000007d000000000000008e000000000000008b000000000000007f00000000",
            INIT_4C => X"0000002b000000000000003f000000000000004d000000000000006700000000",
            INIT_4D => X"0000001a00000000000000110000000000000018000000000000002100000000",
            INIT_4E => X"000000320000000000000048000000000000003e000000000000001f00000000",
            INIT_4F => X"000000880000000000000078000000000000005a000000000000004800000000",
            INIT_50 => X"000000a700000000000000a700000000000000a300000000000000a000000000",
            INIT_51 => X"00000078000000000000008c00000000000000a800000000000000b100000000",
            INIT_52 => X"000000820000000000000076000000000000008f00000000000000ab00000000",
            INIT_53 => X"0000009100000000000000a6000000000000009c000000000000007b00000000",
            INIT_54 => X"0000004e000000000000005b0000000000000069000000000000007c00000000",
            INIT_55 => X"0000004300000000000000380000000000000042000000000000004c00000000",
            INIT_56 => X"0000004900000000000000410000000000000041000000000000004600000000",
            INIT_57 => X"0000006a0000000000000051000000000000007b000000000000006400000000",
            INIT_58 => X"00000093000000000000008c000000000000009f000000000000009c00000000",
            INIT_59 => X"0000007b000000000000009900000000000000aa00000000000000b400000000",
            INIT_5A => X"0000007e0000000000000073000000000000009c000000000000008b00000000",
            INIT_5B => X"000000a200000000000000a8000000000000009e000000000000008300000000",
            INIT_5C => X"00000078000000000000007b0000000000000077000000000000007f00000000",
            INIT_5D => X"0000007700000000000000690000000000000068000000000000007000000000",
            INIT_5E => X"0000006d00000000000000680000000000000069000000000000007400000000",
            INIT_5F => X"00000068000000000000005c0000000000000086000000000000007a00000000",
            INIT_60 => X"0000008b000000000000007b000000000000009e00000000000000a400000000",
            INIT_61 => X"0000008c000000000000008d000000000000009c00000000000000ad00000000",
            INIT_62 => X"000000a100000000000000820000000000000079000000000000008d00000000",
            INIT_63 => X"000000a800000000000000a6000000000000009d000000000000009700000000",
            INIT_64 => X"00000084000000000000008f000000000000008a000000000000009000000000",
            INIT_65 => X"00000094000000000000008a0000000000000085000000000000008100000000",
            INIT_66 => X"0000008400000000000000860000000000000089000000000000008f00000000",
            INIT_67 => X"0000009300000000000000730000000000000064000000000000007800000000",
            INIT_68 => X"000000a800000000000000900000000000000095000000000000008e00000000",
            INIT_69 => X"0000009e000000000000009e00000000000000a100000000000000a700000000",
            INIT_6A => X"000000a90000000000000097000000000000009000000000000000a500000000",
            INIT_6B => X"000000a2000000000000009e00000000000000a000000000000000a100000000",
            INIT_6C => X"0000007f00000000000000890000000000000091000000000000009900000000",
            INIT_6D => X"0000009e00000000000000960000000000000095000000000000008d00000000",
            INIT_6E => X"0000008f00000000000000940000000000000096000000000000009f00000000",
            INIT_6F => X"0000009f000000000000008b0000000000000077000000000000007b00000000",
            INIT_70 => X"000000b900000000000000b300000000000000a6000000000000009800000000",
            INIT_71 => X"000000a800000000000000aa00000000000000a700000000000000a700000000",
            INIT_72 => X"000000b200000000000000ad00000000000000a400000000000000a700000000",
            INIT_73 => X"000000850000000000000089000000000000009d00000000000000a900000000",
            INIT_74 => X"00000088000000000000008c000000000000008f000000000000009200000000",
            INIT_75 => X"0000009d00000000000000980000000000000097000000000000008c00000000",
            INIT_76 => X"000000900000000000000099000000000000009c00000000000000a600000000",
            INIT_77 => X"0000009900000000000000900000000000000083000000000000008500000000",
            INIT_78 => X"000000ab00000000000000b700000000000000b2000000000000009f00000000",
            INIT_79 => X"0000009f0000000000000091000000000000007d000000000000008b00000000",
            INIT_7A => X"0000009c0000000000000095000000000000008b00000000000000a200000000",
            INIT_7B => X"0000007300000000000000830000000000000098000000000000009e00000000",
            INIT_7C => X"0000008f0000000000000094000000000000008e000000000000008400000000",
            INIT_7D => X"000000a1000000000000009c000000000000009d000000000000009000000000",
            INIT_7E => X"0000009c0000000000000094000000000000009f00000000000000a700000000",
            INIT_7F => X"0000009800000000000000990000000000000096000000000000009c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE31;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE32 : if BRAM_NAME = "sampleifmap_layersamples_instance32" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003b00000000000000310000000000000060000000000000007600000000",
            INIT_01 => X"000000530000000000000054000000000000005f000000000000006000000000",
            INIT_02 => X"0000005a00000000000000530000000000000061000000000000005f00000000",
            INIT_03 => X"0000004f000000000000004b0000000000000052000000000000005c00000000",
            INIT_04 => X"00000032000000000000003b0000000000000050000000000000005b00000000",
            INIT_05 => X"0000003300000000000000380000000000000038000000000000003700000000",
            INIT_06 => X"0000003a00000000000000330000000000000038000000000000003c00000000",
            INIT_07 => X"0000002f000000000000002f0000000000000035000000000000004c00000000",
            INIT_08 => X"0000006900000000000000590000000000000058000000000000008200000000",
            INIT_09 => X"00000068000000000000005d0000000000000060000000000000006c00000000",
            INIT_0A => X"0000005b000000000000005a0000000000000062000000000000006500000000",
            INIT_0B => X"00000048000000000000004f0000000000000057000000000000005400000000",
            INIT_0C => X"00000032000000000000003d0000000000000048000000000000005200000000",
            INIT_0D => X"0000003300000000000000370000000000000038000000000000003700000000",
            INIT_0E => X"0000004100000000000000350000000000000028000000000000002b00000000",
            INIT_0F => X"00000039000000000000003a000000000000003d000000000000004b00000000",
            INIT_10 => X"0000007a00000000000000810000000000000068000000000000008400000000",
            INIT_11 => X"0000006a000000000000005f0000000000000059000000000000006c00000000",
            INIT_12 => X"0000005e00000000000000620000000000000069000000000000006200000000",
            INIT_13 => X"0000004c000000000000004f0000000000000050000000000000005500000000",
            INIT_14 => X"0000002a0000000000000036000000000000004c000000000000005500000000",
            INIT_15 => X"00000042000000000000003f000000000000003a000000000000003300000000",
            INIT_16 => X"0000004200000000000000430000000000000042000000000000003c00000000",
            INIT_17 => X"000000390000000000000038000000000000003e000000000000004300000000",
            INIT_18 => X"000000840000000000000088000000000000007f000000000000008100000000",
            INIT_19 => X"000000690000000000000068000000000000005a000000000000007000000000",
            INIT_1A => X"0000006600000000000000650000000000000071000000000000006500000000",
            INIT_1B => X"0000005d0000000000000057000000000000005a000000000000006700000000",
            INIT_1C => X"0000001f0000000000000033000000000000004e000000000000004f00000000",
            INIT_1D => X"0000003e00000000000000390000000000000033000000000000002a00000000",
            INIT_1E => X"0000004a000000000000004b000000000000004d000000000000004600000000",
            INIT_1F => X"0000004500000000000000430000000000000037000000000000003c00000000",
            INIT_20 => X"0000007f0000000000000079000000000000007f000000000000008000000000",
            INIT_21 => X"0000007200000000000000720000000000000063000000000000006d00000000",
            INIT_22 => X"000000710000000000000070000000000000006f000000000000006f00000000",
            INIT_23 => X"0000005c00000000000000590000000000000063000000000000006c00000000",
            INIT_24 => X"0000002c000000000000004e0000000000000059000000000000005e00000000",
            INIT_25 => X"0000002e00000000000000380000000000000034000000000000002700000000",
            INIT_26 => X"0000004900000000000000470000000000000043000000000000003500000000",
            INIT_27 => X"000000470000000000000045000000000000003b000000000000004200000000",
            INIT_28 => X"0000007f00000000000000680000000000000083000000000000008900000000",
            INIT_29 => X"000000740000000000000071000000000000006a000000000000007600000000",
            INIT_2A => X"0000007100000000000000740000000000000075000000000000007300000000",
            INIT_2B => X"00000054000000000000005a0000000000000069000000000000006d00000000",
            INIT_2C => X"0000004f00000000000000670000000000000068000000000000006a00000000",
            INIT_2D => X"0000003d0000000000000052000000000000004d000000000000003a00000000",
            INIT_2E => X"000000460000000000000043000000000000003f000000000000003e00000000",
            INIT_2F => X"0000004b00000000000000460000000000000048000000000000004900000000",
            INIT_30 => X"0000008700000000000000660000000000000077000000000000009800000000",
            INIT_31 => X"0000006f00000000000000730000000000000075000000000000007a00000000",
            INIT_32 => X"00000070000000000000007c000000000000007b000000000000007900000000",
            INIT_33 => X"0000005c00000000000000660000000000000071000000000000007300000000",
            INIT_34 => X"0000006e000000000000006d0000000000000065000000000000006400000000",
            INIT_35 => X"00000043000000000000005b0000000000000057000000000000005c00000000",
            INIT_36 => X"0000003b00000000000000380000000000000040000000000000003e00000000",
            INIT_37 => X"0000004e000000000000004a0000000000000048000000000000004500000000",
            INIT_38 => X"0000007e00000000000000780000000000000059000000000000009300000000",
            INIT_39 => X"0000007900000000000000720000000000000076000000000000007800000000",
            INIT_3A => X"00000073000000000000007c000000000000007a000000000000008000000000",
            INIT_3B => X"00000064000000000000006c000000000000006d000000000000007300000000",
            INIT_3C => X"0000006a000000000000006d0000000000000068000000000000006500000000",
            INIT_3D => X"000000480000000000000057000000000000004b000000000000006600000000",
            INIT_3E => X"00000035000000000000002e000000000000003c000000000000003b00000000",
            INIT_3F => X"0000004b00000000000000490000000000000044000000000000004200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000720000000000000078000000000000006f000000000000007600000000",
            INIT_41 => X"0000007700000000000000750000000000000074000000000000007700000000",
            INIT_42 => X"0000006d000000000000006f000000000000007a000000000000008000000000",
            INIT_43 => X"0000005e00000000000000610000000000000067000000000000007300000000",
            INIT_44 => X"0000006400000000000000610000000000000059000000000000005e00000000",
            INIT_45 => X"000000590000000000000072000000000000005f000000000000006d00000000",
            INIT_46 => X"000000470000000000000040000000000000003a000000000000003e00000000",
            INIT_47 => X"0000004b00000000000000480000000000000048000000000000004600000000",
            INIT_48 => X"0000007800000000000000690000000000000071000000000000007700000000",
            INIT_49 => X"0000006f000000000000007b000000000000007a000000000000007c00000000",
            INIT_4A => X"00000079000000000000007d000000000000007b000000000000007600000000",
            INIT_4B => X"0000006f0000000000000065000000000000006d000000000000007600000000",
            INIT_4C => X"0000006000000000000000520000000000000055000000000000006900000000",
            INIT_4D => X"00000067000000000000007a0000000000000064000000000000006a00000000",
            INIT_4E => X"000000490000000000000047000000000000003e000000000000003d00000000",
            INIT_4F => X"0000004b0000000000000044000000000000004b000000000000004700000000",
            INIT_50 => X"0000007e00000000000000720000000000000048000000000000006400000000",
            INIT_51 => X"0000007e000000000000007c000000000000007f000000000000007800000000",
            INIT_52 => X"0000007b00000000000000800000000000000081000000000000007f00000000",
            INIT_53 => X"0000009000000000000000780000000000000077000000000000007900000000",
            INIT_54 => X"00000058000000000000004f0000000000000063000000000000008300000000",
            INIT_55 => X"0000005b000000000000006c0000000000000061000000000000005f00000000",
            INIT_56 => X"0000003b000000000000003d000000000000003e000000000000002e00000000",
            INIT_57 => X"0000004c00000000000000490000000000000046000000000000004000000000",
            INIT_58 => X"00000069000000000000007f0000000000000034000000000000002200000000",
            INIT_59 => X"000000830000000000000084000000000000007a000000000000005d00000000",
            INIT_5A => X"0000008c00000000000000780000000000000073000000000000008100000000",
            INIT_5B => X"000000850000000000000074000000000000009700000000000000a600000000",
            INIT_5C => X"000000610000000000000056000000000000006e000000000000008d00000000",
            INIT_5D => X"000000310000000000000056000000000000005c000000000000006000000000",
            INIT_5E => X"0000003c000000000000003e000000000000003c000000000000002a00000000",
            INIT_5F => X"0000004a00000000000000450000000000000042000000000000003e00000000",
            INIT_60 => X"0000007d000000000000008e0000000000000040000000000000000400000000",
            INIT_61 => X"00000084000000000000008c000000000000009a000000000000008c00000000",
            INIT_62 => X"0000009c000000000000007b000000000000006b000000000000007f00000000",
            INIT_63 => X"000000530000000000000077000000000000009300000000000000b200000000",
            INIT_64 => X"000000640000000000000053000000000000005b000000000000004000000000",
            INIT_65 => X"00000031000000000000004d000000000000005c000000000000006f00000000",
            INIT_66 => X"000000390000000000000037000000000000002f000000000000002900000000",
            INIT_67 => X"0000004400000000000000420000000000000043000000000000003b00000000",
            INIT_68 => X"0000007b000000000000007a0000000000000048000000000000001800000000",
            INIT_69 => X"0000008d000000000000008f0000000000000096000000000000009c00000000",
            INIT_6A => X"000000a0000000000000008f000000000000006a000000000000007700000000",
            INIT_6B => X"0000007700000000000000800000000000000081000000000000009700000000",
            INIT_6C => X"0000006d00000000000000730000000000000074000000000000004d00000000",
            INIT_6D => X"0000002d0000000000000044000000000000005a000000000000007b00000000",
            INIT_6E => X"000000370000000000000033000000000000002b000000000000002300000000",
            INIT_6F => X"0000003e000000000000003a000000000000003e000000000000003b00000000",
            INIT_70 => X"00000070000000000000004a0000000000000052000000000000004500000000",
            INIT_71 => X"0000008f00000000000000860000000000000091000000000000009600000000",
            INIT_72 => X"0000009c00000000000000a10000000000000084000000000000008300000000",
            INIT_73 => X"0000009700000000000000850000000000000072000000000000007d00000000",
            INIT_74 => X"00000098000000000000009200000000000000a0000000000000009100000000",
            INIT_75 => X"0000002f000000000000004b000000000000005d000000000000008100000000",
            INIT_76 => X"0000004400000000000000380000000000000030000000000000002f00000000",
            INIT_77 => X"000000390000000000000036000000000000003c000000000000003c00000000",
            INIT_78 => X"00000070000000000000003b0000000000000041000000000000005700000000",
            INIT_79 => X"0000007d00000000000000860000000000000096000000000000009800000000",
            INIT_7A => X"000000a500000000000000a7000000000000009b000000000000008f00000000",
            INIT_7B => X"000000a0000000000000008f0000000000000084000000000000009b00000000",
            INIT_7C => X"000000a1000000000000009f000000000000009e00000000000000a200000000",
            INIT_7D => X"0000003900000000000000540000000000000078000000000000008900000000",
            INIT_7E => X"0000005f0000000000000040000000000000002b000000000000003300000000",
            INIT_7F => X"0000003900000000000000360000000000000037000000000000005100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE32;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE33 : if BRAM_NAME = "sampleifmap_layersamples_instance33" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000660000000000000040000000000000004e000000000000005800000000",
            INIT_01 => X"0000006c0000000000000081000000000000008d000000000000009000000000",
            INIT_02 => X"0000009d00000000000000af00000000000000a5000000000000008b00000000",
            INIT_03 => X"0000009f00000000000000860000000000000086000000000000009e00000000",
            INIT_04 => X"0000009800000000000000930000000000000094000000000000009a00000000",
            INIT_05 => X"0000003100000000000000490000000000000087000000000000009a00000000",
            INIT_06 => X"00000067000000000000004b0000000000000023000000000000001e00000000",
            INIT_07 => X"00000039000000000000002c000000000000003d000000000000006f00000000",
            INIT_08 => X"0000007400000000000000570000000000000057000000000000005600000000",
            INIT_09 => X"0000006900000000000000910000000000000093000000000000008f00000000",
            INIT_0A => X"0000006c000000000000008500000000000000b3000000000000008000000000",
            INIT_0B => X"00000079000000000000007a000000000000008b000000000000009100000000",
            INIT_0C => X"00000079000000000000007c0000000000000087000000000000007d00000000",
            INIT_0D => X"00000018000000000000002a0000000000000058000000000000007200000000",
            INIT_0E => X"000000660000000000000049000000000000001d000000000000001300000000",
            INIT_0F => X"0000002e00000000000000270000000000000050000000000000007500000000",
            INIT_10 => X"00000076000000000000004d000000000000005c000000000000005c00000000",
            INIT_11 => X"0000006200000000000000910000000000000099000000000000009c00000000",
            INIT_12 => X"0000007a000000000000007400000000000000aa000000000000005c00000000",
            INIT_13 => X"00000062000000000000004b000000000000008300000000000000a500000000",
            INIT_14 => X"0000004000000000000000550000000000000061000000000000004c00000000",
            INIT_15 => X"0000001b0000000000000011000000000000001b000000000000003600000000",
            INIT_16 => X"0000007500000000000000450000000000000028000000000000001a00000000",
            INIT_17 => X"0000002800000000000000240000000000000064000000000000007f00000000",
            INIT_18 => X"0000006e000000000000003c0000000000000054000000000000005e00000000",
            INIT_19 => X"00000073000000000000009b00000000000000a3000000000000009c00000000",
            INIT_1A => X"000000890000000000000094000000000000007c000000000000002700000000",
            INIT_1B => X"0000009c00000000000000570000000000000071000000000000009500000000",
            INIT_1C => X"00000027000000000000003d0000000000000050000000000000007800000000",
            INIT_1D => X"0000002e00000000000000220000000000000018000000000000002700000000",
            INIT_1E => X"000000780000000000000045000000000000002d000000000000001f00000000",
            INIT_1F => X"000000200000000000000022000000000000007b000000000000009900000000",
            INIT_20 => X"000000720000000000000059000000000000005d000000000000006100000000",
            INIT_21 => X"00000075000000000000009800000000000000a2000000000000009600000000",
            INIT_22 => X"000000740000000000000064000000000000001d000000000000000d00000000",
            INIT_23 => X"0000007c00000000000000490000000000000056000000000000007300000000",
            INIT_24 => X"0000001b000000000000002f000000000000005b000000000000008600000000",
            INIT_25 => X"0000003200000000000000310000000000000032000000000000003100000000",
            INIT_26 => X"0000007d0000000000000042000000000000001e000000000000001900000000",
            INIT_27 => X"000000200000000000000038000000000000009600000000000000a200000000",
            INIT_28 => X"0000006300000000000000570000000000000068000000000000006a00000000",
            INIT_29 => X"0000005700000000000000810000000000000096000000000000008d00000000",
            INIT_2A => X"000000250000000000000016000000000000000b000000000000000f00000000",
            INIT_2B => X"0000003e00000000000000290000000000000039000000000000003600000000",
            INIT_2C => X"0000001a00000000000000360000000000000048000000000000005300000000",
            INIT_2D => X"0000003300000000000000220000000000000023000000000000002000000000",
            INIT_2E => X"00000070000000000000003e000000000000002b000000000000002800000000",
            INIT_2F => X"0000001f000000000000004a000000000000009e000000000000009b00000000",
            INIT_30 => X"0000005a000000000000004f0000000000000068000000000000007000000000",
            INIT_31 => X"0000004200000000000000730000000000000089000000000000007b00000000",
            INIT_32 => X"0000001700000000000000280000000000000042000000000000002f00000000",
            INIT_33 => X"00000045000000000000002c0000000000000026000000000000001b00000000",
            INIT_34 => X"0000001d0000000000000026000000000000001f000000000000003600000000",
            INIT_35 => X"0000001f000000000000000f0000000000000016000000000000001900000000",
            INIT_36 => X"0000004e000000000000003a0000000000000033000000000000003100000000",
            INIT_37 => X"0000001f00000000000000570000000000000094000000000000008600000000",
            INIT_38 => X"0000006000000000000000590000000000000058000000000000006d00000000",
            INIT_39 => X"0000005e00000000000000730000000000000081000000000000006900000000",
            INIT_3A => X"0000003c00000000000000360000000000000047000000000000006100000000",
            INIT_3B => X"0000003c000000000000004b000000000000003e000000000000004200000000",
            INIT_3C => X"0000000e0000000000000009000000000000000a000000000000001a00000000",
            INIT_3D => X"0000000c000000000000000b0000000000000013000000000000001100000000",
            INIT_3E => X"0000003b000000000000003a000000000000001f000000000000001700000000",
            INIT_3F => X"0000002300000000000000690000000000000088000000000000005e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007000000000000000600000000000000046000000000000005b00000000",
            INIT_41 => X"0000009300000000000000890000000000000068000000000000006000000000",
            INIT_42 => X"000000430000000000000045000000000000003a000000000000007500000000",
            INIT_43 => X"00000035000000000000003f0000000000000045000000000000004a00000000",
            INIT_44 => X"0000000d00000000000000130000000000000019000000000000002900000000",
            INIT_45 => X"00000012000000000000000d0000000000000009000000000000000c00000000",
            INIT_46 => X"00000027000000000000003e0000000000000024000000000000000c00000000",
            INIT_47 => X"0000004700000000000000790000000000000068000000000000003400000000",
            INIT_48 => X"000000620000000000000062000000000000005c000000000000005b00000000",
            INIT_49 => X"0000008600000000000000690000000000000056000000000000006100000000",
            INIT_4A => X"00000061000000000000007c000000000000006b000000000000008e00000000",
            INIT_4B => X"00000049000000000000004e0000000000000049000000000000004400000000",
            INIT_4C => X"0000001c0000000000000026000000000000002b000000000000003e00000000",
            INIT_4D => X"00000014000000000000000b000000000000000e000000000000001600000000",
            INIT_4E => X"000000140000000000000030000000000000002a000000000000001400000000",
            INIT_4F => X"0000006400000000000000580000000000000038000000000000002500000000",
            INIT_50 => X"000000620000000000000061000000000000005e000000000000005b00000000",
            INIT_51 => X"0000004c000000000000005b000000000000006f000000000000007100000000",
            INIT_52 => X"000000510000000000000050000000000000006e000000000000008400000000",
            INIT_53 => X"000000540000000000000063000000000000005f000000000000004700000000",
            INIT_54 => X"000000330000000000000038000000000000003d000000000000004800000000",
            INIT_55 => X"0000002b0000000000000020000000000000002b000000000000003500000000",
            INIT_56 => X"0000002800000000000000250000000000000028000000000000002e00000000",
            INIT_57 => X"000000420000000000000030000000000000005a000000000000004000000000",
            INIT_58 => X"0000005200000000000000500000000000000060000000000000005700000000",
            INIT_59 => X"000000480000000000000062000000000000006d000000000000007100000000",
            INIT_5A => X"0000004600000000000000450000000000000073000000000000005c00000000",
            INIT_5B => X"000000580000000000000060000000000000005e000000000000004a00000000",
            INIT_5C => X"0000004a000000000000004c0000000000000047000000000000004500000000",
            INIT_5D => X"0000004b000000000000003d000000000000003c000000000000004200000000",
            INIT_5E => X"00000041000000000000003f0000000000000040000000000000004900000000",
            INIT_5F => X"0000003a0000000000000036000000000000005e000000000000004c00000000",
            INIT_60 => X"0000004c00000000000000430000000000000061000000000000006000000000",
            INIT_61 => X"00000050000000000000004e000000000000005a000000000000006900000000",
            INIT_62 => X"00000062000000000000004c0000000000000048000000000000005700000000",
            INIT_63 => X"0000005a000000000000005d000000000000005c000000000000005700000000",
            INIT_64 => X"0000004600000000000000550000000000000054000000000000004f00000000",
            INIT_65 => X"00000057000000000000004d0000000000000048000000000000004200000000",
            INIT_66 => X"0000004f00000000000000500000000000000052000000000000005300000000",
            INIT_67 => X"0000005e00000000000000460000000000000035000000000000004300000000",
            INIT_68 => X"0000006500000000000000510000000000000054000000000000004900000000",
            INIT_69 => X"0000005b0000000000000058000000000000005b000000000000006100000000",
            INIT_6A => X"00000063000000000000005b0000000000000059000000000000006900000000",
            INIT_6B => X"0000005a000000000000005d000000000000005d000000000000005900000000",
            INIT_6C => X"0000003c00000000000000490000000000000055000000000000005800000000",
            INIT_6D => X"0000005b00000000000000540000000000000052000000000000004900000000",
            INIT_6E => X"0000005500000000000000570000000000000056000000000000005d00000000",
            INIT_6F => X"0000006400000000000000570000000000000044000000000000004300000000",
            INIT_70 => X"00000071000000000000006a0000000000000060000000000000005300000000",
            INIT_71 => X"0000005f0000000000000060000000000000005f000000000000006000000000",
            INIT_72 => X"00000068000000000000006d0000000000000069000000000000006600000000",
            INIT_73 => X"0000004a0000000000000052000000000000005a000000000000005b00000000",
            INIT_74 => X"0000004a000000000000004d000000000000004e000000000000005200000000",
            INIT_75 => X"0000005c00000000000000570000000000000055000000000000004d00000000",
            INIT_76 => X"00000054000000000000005a0000000000000059000000000000006400000000",
            INIT_77 => X"0000005a0000000000000057000000000000004d000000000000004e00000000",
            INIT_78 => X"000000680000000000000071000000000000006b000000000000005c00000000",
            INIT_79 => X"0000005c000000000000004d0000000000000042000000000000005200000000",
            INIT_7A => X"0000005a000000000000005b0000000000000051000000000000005f00000000",
            INIT_7B => X"0000003d000000000000004d000000000000005b000000000000005800000000",
            INIT_7C => X"000000520000000000000056000000000000004d000000000000004600000000",
            INIT_7D => X"00000060000000000000005b000000000000005c000000000000005300000000",
            INIT_7E => X"0000005b0000000000000057000000000000005c000000000000006500000000",
            INIT_7F => X"00000057000000000000005b000000000000005a000000000000005c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE33;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE34 : if BRAM_NAME = "sampleifmap_layersamples_instance34" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000024000000000000001a000000000000003d000000000000005300000000",
            INIT_01 => X"00000036000000000000003a0000000000000043000000000000004100000000",
            INIT_02 => X"0000003b00000000000000340000000000000041000000000000003f00000000",
            INIT_03 => X"00000034000000000000002e0000000000000035000000000000003e00000000",
            INIT_04 => X"00000027000000000000002b0000000000000041000000000000004700000000",
            INIT_05 => X"00000026000000000000002d000000000000002f000000000000002f00000000",
            INIT_06 => X"00000032000000000000002a000000000000002d000000000000002f00000000",
            INIT_07 => X"000000290000000000000029000000000000002e000000000000004500000000",
            INIT_08 => X"00000046000000000000003a0000000000000035000000000000006100000000",
            INIT_09 => X"0000004d00000000000000440000000000000043000000000000004600000000",
            INIT_0A => X"0000003900000000000000380000000000000041000000000000004400000000",
            INIT_0B => X"0000002e00000000000000320000000000000039000000000000003400000000",
            INIT_0C => X"00000026000000000000002b0000000000000034000000000000003c00000000",
            INIT_0D => X"00000028000000000000002c000000000000002f000000000000002f00000000",
            INIT_0E => X"00000038000000000000002b000000000000001e000000000000002000000000",
            INIT_0F => X"0000003100000000000000330000000000000035000000000000004300000000",
            INIT_10 => X"00000051000000000000005c0000000000000047000000000000006400000000",
            INIT_11 => X"0000004e00000000000000440000000000000039000000000000004400000000",
            INIT_12 => X"0000003b000000000000003f0000000000000047000000000000004000000000",
            INIT_13 => X"0000003000000000000000310000000000000030000000000000003400000000",
            INIT_14 => X"0000001e00000000000000210000000000000032000000000000003b00000000",
            INIT_15 => X"0000003800000000000000350000000000000030000000000000002b00000000",
            INIT_16 => X"0000003800000000000000390000000000000038000000000000003300000000",
            INIT_17 => X"00000031000000000000002f0000000000000035000000000000003900000000",
            INIT_18 => X"000000590000000000000061000000000000005f000000000000006000000000",
            INIT_19 => X"0000004800000000000000490000000000000037000000000000004900000000",
            INIT_1A => X"000000420000000000000042000000000000004e000000000000004100000000",
            INIT_1B => X"0000003f00000000000000360000000000000037000000000000004300000000",
            INIT_1C => X"00000012000000000000001a000000000000002e000000000000002f00000000",
            INIT_1D => X"00000035000000000000002f0000000000000029000000000000002200000000",
            INIT_1E => X"0000003e00000000000000400000000000000044000000000000003d00000000",
            INIT_1F => X"0000003c000000000000003a000000000000002d000000000000003000000000",
            INIT_20 => X"0000005700000000000000540000000000000061000000000000005c00000000",
            INIT_21 => X"0000004b000000000000004c000000000000003f000000000000004900000000",
            INIT_22 => X"0000004b000000000000004b000000000000004a000000000000004a00000000",
            INIT_23 => X"0000003b0000000000000035000000000000003b000000000000004300000000",
            INIT_24 => X"0000001e00000000000000330000000000000034000000000000003b00000000",
            INIT_25 => X"00000027000000000000002e0000000000000029000000000000001f00000000",
            INIT_26 => X"0000003d000000000000003d000000000000003b000000000000002e00000000",
            INIT_27 => X"0000003c000000000000003a0000000000000030000000000000003400000000",
            INIT_28 => X"0000005900000000000000470000000000000066000000000000006500000000",
            INIT_29 => X"0000004c000000000000004c0000000000000046000000000000005100000000",
            INIT_2A => X"00000047000000000000004e0000000000000051000000000000004c00000000",
            INIT_2B => X"0000003100000000000000350000000000000043000000000000004400000000",
            INIT_2C => X"0000003900000000000000480000000000000041000000000000004300000000",
            INIT_2D => X"000000320000000000000042000000000000003e000000000000002b00000000",
            INIT_2E => X"0000003a00000000000000380000000000000036000000000000003800000000",
            INIT_2F => X"00000041000000000000003c000000000000003d000000000000003c00000000",
            INIT_30 => X"0000006300000000000000490000000000000059000000000000007800000000",
            INIT_31 => X"0000004b00000000000000510000000000000050000000000000005300000000",
            INIT_32 => X"0000004200000000000000550000000000000057000000000000005100000000",
            INIT_33 => X"000000350000000000000043000000000000004f000000000000004c00000000",
            INIT_34 => X"0000004d000000000000004a0000000000000040000000000000003c00000000",
            INIT_35 => X"0000002f00000000000000410000000000000040000000000000004100000000",
            INIT_36 => X"00000030000000000000002d0000000000000036000000000000003500000000",
            INIT_37 => X"00000042000000000000003f000000000000003d000000000000003a00000000",
            INIT_38 => X"0000005b000000000000005b000000000000003b000000000000007500000000",
            INIT_39 => X"00000054000000000000004f0000000000000051000000000000005100000000",
            INIT_3A => X"0000004800000000000000560000000000000056000000000000005700000000",
            INIT_3B => X"0000003f000000000000004a000000000000004c000000000000004d00000000",
            INIT_3C => X"00000049000000000000004c0000000000000049000000000000004200000000",
            INIT_3D => X"0000002f0000000000000038000000000000002f000000000000004700000000",
            INIT_3E => X"0000002a00000000000000230000000000000031000000000000002c00000000",
            INIT_3F => X"00000040000000000000003e0000000000000039000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000051000000000000005b0000000000000054000000000000005c00000000",
            INIT_41 => X"000000500000000000000050000000000000004f000000000000005300000000",
            INIT_42 => X"0000004600000000000000490000000000000053000000000000005800000000",
            INIT_43 => X"0000003d00000000000000430000000000000048000000000000005100000000",
            INIT_44 => X"0000004600000000000000460000000000000041000000000000004300000000",
            INIT_45 => X"0000003c000000000000004f0000000000000040000000000000004f00000000",
            INIT_46 => X"0000003b0000000000000034000000000000002d000000000000002c00000000",
            INIT_47 => X"00000040000000000000003d000000000000003d000000000000003a00000000",
            INIT_48 => X"0000005a000000000000004c0000000000000058000000000000006100000000",
            INIT_49 => X"0000004700000000000000530000000000000056000000000000005b00000000",
            INIT_4A => X"0000005300000000000000540000000000000052000000000000004f00000000",
            INIT_4B => X"00000055000000000000004d0000000000000053000000000000005800000000",
            INIT_4C => X"000000460000000000000039000000000000003e000000000000005100000000",
            INIT_4D => X"0000004b00000000000000590000000000000048000000000000005000000000",
            INIT_4E => X"0000003c000000000000003a0000000000000031000000000000002b00000000",
            INIT_4F => X"000000400000000000000039000000000000003f000000000000003a00000000",
            INIT_50 => X"0000006200000000000000560000000000000030000000000000005100000000",
            INIT_51 => X"000000540000000000000052000000000000005b000000000000005900000000",
            INIT_52 => X"0000005000000000000000500000000000000054000000000000005b00000000",
            INIT_53 => X"0000007e00000000000000670000000000000065000000000000005e00000000",
            INIT_54 => X"0000004300000000000000370000000000000049000000000000006b00000000",
            INIT_55 => X"000000440000000000000051000000000000004c000000000000004b00000000",
            INIT_56 => X"0000002d000000000000002f0000000000000031000000000000002000000000",
            INIT_57 => X"00000041000000000000003e000000000000003a000000000000003300000000",
            INIT_58 => X"0000004d0000000000000063000000000000001f000000000000001400000000",
            INIT_59 => X"0000005a000000000000005a0000000000000056000000000000004000000000",
            INIT_5A => X"0000005f00000000000000450000000000000045000000000000005f00000000",
            INIT_5B => X"0000007900000000000000670000000000000088000000000000008f00000000",
            INIT_5C => X"00000050000000000000003f0000000000000052000000000000007600000000",
            INIT_5D => X"000000210000000000000042000000000000004d000000000000005200000000",
            INIT_5E => X"0000002e00000000000000300000000000000030000000000000002100000000",
            INIT_5F => X"0000003f000000000000003b0000000000000036000000000000003000000000",
            INIT_60 => X"0000005c00000000000000700000000000000032000000000000000000000000",
            INIT_61 => X"000000620000000000000069000000000000007a000000000000006e00000000",
            INIT_62 => X"0000007700000000000000540000000000000048000000000000006000000000",
            INIT_63 => X"00000049000000000000005f000000000000007d000000000000009d00000000",
            INIT_64 => X"0000005400000000000000410000000000000047000000000000003400000000",
            INIT_65 => X"0000002a0000000000000041000000000000004f000000000000006000000000",
            INIT_66 => X"0000002900000000000000290000000000000025000000000000002500000000",
            INIT_67 => X"0000003a00000000000000390000000000000038000000000000002d00000000",
            INIT_68 => X"0000005c0000000000000061000000000000003c000000000000001400000000",
            INIT_69 => X"0000006f00000000000000700000000000000078000000000000007d00000000",
            INIT_6A => X"00000080000000000000006e000000000000004c000000000000005900000000",
            INIT_6B => X"0000006c00000000000000620000000000000064000000000000007f00000000",
            INIT_6C => X"0000005b00000000000000620000000000000063000000000000004400000000",
            INIT_6D => X"00000029000000000000003a000000000000004c000000000000006a00000000",
            INIT_6E => X"0000002600000000000000250000000000000023000000000000002100000000",
            INIT_6F => X"0000003500000000000000320000000000000034000000000000002e00000000",
            INIT_70 => X"00000058000000000000003a0000000000000046000000000000003b00000000",
            INIT_71 => X"00000073000000000000006a0000000000000075000000000000007b00000000",
            INIT_72 => X"0000007d00000000000000820000000000000067000000000000006600000000",
            INIT_73 => X"0000008900000000000000660000000000000050000000000000005f00000000",
            INIT_74 => X"00000084000000000000007e000000000000008c000000000000008300000000",
            INIT_75 => X"0000002a0000000000000040000000000000004e000000000000006f00000000",
            INIT_76 => X"00000032000000000000002a0000000000000028000000000000002b00000000",
            INIT_77 => X"00000031000000000000002e0000000000000032000000000000002f00000000",
            INIT_78 => X"0000005e00000000000000320000000000000035000000000000004900000000",
            INIT_79 => X"00000062000000000000006c000000000000007c000000000000007e00000000",
            INIT_7A => X"00000088000000000000008a000000000000007d000000000000007200000000",
            INIT_7B => X"0000008c00000000000000710000000000000062000000000000007b00000000",
            INIT_7C => X"0000008c000000000000008a0000000000000089000000000000008f00000000",
            INIT_7D => X"0000003300000000000000490000000000000069000000000000007500000000",
            INIT_7E => X"0000004d00000000000000320000000000000023000000000000002f00000000",
            INIT_7F => X"00000032000000000000002d000000000000002d000000000000004300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE34;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE35 : if BRAM_NAME = "sampleifmap_layersamples_instance35" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000056000000000000003a0000000000000041000000000000004800000000",
            INIT_01 => X"0000005300000000000000690000000000000075000000000000007700000000",
            INIT_02 => X"0000008200000000000000930000000000000089000000000000006e00000000",
            INIT_03 => X"00000087000000000000006d000000000000006b000000000000008200000000",
            INIT_04 => X"00000083000000000000007e000000000000007f000000000000008400000000",
            INIT_05 => X"0000002a000000000000003d0000000000000077000000000000008700000000",
            INIT_06 => X"00000055000000000000003c000000000000001b000000000000001a00000000",
            INIT_07 => X"0000003300000000000000240000000000000033000000000000006100000000",
            INIT_08 => X"0000006600000000000000510000000000000048000000000000004700000000",
            INIT_09 => X"00000050000000000000007a000000000000007c000000000000007800000000",
            INIT_0A => X"00000054000000000000006a0000000000000097000000000000006300000000",
            INIT_0B => X"0000005c00000000000000650000000000000079000000000000007c00000000",
            INIT_0C => X"0000006500000000000000680000000000000073000000000000006300000000",
            INIT_0D => X"00000011000000000000001f0000000000000048000000000000005e00000000",
            INIT_0E => X"00000055000000000000003a0000000000000015000000000000000e00000000",
            INIT_0F => X"00000029000000000000001f0000000000000046000000000000006800000000",
            INIT_10 => X"000000640000000000000044000000000000004e000000000000004f00000000",
            INIT_11 => X"0000004b000000000000007d0000000000000088000000000000008600000000",
            INIT_12 => X"00000061000000000000005b0000000000000093000000000000004700000000",
            INIT_13 => X"0000004800000000000000370000000000000071000000000000008e00000000",
            INIT_14 => X"000000320000000000000045000000000000004f000000000000003500000000",
            INIT_15 => X"00000016000000000000000d0000000000000014000000000000002a00000000",
            INIT_16 => X"0000006000000000000000370000000000000023000000000000001400000000",
            INIT_17 => X"00000023000000000000001e000000000000005b000000000000006f00000000",
            INIT_18 => X"0000005800000000000000320000000000000048000000000000005100000000",
            INIT_19 => X"0000005d000000000000008a0000000000000099000000000000008700000000",
            INIT_1A => X"00000071000000000000007f000000000000006f000000000000001f00000000",
            INIT_1B => X"0000008d0000000000000047000000000000005c000000000000007c00000000",
            INIT_1C => X"0000002100000000000000330000000000000041000000000000006700000000",
            INIT_1D => X"0000002c00000000000000240000000000000019000000000000002400000000",
            INIT_1E => X"000000600000000000000036000000000000002b000000000000001a00000000",
            INIT_1F => X"0000001a000000000000001e0000000000000073000000000000008900000000",
            INIT_20 => X"0000005f000000000000004f0000000000000052000000000000005300000000",
            INIT_21 => X"0000006200000000000000860000000000000096000000000000008200000000",
            INIT_22 => X"0000006300000000000000560000000000000017000000000000000a00000000",
            INIT_23 => X"000000740000000000000042000000000000004c000000000000006500000000",
            INIT_24 => X"000000170000000000000027000000000000004e000000000000007a00000000",
            INIT_25 => X"0000002e000000000000002f000000000000002f000000000000002e00000000",
            INIT_26 => X"000000670000000000000034000000000000001b000000000000001400000000",
            INIT_27 => X"00000019000000000000002f0000000000000089000000000000009200000000",
            INIT_28 => X"00000053000000000000004e000000000000005c000000000000005c00000000",
            INIT_29 => X"00000046000000000000006e0000000000000087000000000000007b00000000",
            INIT_2A => X"0000001d00000000000000100000000000000008000000000000000c00000000",
            INIT_2B => X"0000003800000000000000250000000000000034000000000000002f00000000",
            INIT_2C => X"00000012000000000000002b0000000000000039000000000000004600000000",
            INIT_2D => X"0000002c000000000000001d000000000000001c000000000000001900000000",
            INIT_2E => X"0000005e00000000000000310000000000000026000000000000002100000000",
            INIT_2F => X"00000018000000000000003d000000000000008d000000000000008c00000000",
            INIT_30 => X"0000004e0000000000000046000000000000005d000000000000006100000000",
            INIT_31 => X"0000003000000000000000600000000000000076000000000000006b00000000",
            INIT_32 => X"000000130000000000000022000000000000003a000000000000002500000000",
            INIT_33 => X"0000003b0000000000000026000000000000001f000000000000001300000000",
            INIT_34 => X"00000012000000000000001b0000000000000013000000000000002700000000",
            INIT_35 => X"00000018000000000000000a0000000000000011000000000000001100000000",
            INIT_36 => X"000000400000000000000030000000000000002c000000000000002a00000000",
            INIT_37 => X"0000001800000000000000460000000000000080000000000000007800000000",
            INIT_38 => X"000000580000000000000052000000000000004d000000000000005e00000000",
            INIT_39 => X"0000004b000000000000005f000000000000006b000000000000005b00000000",
            INIT_3A => X"0000003900000000000000300000000000000037000000000000004a00000000",
            INIT_3B => X"0000003300000000000000430000000000000035000000000000003a00000000",
            INIT_3C => X"0000000800000000000000030000000000000004000000000000001000000000",
            INIT_3D => X"0000000600000000000000070000000000000013000000000000000e00000000",
            INIT_3E => X"0000002f00000000000000300000000000000017000000000000001100000000",
            INIT_3F => X"0000001b00000000000000570000000000000073000000000000005100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000690000000000000057000000000000003b000000000000004b00000000",
            INIT_41 => X"0000007e00000000000000750000000000000052000000000000005300000000",
            INIT_42 => X"0000003e00000000000000390000000000000022000000000000005500000000",
            INIT_43 => X"0000002e0000000000000039000000000000003d000000000000004200000000",
            INIT_44 => X"0000000d00000000000000120000000000000017000000000000002400000000",
            INIT_45 => X"0000000e000000000000000c000000000000000e000000000000000f00000000",
            INIT_46 => X"0000001e0000000000000036000000000000001c000000000000000700000000",
            INIT_47 => X"0000003e00000000000000680000000000000055000000000000002800000000",
            INIT_48 => X"000000560000000000000051000000000000004d000000000000004d00000000",
            INIT_49 => X"0000007000000000000000570000000000000045000000000000005500000000",
            INIT_4A => X"0000004f0000000000000064000000000000004f000000000000006f00000000",
            INIT_4B => X"0000003a00000000000000450000000000000043000000000000003b00000000",
            INIT_4C => X"0000001500000000000000200000000000000026000000000000003300000000",
            INIT_4D => X"0000000e0000000000000006000000000000000c000000000000001100000000",
            INIT_4E => X"0000000f00000000000000290000000000000022000000000000000f00000000",
            INIT_4F => X"0000005a000000000000004c000000000000002e000000000000001f00000000",
            INIT_50 => X"0000005500000000000000520000000000000051000000000000004f00000000",
            INIT_51 => X"00000039000000000000004a0000000000000060000000000000006500000000",
            INIT_52 => X"0000003e000000000000003a0000000000000057000000000000006d00000000",
            INIT_53 => X"00000044000000000000005a0000000000000058000000000000003d00000000",
            INIT_54 => X"0000002a000000000000002f0000000000000035000000000000003b00000000",
            INIT_55 => X"0000002300000000000000180000000000000023000000000000002c00000000",
            INIT_56 => X"0000001f000000000000001b000000000000001d000000000000002600000000",
            INIT_57 => X"0000003800000000000000270000000000000052000000000000003900000000",
            INIT_58 => X"0000004a000000000000004a0000000000000057000000000000004c00000000",
            INIT_59 => X"000000390000000000000053000000000000005f000000000000006600000000",
            INIT_5A => X"0000003a00000000000000370000000000000063000000000000004d00000000",
            INIT_5B => X"0000004d00000000000000570000000000000054000000000000003f00000000",
            INIT_5C => X"000000440000000000000043000000000000003c000000000000003900000000",
            INIT_5D => X"0000003f00000000000000310000000000000031000000000000003b00000000",
            INIT_5E => X"0000003300000000000000300000000000000031000000000000003c00000000",
            INIT_5F => X"0000002f000000000000002d0000000000000054000000000000003f00000000",
            INIT_60 => X"000000450000000000000040000000000000005a000000000000005500000000",
            INIT_61 => X"000000440000000000000041000000000000004e000000000000005e00000000",
            INIT_62 => X"0000005a0000000000000042000000000000003c000000000000004c00000000",
            INIT_63 => X"000000510000000000000053000000000000004e000000000000004a00000000",
            INIT_64 => X"00000040000000000000004c0000000000000047000000000000004300000000",
            INIT_65 => X"00000048000000000000003e0000000000000039000000000000003b00000000",
            INIT_66 => X"0000003e00000000000000400000000000000042000000000000004400000000",
            INIT_67 => X"00000053000000000000003d0000000000000029000000000000003200000000",
            INIT_68 => X"0000005c0000000000000049000000000000004b000000000000003d00000000",
            INIT_69 => X"00000050000000000000004e0000000000000051000000000000005700000000",
            INIT_6A => X"000000590000000000000050000000000000004c000000000000005d00000000",
            INIT_6B => X"00000050000000000000004e000000000000004c000000000000004a00000000",
            INIT_6C => X"00000035000000000000003e0000000000000045000000000000004a00000000",
            INIT_6D => X"0000004b00000000000000440000000000000042000000000000004000000000",
            INIT_6E => X"0000004400000000000000480000000000000048000000000000004d00000000",
            INIT_6F => X"00000059000000000000004e0000000000000038000000000000003200000000",
            INIT_70 => X"00000064000000000000005a0000000000000051000000000000004600000000",
            INIT_71 => X"0000005500000000000000570000000000000055000000000000005600000000",
            INIT_72 => X"0000005a000000000000005d0000000000000057000000000000005600000000",
            INIT_73 => X"0000003c000000000000003f0000000000000046000000000000004a00000000",
            INIT_74 => X"0000003e000000000000003e000000000000003c000000000000004200000000",
            INIT_75 => X"0000004c00000000000000470000000000000046000000000000004100000000",
            INIT_76 => X"00000047000000000000004e000000000000004d000000000000005500000000",
            INIT_77 => X"0000004f000000000000004d0000000000000041000000000000003e00000000",
            INIT_78 => X"00000059000000000000005f000000000000005d000000000000004f00000000",
            INIT_79 => X"0000005100000000000000460000000000000039000000000000004600000000",
            INIT_7A => X"0000004700000000000000470000000000000040000000000000005300000000",
            INIT_7B => X"0000002f000000000000003d000000000000004c000000000000004a00000000",
            INIT_7C => X"000000460000000000000048000000000000003f000000000000003800000000",
            INIT_7D => X"00000050000000000000004b000000000000004c000000000000004500000000",
            INIT_7E => X"0000004e0000000000000049000000000000004f000000000000005600000000",
            INIT_7F => X"00000049000000000000004f000000000000004c000000000000004f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE35;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE36 : if BRAM_NAME = "sampleifmap_layersamples_instance36" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d900000000000000d100000000000000b900000000000000a000000000",
            INIT_01 => X"000000f600000000000000f900000000000000f600000000000000e600000000",
            INIT_02 => X"000000dd00000000000000e600000000000000f300000000000000f800000000",
            INIT_03 => X"000000c700000000000000d800000000000000dd00000000000000da00000000",
            INIT_04 => X"000000b400000000000000b800000000000000bb00000000000000bc00000000",
            INIT_05 => X"0000008b0000000000000079000000000000009000000000000000a600000000",
            INIT_06 => X"0000004f00000000000000660000000000000066000000000000006a00000000",
            INIT_07 => X"0000005e000000000000005b0000000000000065000000000000005e00000000",
            INIT_08 => X"000000e600000000000000f200000000000000ef00000000000000e100000000",
            INIT_09 => X"000000eb00000000000000f300000000000000f500000000000000e800000000",
            INIT_0A => X"000000cd00000000000000d800000000000000e600000000000000ed00000000",
            INIT_0B => X"000000ba00000000000000c800000000000000cb00000000000000c900000000",
            INIT_0C => X"0000007f00000000000000a100000000000000ab00000000000000af00000000",
            INIT_0D => X"00000087000000000000007a000000000000008d000000000000008e00000000",
            INIT_0E => X"0000003400000000000000250000000000000052000000000000007600000000",
            INIT_0F => X"000000640000000000000061000000000000006b000000000000005f00000000",
            INIT_10 => X"000000dc00000000000000f100000000000000f900000000000000fc00000000",
            INIT_11 => X"000000d600000000000000df00000000000000e200000000000000d900000000",
            INIT_12 => X"000000b800000000000000c300000000000000cf00000000000000d500000000",
            INIT_13 => X"000000a700000000000000b300000000000000b600000000000000b300000000",
            INIT_14 => X"0000008100000000000000940000000000000098000000000000009f00000000",
            INIT_15 => X"000000720000000000000080000000000000008c000000000000008000000000",
            INIT_16 => X"0000002600000000000000040000000000000028000000000000005700000000",
            INIT_17 => X"0000006900000000000000690000000000000073000000000000006300000000",
            INIT_18 => X"000000d300000000000000de00000000000000e100000000000000e900000000",
            INIT_19 => X"000000c000000000000000c800000000000000cb00000000000000d300000000",
            INIT_1A => X"000000a400000000000000ae00000000000000b700000000000000bb00000000",
            INIT_1B => X"0000009900000000000000a000000000000000a500000000000000a000000000",
            INIT_1C => X"0000008a000000000000008c000000000000008d000000000000009100000000",
            INIT_1D => X"00000069000000000000007f000000000000007d000000000000007d00000000",
            INIT_1E => X"00000037000000000000001a0000000000000025000000000000003b00000000",
            INIT_1F => X"0000006d00000000000000700000000000000078000000000000007000000000",
            INIT_20 => X"000000c900000000000000cf00000000000000c300000000000000cf00000000",
            INIT_21 => X"000000ab00000000000000b300000000000000b400000000000000be00000000",
            INIT_22 => X"000000920000000000000099000000000000009f00000000000000a300000000",
            INIT_23 => X"0000008d00000000000000930000000000000097000000000000009100000000",
            INIT_24 => X"0000008700000000000000830000000000000088000000000000008700000000",
            INIT_25 => X"0000005a0000000000000084000000000000007a000000000000008100000000",
            INIT_26 => X"000000560000000000000030000000000000003d000000000000003a00000000",
            INIT_27 => X"0000006d00000000000000720000000000000078000000000000007500000000",
            INIT_28 => X"000000a200000000000000aa00000000000000ab00000000000000b600000000",
            INIT_29 => X"00000097000000000000009f000000000000009c000000000000009900000000",
            INIT_2A => X"0000008a000000000000008c000000000000008d000000000000009000000000",
            INIT_2B => X"0000008a000000000000008a000000000000008d000000000000008b00000000",
            INIT_2C => X"0000008a0000000000000086000000000000008c000000000000008700000000",
            INIT_2D => X"0000004500000000000000660000000000000089000000000000008c00000000",
            INIT_2E => X"000000740000000000000043000000000000003e000000000000004b00000000",
            INIT_2F => X"0000006e00000000000000700000000000000080000000000000008100000000",
            INIT_30 => X"0000008600000000000000880000000000000088000000000000008d00000000",
            INIT_31 => X"00000085000000000000008c0000000000000086000000000000008800000000",
            INIT_32 => X"0000008d000000000000008b0000000000000089000000000000008700000000",
            INIT_33 => X"00000091000000000000008e0000000000000092000000000000008f00000000",
            INIT_34 => X"0000008f000000000000008a0000000000000091000000000000009100000000",
            INIT_35 => X"00000021000000000000002f000000000000006b000000000000008e00000000",
            INIT_36 => X"0000007f000000000000006c000000000000004b000000000000004800000000",
            INIT_37 => X"00000070000000000000006f0000000000000084000000000000008400000000",
            INIT_38 => X"000000810000000000000080000000000000007d000000000000007600000000",
            INIT_39 => X"00000084000000000000008a0000000000000083000000000000008800000000",
            INIT_3A => X"000000930000000000000090000000000000008c000000000000008800000000",
            INIT_3B => X"00000099000000000000009a000000000000009e000000000000009600000000",
            INIT_3C => X"0000009400000000000000930000000000000095000000000000009200000000",
            INIT_3D => X"00000011000000000000000d0000000000000042000000000000008000000000",
            INIT_3E => X"0000007a00000000000000800000000000000075000000000000005000000000",
            INIT_3F => X"0000007000000000000000720000000000000080000000000000007b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000850000000000000084000000000000007e000000000000007300000000",
            INIT_41 => X"00000089000000000000008f0000000000000087000000000000008b00000000",
            INIT_42 => X"0000009800000000000000950000000000000091000000000000008b00000000",
            INIT_43 => X"000000aa00000000000000a3000000000000009a000000000000009400000000",
            INIT_44 => X"00000094000000000000009d00000000000000a2000000000000009e00000000",
            INIT_45 => X"0000001e000000000000000e000000000000002c000000000000007300000000",
            INIT_46 => X"0000007e0000000000000088000000000000008b000000000000006900000000",
            INIT_47 => X"0000006f0000000000000074000000000000007a000000000000007700000000",
            INIT_48 => X"0000008800000000000000880000000000000080000000000000007600000000",
            INIT_49 => X"0000008d00000000000000910000000000000088000000000000008d00000000",
            INIT_4A => X"000000a5000000000000009a0000000000000093000000000000008d00000000",
            INIT_4B => X"000000a700000000000000a2000000000000009a000000000000009d00000000",
            INIT_4C => X"0000008a00000000000000910000000000000093000000000000009b00000000",
            INIT_4D => X"00000037000000000000002e0000000000000038000000000000006300000000",
            INIT_4E => X"0000007e000000000000007a000000000000007c000000000000006d00000000",
            INIT_4F => X"0000006e00000000000000750000000000000074000000000000007300000000",
            INIT_50 => X"00000089000000000000008b0000000000000084000000000000007d00000000",
            INIT_51 => X"0000008c00000000000000900000000000000088000000000000008e00000000",
            INIT_52 => X"0000009900000000000000960000000000000090000000000000008b00000000",
            INIT_53 => X"000000980000000000000090000000000000008b000000000000008300000000",
            INIT_54 => X"000000d600000000000000d300000000000000ba00000000000000a600000000",
            INIT_55 => X"0000002a0000000000000045000000000000005c000000000000008000000000",
            INIT_56 => X"000000730000000000000063000000000000005f000000000000005500000000",
            INIT_57 => X"0000006b0000000000000071000000000000006f000000000000007000000000",
            INIT_58 => X"0000008a000000000000008e0000000000000089000000000000008500000000",
            INIT_59 => X"0000008a000000000000008e0000000000000088000000000000008d00000000",
            INIT_5A => X"000000840000000000000088000000000000008f000000000000008900000000",
            INIT_5B => X"000000cb00000000000000c900000000000000b6000000000000008e00000000",
            INIT_5C => X"000000c000000000000000cf00000000000000ce00000000000000d200000000",
            INIT_5D => X"0000002a000000000000009200000000000000bd00000000000000a200000000",
            INIT_5E => X"0000007200000000000000670000000000000028000000000000001b00000000",
            INIT_5F => X"00000068000000000000006c000000000000006a000000000000006d00000000",
            INIT_60 => X"0000008b000000000000008f000000000000008b000000000000008c00000000",
            INIT_61 => X"00000089000000000000008a000000000000008c000000000000008f00000000",
            INIT_62 => X"000000a400000000000000900000000000000085000000000000008700000000",
            INIT_63 => X"00000073000000000000008900000000000000a000000000000000ab00000000",
            INIT_64 => X"0000003b000000000000004b000000000000005d000000000000006a00000000",
            INIT_65 => X"0000005f00000000000000c900000000000000dc000000000000006f00000000",
            INIT_66 => X"00000074000000000000003e0000000000000007000000000000000d00000000",
            INIT_67 => X"0000006400000000000000690000000000000065000000000000006300000000",
            INIT_68 => X"0000008c000000000000008f000000000000008a000000000000009000000000",
            INIT_69 => X"0000008700000000000000820000000000000092000000000000009200000000",
            INIT_6A => X"0000006e000000000000008c0000000000000091000000000000008200000000",
            INIT_6B => X"000000130000000000000031000000000000005c000000000000005e00000000",
            INIT_6C => X"0000001200000000000000190000000000000032000000000000001d00000000",
            INIT_6D => X"0000009d00000000000000d200000000000000d1000000000000007800000000",
            INIT_6E => X"0000004400000000000000130000000000000006000000000000002600000000",
            INIT_6F => X"0000005f00000000000000630000000000000052000000000000004500000000",
            INIT_70 => X"0000008e0000000000000092000000000000008b000000000000009100000000",
            INIT_71 => X"000000800000000000000079000000000000008e000000000000009000000000",
            INIT_72 => X"000000440000000000000054000000000000007f000000000000008500000000",
            INIT_73 => X"00000016000000000000002e0000000000000052000000000000005600000000",
            INIT_74 => X"00000041000000000000001e0000000000000032000000000000001300000000",
            INIT_75 => X"000000cb00000000000000cd00000000000000c900000000000000af00000000",
            INIT_76 => X"0000001600000000000000120000000000000010000000000000006600000000",
            INIT_77 => X"00000058000000000000004f0000000000000038000000000000002300000000",
            INIT_78 => X"000000900000000000000094000000000000008b000000000000008f00000000",
            INIT_79 => X"00000083000000000000008b0000000000000084000000000000008a00000000",
            INIT_7A => X"0000005600000000000000480000000000000042000000000000007500000000",
            INIT_7B => X"000000220000000000000028000000000000004e000000000000006a00000000",
            INIT_7C => X"000000b600000000000000730000000000000046000000000000002400000000",
            INIT_7D => X"000000c300000000000000cd00000000000000c500000000000000cb00000000",
            INIT_7E => X"000000120000000000000025000000000000003d000000000000006c00000000",
            INIT_7F => X"000000530000000000000064000000000000004f000000000000001800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE36;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE37 : if BRAM_NAME = "sampleifmap_layersamples_instance37" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000900000000000000093000000000000008b000000000000008e00000000",
            INIT_01 => X"0000007900000000000000840000000000000072000000000000008500000000",
            INIT_02 => X"00000045000000000000003c0000000000000059000000000000005100000000",
            INIT_03 => X"0000009b00000000000000530000000000000044000000000000005500000000",
            INIT_04 => X"000000eb00000000000000ed00000000000000db00000000000000c000000000",
            INIT_05 => X"0000007200000000000000d300000000000000d700000000000000d700000000",
            INIT_06 => X"000000140000000000000035000000000000005d000000000000003000000000",
            INIT_07 => X"00000054000000000000008f000000000000008b000000000000004100000000",
            INIT_08 => X"00000089000000000000008e000000000000008d000000000000008f00000000",
            INIT_09 => X"00000043000000000000003a0000000000000045000000000000007400000000",
            INIT_0A => X"0000001c000000000000001d000000000000004b000000000000005100000000",
            INIT_0B => X"000000f2000000000000008c0000000000000019000000000000002400000000",
            INIT_0C => X"000000dc00000000000000e300000000000000eb00000000000000ec00000000",
            INIT_0D => X"0000003a000000000000009500000000000000df00000000000000db00000000",
            INIT_0E => X"0000004e000000000000004e0000000000000054000000000000003900000000",
            INIT_0F => X"0000005b00000000000000a700000000000000a1000000000000008500000000",
            INIT_10 => X"000000860000000000000088000000000000008c000000000000008f00000000",
            INIT_11 => X"00000034000000000000002d0000000000000047000000000000008d00000000",
            INIT_12 => X"0000001600000000000000170000000000000021000000000000004300000000",
            INIT_13 => X"000000d9000000000000009b0000000000000029000000000000002f00000000",
            INIT_14 => X"000000d000000000000000bf00000000000000be00000000000000c700000000",
            INIT_15 => X"0000006700000000000000ad00000000000000df00000000000000dc00000000",
            INIT_16 => X"0000009500000000000000870000000000000073000000000000005d00000000",
            INIT_17 => X"0000005900000000000000a50000000000000094000000000000009800000000",
            INIT_18 => X"000000b5000000000000007e000000000000008c000000000000008f00000000",
            INIT_19 => X"0000002b0000000000000021000000000000004c00000000000000bd00000000",
            INIT_1A => X"0000001700000000000000100000000000000015000000000000003900000000",
            INIT_1B => X"000000c2000000000000009e0000000000000042000000000000003900000000",
            INIT_1C => X"000000c900000000000000c400000000000000b300000000000000b600000000",
            INIT_1D => X"000000b300000000000000de00000000000000ce00000000000000c200000000",
            INIT_1E => X"000000970000000000000095000000000000009c000000000000009700000000",
            INIT_1F => X"0000004200000000000000880000000000000092000000000000009600000000",
            INIT_20 => X"000000ea000000000000009a0000000000000085000000000000008c00000000",
            INIT_21 => X"0000002a0000000000000026000000000000005a00000000000000b500000000",
            INIT_22 => X"0000000b000000000000000b000000000000000b000000000000003400000000",
            INIT_23 => X"000000ba00000000000000a00000000000000031000000000000001400000000",
            INIT_24 => X"0000007300000000000000b900000000000000b900000000000000b000000000",
            INIT_25 => X"000000c400000000000000a1000000000000005a000000000000004500000000",
            INIT_26 => X"0000009900000000000000a000000000000000aa00000000000000b700000000",
            INIT_27 => X"00000026000000000000004d0000000000000088000000000000009300000000",
            INIT_28 => X"000000a300000000000000a30000000000000080000000000000008200000000",
            INIT_29 => X"0000002e000000000000002d000000000000006a000000000000008b00000000",
            INIT_2A => X"0000000f00000000000000090000000000000003000000000000001c00000000",
            INIT_2B => X"000000b400000000000000a20000000000000036000000000000001e00000000",
            INIT_2C => X"00000015000000000000007100000000000000be00000000000000ac00000000",
            INIT_2D => X"0000009500000000000000300000000000000015000000000000001400000000",
            INIT_2E => X"00000085000000000000008e00000000000000ab00000000000000bb00000000",
            INIT_2F => X"0000002700000000000000150000000000000043000000000000008000000000",
            INIT_30 => X"0000001a00000000000000670000000000000084000000000000007c00000000",
            INIT_31 => X"000000300000000000000034000000000000006c000000000000004800000000",
            INIT_32 => X"0000003b000000000000000b0000000000000007000000000000001200000000",
            INIT_33 => X"000000b000000000000000a50000000000000063000000000000005a00000000",
            INIT_34 => X"0000001d000000000000002a00000000000000a900000000000000b100000000",
            INIT_35 => X"00000046000000000000000e0000000000000026000000000000002f00000000",
            INIT_36 => X"0000007500000000000000750000000000000088000000000000009500000000",
            INIT_37 => X"000000300000000000000015000000000000000e000000000000003c00000000",
            INIT_38 => X"0000001e0000000000000049000000000000007c000000000000007900000000",
            INIT_39 => X"0000001f00000000000000440000000000000072000000000000003b00000000",
            INIT_3A => X"000000480000000000000018000000000000000e000000000000000d00000000",
            INIT_3B => X"000000bb00000000000000bb000000000000006c000000000000004f00000000",
            INIT_3C => X"0000002b000000000000001b000000000000008b00000000000000bf00000000",
            INIT_3D => X"0000001b000000000000001c000000000000001b000000000000001e00000000",
            INIT_3E => X"00000059000000000000007b0000000000000084000000000000006c00000000",
            INIT_3F => X"0000003b000000000000002a0000000000000015000000000000001600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003f00000000000000470000000000000066000000000000006d00000000",
            INIT_41 => X"0000001c000000000000004d0000000000000071000000000000003c00000000",
            INIT_42 => X"000000470000000000000030000000000000001f000000000000001000000000",
            INIT_43 => X"000000b300000000000000bd0000000000000088000000000000004600000000",
            INIT_44 => X"00000036000000000000001f000000000000007400000000000000b400000000",
            INIT_45 => X"0000000e000000000000001b0000000000000029000000000000003500000000",
            INIT_46 => X"0000003c000000000000007c0000000000000085000000000000004800000000",
            INIT_47 => X"0000003b00000000000000320000000000000022000000000000001200000000",
            INIT_48 => X"0000003c000000000000003d0000000000000051000000000000005700000000",
            INIT_49 => X"00000015000000000000004b0000000000000069000000000000003a00000000",
            INIT_4A => X"00000060000000000000004c000000000000002e000000000000001400000000",
            INIT_4B => X"000000a300000000000000a40000000000000091000000000000006100000000",
            INIT_4C => X"000000390000000000000020000000000000007100000000000000aa00000000",
            INIT_4D => X"0000001100000000000000250000000000000031000000000000004700000000",
            INIT_4E => X"000000210000000000000060000000000000006c000000000000002900000000",
            INIT_4F => X"000000320000000000000028000000000000001d000000000000000c00000000",
            INIT_50 => X"0000003c00000000000000400000000000000049000000000000004900000000",
            INIT_51 => X"0000002f0000000000000057000000000000005f000000000000003900000000",
            INIT_52 => X"000000a500000000000000890000000000000062000000000000003d00000000",
            INIT_53 => X"000000b600000000000000b700000000000000b000000000000000a900000000",
            INIT_54 => X"000000360000000000000022000000000000007c00000000000000b600000000",
            INIT_55 => X"0000001b0000000000000033000000000000005c000000000000006000000000",
            INIT_56 => X"0000000c000000000000003b0000000000000046000000000000001100000000",
            INIT_57 => X"00000028000000000000001d0000000000000012000000000000000600000000",
            INIT_58 => X"0000004e00000000000000450000000000000049000000000000004900000000",
            INIT_59 => X"0000002f00000000000000450000000000000059000000000000004100000000",
            INIT_5A => X"00000056000000000000004a000000000000003c000000000000003400000000",
            INIT_5B => X"0000006000000000000000620000000000000060000000000000005b00000000",
            INIT_5C => X"0000003c00000000000000200000000000000053000000000000006200000000",
            INIT_5D => X"00000014000000000000001d000000000000003e000000000000003b00000000",
            INIT_5E => X"00000003000000000000000a0000000000000011000000000000000400000000",
            INIT_5F => X"000000210000000000000011000000000000000a000000000000000700000000",
            INIT_60 => X"0000003600000000000000480000000000000053000000000000004b00000000",
            INIT_61 => X"00000004000000000000000f0000000000000027000000000000002d00000000",
            INIT_62 => X"0000000700000000000000050000000000000002000000000000000300000000",
            INIT_63 => X"0000000b000000000000000a0000000000000008000000000000000700000000",
            INIT_64 => X"000000420000000000000008000000000000000d000000000000000b00000000",
            INIT_65 => X"0000000f0000000000000038000000000000002f000000000000004300000000",
            INIT_66 => X"0000000300000000000000010000000000000002000000000000000200000000",
            INIT_67 => X"00000020000000000000000f000000000000000a000000000000000600000000",
            INIT_68 => X"0000002f00000000000000510000000000000059000000000000005000000000",
            INIT_69 => X"000000190000000000000010000000000000000a000000000000001500000000",
            INIT_6A => X"0000000e000000000000000e000000000000000a000000000000000e00000000",
            INIT_6B => X"0000000c000000000000000e000000000000000e000000000000000e00000000",
            INIT_6C => X"0000001700000000000000060000000000000009000000000000000a00000000",
            INIT_6D => X"00000007000000000000002a0000000000000048000000000000003e00000000",
            INIT_6E => X"0000000500000000000000050000000000000004000000000000000300000000",
            INIT_6F => X"000000210000000000000015000000000000000b000000000000000700000000",
            INIT_70 => X"000000370000000000000049000000000000004f000000000000004900000000",
            INIT_71 => X"0000003a000000000000003b000000000000002f000000000000002e00000000",
            INIT_72 => X"0000001c00000000000000190000000000000011000000000000001a00000000",
            INIT_73 => X"0000001c000000000000001d0000000000000020000000000000001f00000000",
            INIT_74 => X"0000000c00000000000000100000000000000015000000000000001800000000",
            INIT_75 => X"0000000600000000000000080000000000000016000000000000001400000000",
            INIT_76 => X"0000000800000000000000080000000000000007000000000000000800000000",
            INIT_77 => X"0000001f000000000000001b000000000000000f000000000000000b00000000",
            INIT_78 => X"0000004e000000000000004c0000000000000048000000000000004500000000",
            INIT_79 => X"0000003800000000000000480000000000000053000000000000005800000000",
            INIT_7A => X"0000002a000000000000002b0000000000000026000000000000002000000000",
            INIT_7B => X"0000003100000000000000320000000000000033000000000000002f00000000",
            INIT_7C => X"0000001c000000000000001e0000000000000026000000000000002c00000000",
            INIT_7D => X"0000000c00000000000000130000000000000022000000000000002200000000",
            INIT_7E => X"0000000d000000000000000f0000000000000010000000000000000e00000000",
            INIT_7F => X"0000001d000000000000001e000000000000001a000000000000001200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE37;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE38 : if BRAM_NAME = "sampleifmap_layersamples_instance38" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003a00000000000000390000000000000031000000000000002500000000",
            INIT_01 => X"000000510000000000000050000000000000004e000000000000004200000000",
            INIT_02 => X"0000004200000000000000490000000000000052000000000000005600000000",
            INIT_03 => X"0000003800000000000000430000000000000043000000000000004100000000",
            INIT_04 => X"0000007300000000000000400000000000000032000000000000003200000000",
            INIT_05 => X"0000002700000000000000320000000000000038000000000000003400000000",
            INIT_06 => X"00000024000000000000002e0000000000000022000000000000001600000000",
            INIT_07 => X"0000001300000000000000150000000000000012000000000000001d00000000",
            INIT_08 => X"00000044000000000000004d0000000000000048000000000000004300000000",
            INIT_09 => X"000000420000000000000048000000000000004a000000000000004300000000",
            INIT_0A => X"0000003400000000000000390000000000000040000000000000004400000000",
            INIT_0B => X"0000002e00000000000000370000000000000036000000000000003200000000",
            INIT_0C => X"000000290000000000000027000000000000002a000000000000002900000000",
            INIT_0D => X"00000021000000000000001e0000000000000023000000000000002800000000",
            INIT_0E => X"0000001b000000000000001e000000000000002e000000000000002200000000",
            INIT_0F => X"0000001200000000000000160000000000000015000000000000001c00000000",
            INIT_10 => X"0000003e00000000000000480000000000000044000000000000004800000000",
            INIT_11 => X"000000310000000000000038000000000000003d000000000000003a00000000",
            INIT_12 => X"00000028000000000000002b000000000000002d000000000000003000000000",
            INIT_13 => X"00000026000000000000002b000000000000002a000000000000002600000000",
            INIT_14 => X"0000001c000000000000001e0000000000000023000000000000002200000000",
            INIT_15 => X"00000022000000000000001f0000000000000021000000000000002300000000",
            INIT_16 => X"0000000e000000000000000d0000000000000022000000000000003000000000",
            INIT_17 => X"0000001100000000000000130000000000000014000000000000001500000000",
            INIT_18 => X"0000003c000000000000003d0000000000000036000000000000003800000000",
            INIT_19 => X"00000024000000000000002b0000000000000030000000000000003e00000000",
            INIT_1A => X"0000002000000000000000220000000000000023000000000000002300000000",
            INIT_1B => X"0000002000000000000000220000000000000021000000000000001f00000000",
            INIT_1C => X"0000001d000000000000001b000000000000001e000000000000001d00000000",
            INIT_1D => X"00000025000000000000001d000000000000001c000000000000002000000000",
            INIT_1E => X"0000000f000000000000000b0000000000000012000000000000002a00000000",
            INIT_1F => X"0000001100000000000000100000000000000013000000000000001600000000",
            INIT_20 => X"0000003b00000000000000420000000000000039000000000000003900000000",
            INIT_21 => X"0000001b00000000000000200000000000000024000000000000003400000000",
            INIT_22 => X"0000001a000000000000001c000000000000001d000000000000001c00000000",
            INIT_23 => X"0000001e000000000000001c000000000000001a000000000000001a00000000",
            INIT_24 => X"0000001c000000000000001c000000000000001c000000000000001c00000000",
            INIT_25 => X"0000002a00000000000000430000000000000030000000000000001c00000000",
            INIT_26 => X"00000019000000000000000d0000000000000012000000000000001900000000",
            INIT_27 => X"000000110000000000000013000000000000001f000000000000001b00000000",
            INIT_28 => X"00000021000000000000002f000000000000003a000000000000003b00000000",
            INIT_29 => X"000000160000000000000019000000000000001a000000000000001a00000000",
            INIT_2A => X"00000019000000000000001a0000000000000019000000000000001700000000",
            INIT_2B => X"0000001f000000000000001b0000000000000018000000000000001800000000",
            INIT_2C => X"0000001e0000000000000021000000000000001e000000000000001d00000000",
            INIT_2D => X"0000003c000000000000005e000000000000005d000000000000002100000000",
            INIT_2E => X"0000002c000000000000001e000000000000001b000000000000002900000000",
            INIT_2F => X"000000130000000000000018000000000000002d000000000000002b00000000",
            INIT_30 => X"000000140000000000000017000000000000001c000000000000002200000000",
            INIT_31 => X"0000001500000000000000160000000000000017000000000000001600000000",
            INIT_32 => X"0000001a00000000000000190000000000000016000000000000001600000000",
            INIT_33 => X"00000023000000000000001d0000000000000019000000000000001800000000",
            INIT_34 => X"0000001e0000000000000023000000000000001f000000000000002000000000",
            INIT_35 => X"0000002500000000000000370000000000000059000000000000003300000000",
            INIT_36 => X"0000002d000000000000002b0000000000000028000000000000003800000000",
            INIT_37 => X"000000150000000000000017000000000000001e000000000000002400000000",
            INIT_38 => X"0000001200000000000000100000000000000011000000000000001100000000",
            INIT_39 => X"0000001600000000000000160000000000000017000000000000001600000000",
            INIT_3A => X"0000001b000000000000001a0000000000000017000000000000001800000000",
            INIT_3B => X"00000027000000000000001d000000000000001b000000000000001900000000",
            INIT_3C => X"000000300000000000000033000000000000002d000000000000002800000000",
            INIT_3D => X"0000000b00000000000000120000000000000040000000000000004100000000",
            INIT_3E => X"00000020000000000000001f0000000000000025000000000000002200000000",
            INIT_3F => X"0000001500000000000000160000000000000016000000000000001900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001200000000000000120000000000000012000000000000001100000000",
            INIT_41 => X"0000001700000000000000170000000000000016000000000000001500000000",
            INIT_42 => X"0000001e000000000000001c0000000000000018000000000000001900000000",
            INIT_43 => X"0000003b00000000000000330000000000000038000000000000002500000000",
            INIT_44 => X"000000360000000000000037000000000000003a000000000000003b00000000",
            INIT_45 => X"0000001000000000000000110000000000000028000000000000003d00000000",
            INIT_46 => X"0000001b00000000000000180000000000000019000000000000001a00000000",
            INIT_47 => X"0000001400000000000000150000000000000017000000000000001a00000000",
            INIT_48 => X"0000001200000000000000120000000000000012000000000000001300000000",
            INIT_49 => X"0000001800000000000000160000000000000014000000000000001500000000",
            INIT_4A => X"0000003100000000000000200000000000000019000000000000001800000000",
            INIT_4B => X"000000340000000000000039000000000000004c000000000000003e00000000",
            INIT_4C => X"0000003a0000000000000032000000000000002e000000000000003100000000",
            INIT_4D => X"0000002c00000000000000300000000000000031000000000000003800000000",
            INIT_4E => X"0000001900000000000000190000000000000023000000000000002900000000",
            INIT_4F => X"0000001400000000000000140000000000000018000000000000001900000000",
            INIT_50 => X"0000001200000000000000130000000000000012000000000000001400000000",
            INIT_51 => X"0000001700000000000000150000000000000015000000000000001500000000",
            INIT_52 => X"0000003500000000000000240000000000000019000000000000001900000000",
            INIT_53 => X"0000004a000000000000003e0000000000000042000000000000003100000000",
            INIT_54 => X"000000b800000000000000a60000000000000089000000000000006800000000",
            INIT_55 => X"00000021000000000000004b0000000000000068000000000000007c00000000",
            INIT_56 => X"000000190000000000000026000000000000003d000000000000003800000000",
            INIT_57 => X"0000001300000000000000120000000000000019000000000000001800000000",
            INIT_58 => X"0000001300000000000000140000000000000012000000000000001500000000",
            INIT_59 => X"0000001800000000000000160000000000000018000000000000001800000000",
            INIT_5A => X"00000030000000000000001f000000000000001d000000000000001900000000",
            INIT_5B => X"000000be00000000000000b20000000000000097000000000000005500000000",
            INIT_5C => X"000000c500000000000000ca00000000000000cd00000000000000cd00000000",
            INIT_5D => X"00000016000000000000009800000000000000d000000000000000b200000000",
            INIT_5E => X"0000002800000000000000460000000000000025000000000000001800000000",
            INIT_5F => X"0000001100000000000000110000000000000016000000000000001500000000",
            INIT_60 => X"0000001500000000000000160000000000000014000000000000001400000000",
            INIT_61 => X"0000001a00000000000000190000000000000018000000000000001800000000",
            INIT_62 => X"0000007000000000000000420000000000000020000000000000001900000000",
            INIT_63 => X"00000075000000000000008c000000000000009b000000000000009000000000",
            INIT_64 => X"0000003d00000000000000470000000000000058000000000000006400000000",
            INIT_65 => X"0000004e00000000000000d500000000000000e8000000000000007500000000",
            INIT_66 => X"000000460000000000000032000000000000000a000000000000000f00000000",
            INIT_67 => X"0000001000000000000000110000000000000015000000000000001a00000000",
            INIT_68 => X"0000001600000000000000190000000000000016000000000000001400000000",
            INIT_69 => X"0000001a00000000000000190000000000000017000000000000001700000000",
            INIT_6A => X"0000005b00000000000000670000000000000048000000000000001a00000000",
            INIT_6B => X"0000001200000000000000340000000000000056000000000000005000000000",
            INIT_6C => X"00000010000000000000000f0000000000000022000000000000001100000000",
            INIT_6D => X"0000009b00000000000000e000000000000000dd000000000000007c00000000",
            INIT_6E => X"0000003b00000000000000160000000000000007000000000000002400000000",
            INIT_6F => X"0000001000000000000000120000000000000013000000000000002100000000",
            INIT_70 => X"00000016000000000000001b0000000000000017000000000000001800000000",
            INIT_71 => X"0000001500000000000000130000000000000019000000000000001800000000",
            INIT_72 => X"00000029000000000000003a0000000000000055000000000000003700000000",
            INIT_73 => X"000000180000000000000032000000000000004e000000000000003d00000000",
            INIT_74 => X"00000049000000000000001e000000000000002b000000000000000b00000000",
            INIT_75 => X"000000cd00000000000000d100000000000000d800000000000000bf00000000",
            INIT_76 => X"000000170000000000000010000000000000000e000000000000006700000000",
            INIT_77 => X"0000001200000000000000140000000000000016000000000000001b00000000",
            INIT_78 => X"00000017000000000000001a0000000000000016000000000000001a00000000",
            INIT_79 => X"00000034000000000000003c0000000000000025000000000000001900000000",
            INIT_7A => X"0000003b00000000000000380000000000000034000000000000004c00000000",
            INIT_7B => X"00000026000000000000002e000000000000004d000000000000005000000000",
            INIT_7C => X"000000c4000000000000007c0000000000000049000000000000002300000000",
            INIT_7D => X"000000d200000000000000d900000000000000d800000000000000df00000000",
            INIT_7E => X"0000000e00000000000000150000000000000039000000000000007600000000",
            INIT_7F => X"00000011000000000000003e0000000000000047000000000000001f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE38;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE39 : if BRAM_NAME = "sampleifmap_layersamples_instance39" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001700000000000000190000000000000014000000000000001900000000",
            INIT_01 => X"0000005c00000000000000600000000000000035000000000000002100000000",
            INIT_02 => X"00000042000000000000003e000000000000005d000000000000004900000000",
            INIT_03 => X"000000a2000000000000005a0000000000000047000000000000005100000000",
            INIT_04 => X"000000f500000000000000f500000000000000df00000000000000c400000000",
            INIT_05 => X"0000007900000000000000de00000000000000e400000000000000e300000000",
            INIT_06 => X"000000090000000000000011000000000000003b000000000000002500000000",
            INIT_07 => X"000000130000000000000075000000000000008c000000000000004800000000",
            INIT_08 => X"0000001a00000000000000180000000000000015000000000000001900000000",
            INIT_09 => X"000000450000000000000035000000000000002c000000000000002800000000",
            INIT_0A => X"0000002900000000000000250000000000000052000000000000005800000000",
            INIT_0B => X"000000fb00000000000000940000000000000020000000000000003100000000",
            INIT_0C => X"000000e200000000000000e900000000000000f200000000000000f600000000",
            INIT_0D => X"0000001f000000000000008b00000000000000e200000000000000e100000000",
            INIT_0E => X"0000004300000000000000280000000000000019000000000000000b00000000",
            INIT_0F => X"00000022000000000000009700000000000000a2000000000000008500000000",
            INIT_10 => X"0000002600000000000000160000000000000013000000000000001600000000",
            INIT_11 => X"00000036000000000000002e0000000000000046000000000000005d00000000",
            INIT_12 => X"0000001b00000000000000180000000000000026000000000000004b00000000",
            INIT_13 => X"000000e300000000000000a30000000000000031000000000000003800000000",
            INIT_14 => X"000000da00000000000000cb00000000000000cd00000000000000d600000000",
            INIT_15 => X"0000004a00000000000000a300000000000000e400000000000000e500000000",
            INIT_16 => X"000000950000000000000080000000000000005a000000000000003900000000",
            INIT_17 => X"0000003300000000000000a00000000000000096000000000000009700000000",
            INIT_18 => X"0000007c0000000000000026000000000000000f000000000000001300000000",
            INIT_19 => X"0000002a0000000000000024000000000000005a00000000000000af00000000",
            INIT_1A => X"00000015000000000000000b0000000000000017000000000000003f00000000",
            INIT_1B => X"000000d000000000000000aa000000000000004f000000000000004000000000",
            INIT_1C => X"000000d600000000000000d300000000000000c500000000000000c700000000",
            INIT_1D => X"000000b100000000000000e300000000000000d900000000000000ce00000000",
            INIT_1E => X"000000a200000000000000a700000000000000a8000000000000009800000000",
            INIT_1F => X"0000002a00000000000000880000000000000097000000000000009a00000000",
            INIT_20 => X"000000dc0000000000000065000000000000000a000000000000001200000000",
            INIT_21 => X"0000002e000000000000002f000000000000006f00000000000000be00000000",
            INIT_22 => X"0000000e0000000000000009000000000000000a000000000000003900000000",
            INIT_23 => X"000000cc00000000000000b10000000000000042000000000000001f00000000",
            INIT_24 => X"0000007c00000000000000c600000000000000ca00000000000000c200000000",
            INIT_25 => X"000000d300000000000000ac0000000000000066000000000000004f00000000",
            INIT_26 => X"000000a900000000000000b100000000000000b800000000000000c800000000",
            INIT_27 => X"00000011000000000000004a000000000000008c000000000000009c00000000",
            INIT_28 => X"000000a500000000000000840000000000000014000000000000000e00000000",
            INIT_29 => X"0000003400000000000000370000000000000080000000000000009600000000",
            INIT_2A => X"00000016000000000000000a0000000000000003000000000000001e00000000",
            INIT_2B => X"000000c600000000000000b40000000000000048000000000000002d00000000",
            INIT_2C => X"00000019000000000000007b00000000000000cd00000000000000be00000000",
            INIT_2D => X"000000a30000000000000038000000000000001e000000000000001a00000000",
            INIT_2E => X"00000093000000000000009e00000000000000b800000000000000ca00000000",
            INIT_2F => X"00000011000000000000000d0000000000000044000000000000008800000000",
            INIT_30 => X"0000002100000000000000530000000000000023000000000000000a00000000",
            INIT_31 => X"00000035000000000000003e0000000000000082000000000000005300000000",
            INIT_32 => X"0000004800000000000000100000000000000007000000000000001300000000",
            INIT_33 => X"000000c200000000000000b70000000000000075000000000000006c00000000",
            INIT_34 => X"0000001e000000000000002f00000000000000b700000000000000c300000000",
            INIT_35 => X"0000004f0000000000000014000000000000002b000000000000003100000000",
            INIT_36 => X"000000810000000000000084000000000000009400000000000000a100000000",
            INIT_37 => X"000000180000000000000009000000000000000a000000000000004000000000",
            INIT_38 => X"0000002300000000000000370000000000000021000000000000000a00000000",
            INIT_39 => X"00000024000000000000004e0000000000000088000000000000004600000000",
            INIT_3A => X"0000005800000000000000220000000000000011000000000000000f00000000",
            INIT_3B => X"000000cd00000000000000cd000000000000007e000000000000006100000000",
            INIT_3C => X"0000002b0000000000000020000000000000009800000000000000d000000000",
            INIT_3D => X"0000001f0000000000000020000000000000001f000000000000002000000000",
            INIT_3E => X"00000063000000000000008a0000000000000091000000000000007500000000",
            INIT_3F => X"000000210000000000000019000000000000000c000000000000001700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004100000000000000360000000000000015000000000000000a00000000",
            INIT_41 => X"0000002100000000000000570000000000000088000000000000004700000000",
            INIT_42 => X"00000057000000000000003f0000000000000027000000000000001500000000",
            INIT_43 => X"000000c500000000000000cf000000000000009a000000000000005600000000",
            INIT_44 => X"000000380000000000000025000000000000008100000000000000c600000000",
            INIT_45 => X"0000000f000000000000001c000000000000002c000000000000003700000000",
            INIT_46 => X"00000043000000000000008b0000000000000093000000000000004d00000000",
            INIT_47 => X"0000001f000000000000001c0000000000000014000000000000000e00000000",
            INIT_48 => X"0000003e000000000000002f000000000000000e000000000000000700000000",
            INIT_49 => X"0000001c00000000000000560000000000000080000000000000004500000000",
            INIT_4A => X"0000006f000000000000005e000000000000003c000000000000001e00000000",
            INIT_4B => X"000000b400000000000000b600000000000000a2000000000000006f00000000",
            INIT_4C => X"0000003c0000000000000029000000000000007f00000000000000bc00000000",
            INIT_4D => X"0000000f00000000000000230000000000000035000000000000004b00000000",
            INIT_4E => X"00000026000000000000006f000000000000007a000000000000002c00000000",
            INIT_4F => X"000000160000000000000010000000000000000d000000000000000700000000",
            INIT_50 => X"0000003b00000000000000270000000000000011000000000000000b00000000",
            INIT_51 => X"0000003d00000000000000680000000000000075000000000000004600000000",
            INIT_52 => X"000000b7000000000000009f0000000000000079000000000000005100000000",
            INIT_53 => X"000000c700000000000000c900000000000000c300000000000000b900000000",
            INIT_54 => X"0000003c000000000000002a000000000000008800000000000000c600000000",
            INIT_55 => X"0000001c00000000000000340000000000000062000000000000006600000000",
            INIT_56 => X"000000100000000000000045000000000000004f000000000000001500000000",
            INIT_57 => X"00000016000000000000000c0000000000000007000000000000000300000000",
            INIT_58 => X"00000043000000000000001d0000000000000014000000000000001300000000",
            INIT_59 => X"0000003c00000000000000550000000000000067000000000000004900000000",
            INIT_5A => X"00000064000000000000005b0000000000000050000000000000004500000000",
            INIT_5B => X"0000006d00000000000000710000000000000071000000000000006800000000",
            INIT_5C => X"0000004100000000000000250000000000000059000000000000006d00000000",
            INIT_5D => X"00000017000000000000001f0000000000000042000000000000004000000000",
            INIT_5E => X"00000005000000000000000e0000000000000014000000000000000800000000",
            INIT_5F => X"00000018000000000000000b0000000000000006000000000000000600000000",
            INIT_60 => X"00000025000000000000001d000000000000001c000000000000001700000000",
            INIT_61 => X"000000070000000000000016000000000000002c000000000000002c00000000",
            INIT_62 => X"0000000c000000000000000c000000000000000a000000000000000a00000000",
            INIT_63 => X"0000001000000000000000110000000000000010000000000000000d00000000",
            INIT_64 => X"000000430000000000000009000000000000000f000000000000000f00000000",
            INIT_65 => X"0000001000000000000000380000000000000030000000000000004400000000",
            INIT_66 => X"0000000400000000000000030000000000000003000000000000000400000000",
            INIT_67 => X"00000019000000000000000e0000000000000009000000000000000600000000",
            INIT_68 => X"0000002000000000000000270000000000000025000000000000002100000000",
            INIT_69 => X"0000002000000000000000190000000000000012000000000000001700000000",
            INIT_6A => X"0000001700000000000000170000000000000015000000000000001700000000",
            INIT_6B => X"0000000f00000000000000130000000000000015000000000000001700000000",
            INIT_6C => X"000000180000000000000007000000000000000a000000000000000b00000000",
            INIT_6D => X"0000000800000000000000290000000000000047000000000000003e00000000",
            INIT_6E => X"0000000600000000000000050000000000000005000000000000000400000000",
            INIT_6F => X"0000001d0000000000000018000000000000000e000000000000000900000000",
            INIT_70 => X"0000003200000000000000290000000000000025000000000000002300000000",
            INIT_71 => X"0000004d00000000000000510000000000000043000000000000003c00000000",
            INIT_72 => X"00000030000000000000002d0000000000000024000000000000002c00000000",
            INIT_73 => X"000000230000000000000027000000000000002c000000000000003100000000",
            INIT_74 => X"000000100000000000000015000000000000001b000000000000001d00000000",
            INIT_75 => X"00000009000000000000000a0000000000000019000000000000001700000000",
            INIT_76 => X"0000000b000000000000000a0000000000000009000000000000000b00000000",
            INIT_77 => X"0000001e000000000000001f0000000000000014000000000000000e00000000",
            INIT_78 => X"00000057000000000000003b000000000000002a000000000000002a00000000",
            INIT_79 => X"000000520000000000000066000000000000006f000000000000006d00000000",
            INIT_7A => X"000000470000000000000045000000000000003e000000000000003700000000",
            INIT_7B => X"0000004300000000000000460000000000000048000000000000004a00000000",
            INIT_7C => X"00000029000000000000002b0000000000000033000000000000003b00000000",
            INIT_7D => X"000000120000000000000018000000000000002c000000000000002f00000000",
            INIT_7E => X"0000001300000000000000150000000000000016000000000000001400000000",
            INIT_7F => X"0000001e0000000000000020000000000000001c000000000000001600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE39;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE40 : if BRAM_NAME = "sampleifmap_layersamples_instance40" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000a000000000000000e000000000000000b000000000000000d00000000",
            INIT_01 => X"000000020000000000000005000000000000000a000000000000000900000000",
            INIT_02 => X"0000000200000000000000010000000000000003000000000000000300000000",
            INIT_03 => X"0000000000000000000000050000000000000006000000000000000400000000",
            INIT_04 => X"0000005600000000000000230000000000000000000000000000000100000000",
            INIT_05 => X"00000008000000000000001d0000000000000017000000000000001600000000",
            INIT_06 => X"0000001d0000000000000027000000000000001b000000000000000d00000000",
            INIT_07 => X"0000000500000000000000060000000000000008000000000000001300000000",
            INIT_08 => X"00000004000000000000000a000000000000000c000000000000000d00000000",
            INIT_09 => X"0000000000000000000000030000000000000008000000000000000700000000",
            INIT_0A => X"0000000100000000000000010000000000000002000000000000000400000000",
            INIT_0B => X"0000000100000000000000040000000000000004000000000000000200000000",
            INIT_0C => X"0000001300000000000000100000000000000001000000000000000100000000",
            INIT_0D => X"0000000700000000000000060000000000000006000000000000000700000000",
            INIT_0E => X"000000160000000000000017000000000000002e000000000000002100000000",
            INIT_0F => X"0000000600000000000000040000000000000008000000000000001300000000",
            INIT_10 => X"0000000000000000000000030000000000000004000000000000000700000000",
            INIT_11 => X"0000000000000000000000010000000000000004000000000000000400000000",
            INIT_12 => X"0000000400000000000000040000000000000004000000000000000400000000",
            INIT_13 => X"0000000300000000000000050000000000000006000000000000000400000000",
            INIT_14 => X"00000009000000000000000c0000000000000003000000000000000400000000",
            INIT_15 => X"0000000a00000000000000060000000000000007000000000000000400000000",
            INIT_16 => X"0000000c000000000000000d0000000000000023000000000000002800000000",
            INIT_17 => X"0000000600000000000000030000000000000006000000000000000f00000000",
            INIT_18 => X"0000000b00000000000000080000000000000003000000000000000100000000",
            INIT_19 => X"0000000300000000000000030000000000000004000000000000001200000000",
            INIT_1A => X"0000000700000000000000080000000000000006000000000000000500000000",
            INIT_1B => X"0000000600000000000000060000000000000009000000000000000800000000",
            INIT_1C => X"00000009000000000000000a0000000000000005000000000000000700000000",
            INIT_1D => X"000000170000000000000010000000000000000a000000000000000400000000",
            INIT_1E => X"0000000e00000000000000110000000000000016000000000000001e00000000",
            INIT_1F => X"0000000800000000000000050000000000000006000000000000000f00000000",
            INIT_20 => X"0000001a000000000000001d0000000000000013000000000000000c00000000",
            INIT_21 => X"0000000800000000000000070000000000000006000000000000001700000000",
            INIT_22 => X"0000000800000000000000090000000000000008000000000000000700000000",
            INIT_23 => X"000000080000000000000007000000000000000a000000000000000900000000",
            INIT_24 => X"0000000700000000000000080000000000000007000000000000000900000000",
            INIT_25 => X"0000002700000000000000400000000000000025000000000000000800000000",
            INIT_26 => X"00000015000000000000000e0000000000000010000000000000001000000000",
            INIT_27 => X"00000009000000000000000d000000000000000f000000000000000e00000000",
            INIT_28 => X"0000000c0000000000000016000000000000001e000000000000001800000000",
            INIT_29 => X"0000000800000000000000090000000000000006000000000000000900000000",
            INIT_2A => X"0000000a00000000000000090000000000000005000000000000000500000000",
            INIT_2B => X"000000090000000000000007000000000000000a000000000000000b00000000",
            INIT_2C => X"00000007000000000000000b000000000000000b000000000000000a00000000",
            INIT_2D => X"0000003b000000000000005d0000000000000055000000000000001400000000",
            INIT_2E => X"000000200000000000000013000000000000000e000000000000002200000000",
            INIT_2F => X"000000090000000000000010000000000000001b000000000000001700000000",
            INIT_30 => X"00000007000000000000000a000000000000000b000000000000000c00000000",
            INIT_31 => X"00000007000000000000000a0000000000000008000000000000000800000000",
            INIT_32 => X"0000000e000000000000000a0000000000000005000000000000000600000000",
            INIT_33 => X"0000000c000000000000000a000000000000000c000000000000000d00000000",
            INIT_34 => X"00000007000000000000000e000000000000000e000000000000000900000000",
            INIT_35 => X"00000028000000000000003c0000000000000056000000000000002500000000",
            INIT_36 => X"0000001c000000000000001c000000000000001c000000000000003500000000",
            INIT_37 => X"0000000700000000000000060000000000000010000000000000001400000000",
            INIT_38 => X"0000000700000000000000060000000000000006000000000000000300000000",
            INIT_39 => X"00000009000000000000000c000000000000000a000000000000000b00000000",
            INIT_3A => X"0000000e000000000000000c0000000000000008000000000000000900000000",
            INIT_3B => X"0000001300000000000000100000000000000012000000000000000e00000000",
            INIT_3C => X"00000016000000000000001a0000000000000015000000000000001000000000",
            INIT_3D => X"0000000a0000000000000014000000000000003e000000000000003100000000",
            INIT_3E => X"0000000d0000000000000010000000000000001a000000000000001e00000000",
            INIT_3F => X"0000000700000000000000040000000000000008000000000000000900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000080000000000000009000000000000000a000000000000000700000000",
            INIT_41 => X"0000000b000000000000000e000000000000000a000000000000000b00000000",
            INIT_42 => X"0000000f000000000000000e000000000000000c000000000000000d00000000",
            INIT_43 => X"0000002800000000000000220000000000000024000000000000001300000000",
            INIT_44 => X"0000002200000000000000220000000000000020000000000000002400000000",
            INIT_45 => X"00000009000000000000000f000000000000002b000000000000003300000000",
            INIT_46 => X"0000000a0000000000000009000000000000000c000000000000001400000000",
            INIT_47 => X"0000000800000000000000080000000000000008000000000000000800000000",
            INIT_48 => X"00000008000000000000000b000000000000000c000000000000000c00000000",
            INIT_49 => X"0000000d000000000000000e000000000000000a000000000000000c00000000",
            INIT_4A => X"000000220000000000000014000000000000000e000000000000000e00000000",
            INIT_4B => X"0000002600000000000000280000000000000031000000000000002700000000",
            INIT_4C => X"000000320000000000000027000000000000001b000000000000002000000000",
            INIT_4D => X"000000260000000000000034000000000000003b000000000000003600000000",
            INIT_4E => X"0000000c000000000000000b0000000000000015000000000000002300000000",
            INIT_4F => X"0000000a000000000000000b0000000000000009000000000000000600000000",
            INIT_50 => X"00000009000000000000000b000000000000000b000000000000000c00000000",
            INIT_51 => X"0000000d000000000000000d000000000000000a000000000000000c00000000",
            INIT_52 => X"00000028000000000000001b0000000000000010000000000000000d00000000",
            INIT_53 => X"0000003f00000000000000320000000000000032000000000000002000000000",
            INIT_54 => X"000000b400000000000000a10000000000000077000000000000005800000000",
            INIT_55 => X"0000002200000000000000540000000000000071000000000000007900000000",
            INIT_56 => X"00000011000000000000001d0000000000000031000000000000003200000000",
            INIT_57 => X"0000000a000000000000000c000000000000000a000000000000000900000000",
            INIT_58 => X"0000000b000000000000000e000000000000000a000000000000000900000000",
            INIT_59 => X"0000000c000000000000000d000000000000000c000000000000000e00000000",
            INIT_5A => X"0000002700000000000000180000000000000012000000000000000c00000000",
            INIT_5B => X"000000ba00000000000000af0000000000000093000000000000004d00000000",
            INIT_5C => X"000000ca00000000000000d200000000000000c800000000000000c800000000",
            INIT_5D => X"0000001c000000000000009e00000000000000d500000000000000b100000000",
            INIT_5E => X"0000002500000000000000460000000000000022000000000000001300000000",
            INIT_5F => X"00000009000000000000000b0000000000000009000000000000000a00000000",
            INIT_60 => X"0000000d000000000000000f000000000000000a000000000000000800000000",
            INIT_61 => X"0000000e000000000000000d000000000000000e000000000000001000000000",
            INIT_62 => X"0000006c000000000000003e0000000000000018000000000000000c00000000",
            INIT_63 => X"0000007d000000000000009300000000000000a2000000000000008e00000000",
            INIT_64 => X"0000004a0000000000000054000000000000005e000000000000006e00000000",
            INIT_65 => X"0000005400000000000000d700000000000000f1000000000000007e00000000",
            INIT_66 => X"0000004900000000000000340000000000000009000000000000000c00000000",
            INIT_67 => X"000000080000000000000009000000000000000d000000000000001900000000",
            INIT_68 => X"0000000e000000000000000f000000000000000b000000000000000b00000000",
            INIT_69 => X"0000000e000000000000000c0000000000000010000000000000001100000000",
            INIT_6A => X"0000005d00000000000000670000000000000044000000000000001400000000",
            INIT_6B => X"00000019000000000000003d000000000000005f000000000000005600000000",
            INIT_6C => X"0000001700000000000000110000000000000023000000000000001600000000",
            INIT_6D => X"000000a700000000000000eb00000000000000eb000000000000008900000000",
            INIT_6E => X"0000004200000000000000170000000000000007000000000000002a00000000",
            INIT_6F => X"0000000700000000000000090000000000000011000000000000002800000000",
            INIT_70 => X"0000000e0000000000000012000000000000000d000000000000000f00000000",
            INIT_71 => X"00000012000000000000000b0000000000000012000000000000001000000000",
            INIT_72 => X"0000002e000000000000003b0000000000000053000000000000003600000000",
            INIT_73 => X"0000001b00000000000000370000000000000053000000000000004400000000",
            INIT_74 => X"0000004c000000000000001c0000000000000027000000000000000c00000000",
            INIT_75 => X"000000e000000000000000e700000000000000e800000000000000c800000000",
            INIT_76 => X"0000001a00000000000000130000000000000016000000000000007300000000",
            INIT_77 => X"00000008000000000000000d0000000000000016000000000000001f00000000",
            INIT_78 => X"0000000e0000000000000013000000000000000d000000000000001000000000",
            INIT_79 => X"000000370000000000000039000000000000001e000000000000000e00000000",
            INIT_7A => X"0000003c00000000000000390000000000000035000000000000004f00000000",
            INIT_7B => X"000000290000000000000032000000000000004e000000000000005200000000",
            INIT_7C => X"000000c8000000000000007c0000000000000047000000000000002300000000",
            INIT_7D => X"000000dd00000000000000ec00000000000000e600000000000000e700000000",
            INIT_7E => X"0000000e000000000000001a0000000000000044000000000000007e00000000",
            INIT_7F => X"00000009000000000000003f0000000000000049000000000000002000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE40;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE41 : if BRAM_NAME = "sampleifmap_layersamples_instance41" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000110000000000000013000000000000000e000000000000001100000000",
            INIT_01 => X"0000005c000000000000005d000000000000002f000000000000001800000000",
            INIT_02 => X"0000003d000000000000003c0000000000000062000000000000004f00000000",
            INIT_03 => X"000000a6000000000000005e0000000000000047000000000000004c00000000",
            INIT_04 => X"000000fc00000000000000fa00000000000000e200000000000000c600000000",
            INIT_05 => X"0000007c00000000000000e700000000000000f000000000000000ed00000000",
            INIT_06 => X"0000000c000000000000001c000000000000004a000000000000002a00000000",
            INIT_07 => X"00000011000000000000007e0000000000000095000000000000004c00000000",
            INIT_08 => X"0000001500000000000000120000000000000010000000000000001200000000",
            INIT_09 => X"000000480000000000000038000000000000002a000000000000002400000000",
            INIT_0A => X"0000002400000000000000240000000000000058000000000000006000000000",
            INIT_0B => X"00000100000000000000009a0000000000000022000000000000002d00000000",
            INIT_0C => X"000000ed00000000000000f400000000000000f900000000000000fa00000000",
            INIT_0D => X"00000027000000000000009600000000000000ee00000000000000ed00000000",
            INIT_0E => X"0000004d000000000000003b000000000000002e000000000000001500000000",
            INIT_0F => X"0000002600000000000000a300000000000000ae000000000000008e00000000",
            INIT_10 => X"0000002200000000000000100000000000000010000000000000001100000000",
            INIT_11 => X"00000042000000000000003c0000000000000049000000000000005c00000000",
            INIT_12 => X"00000021000000000000001c000000000000002c000000000000005400000000",
            INIT_13 => X"000000f000000000000000ae0000000000000037000000000000003e00000000",
            INIT_14 => X"000000e700000000000000d900000000000000d900000000000000e100000000",
            INIT_15 => X"0000005600000000000000b100000000000000ee00000000000000ef00000000",
            INIT_16 => X"000000a40000000000000092000000000000006a000000000000004500000000",
            INIT_17 => X"0000003700000000000000a900000000000000a100000000000000a400000000",
            INIT_18 => X"0000007d0000000000000020000000000000000a000000000000000d00000000",
            INIT_19 => X"000000380000000000000035000000000000006200000000000000b400000000",
            INIT_1A => X"0000001b000000000000000e000000000000001c000000000000004800000000",
            INIT_1B => X"000000e000000000000000b90000000000000059000000000000004900000000",
            INIT_1C => X"000000e300000000000000e400000000000000d500000000000000d500000000",
            INIT_1D => X"000000c000000000000000f200000000000000e100000000000000d700000000",
            INIT_1E => X"000000b000000000000000b500000000000000b400000000000000a500000000",
            INIT_1F => X"0000002a000000000000008d000000000000009f00000000000000a600000000",
            INIT_20 => X"000000e500000000000000650000000000000007000000000000000c00000000",
            INIT_21 => X"00000039000000000000003e000000000000007b00000000000000c900000000",
            INIT_22 => X"0000000f0000000000000009000000000000000f000000000000004100000000",
            INIT_23 => X"000000da00000000000000bf000000000000004f000000000000002600000000",
            INIT_24 => X"0000008a00000000000000d800000000000000db00000000000000d000000000",
            INIT_25 => X"000000e400000000000000b8000000000000006d000000000000005800000000",
            INIT_26 => X"000000b500000000000000bf00000000000000c900000000000000da00000000",
            INIT_27 => X"0000000e000000000000004d000000000000009300000000000000a600000000",
            INIT_28 => X"000000b3000000000000008b0000000000000018000000000000000d00000000",
            INIT_29 => X"0000003d0000000000000045000000000000008d00000000000000a200000000",
            INIT_2A => X"0000001b000000000000000b0000000000000004000000000000002300000000",
            INIT_2B => X"000000d400000000000000c20000000000000056000000000000003600000000",
            INIT_2C => X"00000024000000000000008800000000000000db00000000000000cc00000000",
            INIT_2D => X"000000b100000000000000400000000000000022000000000000002000000000",
            INIT_2E => X"0000009f00000000000000ad00000000000000cc00000000000000dd00000000",
            INIT_2F => X"0000000d000000000000000f0000000000000049000000000000009000000000",
            INIT_30 => X"00000031000000000000005b0000000000000027000000000000000900000000",
            INIT_31 => X"0000003e000000000000004c000000000000008f000000000000006000000000",
            INIT_32 => X"0000005100000000000000150000000000000007000000000000001500000000",
            INIT_33 => X"000000d000000000000000c50000000000000083000000000000007900000000",
            INIT_34 => X"00000026000000000000003800000000000000c100000000000000d100000000",
            INIT_35 => X"000000590000000000000019000000000000002e000000000000003700000000",
            INIT_36 => X"0000008d000000000000009500000000000000a900000000000000b200000000",
            INIT_37 => X"000000140000000000000008000000000000000e000000000000004800000000",
            INIT_38 => X"00000030000000000000003b0000000000000022000000000000000500000000",
            INIT_39 => X"0000002d000000000000005c0000000000000095000000000000005300000000",
            INIT_3A => X"00000064000000000000002a0000000000000013000000000000000f00000000",
            INIT_3B => X"000000db00000000000000db000000000000008c000000000000006f00000000",
            INIT_3C => X"00000033000000000000002600000000000000a000000000000000de00000000",
            INIT_3D => X"0000002700000000000000240000000000000023000000000000002500000000",
            INIT_3E => X"0000006e000000000000009b00000000000000a4000000000000008200000000",
            INIT_3F => X"0000001e0000000000000016000000000000000c000000000000001d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004d000000000000003a0000000000000017000000000000000700000000",
            INIT_41 => X"0000002a00000000000000650000000000000094000000000000005400000000",
            INIT_42 => X"00000065000000000000004a000000000000002b000000000000001600000000",
            INIT_43 => X"000000d300000000000000dd00000000000000a8000000000000006400000000",
            INIT_44 => X"00000040000000000000002b000000000000008900000000000000d400000000",
            INIT_45 => X"0000001500000000000000230000000000000034000000000000003f00000000",
            INIT_46 => X"0000004e000000000000009a00000000000000a2000000000000005600000000",
            INIT_47 => X"0000001c00000000000000180000000000000012000000000000001300000000",
            INIT_48 => X"0000004c00000000000000370000000000000015000000000000000900000000",
            INIT_49 => X"000000250000000000000065000000000000008c000000000000005200000000",
            INIT_4A => X"0000007f000000000000006c0000000000000043000000000000002100000000",
            INIT_4B => X"000000c200000000000000c300000000000000b0000000000000007e00000000",
            INIT_4C => X"000000460000000000000030000000000000008700000000000000c900000000",
            INIT_4D => X"00000015000000000000002e0000000000000041000000000000005600000000",
            INIT_4E => X"00000031000000000000007b0000000000000083000000000000003200000000",
            INIT_4F => X"00000014000000000000000b000000000000000a000000000000000b00000000",
            INIT_50 => X"0000004900000000000000310000000000000017000000000000000b00000000",
            INIT_51 => X"0000004b00000000000000780000000000000084000000000000005700000000",
            INIT_52 => X"000000c800000000000000b10000000000000086000000000000005d00000000",
            INIT_53 => X"000000d500000000000000d400000000000000cf00000000000000c800000000",
            INIT_54 => X"000000480000000000000035000000000000009400000000000000d600000000",
            INIT_55 => X"000000220000000000000040000000000000006e000000000000007100000000",
            INIT_56 => X"00000016000000000000004c0000000000000055000000000000001800000000",
            INIT_57 => X"00000016000000000000000d0000000000000009000000000000000700000000",
            INIT_58 => X"0000004e00000000000000250000000000000016000000000000000f00000000",
            INIT_59 => X"0000004800000000000000600000000000000073000000000000005700000000",
            INIT_5A => X"000000720000000000000069000000000000005d000000000000005200000000",
            INIT_5B => X"0000007b000000000000007e000000000000007d000000000000007700000000",
            INIT_5C => X"0000004c00000000000000300000000000000066000000000000007c00000000",
            INIT_5D => X"0000001b0000000000000029000000000000004e000000000000004b00000000",
            INIT_5E => X"0000000600000000000000100000000000000018000000000000000900000000",
            INIT_5F => X"00000019000000000000000f000000000000000a000000000000000800000000",
            INIT_60 => X"0000002b0000000000000023000000000000001f000000000000001500000000",
            INIT_61 => X"0000000c00000000000000190000000000000030000000000000003200000000",
            INIT_62 => X"000000110000000000000011000000000000000e000000000000000e00000000",
            INIT_63 => X"00000019000000000000001a0000000000000018000000000000001400000000",
            INIT_64 => X"0000004a000000000000000d0000000000000014000000000000001800000000",
            INIT_65 => X"000000120000000000000041000000000000003b000000000000004e00000000",
            INIT_66 => X"0000000300000000000000040000000000000005000000000000000300000000",
            INIT_67 => X"0000001a000000000000000d0000000000000009000000000000000500000000",
            INIT_68 => X"00000025000000000000002c0000000000000028000000000000002100000000",
            INIT_69 => X"00000025000000000000001e0000000000000017000000000000001e00000000",
            INIT_6A => X"0000001c000000000000001c0000000000000019000000000000001c00000000",
            INIT_6B => X"0000001300000000000000170000000000000018000000000000001b00000000",
            INIT_6C => X"0000001c00000000000000060000000000000009000000000000000f00000000",
            INIT_6D => X"00000008000000000000002f0000000000000053000000000000004700000000",
            INIT_6E => X"0000000400000000000000050000000000000005000000000000000200000000",
            INIT_6F => X"0000001c0000000000000015000000000000000b000000000000000600000000",
            INIT_70 => X"0000003b00000000000000300000000000000029000000000000002500000000",
            INIT_71 => X"00000059000000000000005c000000000000004f000000000000004900000000",
            INIT_72 => X"0000003b0000000000000038000000000000002f000000000000003800000000",
            INIT_73 => X"00000028000000000000002b0000000000000030000000000000003900000000",
            INIT_74 => X"000000150000000000000015000000000000001b000000000000002300000000",
            INIT_75 => X"0000000800000000000000100000000000000025000000000000002100000000",
            INIT_76 => X"0000000a000000000000000a0000000000000009000000000000000800000000",
            INIT_77 => X"0000001c000000000000001d0000000000000012000000000000000d00000000",
            INIT_78 => X"0000006500000000000000460000000000000031000000000000002c00000000",
            INIT_79 => X"0000006300000000000000760000000000000080000000000000008000000000",
            INIT_7A => X"000000550000000000000054000000000000004e000000000000004700000000",
            INIT_7B => X"0000004f00000000000000510000000000000053000000000000005700000000",
            INIT_7C => X"000000310000000000000031000000000000003c000000000000004700000000",
            INIT_7D => X"0000001300000000000000200000000000000038000000000000003a00000000",
            INIT_7E => X"0000001500000000000000180000000000000018000000000000001300000000",
            INIT_7F => X"0000001c0000000000000022000000000000001f000000000000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE41;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE42 : if BRAM_NAME = "sampleifmap_layersamples_instance42" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004d00000000000000510000000000000052000000000000005300000000",
            INIT_01 => X"0000005c000000000000005b0000000000000055000000000000005100000000",
            INIT_02 => X"0000005c0000000000000065000000000000005f000000000000005c00000000",
            INIT_03 => X"0000004c00000000000000500000000000000052000000000000005700000000",
            INIT_04 => X"0000003e000000000000003f0000000000000041000000000000004400000000",
            INIT_05 => X"0000002f00000000000000340000000000000038000000000000003c00000000",
            INIT_06 => X"0000002200000000000000230000000000000025000000000000002a00000000",
            INIT_07 => X"000000150000000000000019000000000000001d000000000000002400000000",
            INIT_08 => X"0000004d00000000000000530000000000000053000000000000005400000000",
            INIT_09 => X"0000005d000000000000005a0000000000000054000000000000005000000000",
            INIT_0A => X"00000061000000000000005f0000000000000058000000000000005a00000000",
            INIT_0B => X"0000004c000000000000004e0000000000000052000000000000005800000000",
            INIT_0C => X"0000004200000000000000400000000000000044000000000000004700000000",
            INIT_0D => X"0000002e00000000000000340000000000000036000000000000003d00000000",
            INIT_0E => X"0000002300000000000000240000000000000026000000000000002a00000000",
            INIT_0F => X"0000001f000000000000001d000000000000001e000000000000002400000000",
            INIT_10 => X"0000004b00000000000000500000000000000051000000000000005200000000",
            INIT_11 => X"0000004c00000000000000580000000000000054000000000000004b00000000",
            INIT_12 => X"0000006300000000000000570000000000000056000000000000005200000000",
            INIT_13 => X"0000004c000000000000004d0000000000000058000000000000006500000000",
            INIT_14 => X"0000004000000000000000400000000000000044000000000000004900000000",
            INIT_15 => X"0000002d00000000000000340000000000000037000000000000003a00000000",
            INIT_16 => X"0000002c00000000000000290000000000000028000000000000002b00000000",
            INIT_17 => X"0000003500000000000000310000000000000030000000000000003100000000",
            INIT_18 => X"0000004e00000000000000500000000000000051000000000000005300000000",
            INIT_19 => X"0000003200000000000000500000000000000057000000000000004a00000000",
            INIT_1A => X"0000005b00000000000000570000000000000061000000000000005500000000",
            INIT_1B => X"0000005000000000000000580000000000000066000000000000006800000000",
            INIT_1C => X"0000003f000000000000003f0000000000000040000000000000004900000000",
            INIT_1D => X"0000003a00000000000000390000000000000038000000000000003b00000000",
            INIT_1E => X"000000470000000000000044000000000000003f000000000000003d00000000",
            INIT_1F => X"0000004500000000000000450000000000000047000000000000004900000000",
            INIT_20 => X"0000004f000000000000004f000000000000004f000000000000004f00000000",
            INIT_21 => X"00000037000000000000004c0000000000000053000000000000004a00000000",
            INIT_22 => X"0000004b000000000000004b0000000000000054000000000000005300000000",
            INIT_23 => X"00000057000000000000005a0000000000000059000000000000004e00000000",
            INIT_24 => X"0000004600000000000000430000000000000042000000000000005300000000",
            INIT_25 => X"0000005700000000000000540000000000000050000000000000004e00000000",
            INIT_26 => X"0000005900000000000000590000000000000056000000000000005700000000",
            INIT_27 => X"00000049000000000000004f0000000000000054000000000000005800000000",
            INIT_28 => X"0000004d000000000000004b000000000000004a000000000000004c00000000",
            INIT_29 => X"0000004600000000000000460000000000000049000000000000004900000000",
            INIT_2A => X"0000004900000000000000470000000000000045000000000000004600000000",
            INIT_2B => X"00000051000000000000004e000000000000004e000000000000004b00000000",
            INIT_2C => X"0000006200000000000000600000000000000059000000000000005a00000000",
            INIT_2D => X"0000006800000000000000660000000000000068000000000000006400000000",
            INIT_2E => X"0000005e0000000000000061000000000000005f000000000000006300000000",
            INIT_2F => X"0000004200000000000000490000000000000050000000000000005700000000",
            INIT_30 => X"0000004900000000000000470000000000000048000000000000004a00000000",
            INIT_31 => X"00000033000000000000002b000000000000003e000000000000004a00000000",
            INIT_32 => X"0000004700000000000000440000000000000040000000000000004400000000",
            INIT_33 => X"0000005e0000000000000051000000000000004a000000000000004b00000000",
            INIT_34 => X"00000072000000000000006e0000000000000062000000000000006000000000",
            INIT_35 => X"0000006d00000000000000680000000000000064000000000000006600000000",
            INIT_36 => X"000000500000000000000055000000000000005b000000000000006300000000",
            INIT_37 => X"0000004300000000000000460000000000000049000000000000004c00000000",
            INIT_38 => X"0000004800000000000000470000000000000048000000000000004700000000",
            INIT_39 => X"00000029000000000000002a000000000000003a000000000000004700000000",
            INIT_3A => X"0000003f000000000000003a0000000000000036000000000000003900000000",
            INIT_3B => X"0000006000000000000000520000000000000047000000000000004100000000",
            INIT_3C => X"00000067000000000000005d000000000000005e000000000000006900000000",
            INIT_3D => X"00000061000000000000006c000000000000006a000000000000006700000000",
            INIT_3E => X"000000500000000000000054000000000000005b000000000000005d00000000",
            INIT_3F => X"0000004d000000000000004f0000000000000050000000000000005000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000052000000000000004b0000000000000049000000000000004900000000",
            INIT_41 => X"0000002e00000000000000570000000000000067000000000000005800000000",
            INIT_42 => X"0000005200000000000000450000000000000038000000000000003800000000",
            INIT_43 => X"00000057000000000000005a0000000000000057000000000000005100000000",
            INIT_44 => X"0000005b000000000000005e0000000000000063000000000000006200000000",
            INIT_45 => X"00000066000000000000006a0000000000000066000000000000006100000000",
            INIT_46 => X"0000005c00000000000000610000000000000063000000000000005e00000000",
            INIT_47 => X"0000005f000000000000005b0000000000000059000000000000005900000000",
            INIT_48 => X"0000007b000000000000006d000000000000005f000000000000005600000000",
            INIT_49 => X"0000003300000000000000680000000000000099000000000000008800000000",
            INIT_4A => X"000000610000000000000049000000000000003b000000000000003c00000000",
            INIT_4B => X"0000005a0000000000000066000000000000006c000000000000006500000000",
            INIT_4C => X"0000005d00000000000000610000000000000061000000000000005f00000000",
            INIT_4D => X"0000006e00000000000000690000000000000063000000000000005d00000000",
            INIT_4E => X"0000006c000000000000006c0000000000000069000000000000006700000000",
            INIT_4F => X"0000006e000000000000006e000000000000006e000000000000006d00000000",
            INIT_50 => X"0000009d0000000000000096000000000000008b000000000000007f00000000",
            INIT_51 => X"00000032000000000000005700000000000000a200000000000000a000000000",
            INIT_52 => X"0000005800000000000000350000000000000038000000000000004300000000",
            INIT_53 => X"0000005a000000000000006b0000000000000070000000000000006500000000",
            INIT_54 => X"00000060000000000000005e0000000000000060000000000000005e00000000",
            INIT_55 => X"000000650000000000000060000000000000005f000000000000006000000000",
            INIT_56 => X"0000007e000000000000007d0000000000000071000000000000006800000000",
            INIT_57 => X"0000007000000000000000740000000000000077000000000000007b00000000",
            INIT_58 => X"000000a2000000000000009f000000000000009d000000000000009800000000",
            INIT_59 => X"0000002c000000000000005a000000000000009f00000000000000a000000000",
            INIT_5A => X"00000056000000000000003a0000000000000045000000000000004800000000",
            INIT_5B => X"0000005c0000000000000061000000000000005a000000000000006700000000",
            INIT_5C => X"0000005e000000000000005f0000000000000060000000000000005a00000000",
            INIT_5D => X"0000005c00000000000000570000000000000062000000000000006300000000",
            INIT_5E => X"0000008300000000000000830000000000000070000000000000006100000000",
            INIT_5F => X"0000006c00000000000000740000000000000079000000000000007f00000000",
            INIT_60 => X"0000009d00000000000000a0000000000000009e000000000000009b00000000",
            INIT_61 => X"0000003000000000000000720000000000000094000000000000009800000000",
            INIT_62 => X"00000067000000000000005e0000000000000058000000000000004400000000",
            INIT_63 => X"0000005d00000000000000580000000000000060000000000000007300000000",
            INIT_64 => X"0000005e00000000000000620000000000000065000000000000005900000000",
            INIT_65 => X"0000005500000000000000540000000000000065000000000000006300000000",
            INIT_66 => X"00000084000000000000007d000000000000006e000000000000006900000000",
            INIT_67 => X"0000005f000000000000006b0000000000000076000000000000007f00000000",
            INIT_68 => X"0000009200000000000000950000000000000094000000000000009400000000",
            INIT_69 => X"000000500000000000000088000000000000008e000000000000009000000000",
            INIT_6A => X"00000068000000000000005e0000000000000048000000000000002f00000000",
            INIT_6B => X"0000005e000000000000005c0000000000000071000000000000007200000000",
            INIT_6C => X"0000005d00000000000000610000000000000067000000000000005d00000000",
            INIT_6D => X"0000005200000000000000550000000000000061000000000000006000000000",
            INIT_6E => X"00000079000000000000006f000000000000006b000000000000006b00000000",
            INIT_6F => X"0000004d00000000000000570000000000000064000000000000007000000000",
            INIT_70 => X"0000008c000000000000008a0000000000000087000000000000008600000000",
            INIT_71 => X"0000008900000000000000970000000000000093000000000000008e00000000",
            INIT_72 => X"0000003e00000000000000320000000000000049000000000000005d00000000",
            INIT_73 => X"00000062000000000000005a000000000000005e000000000000005900000000",
            INIT_74 => X"0000006100000000000000670000000000000069000000000000006600000000",
            INIT_75 => X"000000530000000000000056000000000000005e000000000000005e00000000",
            INIT_76 => X"00000066000000000000005c0000000000000065000000000000005f00000000",
            INIT_77 => X"0000004b000000000000004a0000000000000052000000000000005f00000000",
            INIT_78 => X"00000090000000000000008b0000000000000086000000000000008300000000",
            INIT_79 => X"00000098000000000000009a000000000000009f000000000000009800000000",
            INIT_7A => X"0000003900000000000000350000000000000076000000000000009e00000000",
            INIT_7B => X"00000066000000000000005f0000000000000064000000000000006700000000",
            INIT_7C => X"0000006a000000000000006f0000000000000074000000000000006e00000000",
            INIT_7D => X"000000550000000000000057000000000000005b000000000000006100000000",
            INIT_7E => X"0000005300000000000000550000000000000062000000000000005400000000",
            INIT_7F => X"0000005f000000000000005a0000000000000055000000000000005300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE42;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE43 : if BRAM_NAME = "sampleifmap_layersamples_instance43" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a000000000000000980000000000000090000000000000008700000000",
            INIT_01 => X"00000073000000000000008900000000000000a100000000000000a400000000",
            INIT_02 => X"0000006e00000000000000800000000000000091000000000000009d00000000",
            INIT_03 => X"000000670000000000000068000000000000007a000000000000007b00000000",
            INIT_04 => X"00000068000000000000006c000000000000006d000000000000006900000000",
            INIT_05 => X"000000570000000000000058000000000000005a000000000000006100000000",
            INIT_06 => X"000000550000000000000057000000000000005c000000000000004f00000000",
            INIT_07 => X"0000005e00000000000000690000000000000069000000000000006500000000",
            INIT_08 => X"000000a4000000000000009f000000000000009a000000000000009400000000",
            INIT_09 => X"0000007f00000000000000b000000000000000b300000000000000aa00000000",
            INIT_0A => X"00000098000000000000009d00000000000000c500000000000000b000000000",
            INIT_0B => X"0000006700000000000000800000000000000091000000000000007100000000",
            INIT_0C => X"0000006600000000000000680000000000000065000000000000006700000000",
            INIT_0D => X"00000059000000000000005b000000000000005f000000000000006100000000",
            INIT_0E => X"0000005b000000000000005b0000000000000056000000000000004f00000000",
            INIT_0F => X"0000004600000000000000560000000000000068000000000000006d00000000",
            INIT_10 => X"000000c500000000000000b200000000000000a4000000000000009b00000000",
            INIT_11 => X"000000c400000000000000f800000000000000ee00000000000000dd00000000",
            INIT_12 => X"000000b800000000000000b000000000000000c8000000000000009c00000000",
            INIT_13 => X"0000006a0000000000000089000000000000008e000000000000006c00000000",
            INIT_14 => X"0000006500000000000000640000000000000063000000000000006400000000",
            INIT_15 => X"00000059000000000000005f0000000000000063000000000000006500000000",
            INIT_16 => X"00000053000000000000005c0000000000000051000000000000005000000000",
            INIT_17 => X"0000004700000000000000490000000000000052000000000000005800000000",
            INIT_18 => X"000000f900000000000000eb00000000000000d600000000000000bf00000000",
            INIT_19 => X"000000f400000000000000fb00000000000000f600000000000000fd00000000",
            INIT_1A => X"000000c300000000000000ac000000000000009e00000000000000a000000000",
            INIT_1B => X"0000006e000000000000008b0000000000000072000000000000007100000000",
            INIT_1C => X"0000006300000000000000610000000000000062000000000000006200000000",
            INIT_1D => X"0000005c00000000000000660000000000000068000000000000006700000000",
            INIT_1E => X"000000490000000000000055000000000000004e000000000000005300000000",
            INIT_1F => X"00000048000000000000004a0000000000000050000000000000004b00000000",
            INIT_20 => X"000000fe00000000000000fd00000000000000fc00000000000000f500000000",
            INIT_21 => X"000000c900000000000000ba00000000000000bb00000000000000f300000000",
            INIT_22 => X"0000009c00000000000000970000000000000080000000000000009100000000",
            INIT_23 => X"000000720000000000000080000000000000006a000000000000007400000000",
            INIT_24 => X"0000006700000000000000650000000000000067000000000000006800000000",
            INIT_25 => X"0000005c0000000000000069000000000000006e000000000000006c00000000",
            INIT_26 => X"000000550000000000000054000000000000004c000000000000005200000000",
            INIT_27 => X"00000049000000000000004d0000000000000053000000000000004e00000000",
            INIT_28 => X"0000010000000000000000fc00000000000000fc00000000000000fb00000000",
            INIT_29 => X"00000072000000000000006b000000000000007e00000000000000e900000000",
            INIT_2A => X"0000006e00000000000000780000000000000073000000000000006900000000",
            INIT_2B => X"0000006700000000000000680000000000000063000000000000006300000000",
            INIT_2C => X"0000006b000000000000006b000000000000006e000000000000006d00000000",
            INIT_2D => X"000000560000000000000060000000000000006e000000000000007000000000",
            INIT_2E => X"00000068000000000000005a000000000000004c000000000000004e00000000",
            INIT_2F => X"0000004f00000000000000520000000000000052000000000000005b00000000",
            INIT_30 => X"000000eb00000000000000f600000000000000f800000000000000f800000000",
            INIT_31 => X"000000760000000000000072000000000000007c00000000000000c800000000",
            INIT_32 => X"0000004f00000000000000530000000000000057000000000000005d00000000",
            INIT_33 => X"00000044000000000000004b0000000000000056000000000000005000000000",
            INIT_34 => X"0000006100000000000000620000000000000064000000000000005f00000000",
            INIT_35 => X"0000006100000000000000610000000000000061000000000000006200000000",
            INIT_36 => X"0000006f000000000000005b0000000000000057000000000000005b00000000",
            INIT_37 => X"0000005200000000000000520000000000000055000000000000006e00000000",
            INIT_38 => X"0000009600000000000000b500000000000000d600000000000000eb00000000",
            INIT_39 => X"0000008400000000000000850000000000000088000000000000008a00000000",
            INIT_3A => X"0000003c0000000000000039000000000000003d000000000000006400000000",
            INIT_3B => X"0000003a00000000000000600000000000000059000000000000004300000000",
            INIT_3C => X"0000005000000000000000470000000000000045000000000000003300000000",
            INIT_3D => X"0000006500000000000000680000000000000065000000000000005e00000000",
            INIT_3E => X"0000006d000000000000005e0000000000000057000000000000005d00000000",
            INIT_3F => X"0000005100000000000000510000000000000062000000000000007700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000078000000000000007a0000000000000082000000000000009900000000",
            INIT_41 => X"00000067000000000000006f000000000000007a000000000000007c00000000",
            INIT_42 => X"000000340000000000000039000000000000005a000000000000006a00000000",
            INIT_43 => X"00000053000000000000006a0000000000000066000000000000004500000000",
            INIT_44 => X"00000055000000000000004d0000000000000047000000000000004000000000",
            INIT_45 => X"0000006d00000000000000660000000000000067000000000000006400000000",
            INIT_46 => X"00000063000000000000005d0000000000000057000000000000006a00000000",
            INIT_47 => X"00000050000000000000005c0000000000000073000000000000007100000000",
            INIT_48 => X"0000006d0000000000000072000000000000006f000000000000006d00000000",
            INIT_49 => X"0000006d00000000000000660000000000000061000000000000006500000000",
            INIT_4A => X"0000005500000000000000670000000000000078000000000000007500000000",
            INIT_4B => X"00000059000000000000005f0000000000000065000000000000005d00000000",
            INIT_4C => X"0000005a0000000000000052000000000000004b000000000000004a00000000",
            INIT_4D => X"0000006600000000000000690000000000000077000000000000007200000000",
            INIT_4E => X"00000062000000000000005e000000000000006b000000000000006f00000000",
            INIT_4F => X"0000004f000000000000006b0000000000000075000000000000006500000000",
            INIT_50 => X"0000005b000000000000005d0000000000000062000000000000006900000000",
            INIT_51 => X"00000071000000000000006f000000000000006a000000000000006300000000",
            INIT_52 => X"0000005f00000000000000610000000000000068000000000000007000000000",
            INIT_53 => X"0000005c0000000000000054000000000000004c000000000000005000000000",
            INIT_54 => X"00000059000000000000004f0000000000000048000000000000005100000000",
            INIT_55 => X"0000005e0000000000000069000000000000007b000000000000007500000000",
            INIT_56 => X"0000006500000000000000670000000000000067000000000000006000000000",
            INIT_57 => X"0000005a000000000000006f0000000000000069000000000000006000000000",
            INIT_58 => X"00000065000000000000005e0000000000000057000000000000005700000000",
            INIT_59 => X"00000064000000000000006b000000000000006e000000000000006c00000000",
            INIT_5A => X"0000006800000000000000560000000000000051000000000000005b00000000",
            INIT_5B => X"0000005c000000000000004c0000000000000049000000000000005d00000000",
            INIT_5C => X"0000004f000000000000004f000000000000004d000000000000005800000000",
            INIT_5D => X"00000056000000000000005d0000000000000064000000000000005b00000000",
            INIT_5E => X"000000600000000000000061000000000000005c000000000000005700000000",
            INIT_5F => X"0000006500000000000000660000000000000060000000000000006000000000",
            INIT_60 => X"0000006900000000000000670000000000000060000000000000005a00000000",
            INIT_61 => X"000000500000000000000056000000000000005f000000000000006500000000",
            INIT_62 => X"0000006a00000000000000600000000000000055000000000000005100000000",
            INIT_63 => X"0000005d00000000000000600000000000000055000000000000006200000000",
            INIT_64 => X"0000004c000000000000004f0000000000000051000000000000005800000000",
            INIT_65 => X"0000005b0000000000000054000000000000004c000000000000004700000000",
            INIT_66 => X"0000005a00000000000000530000000000000056000000000000005c00000000",
            INIT_67 => X"00000060000000000000005b0000000000000060000000000000006200000000",
            INIT_68 => X"00000056000000000000005f0000000000000063000000000000006400000000",
            INIT_69 => X"0000004f000000000000004f000000000000004f000000000000005000000000",
            INIT_6A => X"0000006c00000000000000620000000000000053000000000000005200000000",
            INIT_6B => X"0000005900000000000000610000000000000060000000000000006300000000",
            INIT_6C => X"00000051000000000000004f0000000000000054000000000000005c00000000",
            INIT_6D => X"000000590000000000000052000000000000004a000000000000004c00000000",
            INIT_6E => X"0000005600000000000000520000000000000055000000000000005a00000000",
            INIT_6F => X"000000530000000000000053000000000000005c000000000000005d00000000",
            INIT_70 => X"000000470000000000000049000000000000004e000000000000005700000000",
            INIT_71 => X"0000005300000000000000590000000000000057000000000000004d00000000",
            INIT_72 => X"0000006a0000000000000061000000000000004f000000000000005100000000",
            INIT_73 => X"0000005c00000000000000590000000000000067000000000000006400000000",
            INIT_74 => X"0000005900000000000000580000000000000057000000000000006000000000",
            INIT_75 => X"000000530000000000000054000000000000004f000000000000005200000000",
            INIT_76 => X"000000530000000000000056000000000000005a000000000000005600000000",
            INIT_77 => X"00000049000000000000004f0000000000000056000000000000005600000000",
            INIT_78 => X"000000490000000000000046000000000000003f000000000000003e00000000",
            INIT_79 => X"0000005100000000000000530000000000000056000000000000005400000000",
            INIT_7A => X"0000006b000000000000005e000000000000004a000000000000004e00000000",
            INIT_7B => X"00000058000000000000005b0000000000000068000000000000005f00000000",
            INIT_7C => X"0000005900000000000000580000000000000058000000000000005b00000000",
            INIT_7D => X"0000005300000000000000550000000000000050000000000000005500000000",
            INIT_7E => X"0000005000000000000000560000000000000059000000000000005400000000",
            INIT_7F => X"00000048000000000000004c000000000000004d000000000000004c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE43;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE44 : if BRAM_NAME = "sampleifmap_layersamples_instance44" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000059000000000000005d000000000000005e000000000000005e00000000",
            INIT_01 => X"000000600000000000000060000000000000005a000000000000005a00000000",
            INIT_02 => X"00000065000000000000006e0000000000000066000000000000006100000000",
            INIT_03 => X"0000005200000000000000550000000000000058000000000000005e00000000",
            INIT_04 => X"000000480000000000000049000000000000004b000000000000004e00000000",
            INIT_05 => X"00000038000000000000003d0000000000000041000000000000004500000000",
            INIT_06 => X"000000270000000000000029000000000000002e000000000000003300000000",
            INIT_07 => X"00000019000000000000001d0000000000000022000000000000002800000000",
            INIT_08 => X"00000059000000000000005f000000000000005f000000000000006000000000",
            INIT_09 => X"00000062000000000000005f0000000000000059000000000000005900000000",
            INIT_0A => X"0000006b000000000000006a0000000000000060000000000000006100000000",
            INIT_0B => X"0000005200000000000000550000000000000059000000000000006000000000",
            INIT_0C => X"000000490000000000000047000000000000004b000000000000004f00000000",
            INIT_0D => X"00000035000000000000003b000000000000003d000000000000004400000000",
            INIT_0E => X"000000250000000000000027000000000000002c000000000000003100000000",
            INIT_0F => X"0000001f000000000000001f0000000000000020000000000000002600000000",
            INIT_10 => X"00000057000000000000005c000000000000005c000000000000005e00000000",
            INIT_11 => X"00000051000000000000005d000000000000005a000000000000005400000000",
            INIT_12 => X"0000006e00000000000000630000000000000060000000000000005900000000",
            INIT_13 => X"0000005400000000000000560000000000000062000000000000007000000000",
            INIT_14 => X"0000004600000000000000440000000000000049000000000000004f00000000",
            INIT_15 => X"000000300000000000000036000000000000003a000000000000003f00000000",
            INIT_16 => X"0000002b0000000000000029000000000000002b000000000000002e00000000",
            INIT_17 => X"000000310000000000000030000000000000002e000000000000002f00000000",
            INIT_18 => X"0000005a000000000000005c000000000000005d000000000000005f00000000",
            INIT_19 => X"000000390000000000000056000000000000005d000000000000005300000000",
            INIT_1A => X"000000680000000000000063000000000000006b000000000000005d00000000",
            INIT_1B => X"0000005a00000000000000650000000000000072000000000000007400000000",
            INIT_1C => X"0000004200000000000000420000000000000043000000000000004e00000000",
            INIT_1D => X"0000003900000000000000380000000000000038000000000000003e00000000",
            INIT_1E => X"000000420000000000000041000000000000003e000000000000003c00000000",
            INIT_1F => X"0000003d000000000000003f0000000000000041000000000000004300000000",
            INIT_20 => X"0000005b000000000000005b000000000000005b000000000000005c00000000",
            INIT_21 => X"0000003e00000000000000520000000000000059000000000000005300000000",
            INIT_22 => X"000000580000000000000058000000000000005f000000000000005c00000000",
            INIT_23 => X"0000006400000000000000690000000000000068000000000000005c00000000",
            INIT_24 => X"0000004800000000000000450000000000000046000000000000005b00000000",
            INIT_25 => X"000000530000000000000050000000000000004d000000000000005000000000",
            INIT_26 => X"0000005000000000000000510000000000000051000000000000005300000000",
            INIT_27 => X"0000003f0000000000000046000000000000004b000000000000004f00000000",
            INIT_28 => X"0000005900000000000000570000000000000056000000000000005800000000",
            INIT_29 => X"0000004d000000000000004c000000000000004f000000000000005200000000",
            INIT_2A => X"0000005700000000000000550000000000000052000000000000005000000000",
            INIT_2B => X"0000005f000000000000005e000000000000005e000000000000005a00000000",
            INIT_2C => X"000000630000000000000062000000000000005e000000000000006300000000",
            INIT_2D => X"0000006200000000000000600000000000000064000000000000006400000000",
            INIT_2E => X"0000005300000000000000580000000000000058000000000000005d00000000",
            INIT_2F => X"00000037000000000000003e0000000000000045000000000000004c00000000",
            INIT_30 => X"0000005400000000000000520000000000000054000000000000005500000000",
            INIT_31 => X"00000037000000000000002a000000000000003d000000000000005100000000",
            INIT_32 => X"0000005900000000000000580000000000000057000000000000005300000000",
            INIT_33 => X"00000065000000000000005d0000000000000057000000000000005b00000000",
            INIT_34 => X"0000007300000000000000700000000000000064000000000000006200000000",
            INIT_35 => X"0000006700000000000000670000000000000067000000000000006900000000",
            INIT_36 => X"0000004a000000000000004e0000000000000050000000000000005b00000000",
            INIT_37 => X"000000360000000000000039000000000000003f000000000000004400000000",
            INIT_38 => X"0000005400000000000000520000000000000053000000000000005200000000",
            INIT_39 => X"0000002c00000000000000260000000000000037000000000000004c00000000",
            INIT_3A => X"0000005100000000000000520000000000000055000000000000004c00000000",
            INIT_3B => X"00000063000000000000005b0000000000000053000000000000005000000000",
            INIT_3C => X"0000006c00000000000000610000000000000060000000000000006700000000",
            INIT_3D => X"0000005e00000000000000710000000000000072000000000000006d00000000",
            INIT_3E => X"0000004b000000000000004d000000000000004d000000000000005200000000",
            INIT_3F => X"0000003b00000000000000400000000000000044000000000000004700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005b00000000000000540000000000000052000000000000005100000000",
            INIT_41 => X"0000003100000000000000550000000000000068000000000000005e00000000",
            INIT_42 => X"00000063000000000000005b0000000000000054000000000000004900000000",
            INIT_43 => X"0000005e00000000000000650000000000000064000000000000006100000000",
            INIT_44 => X"0000006200000000000000650000000000000068000000000000006500000000",
            INIT_45 => X"000000670000000000000072000000000000006f000000000000006a00000000",
            INIT_46 => X"0000004e00000000000000520000000000000055000000000000005700000000",
            INIT_47 => X"0000004800000000000000470000000000000046000000000000004a00000000",
            INIT_48 => X"0000008000000000000000730000000000000065000000000000005c00000000",
            INIT_49 => X"000000360000000000000068000000000000009d000000000000008e00000000",
            INIT_4A => X"00000071000000000000005d0000000000000054000000000000004b00000000",
            INIT_4B => X"000000650000000000000075000000000000007c000000000000007500000000",
            INIT_4C => X"00000067000000000000006b000000000000006a000000000000006700000000",
            INIT_4D => X"000000760000000000000074000000000000006e000000000000006800000000",
            INIT_4E => X"000000540000000000000055000000000000005a000000000000006400000000",
            INIT_4F => X"0000005200000000000000550000000000000055000000000000005500000000",
            INIT_50 => X"000000a00000000000000099000000000000008e000000000000008200000000",
            INIT_51 => X"00000035000000000000005900000000000000aa00000000000000a600000000",
            INIT_52 => X"000000680000000000000046000000000000004d000000000000005000000000",
            INIT_53 => X"0000006b000000000000007f0000000000000082000000000000007700000000",
            INIT_54 => X"0000006a0000000000000069000000000000006c000000000000006a00000000",
            INIT_55 => X"00000072000000000000006e0000000000000069000000000000006a00000000",
            INIT_56 => X"0000006000000000000000620000000000000062000000000000006900000000",
            INIT_57 => X"000000550000000000000059000000000000005b000000000000005e00000000",
            INIT_58 => X"000000a400000000000000a2000000000000009f000000000000009a00000000",
            INIT_59 => X"0000002e000000000000005d00000000000000a900000000000000a700000000",
            INIT_5A => X"00000067000000000000004a0000000000000056000000000000005100000000",
            INIT_5B => X"00000072000000000000007a0000000000000070000000000000007b00000000",
            INIT_5C => X"00000067000000000000006a000000000000006d000000000000006a00000000",
            INIT_5D => X"0000006e00000000000000670000000000000069000000000000006b00000000",
            INIT_5E => X"0000006300000000000000650000000000000061000000000000006600000000",
            INIT_5F => X"00000055000000000000005a000000000000005e000000000000006000000000",
            INIT_60 => X"0000009e00000000000000a1000000000000009f000000000000009d00000000",
            INIT_61 => X"000000300000000000000075000000000000009f000000000000009e00000000",
            INIT_62 => X"00000078000000000000006c0000000000000065000000000000004900000000",
            INIT_63 => X"0000007500000000000000740000000000000078000000000000008700000000",
            INIT_64 => X"00000066000000000000006c0000000000000073000000000000006b00000000",
            INIT_65 => X"000000690000000000000064000000000000006a000000000000006900000000",
            INIT_66 => X"0000006500000000000000600000000000000060000000000000007000000000",
            INIT_67 => X"0000004c0000000000000055000000000000005d000000000000006200000000",
            INIT_68 => X"0000009300000000000000970000000000000098000000000000009900000000",
            INIT_69 => X"0000004c00000000000000870000000000000093000000000000009300000000",
            INIT_6A => X"0000007500000000000000670000000000000049000000000000002c00000000",
            INIT_6B => X"0000007100000000000000730000000000000085000000000000008300000000",
            INIT_6C => X"0000006b00000000000000710000000000000077000000000000006c00000000",
            INIT_6D => X"000000640000000000000065000000000000006a000000000000006a00000000",
            INIT_6E => X"00000062000000000000005d0000000000000069000000000000007500000000",
            INIT_6F => X"00000040000000000000004a0000000000000055000000000000005d00000000",
            INIT_70 => X"0000008e000000000000008e000000000000008e000000000000008f00000000",
            INIT_71 => X"0000008300000000000000950000000000000094000000000000008f00000000",
            INIT_72 => X"0000004600000000000000350000000000000041000000000000005400000000",
            INIT_73 => X"0000006d0000000000000068000000000000006b000000000000006300000000",
            INIT_74 => X"00000075000000000000007d000000000000007c000000000000007200000000",
            INIT_75 => X"000000620000000000000065000000000000006c000000000000006e00000000",
            INIT_76 => X"0000005a0000000000000058000000000000006f000000000000006c00000000",
            INIT_77 => X"0000003f00000000000000410000000000000048000000000000005500000000",
            INIT_78 => X"00000091000000000000008e000000000000008d000000000000008c00000000",
            INIT_79 => X"00000093000000000000009900000000000000a0000000000000009900000000",
            INIT_7A => X"0000003a0000000000000034000000000000006f000000000000009700000000",
            INIT_7B => X"0000006e00000000000000650000000000000068000000000000006a00000000",
            INIT_7C => X"0000008000000000000000870000000000000089000000000000007b00000000",
            INIT_7D => X"000000650000000000000068000000000000006c000000000000007300000000",
            INIT_7E => X"0000004e0000000000000059000000000000006f000000000000006300000000",
            INIT_7F => X"0000004d000000000000004a0000000000000048000000000000004a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE44;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE45 : if BRAM_NAME = "sampleifmap_layersamples_instance45" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009f000000000000009b0000000000000095000000000000008f00000000",
            INIT_01 => X"00000072000000000000008800000000000000a000000000000000a400000000",
            INIT_02 => X"00000068000000000000007a000000000000008f000000000000009b00000000",
            INIT_03 => X"0000006c00000000000000660000000000000077000000000000007600000000",
            INIT_04 => X"0000008000000000000000850000000000000084000000000000007800000000",
            INIT_05 => X"0000006a000000000000006b000000000000006d000000000000007500000000",
            INIT_06 => X"000000560000000000000062000000000000006c000000000000006100000000",
            INIT_07 => X"00000044000000000000004f0000000000000054000000000000005a00000000",
            INIT_08 => X"000000a1000000000000009f000000000000009d000000000000009a00000000",
            INIT_09 => X"0000008100000000000000b000000000000000b100000000000000a700000000",
            INIT_0A => X"0000008e000000000000009700000000000000c700000000000000b300000000",
            INIT_0B => X"0000006c000000000000007b0000000000000089000000000000006800000000",
            INIT_0C => X"000000800000000000000083000000000000007e000000000000007900000000",
            INIT_0D => X"0000006e00000000000000700000000000000073000000000000007700000000",
            INIT_0E => X"0000005e000000000000006a0000000000000069000000000000006300000000",
            INIT_0F => X"000000270000000000000034000000000000004a000000000000005c00000000",
            INIT_10 => X"000000c100000000000000b000000000000000a4000000000000009d00000000",
            INIT_11 => X"000000c700000000000000f700000000000000ec00000000000000da00000000",
            INIT_12 => X"000000b100000000000000ad00000000000000ce00000000000000a300000000",
            INIT_13 => X"0000007100000000000000860000000000000088000000000000006500000000",
            INIT_14 => X"000000810000000000000082000000000000007e000000000000007700000000",
            INIT_15 => X"000000710000000000000076000000000000007a000000000000007d00000000",
            INIT_16 => X"00000050000000000000006a0000000000000067000000000000006800000000",
            INIT_17 => X"000000270000000000000025000000000000002c000000000000003e00000000",
            INIT_18 => X"000000f600000000000000e800000000000000d400000000000000c000000000",
            INIT_19 => X"000000f700000000000000fa00000000000000f200000000000000fa00000000",
            INIT_1A => X"000000c100000000000000ae00000000000000aa00000000000000a900000000",
            INIT_1B => X"00000078000000000000008b0000000000000070000000000000006e00000000",
            INIT_1C => X"000000800000000000000080000000000000007e000000000000007600000000",
            INIT_1D => X"00000074000000000000007e000000000000007f000000000000008000000000",
            INIT_1E => X"0000003e00000000000000600000000000000066000000000000006c00000000",
            INIT_1F => X"0000002b00000000000000270000000000000025000000000000002a00000000",
            INIT_20 => X"000000fb00000000000000fa00000000000000fb00000000000000f500000000",
            INIT_21 => X"000000d200000000000000be00000000000000ba00000000000000f100000000",
            INIT_22 => X"000000a0000000000000009c000000000000009200000000000000a100000000",
            INIT_23 => X"0000007a00000000000000870000000000000073000000000000007d00000000",
            INIT_24 => X"000000800000000000000081000000000000007f000000000000007800000000",
            INIT_25 => X"00000074000000000000007d000000000000007f000000000000007f00000000",
            INIT_26 => X"0000004200000000000000570000000000000062000000000000006a00000000",
            INIT_27 => X"000000290000000000000029000000000000002a000000000000002d00000000",
            INIT_28 => X"000000fe00000000000000fb00000000000000fb00000000000000fb00000000",
            INIT_29 => X"000000820000000000000074000000000000008300000000000000ea00000000",
            INIT_2A => X"0000007c0000000000000082000000000000008a000000000000007f00000000",
            INIT_2B => X"0000006b00000000000000720000000000000077000000000000007a00000000",
            INIT_2C => X"0000007f00000000000000820000000000000080000000000000007600000000",
            INIT_2D => X"0000006c000000000000006f0000000000000077000000000000007d00000000",
            INIT_2E => X"000000500000000000000052000000000000005a000000000000006300000000",
            INIT_2F => X"00000029000000000000002c000000000000002f000000000000003d00000000",
            INIT_30 => X"000000ef00000000000000f900000000000000fc00000000000000fc00000000",
            INIT_31 => X"00000083000000000000007b000000000000008000000000000000cb00000000",
            INIT_32 => X"000000670000000000000066000000000000006c000000000000006f00000000",
            INIT_33 => X"0000004400000000000000510000000000000069000000000000006a00000000",
            INIT_34 => X"0000007400000000000000780000000000000075000000000000006600000000",
            INIT_35 => X"000000730000000000000070000000000000006b000000000000006e00000000",
            INIT_36 => X"00000054000000000000004b0000000000000059000000000000006800000000",
            INIT_37 => X"0000002d000000000000002d0000000000000034000000000000005100000000",
            INIT_38 => X"000000a000000000000000bf00000000000000df00000000000000f500000000",
            INIT_39 => X"0000008a00000000000000890000000000000089000000000000009000000000",
            INIT_3A => X"000000570000000000000051000000000000004b000000000000006d00000000",
            INIT_3B => X"0000003a00000000000000630000000000000066000000000000005a00000000",
            INIT_3C => X"00000065000000000000005f0000000000000056000000000000003a00000000",
            INIT_3D => X"00000074000000000000007a0000000000000074000000000000006d00000000",
            INIT_3E => X"000000500000000000000046000000000000004d000000000000006100000000",
            INIT_3F => X"0000002f000000000000002f0000000000000042000000000000005900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000840000000000000086000000000000008d00000000000000a500000000",
            INIT_41 => X"000000690000000000000070000000000000007b000000000000008200000000",
            INIT_42 => X"00000047000000000000004a000000000000005e000000000000006b00000000",
            INIT_43 => X"00000056000000000000006f000000000000006e000000000000005300000000",
            INIT_44 => X"0000006c0000000000000066000000000000005a000000000000004800000000",
            INIT_45 => X"0000007c000000000000007b000000000000007b000000000000007600000000",
            INIT_46 => X"0000004400000000000000420000000000000049000000000000006c00000000",
            INIT_47 => X"00000030000000000000003d0000000000000054000000000000005200000000",
            INIT_48 => X"00000075000000000000007a0000000000000078000000000000007500000000",
            INIT_49 => X"0000006a00000000000000650000000000000061000000000000006a00000000",
            INIT_4A => X"00000057000000000000006a0000000000000073000000000000007000000000",
            INIT_4B => X"0000006100000000000000680000000000000068000000000000005c00000000",
            INIT_4C => X"00000072000000000000006c000000000000005f000000000000005400000000",
            INIT_4D => X"0000007a0000000000000082000000000000008e000000000000008600000000",
            INIT_4E => X"0000004000000000000000450000000000000064000000000000007700000000",
            INIT_4F => X"00000032000000000000004f0000000000000057000000000000004500000000",
            INIT_50 => X"0000005e00000000000000600000000000000066000000000000006c00000000",
            INIT_51 => X"0000006b000000000000006e000000000000006b000000000000006500000000",
            INIT_52 => X"000000510000000000000056000000000000005d000000000000006700000000",
            INIT_53 => X"00000068000000000000005d0000000000000048000000000000004200000000",
            INIT_54 => X"00000071000000000000006b000000000000005f000000000000005e00000000",
            INIT_55 => X"0000007a00000000000000850000000000000094000000000000008900000000",
            INIT_56 => X"000000420000000000000051000000000000006b000000000000007200000000",
            INIT_57 => X"0000003f0000000000000055000000000000004b000000000000004000000000",
            INIT_58 => X"00000063000000000000005d0000000000000057000000000000005800000000",
            INIT_59 => X"000000570000000000000065000000000000006c000000000000006b00000000",
            INIT_5A => X"000000530000000000000041000000000000003c000000000000004900000000",
            INIT_5B => X"0000005e000000000000004e000000000000003f000000000000004a00000000",
            INIT_5C => X"0000005d000000000000005f0000000000000057000000000000005900000000",
            INIT_5D => X"00000072000000000000007a000000000000007b000000000000006900000000",
            INIT_5E => X"0000003b000000000000004e0000000000000068000000000000006d00000000",
            INIT_5F => X"0000004b000000000000004a000000000000003f000000000000003c00000000",
            INIT_60 => X"0000005f0000000000000061000000000000005f000000000000005d00000000",
            INIT_61 => X"0000003800000000000000450000000000000054000000000000005b00000000",
            INIT_62 => X"0000005500000000000000420000000000000031000000000000003200000000",
            INIT_63 => X"0000004800000000000000550000000000000049000000000000005300000000",
            INIT_64 => X"000000440000000000000043000000000000003e000000000000003e00000000",
            INIT_65 => X"0000006800000000000000640000000000000058000000000000004500000000",
            INIT_66 => X"000000330000000000000040000000000000005a000000000000006500000000",
            INIT_67 => X"00000045000000000000003a0000000000000036000000000000003500000000",
            INIT_68 => X"000000440000000000000051000000000000005b000000000000006000000000",
            INIT_69 => X"0000003000000000000000340000000000000037000000000000003b00000000",
            INIT_6A => X"000000520000000000000040000000000000002e000000000000002f00000000",
            INIT_6B => X"00000039000000000000004d000000000000004f000000000000005200000000",
            INIT_6C => X"0000003a00000000000000340000000000000032000000000000003500000000",
            INIT_6D => X"0000004a0000000000000047000000000000003f000000000000003a00000000",
            INIT_6E => X"0000002e00000000000000340000000000000041000000000000004800000000",
            INIT_6F => X"0000003600000000000000300000000000000031000000000000003000000000",
            INIT_70 => X"0000002b0000000000000031000000000000003c000000000000004900000000",
            INIT_71 => X"0000003000000000000000340000000000000030000000000000002c00000000",
            INIT_72 => X"00000049000000000000003a000000000000002c000000000000003000000000",
            INIT_73 => X"00000035000000000000003e000000000000004f000000000000004b00000000",
            INIT_74 => X"000000390000000000000034000000000000002e000000000000003200000000",
            INIT_75 => X"0000002f0000000000000033000000000000002f000000000000003400000000",
            INIT_76 => X"0000002a000000000000002e0000000000000031000000000000002f00000000",
            INIT_77 => X"0000002a000000000000002b000000000000002d000000000000002b00000000",
            INIT_78 => X"0000002500000000000000270000000000000025000000000000002900000000",
            INIT_79 => X"0000002d00000000000000290000000000000029000000000000002a00000000",
            INIT_7A => X"000000470000000000000036000000000000002b000000000000002f00000000",
            INIT_7B => X"0000002e000000000000003b000000000000004c000000000000004300000000",
            INIT_7C => X"00000030000000000000002d000000000000002a000000000000002b00000000",
            INIT_7D => X"0000002d0000000000000031000000000000002d000000000000002f00000000",
            INIT_7E => X"00000027000000000000002a000000000000002d000000000000002b00000000",
            INIT_7F => X"0000002600000000000000280000000000000028000000000000002500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE45;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE46 : if BRAM_NAME = "sampleifmap_layersamples_instance46" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004f00000000000000530000000000000054000000000000005500000000",
            INIT_01 => X"0000005f000000000000005d0000000000000052000000000000005000000000",
            INIT_02 => X"00000048000000000000004f0000000000000055000000000000005a00000000",
            INIT_03 => X"0000004f0000000000000054000000000000004e000000000000004b00000000",
            INIT_04 => X"0000003d000000000000003c000000000000003e000000000000004400000000",
            INIT_05 => X"000000330000000000000038000000000000003b000000000000003c00000000",
            INIT_06 => X"0000002300000000000000250000000000000029000000000000002e00000000",
            INIT_07 => X"000000150000000000000019000000000000001e000000000000002400000000",
            INIT_08 => X"0000004f00000000000000550000000000000055000000000000005600000000",
            INIT_09 => X"0000005d000000000000005a0000000000000050000000000000004e00000000",
            INIT_0A => X"0000004700000000000000460000000000000049000000000000005400000000",
            INIT_0B => X"0000004800000000000000470000000000000045000000000000004400000000",
            INIT_0C => X"0000003e000000000000003e0000000000000043000000000000004600000000",
            INIT_0D => X"0000002e00000000000000340000000000000035000000000000003800000000",
            INIT_0E => X"0000002000000000000000220000000000000025000000000000002900000000",
            INIT_0F => X"0000001b000000000000001a000000000000001b000000000000002100000000",
            INIT_10 => X"0000004e00000000000000520000000000000053000000000000005400000000",
            INIT_11 => X"0000004800000000000000560000000000000050000000000000004900000000",
            INIT_12 => X"0000004300000000000000380000000000000041000000000000004600000000",
            INIT_13 => X"0000003c0000000000000036000000000000003f000000000000004800000000",
            INIT_14 => X"0000003a000000000000003d0000000000000041000000000000004200000000",
            INIT_15 => X"00000026000000000000002d000000000000002f000000000000003000000000",
            INIT_16 => X"0000002500000000000000220000000000000021000000000000002400000000",
            INIT_17 => X"0000002c000000000000002a0000000000000029000000000000002a00000000",
            INIT_18 => X"0000005000000000000000520000000000000053000000000000005500000000",
            INIT_19 => X"0000002b000000000000004d0000000000000052000000000000004800000000",
            INIT_1A => X"0000003400000000000000320000000000000045000000000000004300000000",
            INIT_1B => X"0000002f0000000000000032000000000000003f000000000000004100000000",
            INIT_1C => X"0000003600000000000000390000000000000034000000000000003200000000",
            INIT_1D => X"0000002c000000000000002b000000000000002b000000000000002d00000000",
            INIT_1E => X"0000003b00000000000000380000000000000032000000000000002f00000000",
            INIT_1F => X"000000370000000000000038000000000000003b000000000000003c00000000",
            INIT_20 => X"0000005100000000000000510000000000000051000000000000005200000000",
            INIT_21 => X"0000002c0000000000000046000000000000004c000000000000004800000000",
            INIT_22 => X"0000001d00000000000000220000000000000033000000000000003d00000000",
            INIT_23 => X"0000002300000000000000260000000000000027000000000000001f00000000",
            INIT_24 => X"0000003b0000000000000039000000000000002b000000000000002900000000",
            INIT_25 => X"000000440000000000000041000000000000003d000000000000003d00000000",
            INIT_26 => X"0000004800000000000000470000000000000042000000000000004400000000",
            INIT_27 => X"00000038000000000000003e0000000000000043000000000000004700000000",
            INIT_28 => X"0000004f000000000000004c000000000000004c000000000000004d00000000",
            INIT_29 => X"00000038000000000000003e0000000000000042000000000000004700000000",
            INIT_2A => X"00000017000000000000001a0000000000000021000000000000002c00000000",
            INIT_2B => X"0000000e000000000000000f0000000000000014000000000000001600000000",
            INIT_2C => X"00000054000000000000004f0000000000000035000000000000001f00000000",
            INIT_2D => X"00000050000000000000004e0000000000000052000000000000005300000000",
            INIT_2E => X"0000004b000000000000004d0000000000000048000000000000004c00000000",
            INIT_2F => X"0000002e0000000000000035000000000000003c000000000000004400000000",
            INIT_30 => X"0000004800000000000000460000000000000047000000000000004900000000",
            INIT_31 => X"0000002000000000000000200000000000000037000000000000004700000000",
            INIT_32 => X"0000001300000000000000140000000000000018000000000000002600000000",
            INIT_33 => X"00000015000000000000000e000000000000000b000000000000001200000000",
            INIT_34 => X"0000005900000000000000460000000000000029000000000000001800000000",
            INIT_35 => X"00000052000000000000004f0000000000000050000000000000005600000000",
            INIT_36 => X"0000004300000000000000480000000000000048000000000000004b00000000",
            INIT_37 => X"0000002a000000000000002d0000000000000034000000000000003b00000000",
            INIT_38 => X"0000004500000000000000440000000000000045000000000000004400000000",
            INIT_39 => X"00000011000000000000001c0000000000000033000000000000004300000000",
            INIT_3A => X"0000000b000000000000000a000000000000000c000000000000001700000000",
            INIT_3B => X"000000180000000000000011000000000000000b000000000000000900000000",
            INIT_3C => X"0000003f00000000000000210000000000000016000000000000001c00000000",
            INIT_3D => X"00000040000000000000004d000000000000004f000000000000004d00000000",
            INIT_3E => X"0000004200000000000000480000000000000049000000000000004100000000",
            INIT_3F => X"0000002b000000000000002f0000000000000036000000000000003c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004e00000000000000470000000000000045000000000000004400000000",
            INIT_41 => X"000000130000000000000046000000000000005d000000000000005200000000",
            INIT_42 => X"000000250000000000000019000000000000000c000000000000001200000000",
            INIT_43 => X"0000001400000000000000210000000000000021000000000000002000000000",
            INIT_44 => X"0000002100000000000000190000000000000018000000000000001600000000",
            INIT_45 => X"0000003b000000000000003c0000000000000038000000000000003100000000",
            INIT_46 => X"0000003f0000000000000049000000000000004b000000000000003b00000000",
            INIT_47 => X"0000003500000000000000340000000000000034000000000000003900000000",
            INIT_48 => X"0000007500000000000000670000000000000059000000000000005000000000",
            INIT_49 => X"000000160000000000000055000000000000008d000000000000008000000000",
            INIT_4A => X"000000380000000000000021000000000000000f000000000000001500000000",
            INIT_4B => X"0000001c0000000000000035000000000000003d000000000000003900000000",
            INIT_4C => X"0000001400000000000000160000000000000016000000000000001500000000",
            INIT_4D => X"0000003a000000000000002d0000000000000023000000000000001800000000",
            INIT_4E => X"0000004100000000000000460000000000000048000000000000003d00000000",
            INIT_4F => X"0000003d000000000000003f0000000000000040000000000000004100000000",
            INIT_50 => X"00000095000000000000008e0000000000000083000000000000007700000000",
            INIT_51 => X"0000001800000000000000470000000000000098000000000000009800000000",
            INIT_52 => X"0000003100000000000000150000000000000011000000000000001e00000000",
            INIT_53 => X"00000021000000000000003f0000000000000044000000000000003c00000000",
            INIT_54 => X"000000110000000000000015000000000000001b000000000000001900000000",
            INIT_55 => X"0000002b000000000000001c0000000000000014000000000000000f00000000",
            INIT_56 => X"0000004a000000000000004d0000000000000046000000000000003700000000",
            INIT_57 => X"0000004100000000000000440000000000000047000000000000004900000000",
            INIT_58 => X"0000009900000000000000960000000000000094000000000000008f00000000",
            INIT_59 => X"00000017000000000000004f0000000000000099000000000000009900000000",
            INIT_5A => X"0000002e00000000000000190000000000000022000000000000002800000000",
            INIT_5B => X"0000002700000000000000370000000000000030000000000000003d00000000",
            INIT_5C => X"00000015000000000000001f0000000000000024000000000000001d00000000",
            INIT_5D => X"0000001f00000000000000120000000000000015000000000000001300000000",
            INIT_5E => X"0000004d000000000000004c000000000000003b000000000000002a00000000",
            INIT_5F => X"00000045000000000000004a000000000000004c000000000000004d00000000",
            INIT_60 => X"0000009400000000000000970000000000000095000000000000009200000000",
            INIT_61 => X"00000020000000000000006b0000000000000092000000000000009200000000",
            INIT_62 => X"0000003b00000000000000340000000000000037000000000000002b00000000",
            INIT_63 => X"00000029000000000000002c0000000000000034000000000000004700000000",
            INIT_64 => X"0000001e000000000000002c0000000000000032000000000000002200000000",
            INIT_65 => X"000000190000000000000012000000000000001c000000000000001a00000000",
            INIT_66 => X"0000005100000000000000450000000000000032000000000000002e00000000",
            INIT_67 => X"000000420000000000000049000000000000004f000000000000005100000000",
            INIT_68 => X"0000008b000000000000008f000000000000008f000000000000009000000000",
            INIT_69 => X"00000040000000000000007e0000000000000089000000000000008a00000000",
            INIT_6A => X"00000041000000000000003d000000000000002e000000000000001a00000000",
            INIT_6B => X"0000002400000000000000280000000000000040000000000000004600000000",
            INIT_6C => X"0000002800000000000000330000000000000036000000000000002400000000",
            INIT_6D => X"000000130000000000000012000000000000001d000000000000002100000000",
            INIT_6E => X"0000004e000000000000003c0000000000000033000000000000002f00000000",
            INIT_6F => X"000000370000000000000040000000000000004a000000000000004f00000000",
            INIT_70 => X"0000008600000000000000860000000000000084000000000000008500000000",
            INIT_71 => X"0000007700000000000000890000000000000088000000000000008600000000",
            INIT_72 => X"00000021000000000000001b0000000000000031000000000000004700000000",
            INIT_73 => X"000000220000000000000020000000000000002a000000000000002e00000000",
            INIT_74 => X"00000032000000000000003d0000000000000039000000000000002800000000",
            INIT_75 => X"000000110000000000000011000000000000001c000000000000002700000000",
            INIT_76 => X"0000004100000000000000300000000000000033000000000000002400000000",
            INIT_77 => X"000000320000000000000036000000000000003e000000000000004600000000",
            INIT_78 => X"000000850000000000000081000000000000007f000000000000007d00000000",
            INIT_79 => X"0000008100000000000000880000000000000091000000000000008c00000000",
            INIT_7A => X"0000001e000000000000001e000000000000005a000000000000008400000000",
            INIT_7B => X"0000002700000000000000270000000000000033000000000000004000000000",
            INIT_7C => X"0000003d00000000000000450000000000000045000000000000003100000000",
            INIT_7D => X"000000130000000000000014000000000000001c000000000000002c00000000",
            INIT_7E => X"0000002d00000000000000290000000000000030000000000000001900000000",
            INIT_7F => X"0000003d000000000000003c0000000000000039000000000000003500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE46;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE47 : if BRAM_NAME = "sampleifmap_layersamples_instance47" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000091000000000000008b0000000000000084000000000000007d00000000",
            INIT_01 => X"0000005a00000000000000750000000000000091000000000000009500000000",
            INIT_02 => X"0000005000000000000000620000000000000072000000000000008000000000",
            INIT_03 => X"000000280000000000000031000000000000004d000000000000005700000000",
            INIT_04 => X"0000003c0000000000000044000000000000003f000000000000002e00000000",
            INIT_05 => X"000000170000000000000019000000000000001f000000000000002d00000000",
            INIT_06 => X"0000002d000000000000002b000000000000002a000000000000001500000000",
            INIT_07 => X"00000032000000000000003e0000000000000042000000000000004000000000",
            INIT_08 => X"000000930000000000000090000000000000008c000000000000008800000000",
            INIT_09 => X"00000068000000000000009e00000000000000a4000000000000009a00000000",
            INIT_0A => X"00000077000000000000007a00000000000000a6000000000000009500000000",
            INIT_0B => X"00000029000000000000004b0000000000000067000000000000005000000000",
            INIT_0C => X"0000003c00000000000000410000000000000038000000000000002d00000000",
            INIT_0D => X"0000001b000000000000001f0000000000000028000000000000003000000000",
            INIT_0E => X"00000032000000000000002f0000000000000023000000000000001500000000",
            INIT_0F => X"0000001400000000000000230000000000000039000000000000004100000000",
            INIT_10 => X"000000b600000000000000a40000000000000097000000000000009000000000",
            INIT_11 => X"000000b200000000000000eb00000000000000e600000000000000d200000000",
            INIT_12 => X"00000095000000000000008a00000000000000ab000000000000008500000000",
            INIT_13 => X"0000002d00000000000000550000000000000067000000000000004d00000000",
            INIT_14 => X"0000003c000000000000003f0000000000000038000000000000002b00000000",
            INIT_15 => X"0000001d00000000000000270000000000000030000000000000003500000000",
            INIT_16 => X"00000027000000000000002f000000000000001d000000000000001700000000",
            INIT_17 => X"000000150000000000000016000000000000001f000000000000002700000000",
            INIT_18 => X"000000f000000000000000e100000000000000cd00000000000000b700000000",
            INIT_19 => X"000000e600000000000000f200000000000000f200000000000000f800000000",
            INIT_1A => X"0000009f00000000000000840000000000000084000000000000008d00000000",
            INIT_1B => X"000000310000000000000056000000000000004d000000000000005300000000",
            INIT_1C => X"0000003a000000000000003c0000000000000037000000000000002a00000000",
            INIT_1D => X"00000021000000000000002f0000000000000037000000000000003900000000",
            INIT_1E => X"0000001c0000000000000027000000000000001a000000000000001900000000",
            INIT_1F => X"0000001b000000000000001c000000000000001d000000000000001900000000",
            INIT_20 => X"000000f900000000000000f700000000000000f800000000000000f100000000",
            INIT_21 => X"000000b500000000000000ab00000000000000b000000000000000ec00000000",
            INIT_22 => X"0000007600000000000000720000000000000062000000000000007800000000",
            INIT_23 => X"000000340000000000000047000000000000003c000000000000004d00000000",
            INIT_24 => X"0000003a00000000000000390000000000000036000000000000002e00000000",
            INIT_25 => X"0000002000000000000000300000000000000039000000000000003b00000000",
            INIT_26 => X"0000002500000000000000250000000000000017000000000000001800000000",
            INIT_27 => X"0000001a000000000000001f0000000000000020000000000000001c00000000",
            INIT_28 => X"000000fd00000000000000f900000000000000f900000000000000f800000000",
            INIT_29 => X"000000550000000000000053000000000000006a00000000000000e000000000",
            INIT_2A => X"000000410000000000000051000000000000004e000000000000004700000000",
            INIT_2B => X"000000310000000000000034000000000000002e000000000000003000000000",
            INIT_2C => X"0000003900000000000000360000000000000037000000000000003300000000",
            INIT_2D => X"0000001b00000000000000240000000000000033000000000000003d00000000",
            INIT_2E => X"0000003600000000000000270000000000000016000000000000001500000000",
            INIT_2F => X"0000001c000000000000001f000000000000001f000000000000002800000000",
            INIT_30 => X"000000eb00000000000000f500000000000000f800000000000000f700000000",
            INIT_31 => X"0000005e0000000000000060000000000000006d00000000000000c200000000",
            INIT_32 => X"0000001900000000000000230000000000000035000000000000004100000000",
            INIT_33 => X"00000020000000000000002d000000000000002b000000000000001c00000000",
            INIT_34 => X"0000002f000000000000002f0000000000000033000000000000002e00000000",
            INIT_35 => X"00000029000000000000002b000000000000002d000000000000003000000000",
            INIT_36 => X"0000003a0000000000000024000000000000001e000000000000002200000000",
            INIT_37 => X"0000001e000000000000001d0000000000000021000000000000003900000000",
            INIT_38 => X"0000009800000000000000b600000000000000d700000000000000ec00000000",
            INIT_39 => X"00000074000000000000007a0000000000000081000000000000008800000000",
            INIT_3A => X"00000009000000000000000d0000000000000023000000000000005100000000",
            INIT_3B => X"0000002200000000000000490000000000000034000000000000001400000000",
            INIT_3C => X"00000020000000000000001a000000000000001c000000000000001100000000",
            INIT_3D => X"00000031000000000000003b000000000000003b000000000000002f00000000",
            INIT_3E => X"000000340000000000000022000000000000001a000000000000002300000000",
            INIT_3F => X"0000001d000000000000001c000000000000002c000000000000003f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000078000000000000007a0000000000000082000000000000009a00000000",
            INIT_41 => X"0000005c00000000000000680000000000000076000000000000007b00000000",
            INIT_42 => X"00000012000000000000001f0000000000000046000000000000005a00000000",
            INIT_43 => X"000000340000000000000045000000000000003d000000000000001d00000000",
            INIT_44 => X"0000002800000000000000240000000000000024000000000000002200000000",
            INIT_45 => X"0000003d00000000000000410000000000000047000000000000003a00000000",
            INIT_46 => X"00000028000000000000001f0000000000000017000000000000003000000000",
            INIT_47 => X"0000001c0000000000000027000000000000003c000000000000003800000000",
            INIT_48 => X"00000068000000000000006d000000000000006b000000000000006900000000",
            INIT_49 => X"0000005d000000000000005b0000000000000058000000000000005f00000000",
            INIT_4A => X"0000003e00000000000000560000000000000062000000000000006000000000",
            INIT_4B => X"00000031000000000000002f0000000000000038000000000000003800000000",
            INIT_4C => X"00000030000000000000002a0000000000000025000000000000002800000000",
            INIT_4D => X"000000390000000000000048000000000000005b000000000000004c00000000",
            INIT_4E => X"00000023000000000000001d000000000000002c000000000000003600000000",
            INIT_4F => X"0000001d0000000000000037000000000000003d000000000000002a00000000",
            INIT_50 => X"0000005100000000000000530000000000000059000000000000005f00000000",
            INIT_51 => X"00000058000000000000005b0000000000000058000000000000005600000000",
            INIT_52 => X"0000003e00000000000000440000000000000049000000000000005300000000",
            INIT_53 => X"00000034000000000000002c0000000000000023000000000000002800000000",
            INIT_54 => X"000000310000000000000027000000000000001e000000000000002800000000",
            INIT_55 => X"000000320000000000000047000000000000005f000000000000005100000000",
            INIT_56 => X"000000230000000000000025000000000000002a000000000000002900000000",
            INIT_57 => X"00000028000000000000003a0000000000000030000000000000002200000000",
            INIT_58 => X"00000055000000000000004f0000000000000049000000000000004b00000000",
            INIT_59 => X"00000040000000000000004c0000000000000053000000000000005700000000",
            INIT_5A => X"0000003b000000000000002a0000000000000027000000000000003300000000",
            INIT_5B => X"0000003100000000000000290000000000000022000000000000003200000000",
            INIT_5C => X"000000270000000000000024000000000000001e000000000000002600000000",
            INIT_5D => X"0000002d000000000000003c0000000000000045000000000000003700000000",
            INIT_5E => X"0000001d00000000000000220000000000000026000000000000002600000000",
            INIT_5F => X"0000003300000000000000300000000000000024000000000000002000000000",
            INIT_60 => X"0000004d000000000000004f000000000000004e000000000000004c00000000",
            INIT_61 => X"00000021000000000000002c0000000000000039000000000000004400000000",
            INIT_62 => X"0000003d000000000000002e000000000000001e000000000000001d00000000",
            INIT_63 => X"0000002600000000000000320000000000000029000000000000003700000000",
            INIT_64 => X"0000001e000000000000001d000000000000001a000000000000001d00000000",
            INIT_65 => X"00000030000000000000002e0000000000000025000000000000001d00000000",
            INIT_66 => X"0000001800000000000000190000000000000025000000000000002e00000000",
            INIT_67 => X"0000002f00000000000000240000000000000020000000000000001e00000000",
            INIT_68 => X"000000320000000000000040000000000000004a000000000000005000000000",
            INIT_69 => X"0000001b000000000000001e0000000000000020000000000000002600000000",
            INIT_6A => X"0000003c000000000000002d000000000000001b000000000000001b00000000",
            INIT_6B => X"0000001d000000000000002c000000000000002f000000000000003500000000",
            INIT_6C => X"0000001c00000000000000170000000000000017000000000000001c00000000",
            INIT_6D => X"0000002500000000000000200000000000000018000000000000001900000000",
            INIT_6E => X"000000150000000000000015000000000000001d000000000000002300000000",
            INIT_6F => X"00000022000000000000001c000000000000001e000000000000001a00000000",
            INIT_70 => X"0000001a0000000000000021000000000000002d000000000000003a00000000",
            INIT_71 => X"0000001c0000000000000021000000000000001d000000000000001a00000000",
            INIT_72 => X"0000003300000000000000270000000000000018000000000000001b00000000",
            INIT_73 => X"0000001c00000000000000210000000000000032000000000000003100000000",
            INIT_74 => X"0000001d00000000000000190000000000000015000000000000001b00000000",
            INIT_75 => X"0000001700000000000000190000000000000015000000000000001800000000",
            INIT_76 => X"000000120000000000000016000000000000001a000000000000001700000000",
            INIT_77 => X"000000170000000000000019000000000000001a000000000000001500000000",
            INIT_78 => X"0000001500000000000000180000000000000017000000000000001b00000000",
            INIT_79 => X"0000001900000000000000180000000000000019000000000000001a00000000",
            INIT_7A => X"0000003000000000000000210000000000000016000000000000001a00000000",
            INIT_7B => X"0000001800000000000000230000000000000033000000000000002a00000000",
            INIT_7C => X"0000001800000000000000150000000000000014000000000000001500000000",
            INIT_7D => X"00000019000000000000001d0000000000000017000000000000001700000000",
            INIT_7E => X"000000120000000000000016000000000000001b000000000000001800000000",
            INIT_7F => X"0000001600000000000000180000000000000016000000000000001100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE47;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE48 : if BRAM_NAME = "sampleifmap_layersamples_instance48" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004100000000000000150000000000000013000000000000001700000000",
            INIT_01 => X"000000b200000000000000b700000000000000bc00000000000000a400000000",
            INIT_02 => X"000000ba00000000000000ba00000000000000ac00000000000000aa00000000",
            INIT_03 => X"000000b700000000000000b600000000000000b700000000000000b800000000",
            INIT_04 => X"0000005c000000000000007f00000000000000a400000000000000b400000000",
            INIT_05 => X"000000c20000000000000099000000000000006e000000000000006b00000000",
            INIT_06 => X"000000c600000000000000c500000000000000c900000000000000c300000000",
            INIT_07 => X"000000c500000000000000c700000000000000c800000000000000c900000000",
            INIT_08 => X"0000002e00000000000000150000000000000013000000000000001700000000",
            INIT_09 => X"000000b200000000000000bf00000000000000ca000000000000009900000000",
            INIT_0A => X"000000b700000000000000a9000000000000009e00000000000000a400000000",
            INIT_0B => X"000000b200000000000000b400000000000000b800000000000000ba00000000",
            INIT_0C => X"00000056000000000000008a00000000000000ad00000000000000b400000000",
            INIT_0D => X"000000ce00000000000000b4000000000000006a000000000000004a00000000",
            INIT_0E => X"000000ce00000000000000d000000000000000d500000000000000cf00000000",
            INIT_0F => X"000000ca00000000000000cc00000000000000cd00000000000000cf00000000",
            INIT_10 => X"0000001f00000000000000170000000000000014000000000000001700000000",
            INIT_11 => X"000000a800000000000000b900000000000000c8000000000000007f00000000",
            INIT_12 => X"000000a2000000000000009a000000000000009e000000000000009f00000000",
            INIT_13 => X"000000b200000000000000b300000000000000b200000000000000b200000000",
            INIT_14 => X"0000007d00000000000000b600000000000000be00000000000000b500000000",
            INIT_15 => X"000000d100000000000000c50000000000000072000000000000004700000000",
            INIT_16 => X"000000d300000000000000d500000000000000d800000000000000d500000000",
            INIT_17 => X"000000ce00000000000000d000000000000000d300000000000000d400000000",
            INIT_18 => X"0000001700000000000000180000000000000015000000000000001700000000",
            INIT_19 => X"000000a000000000000000af00000000000000bd000000000000006300000000",
            INIT_1A => X"0000009500000000000000a600000000000000a800000000000000a800000000",
            INIT_1B => X"000000c300000000000000bf00000000000000ba00000000000000aa00000000",
            INIT_1C => X"0000008d00000000000000bc00000000000000c800000000000000c300000000",
            INIT_1D => X"000000d600000000000000d20000000000000092000000000000006300000000",
            INIT_1E => X"000000d500000000000000d400000000000000d400000000000000d500000000",
            INIT_1F => X"000000d600000000000000d700000000000000d900000000000000d900000000",
            INIT_20 => X"0000001500000000000000170000000000000017000000000000001900000000",
            INIT_21 => X"0000009700000000000000a500000000000000aa000000000000004800000000",
            INIT_22 => X"0000009b00000000000000b900000000000000b700000000000000af00000000",
            INIT_23 => X"000000bc00000000000000a9000000000000009d000000000000009200000000",
            INIT_24 => X"0000008d00000000000000b200000000000000c400000000000000c500000000",
            INIT_25 => X"000000db00000000000000d300000000000000ac000000000000007900000000",
            INIT_26 => X"000000d900000000000000d900000000000000d900000000000000dd00000000",
            INIT_27 => X"000000ce00000000000000d100000000000000d400000000000000d600000000",
            INIT_28 => X"00000017000000000000001a000000000000001b000000000000001a00000000",
            INIT_29 => X"0000009a00000000000000a4000000000000008f000000000000003100000000",
            INIT_2A => X"000000a600000000000000c800000000000000c200000000000000a900000000",
            INIT_2B => X"000000970000000000000080000000000000007d000000000000008200000000",
            INIT_2C => X"0000008f000000000000009400000000000000a500000000000000a500000000",
            INIT_2D => X"000000c900000000000000bc00000000000000b6000000000000009300000000",
            INIT_2E => X"000000db00000000000000d500000000000000d900000000000000d400000000",
            INIT_2F => X"000000d300000000000000d700000000000000d700000000000000dc00000000",
            INIT_30 => X"00000019000000000000001b000000000000001a000000000000001e00000000",
            INIT_31 => X"000000ab00000000000000b4000000000000007d000000000000002500000000",
            INIT_32 => X"000000b300000000000000ca00000000000000c500000000000000a900000000",
            INIT_33 => X"00000082000000000000007a0000000000000071000000000000008b00000000",
            INIT_34 => X"0000008c000000000000007a0000000000000085000000000000007700000000",
            INIT_35 => X"000000c900000000000000bf00000000000000cb00000000000000b900000000",
            INIT_36 => X"000000db00000000000000d700000000000000da00000000000000d700000000",
            INIT_37 => X"000000e000000000000000dc00000000000000da00000000000000dc00000000",
            INIT_38 => X"00000024000000000000001f0000000000000030000000000000005e00000000",
            INIT_39 => X"000000a800000000000000c100000000000000af000000000000006400000000",
            INIT_3A => X"000000c300000000000000c600000000000000c000000000000000a300000000",
            INIT_3B => X"00000084000000000000008e000000000000009100000000000000ae00000000",
            INIT_3C => X"0000008b000000000000007a0000000000000079000000000000006a00000000",
            INIT_3D => X"000000d500000000000000bd00000000000000d100000000000000c000000000",
            INIT_3E => X"000000e800000000000000ef00000000000000ed00000000000000f200000000",
            INIT_3F => X"000000e500000000000000de00000000000000d500000000000000d000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007a0000000000000072000000000000009e00000000000000b400000000",
            INIT_41 => X"000000a000000000000000be00000000000000be00000000000000b100000000",
            INIT_42 => X"000000c800000000000000c500000000000000ad000000000000008500000000",
            INIT_43 => X"0000009200000000000000a700000000000000b900000000000000c200000000",
            INIT_44 => X"0000008d00000000000000850000000000000081000000000000008100000000",
            INIT_45 => X"000000dc00000000000000bd00000000000000c900000000000000b100000000",
            INIT_46 => X"000000d500000000000000e800000000000000eb00000000000000f100000000",
            INIT_47 => X"000000ea00000000000000e100000000000000c700000000000000bd00000000",
            INIT_48 => X"000000ba00000000000000b200000000000000c000000000000000c500000000",
            INIT_49 => X"0000009d00000000000000c500000000000000c300000000000000c100000000",
            INIT_4A => X"000000bf00000000000000b900000000000000a3000000000000008000000000",
            INIT_4B => X"0000009700000000000000b200000000000000c300000000000000c100000000",
            INIT_4C => X"0000008600000000000000830000000000000081000000000000007200000000",
            INIT_4D => X"000000ea00000000000000d000000000000000c200000000000000aa00000000",
            INIT_4E => X"000000c900000000000000eb00000000000000f000000000000000ec00000000",
            INIT_4F => X"000000eb00000000000000d000000000000000bb00000000000000b900000000",
            INIT_50 => X"000000c000000000000000bb00000000000000c400000000000000ca00000000",
            INIT_51 => X"0000009700000000000000c500000000000000cd00000000000000c800000000",
            INIT_52 => X"000000bd00000000000000b800000000000000af000000000000009500000000",
            INIT_53 => X"0000008800000000000000a800000000000000bb00000000000000c100000000",
            INIT_54 => X"0000008100000000000000800000000000000080000000000000007500000000",
            INIT_55 => X"000000f000000000000000cd00000000000000b500000000000000a700000000",
            INIT_56 => X"000000ce00000000000000ee00000000000000f300000000000000f300000000",
            INIT_57 => X"000000dd00000000000000c100000000000000bb00000000000000ba00000000",
            INIT_58 => X"000000c000000000000000c500000000000000cd00000000000000cd00000000",
            INIT_59 => X"000000a000000000000000c200000000000000d000000000000000cb00000000",
            INIT_5A => X"000000bf00000000000000c100000000000000bf00000000000000a800000000",
            INIT_5B => X"00000077000000000000009200000000000000ac00000000000000c100000000",
            INIT_5C => X"000000870000000000000085000000000000008e000000000000007c00000000",
            INIT_5D => X"000000ea00000000000000bf00000000000000b000000000000000a700000000",
            INIT_5E => X"000000d700000000000000ec00000000000000f100000000000000f300000000",
            INIT_5F => X"000000c400000000000000b900000000000000b800000000000000ba00000000",
            INIT_60 => X"000000c100000000000000c800000000000000cc00000000000000ce00000000",
            INIT_61 => X"000000b400000000000000bf00000000000000c700000000000000c500000000",
            INIT_62 => X"000000ad00000000000000b700000000000000b300000000000000ac00000000",
            INIT_63 => X"00000083000000000000009800000000000000ae00000000000000ae00000000",
            INIT_64 => X"0000009a000000000000008e00000000000000a6000000000000008d00000000",
            INIT_65 => X"000000e600000000000000bf00000000000000ac00000000000000a900000000",
            INIT_66 => X"000000e400000000000000ef00000000000000f100000000000000f000000000",
            INIT_67 => X"000000c000000000000000b800000000000000ba00000000000000c800000000",
            INIT_68 => X"000000bf00000000000000c600000000000000ca00000000000000d200000000",
            INIT_69 => X"000000ca00000000000000b100000000000000b400000000000000c900000000",
            INIT_6A => X"0000008e000000000000008e000000000000009a00000000000000ab00000000",
            INIT_6B => X"0000009c000000000000009300000000000000a800000000000000a800000000",
            INIT_6C => X"000000a4000000000000009600000000000000a900000000000000af00000000",
            INIT_6D => X"000000e600000000000000c500000000000000a0000000000000009e00000000",
            INIT_6E => X"000000f200000000000000f400000000000000f100000000000000f100000000",
            INIT_6F => X"000000d700000000000000c300000000000000bf00000000000000e200000000",
            INIT_70 => X"000000c000000000000000c700000000000000c900000000000000d300000000",
            INIT_71 => X"000000d700000000000000a100000000000000aa00000000000000cf00000000",
            INIT_72 => X"000000ac00000000000000ad00000000000000ba00000000000000bd00000000",
            INIT_73 => X"0000007f000000000000008900000000000000b100000000000000be00000000",
            INIT_74 => X"000000a0000000000000009600000000000000ae00000000000000b400000000",
            INIT_75 => X"000000ec00000000000000c100000000000000b000000000000000af00000000",
            INIT_76 => X"000000fb00000000000000f300000000000000f200000000000000f500000000",
            INIT_77 => X"000000e100000000000000d400000000000000c900000000000000ef00000000",
            INIT_78 => X"000000c100000000000000c500000000000000c400000000000000d300000000",
            INIT_79 => X"000000d9000000000000009a00000000000000b500000000000000d100000000",
            INIT_7A => X"000000b900000000000000c300000000000000c500000000000000ce00000000",
            INIT_7B => X"0000009800000000000000a600000000000000ad00000000000000aa00000000",
            INIT_7C => X"0000009800000000000000a600000000000000b800000000000000a300000000",
            INIT_7D => X"000000cc00000000000000af00000000000000b500000000000000c000000000",
            INIT_7E => X"000000f700000000000000f400000000000000f300000000000000ee00000000",
            INIT_7F => X"000000e200000000000000e200000000000000d500000000000000df00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE48;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE49 : if BRAM_NAME = "sampleifmap_layersamples_instance49" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b500000000000000b400000000000000c200000000000000d600000000",
            INIT_01 => X"000000c6000000000000009b00000000000000c400000000000000c500000000",
            INIT_02 => X"000000b700000000000000ae00000000000000c000000000000000d600000000",
            INIT_03 => X"000000b200000000000000ae00000000000000a100000000000000ad00000000",
            INIT_04 => X"0000009300000000000000bd00000000000000a4000000000000008000000000",
            INIT_05 => X"00000076000000000000009c00000000000000b400000000000000a700000000",
            INIT_06 => X"000000eb00000000000000ef00000000000000d7000000000000009d00000000",
            INIT_07 => X"000000e400000000000000ea00000000000000d600000000000000ce00000000",
            INIT_08 => X"000000a300000000000000a600000000000000c600000000000000d700000000",
            INIT_09 => X"000000b900000000000000be00000000000000ca00000000000000b400000000",
            INIT_0A => X"000000d600000000000000cd00000000000000d200000000000000cf00000000",
            INIT_0B => X"000000ad00000000000000b000000000000000ae00000000000000c100000000",
            INIT_0C => X"0000009900000000000000bf0000000000000089000000000000008100000000",
            INIT_0D => X"0000008700000000000000ab00000000000000c800000000000000a300000000",
            INIT_0E => X"000000c100000000000000b80000000000000090000000000000007400000000",
            INIT_0F => X"000000eb00000000000000ef00000000000000d200000000000000bb00000000",
            INIT_10 => X"000000a400000000000000ae00000000000000cd00000000000000d800000000",
            INIT_11 => X"000000c200000000000000d200000000000000cb00000000000000b900000000",
            INIT_12 => X"000000e200000000000000da00000000000000d300000000000000bf00000000",
            INIT_13 => X"000000b300000000000000be00000000000000cb00000000000000e100000000",
            INIT_14 => X"0000009e00000000000000a80000000000000079000000000000009700000000",
            INIT_15 => X"000000ac00000000000000aa00000000000000c200000000000000a700000000",
            INIT_16 => X"000000a900000000000000990000000000000083000000000000009a00000000",
            INIT_17 => X"000000ec00000000000000de00000000000000b800000000000000a200000000",
            INIT_18 => X"000000b400000000000000c000000000000000d000000000000000d800000000",
            INIT_19 => X"000000d200000000000000d100000000000000ca00000000000000c500000000",
            INIT_1A => X"000000cc00000000000000c500000000000000bd00000000000000ba00000000",
            INIT_1B => X"000000b500000000000000cf00000000000000d500000000000000d100000000",
            INIT_1C => X"000000af0000000000000092000000000000009500000000000000b200000000",
            INIT_1D => X"000000ab000000000000009c00000000000000ae00000000000000b700000000",
            INIT_1E => X"000000b400000000000000a9000000000000009400000000000000a300000000",
            INIT_1F => X"000000cc00000000000000ac00000000000000a000000000000000a600000000",
            INIT_20 => X"000000b600000000000000ca00000000000000d500000000000000da00000000",
            INIT_21 => X"000000ca00000000000000c900000000000000cb00000000000000bf00000000",
            INIT_22 => X"000000c000000000000000c100000000000000c300000000000000ca00000000",
            INIT_23 => X"000000c700000000000000cf00000000000000c600000000000000b200000000",
            INIT_24 => X"000000bb00000000000000a600000000000000cb00000000000000d300000000",
            INIT_25 => X"000000a60000000000000093000000000000009b00000000000000b100000000",
            INIT_26 => X"000000af00000000000000b600000000000000ab00000000000000a700000000",
            INIT_27 => X"000000a7000000000000009f000000000000009c000000000000009c00000000",
            INIT_28 => X"000000ba00000000000000d100000000000000d700000000000000d900000000",
            INIT_29 => X"000000c800000000000000d000000000000000c800000000000000b300000000",
            INIT_2A => X"000000ba00000000000000d200000000000000d700000000000000d100000000",
            INIT_2B => X"000000c200000000000000c400000000000000b600000000000000a100000000",
            INIT_2C => X"000000b900000000000000be00000000000000cf00000000000000cb00000000",
            INIT_2D => X"000000a6000000000000009b000000000000008e000000000000009b00000000",
            INIT_2E => X"0000009f00000000000000ad00000000000000b300000000000000ac00000000",
            INIT_2F => X"0000008f000000000000009e000000000000009e000000000000009600000000",
            INIT_30 => X"000000c000000000000000d600000000000000d500000000000000d600000000",
            INIT_31 => X"000000d900000000000000da00000000000000c500000000000000a900000000",
            INIT_32 => X"000000c300000000000000d400000000000000d900000000000000d700000000",
            INIT_33 => X"000000bf00000000000000c300000000000000b300000000000000aa00000000",
            INIT_34 => X"000000aa00000000000000c000000000000000c000000000000000be00000000",
            INIT_35 => X"000000aa00000000000000a7000000000000008e000000000000008400000000",
            INIT_36 => X"0000009d00000000000000ad00000000000000b300000000000000aa00000000",
            INIT_37 => X"0000007d00000000000000860000000000000093000000000000009d00000000",
            INIT_38 => X"000000ca00000000000000d300000000000000d100000000000000d500000000",
            INIT_39 => X"000000de00000000000000d800000000000000c100000000000000a800000000",
            INIT_3A => X"000000cd00000000000000d300000000000000de00000000000000df00000000",
            INIT_3B => X"000000c600000000000000c900000000000000c200000000000000c200000000",
            INIT_3C => X"0000009900000000000000bc00000000000000c400000000000000c600000000",
            INIT_3D => X"000000a700000000000000ab000000000000009b000000000000008600000000",
            INIT_3E => X"000000a500000000000000b200000000000000bd00000000000000a600000000",
            INIT_3F => X"000000890000000000000085000000000000008e00000000000000a300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ca00000000000000ce00000000000000ce00000000000000d300000000",
            INIT_41 => X"000000d500000000000000d300000000000000bf00000000000000af00000000",
            INIT_42 => X"000000ab00000000000000c600000000000000d800000000000000d600000000",
            INIT_43 => X"000000c900000000000000c900000000000000ce00000000000000c200000000",
            INIT_44 => X"0000009600000000000000b100000000000000c500000000000000c800000000",
            INIT_45 => X"0000009d00000000000000a7000000000000009e000000000000009000000000",
            INIT_46 => X"000000a800000000000000b000000000000000b5000000000000009f00000000",
            INIT_47 => X"0000009000000000000000950000000000000096000000000000009800000000",
            INIT_48 => X"000000c100000000000000c900000000000000cc00000000000000d200000000",
            INIT_49 => X"000000d200000000000000d000000000000000bc00000000000000b500000000",
            INIT_4A => X"0000007a00000000000000a000000000000000ce00000000000000cd00000000",
            INIT_4B => X"000000c200000000000000c600000000000000d000000000000000b100000000",
            INIT_4C => X"0000009600000000000000a600000000000000b800000000000000c100000000",
            INIT_4D => X"0000009900000000000000a0000000000000009c000000000000008b00000000",
            INIT_4E => X"0000009b000000000000009f00000000000000a0000000000000009b00000000",
            INIT_4F => X"00000083000000000000008c0000000000000098000000000000009800000000",
            INIT_50 => X"000000bb00000000000000c600000000000000ca00000000000000d200000000",
            INIT_51 => X"000000d600000000000000cd00000000000000b200000000000000ae00000000",
            INIT_52 => X"0000008300000000000000a400000000000000cb00000000000000d100000000",
            INIT_53 => X"000000b600000000000000bb00000000000000ca00000000000000b400000000",
            INIT_54 => X"0000008b000000000000009d00000000000000a900000000000000b600000000",
            INIT_55 => X"00000090000000000000009a0000000000000099000000000000008600000000",
            INIT_56 => X"0000008d0000000000000083000000000000008d000000000000009700000000",
            INIT_57 => X"000000930000000000000096000000000000009b000000000000009d00000000",
            INIT_58 => X"000000b500000000000000c200000000000000c800000000000000d200000000",
            INIT_59 => X"000000d700000000000000c400000000000000a800000000000000a800000000",
            INIT_5A => X"000000b800000000000000bd00000000000000c700000000000000d400000000",
            INIT_5B => X"000000ac00000000000000ad00000000000000b900000000000000cb00000000",
            INIT_5C => X"000000760000000000000093000000000000009b00000000000000a300000000",
            INIT_5D => X"0000008d00000000000000910000000000000094000000000000008300000000",
            INIT_5E => X"00000085000000000000007f0000000000000084000000000000009000000000",
            INIT_5F => X"0000009c00000000000000a200000000000000a3000000000000009500000000",
            INIT_60 => X"000000b400000000000000bd00000000000000c200000000000000d000000000",
            INIT_61 => X"000000d300000000000000bd000000000000009e00000000000000a200000000",
            INIT_62 => X"000000c700000000000000c200000000000000c500000000000000d300000000",
            INIT_63 => X"000000a400000000000000a300000000000000ac00000000000000bf00000000",
            INIT_64 => X"0000006d00000000000000820000000000000093000000000000009e00000000",
            INIT_65 => X"0000009100000000000000900000000000000090000000000000008900000000",
            INIT_66 => X"00000086000000000000007c0000000000000084000000000000009000000000",
            INIT_67 => X"00000093000000000000009f00000000000000a2000000000000009700000000",
            INIT_68 => X"000000b500000000000000b000000000000000b100000000000000c200000000",
            INIT_69 => X"000000cd00000000000000b3000000000000008f000000000000009f00000000",
            INIT_6A => X"000000be00000000000000c200000000000000c700000000000000d000000000",
            INIT_6B => X"000000a1000000000000009c00000000000000a500000000000000b500000000",
            INIT_6C => X"0000007200000000000000700000000000000088000000000000009500000000",
            INIT_6D => X"00000092000000000000008a0000000000000085000000000000008900000000",
            INIT_6E => X"0000009000000000000000830000000000000083000000000000009200000000",
            INIT_6F => X"0000008d00000000000000940000000000000095000000000000009600000000",
            INIT_70 => X"000000b200000000000000a5000000000000009d00000000000000ac00000000",
            INIT_71 => X"000000c7000000000000009c000000000000008500000000000000a700000000",
            INIT_72 => X"000000c200000000000000c700000000000000c700000000000000ce00000000",
            INIT_73 => X"0000008b0000000000000084000000000000008500000000000000a000000000",
            INIT_74 => X"0000007e000000000000006b000000000000007e000000000000008c00000000",
            INIT_75 => X"00000095000000000000008a0000000000000081000000000000008200000000",
            INIT_76 => X"0000008e0000000000000091000000000000008c000000000000008d00000000",
            INIT_77 => X"000000980000000000000095000000000000008c000000000000008800000000",
            INIT_78 => X"0000009b00000000000000900000000000000086000000000000009700000000",
            INIT_79 => X"000000b70000000000000082000000000000007d000000000000009e00000000",
            INIT_7A => X"000000a500000000000000b700000000000000bf00000000000000c500000000",
            INIT_7B => X"00000069000000000000005e0000000000000067000000000000008000000000",
            INIT_7C => X"0000007c00000000000000750000000000000070000000000000007700000000",
            INIT_7D => X"0000008f000000000000008b000000000000007d000000000000007900000000",
            INIT_7E => X"0000007d0000000000000081000000000000008c000000000000008b00000000",
            INIT_7F => X"00000096000000000000009b0000000000000095000000000000008400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE49;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE50 : if BRAM_NAME = "sampleifmap_layersamples_instance50" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002f00000000000000100000000000000015000000000000001300000000",
            INIT_01 => X"0000008e00000000000000930000000000000093000000000000008300000000",
            INIT_02 => X"0000008e00000000000000900000000000000089000000000000008700000000",
            INIT_03 => X"0000008f000000000000008c000000000000008c000000000000008d00000000",
            INIT_04 => X"000000490000000000000060000000000000007e000000000000008c00000000",
            INIT_05 => X"000000a40000000000000082000000000000005d000000000000005f00000000",
            INIT_06 => X"0000009d000000000000009b000000000000009c000000000000009b00000000",
            INIT_07 => X"000000970000000000000098000000000000009b000000000000009e00000000",
            INIT_08 => X"0000001f00000000000000110000000000000014000000000000001400000000",
            INIT_09 => X"00000092000000000000009b00000000000000a1000000000000007a00000000",
            INIT_0A => X"00000095000000000000008b0000000000000088000000000000008a00000000",
            INIT_0B => X"0000009700000000000000920000000000000096000000000000009800000000",
            INIT_0C => X"0000004900000000000000750000000000000096000000000000009f00000000",
            INIT_0D => X"000000af000000000000009c0000000000000058000000000000004100000000",
            INIT_0E => X"000000ad00000000000000ab00000000000000a900000000000000a800000000",
            INIT_0F => X"000000a300000000000000a400000000000000a800000000000000ac00000000",
            INIT_10 => X"0000001500000000000000140000000000000014000000000000001400000000",
            INIT_11 => X"0000008c000000000000009700000000000000a2000000000000006600000000",
            INIT_12 => X"0000008b00000000000000880000000000000095000000000000008d00000000",
            INIT_13 => X"0000009f00000000000000980000000000000099000000000000009a00000000",
            INIT_14 => X"0000006d00000000000000a100000000000000ab00000000000000a600000000",
            INIT_15 => X"000000b700000000000000b10000000000000061000000000000003a00000000",
            INIT_16 => X"000000b200000000000000b100000000000000b200000000000000b300000000",
            INIT_17 => X"000000a600000000000000a900000000000000ad00000000000000b100000000",
            INIT_18 => X"0000001100000000000000150000000000000014000000000000001400000000",
            INIT_19 => X"00000082000000000000008c0000000000000099000000000000004f00000000",
            INIT_1A => X"00000087000000000000009d00000000000000a4000000000000009700000000",
            INIT_1B => X"000000b000000000000000a900000000000000a6000000000000009900000000",
            INIT_1C => X"0000007600000000000000a100000000000000af00000000000000b000000000",
            INIT_1D => X"000000c300000000000000c40000000000000085000000000000005200000000",
            INIT_1E => X"000000b300000000000000b400000000000000b700000000000000bd00000000",
            INIT_1F => X"000000ab00000000000000ad00000000000000b100000000000000b300000000",
            INIT_20 => X"0000001300000000000000150000000000000014000000000000001500000000",
            INIT_21 => X"0000007700000000000000820000000000000089000000000000003800000000",
            INIT_22 => X"0000009200000000000000b300000000000000b2000000000000009c00000000",
            INIT_23 => X"000000a70000000000000094000000000000008b000000000000008400000000",
            INIT_24 => X"00000078000000000000009800000000000000a900000000000000af00000000",
            INIT_25 => X"000000d200000000000000ce00000000000000a7000000000000006d00000000",
            INIT_26 => X"000000bf00000000000000c300000000000000c900000000000000d100000000",
            INIT_27 => X"000000ac00000000000000b100000000000000b600000000000000ba00000000",
            INIT_28 => X"0000001600000000000000170000000000000016000000000000001600000000",
            INIT_29 => X"0000007800000000000000820000000000000073000000000000002600000000",
            INIT_2A => X"0000009e00000000000000c300000000000000b9000000000000009200000000",
            INIT_2B => X"00000084000000000000006b000000000000006c000000000000007600000000",
            INIT_2C => X"000000840000000000000081000000000000008f000000000000009200000000",
            INIT_2D => X"000000c700000000000000be00000000000000b7000000000000008f00000000",
            INIT_2E => X"000000d100000000000000cc00000000000000d100000000000000cf00000000",
            INIT_2F => X"000000c200000000000000c700000000000000ca00000000000000d100000000",
            INIT_30 => X"0000001400000000000000150000000000000013000000000000001800000000",
            INIT_31 => X"0000009400000000000000a10000000000000071000000000000001e00000000",
            INIT_32 => X"000000aa00000000000000c200000000000000ba000000000000009700000000",
            INIT_33 => X"0000007100000000000000690000000000000062000000000000008000000000",
            INIT_34 => X"00000080000000000000006b0000000000000074000000000000006800000000",
            INIT_35 => X"000000c500000000000000c000000000000000ca00000000000000b200000000",
            INIT_36 => X"000000d700000000000000d100000000000000cf00000000000000ce00000000",
            INIT_37 => X"000000da00000000000000d700000000000000d600000000000000d800000000",
            INIT_38 => X"0000001d00000000000000180000000000000029000000000000005800000000",
            INIT_39 => X"0000009c00000000000000ba00000000000000ae000000000000006000000000",
            INIT_3A => X"000000ba00000000000000bd00000000000000b5000000000000009500000000",
            INIT_3B => X"000000760000000000000081000000000000008400000000000000a400000000",
            INIT_3C => X"0000007c000000000000006c000000000000006b000000000000005c00000000",
            INIT_3D => X"000000ce00000000000000bb00000000000000cc00000000000000b400000000",
            INIT_3E => X"000000e400000000000000e700000000000000e000000000000000e600000000",
            INIT_3F => X"000000e200000000000000dc00000000000000d300000000000000cd00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000075000000000000006d000000000000009900000000000000b100000000",
            INIT_41 => X"0000009300000000000000b700000000000000bd00000000000000af00000000",
            INIT_42 => X"000000c000000000000000bc00000000000000a1000000000000007800000000",
            INIT_43 => X"00000083000000000000009a00000000000000ad00000000000000b800000000",
            INIT_44 => X"0000007f00000000000000770000000000000073000000000000007300000000",
            INIT_45 => X"000000d800000000000000bc00000000000000c500000000000000a600000000",
            INIT_46 => X"000000d300000000000000e300000000000000e200000000000000e900000000",
            INIT_47 => X"000000e800000000000000e000000000000000c600000000000000bc00000000",
            INIT_48 => X"000000b600000000000000af00000000000000bc00000000000000c200000000",
            INIT_49 => X"0000009000000000000000be00000000000000c200000000000000bf00000000",
            INIT_4A => X"000000b600000000000000b10000000000000098000000000000007300000000",
            INIT_4B => X"0000008a00000000000000a400000000000000b600000000000000b700000000",
            INIT_4C => X"0000007b00000000000000770000000000000076000000000000006600000000",
            INIT_4D => X"000000e900000000000000d000000000000000bd00000000000000a000000000",
            INIT_4E => X"000000cb00000000000000ea00000000000000eb00000000000000e800000000",
            INIT_4F => X"000000eb00000000000000d100000000000000bd00000000000000bb00000000",
            INIT_50 => X"000000bb00000000000000b700000000000000c000000000000000c700000000",
            INIT_51 => X"0000008a00000000000000bf00000000000000cd00000000000000c600000000",
            INIT_52 => X"000000b500000000000000b000000000000000a5000000000000008800000000",
            INIT_53 => X"0000007c000000000000009a00000000000000af00000000000000b800000000",
            INIT_54 => X"0000007800000000000000770000000000000076000000000000006b00000000",
            INIT_55 => X"000000f000000000000000cd00000000000000b0000000000000009e00000000",
            INIT_56 => X"000000d400000000000000f200000000000000f400000000000000f300000000",
            INIT_57 => X"000000e000000000000000c600000000000000c000000000000000c000000000",
            INIT_58 => X"000000bb00000000000000c100000000000000c900000000000000c900000000",
            INIT_59 => X"0000009200000000000000bc00000000000000d100000000000000c900000000",
            INIT_5A => X"000000b700000000000000b900000000000000b6000000000000009b00000000",
            INIT_5B => X"0000006b0000000000000084000000000000009f00000000000000b700000000",
            INIT_5C => X"0000007e000000000000007c0000000000000085000000000000007300000000",
            INIT_5D => X"000000eb00000000000000bd00000000000000aa000000000000009e00000000",
            INIT_5E => X"000000de00000000000000f200000000000000f600000000000000f600000000",
            INIT_5F => X"000000ca00000000000000c000000000000000c000000000000000c200000000",
            INIT_60 => X"000000bd00000000000000c500000000000000c900000000000000cb00000000",
            INIT_61 => X"000000a500000000000000b700000000000000c600000000000000c400000000",
            INIT_62 => X"000000a500000000000000b000000000000000aa000000000000009f00000000",
            INIT_63 => X"00000078000000000000008a00000000000000a200000000000000a400000000",
            INIT_64 => X"000000920000000000000087000000000000009f000000000000008500000000",
            INIT_65 => X"000000e700000000000000bd00000000000000a500000000000000a100000000",
            INIT_66 => X"000000ea00000000000000f700000000000000f800000000000000f400000000",
            INIT_67 => X"000000c700000000000000c100000000000000c300000000000000d000000000",
            INIT_68 => X"000000b900000000000000c400000000000000ca00000000000000d000000000",
            INIT_69 => X"000000b9000000000000009c00000000000000a700000000000000c100000000",
            INIT_6A => X"000000870000000000000087000000000000009100000000000000a100000000",
            INIT_6B => X"0000008f0000000000000089000000000000009e00000000000000a100000000",
            INIT_6C => X"000000a2000000000000009500000000000000a400000000000000a400000000",
            INIT_6D => X"000000e400000000000000c3000000000000009d000000000000009900000000",
            INIT_6E => X"000000f500000000000000f900000000000000f700000000000000f200000000",
            INIT_6F => X"000000de00000000000000cc00000000000000c700000000000000e800000000",
            INIT_70 => X"000000b600000000000000c500000000000000cc00000000000000d200000000",
            INIT_71 => X"000000c1000000000000007d000000000000008e00000000000000bf00000000",
            INIT_72 => X"000000a700000000000000a600000000000000b100000000000000b500000000",
            INIT_73 => X"00000072000000000000008200000000000000aa00000000000000b800000000",
            INIT_74 => X"0000009e000000000000009800000000000000aa00000000000000a500000000",
            INIT_75 => X"000000e700000000000000bd00000000000000ae00000000000000ab00000000",
            INIT_76 => X"000000fb00000000000000f500000000000000f400000000000000f200000000",
            INIT_77 => X"000000e900000000000000dd00000000000000cf00000000000000f200000000",
            INIT_78 => X"000000b900000000000000c500000000000000c800000000000000d400000000",
            INIT_79 => X"000000c00000000000000070000000000000009100000000000000bd00000000",
            INIT_7A => X"000000b400000000000000bd00000000000000be00000000000000c700000000",
            INIT_7B => X"0000008900000000000000a000000000000000a700000000000000a400000000",
            INIT_7C => X"0000009100000000000000a200000000000000b0000000000000009200000000",
            INIT_7D => X"000000c300000000000000a800000000000000b100000000000000b800000000",
            INIT_7E => X"000000f900000000000000f500000000000000f100000000000000e800000000",
            INIT_7F => X"000000eb00000000000000ec00000000000000dd00000000000000e400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE50;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE51 : if BRAM_NAME = "sampleifmap_layersamples_instance51" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ae00000000000000b600000000000000c700000000000000d800000000",
            INIT_01 => X"000000ad000000000000006e000000000000009b00000000000000b000000000",
            INIT_02 => X"000000b200000000000000a800000000000000ba00000000000000d000000000",
            INIT_03 => X"000000a400000000000000a7000000000000009b00000000000000a800000000",
            INIT_04 => X"0000008600000000000000b10000000000000096000000000000006e00000000",
            INIT_05 => X"00000068000000000000009000000000000000ab000000000000009a00000000",
            INIT_06 => X"000000ed00000000000000ee00000000000000d1000000000000009100000000",
            INIT_07 => X"000000ed00000000000000f300000000000000dd00000000000000d200000000",
            INIT_08 => X"0000009e00000000000000a900000000000000ce00000000000000db00000000",
            INIT_09 => X"000000a2000000000000009500000000000000a700000000000000a300000000",
            INIT_0A => X"000000d100000000000000c800000000000000cd00000000000000ca00000000",
            INIT_0B => X"000000a100000000000000aa00000000000000a800000000000000bc00000000",
            INIT_0C => X"0000008700000000000000ad0000000000000078000000000000007000000000",
            INIT_0D => X"00000073000000000000009b00000000000000ba000000000000009300000000",
            INIT_0E => X"000000bc00000000000000b20000000000000084000000000000006200000000",
            INIT_0F => X"000000ef00000000000000f300000000000000d400000000000000b900000000",
            INIT_10 => X"000000a100000000000000b300000000000000d600000000000000dd00000000",
            INIT_11 => X"000000b100000000000000b300000000000000b500000000000000af00000000",
            INIT_12 => X"000000dd00000000000000d400000000000000cf00000000000000bd00000000",
            INIT_13 => X"000000ab00000000000000b800000000000000c500000000000000dc00000000",
            INIT_14 => X"0000008c00000000000000950000000000000067000000000000008b00000000",
            INIT_15 => X"00000093000000000000009400000000000000b1000000000000009700000000",
            INIT_16 => X"0000009c000000000000008a0000000000000070000000000000008300000000",
            INIT_17 => X"000000ea00000000000000d900000000000000b1000000000000009700000000",
            INIT_18 => X"000000b200000000000000c600000000000000da00000000000000df00000000",
            INIT_19 => X"000000c800000000000000be00000000000000c200000000000000c200000000",
            INIT_1A => X"000000c700000000000000bf00000000000000b800000000000000ba00000000",
            INIT_1B => X"000000b100000000000000c800000000000000d000000000000000cb00000000",
            INIT_1C => X"0000009e000000000000007f000000000000008700000000000000ab00000000",
            INIT_1D => X"0000008f0000000000000083000000000000009b00000000000000a800000000",
            INIT_1E => X"0000009f0000000000000094000000000000007e000000000000008900000000",
            INIT_1F => X"000000c5000000000000009e0000000000000090000000000000009300000000",
            INIT_20 => X"000000b700000000000000d000000000000000dd00000000000000e100000000",
            INIT_21 => X"000000c200000000000000be00000000000000c700000000000000bf00000000",
            INIT_22 => X"000000ba00000000000000be00000000000000bc00000000000000c600000000",
            INIT_23 => X"000000bf00000000000000c600000000000000c100000000000000ab00000000",
            INIT_24 => X"000000a9000000000000009400000000000000bf00000000000000cf00000000",
            INIT_25 => X"0000008d000000000000007b000000000000008700000000000000a000000000",
            INIT_26 => X"00000098000000000000009f0000000000000095000000000000008e00000000",
            INIT_27 => X"0000009a000000000000008c0000000000000088000000000000008700000000",
            INIT_28 => X"000000be00000000000000d600000000000000dd00000000000000de00000000",
            INIT_29 => X"000000be00000000000000c800000000000000c300000000000000b300000000",
            INIT_2A => X"000000b200000000000000d100000000000000cd00000000000000c600000000",
            INIT_2B => X"000000b500000000000000b600000000000000b3000000000000009700000000",
            INIT_2C => X"000000a500000000000000ae00000000000000c400000000000000c500000000",
            INIT_2D => X"000000930000000000000089000000000000007c000000000000008600000000",
            INIT_2E => X"0000008b000000000000009900000000000000a1000000000000009900000000",
            INIT_2F => X"0000007d000000000000008b000000000000008b000000000000008300000000",
            INIT_30 => X"000000c600000000000000db00000000000000da00000000000000db00000000",
            INIT_31 => X"000000cf00000000000000d200000000000000bf00000000000000aa00000000",
            INIT_32 => X"000000b400000000000000cf00000000000000ce00000000000000cb00000000",
            INIT_33 => X"000000b000000000000000b400000000000000ae000000000000009c00000000",
            INIT_34 => X"0000009600000000000000b000000000000000b500000000000000b600000000",
            INIT_35 => X"000000980000000000000096000000000000007d000000000000006f00000000",
            INIT_36 => X"0000008a000000000000009a00000000000000a1000000000000009800000000",
            INIT_37 => X"0000006a00000000000000730000000000000080000000000000008a00000000",
            INIT_38 => X"000000cf00000000000000d900000000000000d600000000000000da00000000",
            INIT_39 => X"000000d500000000000000d200000000000000bc00000000000000aa00000000",
            INIT_3A => X"000000b600000000000000c700000000000000d300000000000000d400000000",
            INIT_3B => X"000000b500000000000000ba00000000000000ba00000000000000ae00000000",
            INIT_3C => X"0000008500000000000000ab00000000000000b600000000000000ba00000000",
            INIT_3D => X"00000095000000000000009a0000000000000089000000000000007200000000",
            INIT_3E => X"00000092000000000000009f00000000000000ab000000000000009400000000",
            INIT_3F => X"000000760000000000000073000000000000007b000000000000009000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d100000000000000d400000000000000d400000000000000d800000000",
            INIT_41 => X"000000cd00000000000000cf00000000000000bd00000000000000b300000000",
            INIT_42 => X"0000008a00000000000000b100000000000000cd00000000000000cd00000000",
            INIT_43 => X"000000b600000000000000bb00000000000000c300000000000000a700000000",
            INIT_44 => X"00000082000000000000009e00000000000000b500000000000000b900000000",
            INIT_45 => X"0000008c0000000000000096000000000000008d000000000000007d00000000",
            INIT_46 => X"00000095000000000000009d00000000000000a3000000000000008d00000000",
            INIT_47 => X"0000007c00000000000000820000000000000083000000000000008500000000",
            INIT_48 => X"000000c800000000000000d000000000000000d200000000000000d700000000",
            INIT_49 => X"000000cc00000000000000ce00000000000000be00000000000000bb00000000",
            INIT_4A => X"00000050000000000000008300000000000000c400000000000000c600000000",
            INIT_4B => X"000000ae00000000000000b800000000000000c2000000000000009100000000",
            INIT_4C => X"00000083000000000000009300000000000000a500000000000000ae00000000",
            INIT_4D => X"00000088000000000000008f000000000000008b000000000000007800000000",
            INIT_4E => X"00000088000000000000008c000000000000008e000000000000008900000000",
            INIT_4F => X"0000007000000000000000790000000000000085000000000000008500000000",
            INIT_50 => X"000000c200000000000000cd00000000000000d000000000000000d700000000",
            INIT_51 => X"000000d100000000000000cd00000000000000b700000000000000b500000000",
            INIT_52 => X"00000051000000000000008100000000000000c200000000000000cc00000000",
            INIT_53 => X"000000a100000000000000ab00000000000000ba000000000000008e00000000",
            INIT_54 => X"000000780000000000000089000000000000009500000000000000a100000000",
            INIT_55 => X"0000007e00000000000000890000000000000087000000000000007300000000",
            INIT_56 => X"0000007a0000000000000070000000000000007b000000000000008500000000",
            INIT_57 => X"0000008000000000000000830000000000000088000000000000008a00000000",
            INIT_58 => X"000000bc00000000000000c800000000000000cd00000000000000d600000000",
            INIT_59 => X"000000d400000000000000c600000000000000af00000000000000b000000000",
            INIT_5A => X"0000008e00000000000000a000000000000000c000000000000000d000000000",
            INIT_5B => X"00000095000000000000009b00000000000000a800000000000000aa00000000",
            INIT_5C => X"00000064000000000000007f0000000000000085000000000000008d00000000",
            INIT_5D => X"0000007b00000000000000800000000000000083000000000000007100000000",
            INIT_5E => X"00000072000000000000006c0000000000000072000000000000007e00000000",
            INIT_5F => X"0000008900000000000000900000000000000090000000000000008200000000",
            INIT_60 => X"000000b700000000000000c000000000000000c400000000000000d200000000",
            INIT_61 => X"000000d200000000000000c000000000000000a600000000000000a900000000",
            INIT_62 => X"000000b400000000000000b600000000000000c000000000000000d100000000",
            INIT_63 => X"0000008c000000000000008d000000000000009900000000000000ab00000000",
            INIT_64 => X"0000005c000000000000006f000000000000007d000000000000008600000000",
            INIT_65 => X"0000007f000000000000007e000000000000007e000000000000007800000000",
            INIT_66 => X"0000007400000000000000690000000000000072000000000000007e00000000",
            INIT_67 => X"00000081000000000000008d0000000000000090000000000000008500000000",
            INIT_68 => X"000000b900000000000000b300000000000000b300000000000000c400000000",
            INIT_69 => X"000000cc00000000000000b5000000000000009700000000000000a600000000",
            INIT_6A => X"000000b300000000000000ba00000000000000c200000000000000cd00000000",
            INIT_6B => X"000000880000000000000085000000000000009200000000000000a600000000",
            INIT_6C => X"00000061000000000000005d0000000000000072000000000000007e00000000",
            INIT_6D => X"0000008000000000000000780000000000000073000000000000007800000000",
            INIT_6E => X"0000007e00000000000000710000000000000071000000000000008000000000",
            INIT_6F => X"0000007b00000000000000820000000000000083000000000000008400000000",
            INIT_70 => X"000000b800000000000000aa00000000000000a100000000000000b100000000",
            INIT_71 => X"000000c3000000000000009c000000000000008c00000000000000ae00000000",
            INIT_72 => X"000000b600000000000000bf00000000000000c100000000000000c900000000",
            INIT_73 => X"00000073000000000000006c0000000000000071000000000000009100000000",
            INIT_74 => X"0000006e0000000000000059000000000000006a000000000000007600000000",
            INIT_75 => X"0000008300000000000000780000000000000070000000000000007200000000",
            INIT_76 => X"0000007c000000000000007f000000000000007a000000000000007b00000000",
            INIT_77 => X"000000860000000000000082000000000000007a000000000000007500000000",
            INIT_78 => X"000000a10000000000000097000000000000008c000000000000009d00000000",
            INIT_79 => X"000000b10000000000000080000000000000008200000000000000a600000000",
            INIT_7A => X"0000009a00000000000000af00000000000000b700000000000000bf00000000",
            INIT_7B => X"0000005300000000000000470000000000000053000000000000007000000000",
            INIT_7C => X"0000006e0000000000000065000000000000005e000000000000006300000000",
            INIT_7D => X"0000007e0000000000000079000000000000006c000000000000006c00000000",
            INIT_7E => X"0000006b000000000000006f000000000000007a000000000000007900000000",
            INIT_7F => X"0000008400000000000000890000000000000084000000000000007300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE51;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE52 : if BRAM_NAME = "sampleifmap_layersamples_instance52" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000280000000000000013000000000000001c000000000000001700000000",
            INIT_01 => X"00000074000000000000006d0000000000000073000000000000007100000000",
            INIT_02 => X"00000069000000000000006a0000000000000067000000000000007100000000",
            INIT_03 => X"0000006b00000000000000690000000000000069000000000000006900000000",
            INIT_04 => X"0000003a000000000000004c0000000000000063000000000000006a00000000",
            INIT_05 => X"0000008900000000000000720000000000000056000000000000005400000000",
            INIT_06 => X"0000007d000000000000007c000000000000007d000000000000007c00000000",
            INIT_07 => X"00000078000000000000007a000000000000007d000000000000007f00000000",
            INIT_08 => X"0000001a0000000000000014000000000000001b000000000000001800000000",
            INIT_09 => X"0000007c00000000000000760000000000000082000000000000006a00000000",
            INIT_0A => X"00000075000000000000006d0000000000000072000000000000007d00000000",
            INIT_0B => X"0000007900000000000000720000000000000076000000000000007800000000",
            INIT_0C => X"00000044000000000000006a0000000000000083000000000000008500000000",
            INIT_0D => X"00000096000000000000008c0000000000000051000000000000003e00000000",
            INIT_0E => X"000000880000000000000089000000000000008c000000000000008a00000000",
            INIT_0F => X"0000008000000000000000810000000000000085000000000000008800000000",
            INIT_10 => X"000000120000000000000017000000000000001a000000000000001800000000",
            INIT_11 => X"0000007b00000000000000740000000000000083000000000000005800000000",
            INIT_12 => X"000000740000000000000074000000000000008d000000000000008b00000000",
            INIT_13 => X"00000084000000000000007d000000000000007f000000000000008100000000",
            INIT_14 => X"000000690000000000000098000000000000009a000000000000008e00000000",
            INIT_15 => X"0000009e000000000000009f0000000000000059000000000000003700000000",
            INIT_16 => X"0000008e00000000000000920000000000000097000000000000009700000000",
            INIT_17 => X"000000840000000000000088000000000000008b000000000000008e00000000",
            INIT_18 => X"0000001200000000000000190000000000000019000000000000001800000000",
            INIT_19 => X"00000073000000000000006a000000000000007c000000000000004500000000",
            INIT_1A => X"00000078000000000000009200000000000000a6000000000000009c00000000",
            INIT_1B => X"0000009700000000000000950000000000000094000000000000008900000000",
            INIT_1C => X"0000006d0000000000000094000000000000009c000000000000009600000000",
            INIT_1D => X"000000a900000000000000b1000000000000007a000000000000004a00000000",
            INIT_1E => X"000000950000000000000098000000000000009d00000000000000a100000000",
            INIT_1F => X"0000008e00000000000000910000000000000094000000000000009600000000",
            INIT_20 => X"0000001700000000000000190000000000000018000000000000001900000000",
            INIT_21 => X"000000680000000000000060000000000000006d000000000000003300000000",
            INIT_22 => X"0000008d00000000000000b200000000000000b800000000000000a100000000",
            INIT_23 => X"0000009300000000000000860000000000000080000000000000007c00000000",
            INIT_24 => X"0000006c00000000000000890000000000000096000000000000009700000000",
            INIT_25 => X"000000b500000000000000b70000000000000098000000000000006000000000",
            INIT_26 => X"000000a400000000000000a800000000000000ae00000000000000b300000000",
            INIT_27 => X"000000930000000000000098000000000000009c00000000000000a000000000",
            INIT_28 => X"0000001c000000000000001b000000000000001a000000000000001a00000000",
            INIT_29 => X"00000066000000000000005f0000000000000059000000000000002300000000",
            INIT_2A => X"0000009f00000000000000c700000000000000c1000000000000009600000000",
            INIT_2B => X"0000007600000000000000620000000000000066000000000000007400000000",
            INIT_2C => X"0000007a00000000000000770000000000000083000000000000008200000000",
            INIT_2D => X"000000aa00000000000000a600000000000000a7000000000000008400000000",
            INIT_2E => X"000000b700000000000000b300000000000000b700000000000000b200000000",
            INIT_2F => X"000000a900000000000000af00000000000000b100000000000000b700000000",
            INIT_30 => X"0000001a00000000000000190000000000000016000000000000001a00000000",
            INIT_31 => X"0000007b0000000000000080000000000000005c000000000000001d00000000",
            INIT_32 => X"000000ab00000000000000c700000000000000c3000000000000009300000000",
            INIT_33 => X"0000006a0000000000000063000000000000005e000000000000007e00000000",
            INIT_34 => X"0000007a0000000000000065000000000000006d000000000000006000000000",
            INIT_35 => X"000000b000000000000000aa00000000000000c000000000000000ac00000000",
            INIT_36 => X"000000ca00000000000000c500000000000000c400000000000000c300000000",
            INIT_37 => X"000000c200000000000000bf00000000000000bf00000000000000c500000000",
            INIT_38 => X"0000001900000000000000110000000000000021000000000000004d00000000",
            INIT_39 => X"0000007e000000000000009b000000000000009a000000000000005800000000",
            INIT_3A => X"000000b900000000000000c100000000000000be000000000000008c00000000",
            INIT_3B => X"00000071000000000000007b000000000000008100000000000000a300000000",
            INIT_3C => X"0000007900000000000000680000000000000067000000000000005800000000",
            INIT_3D => X"000000bd00000000000000a500000000000000c600000000000000b100000000",
            INIT_3E => X"000000da00000000000000e000000000000000db00000000000000e400000000",
            INIT_3F => X"000000cd00000000000000c400000000000000bb00000000000000ba00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006000000000000000560000000000000080000000000000009500000000",
            INIT_41 => X"00000077000000000000009900000000000000a7000000000000009b00000000",
            INIT_42 => X"000000bf00000000000000bf00000000000000a8000000000000006f00000000",
            INIT_43 => X"0000007f000000000000009400000000000000aa00000000000000b700000000",
            INIT_44 => X"0000007c00000000000000740000000000000070000000000000007000000000",
            INIT_45 => X"000000c100000000000000a200000000000000bb00000000000000a300000000",
            INIT_46 => X"000000bb00000000000000cf00000000000000d500000000000000df00000000",
            INIT_47 => X"000000d200000000000000c400000000000000a6000000000000009d00000000",
            INIT_48 => X"0000009b0000000000000092000000000000009e00000000000000a100000000",
            INIT_49 => X"00000075000000000000009f00000000000000a900000000000000a700000000",
            INIT_4A => X"000000b500000000000000b3000000000000009b000000000000006800000000",
            INIT_4B => X"00000087000000000000009f00000000000000b400000000000000b600000000",
            INIT_4C => X"0000007900000000000000750000000000000074000000000000006400000000",
            INIT_4D => X"000000cc00000000000000b200000000000000b2000000000000009e00000000",
            INIT_4E => X"000000a700000000000000cb00000000000000d600000000000000d800000000",
            INIT_4F => X"000000cf00000000000000b00000000000000096000000000000009300000000",
            INIT_50 => X"000000a5000000000000009e00000000000000a500000000000000aa00000000",
            INIT_51 => X"0000007000000000000000a000000000000000b000000000000000af00000000",
            INIT_52 => X"000000b400000000000000b100000000000000a4000000000000007b00000000",
            INIT_53 => X"00000079000000000000009500000000000000ac00000000000000b600000000",
            INIT_54 => X"0000007600000000000000750000000000000074000000000000006a00000000",
            INIT_55 => X"000000d100000000000000af00000000000000a6000000000000009c00000000",
            INIT_56 => X"000000a900000000000000cd00000000000000d800000000000000de00000000",
            INIT_57 => X"000000ba000000000000009f0000000000000093000000000000009100000000",
            INIT_58 => X"000000a600000000000000a900000000000000ae00000000000000ac00000000",
            INIT_59 => X"0000007a000000000000009d00000000000000b000000000000000b000000000",
            INIT_5A => X"000000b600000000000000b900000000000000b1000000000000008d00000000",
            INIT_5B => X"00000068000000000000007f000000000000009d00000000000000b600000000",
            INIT_5C => X"0000007d000000000000007b0000000000000084000000000000007300000000",
            INIT_5D => X"000000ce00000000000000a300000000000000a4000000000000009f00000000",
            INIT_5E => X"000000b500000000000000cd00000000000000d900000000000000e000000000",
            INIT_5F => X"0000009c0000000000000093000000000000008e000000000000009200000000",
            INIT_60 => X"000000a000000000000000a500000000000000a700000000000000a700000000",
            INIT_61 => X"0000008f000000000000009900000000000000a400000000000000a500000000",
            INIT_62 => X"000000a400000000000000ae00000000000000a3000000000000009100000000",
            INIT_63 => X"000000760000000000000085000000000000009f00000000000000a300000000",
            INIT_64 => X"000000920000000000000087000000000000009f000000000000008600000000",
            INIT_65 => X"000000cd00000000000000a800000000000000a300000000000000a300000000",
            INIT_66 => X"000000c700000000000000d600000000000000dc00000000000000df00000000",
            INIT_67 => X"000000980000000000000090000000000000009000000000000000a300000000",
            INIT_68 => X"0000009b00000000000000a000000000000000a200000000000000a900000000",
            INIT_69 => X"000000a40000000000000083000000000000008800000000000000a300000000",
            INIT_6A => X"0000008500000000000000840000000000000088000000000000009200000000",
            INIT_6B => X"000000920000000000000087000000000000009e000000000000009f00000000",
            INIT_6C => X"0000009e000000000000009000000000000000a200000000000000a700000000",
            INIT_6D => X"000000cb00000000000000b00000000000000098000000000000009800000000",
            INIT_6E => X"000000da00000000000000dd00000000000000d800000000000000d700000000",
            INIT_6F => X"000000b600000000000000a2000000000000009f00000000000000c500000000",
            INIT_70 => X"0000009d00000000000000a200000000000000a400000000000000ae00000000",
            INIT_71 => X"000000b2000000000000006d000000000000007800000000000000a800000000",
            INIT_72 => X"000000a300000000000000a100000000000000a700000000000000a600000000",
            INIT_73 => X"00000078000000000000008400000000000000ab00000000000000b600000000",
            INIT_74 => X"00000095000000000000008c00000000000000a300000000000000a900000000",
            INIT_75 => X"000000cc00000000000000aa00000000000000a400000000000000a600000000",
            INIT_76 => X"000000e400000000000000da00000000000000d500000000000000d300000000",
            INIT_77 => X"000000c700000000000000bb00000000000000b000000000000000d600000000",
            INIT_78 => X"0000009f00000000000000a100000000000000a000000000000000af00000000",
            INIT_79 => X"000000b70000000000000068000000000000008400000000000000aa00000000",
            INIT_7A => X"000000b000000000000000b800000000000000b600000000000000bc00000000",
            INIT_7B => X"0000008d00000000000000a300000000000000a800000000000000a200000000",
            INIT_7C => X"00000085000000000000009200000000000000a5000000000000009100000000",
            INIT_7D => X"000000a9000000000000009600000000000000a500000000000000af00000000",
            INIT_7E => X"000000dd00000000000000d900000000000000d400000000000000ca00000000",
            INIT_7F => X"000000c700000000000000c700000000000000ba00000000000000c400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE52;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE53 : if BRAM_NAME = "sampleifmap_layersamples_instance53" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000940000000000000092000000000000009f00000000000000b300000000",
            INIT_01 => X"000000a8000000000000006d000000000000009700000000000000a100000000",
            INIT_02 => X"000000ae00000000000000a400000000000000b500000000000000c700000000",
            INIT_03 => X"000000a600000000000000aa000000000000009c00000000000000a500000000",
            INIT_04 => X"00000077000000000000009f0000000000000088000000000000006900000000",
            INIT_05 => X"00000050000000000000007e000000000000009e000000000000008f00000000",
            INIT_06 => X"000000cd00000000000000d100000000000000b7000000000000007600000000",
            INIT_07 => X"000000c500000000000000c900000000000000b700000000000000af00000000",
            INIT_08 => X"00000083000000000000008500000000000000a400000000000000b500000000",
            INIT_09 => X"0000009f000000000000009700000000000000a5000000000000009500000000",
            INIT_0A => X"000000cd00000000000000c400000000000000c700000000000000c200000000",
            INIT_0B => X"000000a200000000000000ac00000000000000a800000000000000b900000000",
            INIT_0C => X"00000077000000000000009b0000000000000069000000000000006800000000",
            INIT_0D => X"0000005c000000000000008800000000000000ad000000000000008600000000",
            INIT_0E => X"0000009e0000000000000098000000000000006f000000000000004b00000000",
            INIT_0F => X"000000c800000000000000cb00000000000000b0000000000000009800000000",
            INIT_10 => X"00000085000000000000008e00000000000000ac00000000000000b700000000",
            INIT_11 => X"000000aa00000000000000b100000000000000b0000000000000009f00000000",
            INIT_12 => X"000000d900000000000000cf00000000000000c500000000000000b100000000",
            INIT_13 => X"000000aa00000000000000bb00000000000000c600000000000000d900000000",
            INIT_14 => X"0000007e0000000000000085000000000000005a000000000000008300000000",
            INIT_15 => X"0000007e000000000000008200000000000000a2000000000000008b00000000",
            INIT_16 => X"0000008400000000000000760000000000000060000000000000006f00000000",
            INIT_17 => X"000000c700000000000000b80000000000000092000000000000007c00000000",
            INIT_18 => X"0000009500000000000000a100000000000000b000000000000000b900000000",
            INIT_19 => X"000000bc00000000000000b600000000000000b700000000000000af00000000",
            INIT_1A => X"000000c200000000000000b900000000000000aa00000000000000aa00000000",
            INIT_1B => X"000000af00000000000000ca00000000000000d000000000000000c900000000",
            INIT_1C => X"000000910000000000000071000000000000007b00000000000000a400000000",
            INIT_1D => X"0000007b0000000000000071000000000000008c000000000000009d00000000",
            INIT_1E => X"0000008e00000000000000860000000000000070000000000000007700000000",
            INIT_1F => X"000000a600000000000000840000000000000079000000000000007f00000000",
            INIT_20 => X"0000009b00000000000000ad00000000000000b700000000000000bd00000000",
            INIT_21 => X"000000b200000000000000b100000000000000ba00000000000000ab00000000",
            INIT_22 => X"000000b100000000000000b200000000000000ac00000000000000b400000000",
            INIT_23 => X"000000bd00000000000000c300000000000000bc00000000000000a400000000",
            INIT_24 => X"0000009d000000000000008800000000000000b600000000000000c900000000",
            INIT_25 => X"0000007c000000000000006a0000000000000078000000000000009300000000",
            INIT_26 => X"0000008a0000000000000094000000000000008a000000000000008000000000",
            INIT_27 => X"00000082000000000000007a0000000000000077000000000000007800000000",
            INIT_28 => X"000000a100000000000000b700000000000000bc00000000000000bd00000000",
            INIT_29 => X"000000b000000000000000bb00000000000000b7000000000000009e00000000",
            INIT_2A => X"000000a400000000000000c000000000000000bf00000000000000b800000000",
            INIT_2B => X"000000b100000000000000ad00000000000000a6000000000000008b00000000",
            INIT_2C => X"0000009600000000000000a200000000000000bc00000000000000c000000000",
            INIT_2D => X"000000850000000000000079000000000000006b000000000000007600000000",
            INIT_2E => X"0000007d000000000000008d0000000000000096000000000000008e00000000",
            INIT_2F => X"0000006c000000000000007d000000000000007c000000000000007500000000",
            INIT_30 => X"000000a600000000000000bb00000000000000ba00000000000000ba00000000",
            INIT_31 => X"000000c500000000000000c700000000000000b4000000000000009400000000",
            INIT_32 => X"000000a800000000000000c000000000000000c300000000000000c100000000",
            INIT_33 => X"000000aa00000000000000a9000000000000009f000000000000009100000000",
            INIT_34 => X"0000008600000000000000a300000000000000ac00000000000000af00000000",
            INIT_35 => X"0000008b0000000000000086000000000000006c000000000000005d00000000",
            INIT_36 => X"0000007c000000000000008e0000000000000097000000000000008d00000000",
            INIT_37 => X"0000005b00000000000000650000000000000072000000000000007c00000000",
            INIT_38 => X"000000ac00000000000000b700000000000000b500000000000000ba00000000",
            INIT_39 => X"000000cf00000000000000c900000000000000b0000000000000008f00000000",
            INIT_3A => X"000000af00000000000000bd00000000000000cb00000000000000ce00000000",
            INIT_3B => X"000000ac00000000000000ae00000000000000ab00000000000000a500000000",
            INIT_3C => X"00000075000000000000009e00000000000000ab00000000000000b200000000",
            INIT_3D => X"00000088000000000000008a0000000000000078000000000000006100000000",
            INIT_3E => X"00000084000000000000009200000000000000a1000000000000008a00000000",
            INIT_3F => X"000000680000000000000064000000000000006d000000000000008200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a900000000000000af00000000000000b200000000000000b800000000",
            INIT_41 => X"000000ca00000000000000c600000000000000aa000000000000009200000000",
            INIT_42 => X"0000008800000000000000ab00000000000000c500000000000000c800000000",
            INIT_43 => X"000000aa00000000000000ab00000000000000b400000000000000a100000000",
            INIT_44 => X"00000073000000000000009000000000000000a800000000000000ad00000000",
            INIT_45 => X"0000007e0000000000000086000000000000007c000000000000006c00000000",
            INIT_46 => X"0000008700000000000000910000000000000099000000000000008200000000",
            INIT_47 => X"0000006f00000000000000740000000000000075000000000000007700000000",
            INIT_48 => X"0000009d00000000000000a800000000000000b000000000000000b800000000",
            INIT_49 => X"000000c800000000000000c000000000000000a2000000000000009300000000",
            INIT_4A => X"00000052000000000000008100000000000000b900000000000000bf00000000",
            INIT_4B => X"0000009f00000000000000a600000000000000b3000000000000008d00000000",
            INIT_4C => X"0000007400000000000000840000000000000096000000000000009f00000000",
            INIT_4D => X"0000007a000000000000007f000000000000007a000000000000006900000000",
            INIT_4E => X"0000007a00000000000000800000000000000084000000000000007f00000000",
            INIT_4F => X"00000062000000000000006b0000000000000077000000000000007700000000",
            INIT_50 => X"0000009400000000000000a300000000000000ac00000000000000b800000000",
            INIT_51 => X"000000ca00000000000000ba0000000000000092000000000000008600000000",
            INIT_52 => X"00000058000000000000008200000000000000b200000000000000c000000000",
            INIT_53 => X"00000090000000000000009800000000000000ac000000000000008c00000000",
            INIT_54 => X"00000069000000000000007a0000000000000084000000000000009100000000",
            INIT_55 => X"0000007000000000000000790000000000000077000000000000006400000000",
            INIT_56 => X"0000006c00000000000000640000000000000071000000000000007a00000000",
            INIT_57 => X"000000720000000000000075000000000000007a000000000000007c00000000",
            INIT_58 => X"0000008e000000000000009e00000000000000a900000000000000b700000000",
            INIT_59 => X"000000cc00000000000000b20000000000000084000000000000007e00000000",
            INIT_5A => X"00000090000000000000009d00000000000000af00000000000000c300000000",
            INIT_5B => X"000000830000000000000087000000000000009800000000000000a400000000",
            INIT_5C => X"00000054000000000000006f0000000000000074000000000000007c00000000",
            INIT_5D => X"0000006d00000000000000710000000000000073000000000000006100000000",
            INIT_5E => X"00000064000000000000005f0000000000000066000000000000007200000000",
            INIT_5F => X"0000007b00000000000000820000000000000082000000000000007400000000",
            INIT_60 => X"0000008e000000000000009900000000000000a100000000000000b100000000",
            INIT_61 => X"000000cc00000000000000b2000000000000007a000000000000007700000000",
            INIT_62 => X"000000a800000000000000aa00000000000000b400000000000000c500000000",
            INIT_63 => X"0000007b000000000000007a0000000000000087000000000000009d00000000",
            INIT_64 => X"0000004b000000000000005e000000000000006d000000000000007700000000",
            INIT_65 => X"000000710000000000000070000000000000006f000000000000006800000000",
            INIT_66 => X"00000066000000000000005c0000000000000064000000000000007000000000",
            INIT_67 => X"00000073000000000000007e0000000000000082000000000000007700000000",
            INIT_68 => X"00000091000000000000008d000000000000009000000000000000a300000000",
            INIT_69 => X"000000c800000000000000a9000000000000006b000000000000007400000000",
            INIT_6A => X"000000a300000000000000ac00000000000000b700000000000000c200000000",
            INIT_6B => X"0000007900000000000000730000000000000081000000000000009600000000",
            INIT_6C => X"00000051000000000000004e0000000000000064000000000000007000000000",
            INIT_6D => X"00000072000000000000006a0000000000000065000000000000006800000000",
            INIT_6E => X"0000007000000000000000630000000000000063000000000000007200000000",
            INIT_6F => X"0000006e00000000000000740000000000000075000000000000007600000000",
            INIT_70 => X"0000008f0000000000000083000000000000007e000000000000008e00000000",
            INIT_71 => X"000000c00000000000000091000000000000005f000000000000007c00000000",
            INIT_72 => X"000000a800000000000000b200000000000000b700000000000000be00000000",
            INIT_73 => X"00000065000000000000005c0000000000000062000000000000008200000000",
            INIT_74 => X"0000005f000000000000004b000000000000005c000000000000006800000000",
            INIT_75 => X"00000074000000000000006a0000000000000061000000000000006300000000",
            INIT_76 => X"0000006e0000000000000071000000000000006c000000000000006d00000000",
            INIT_77 => X"000000770000000000000074000000000000006c000000000000006700000000",
            INIT_78 => X"0000007800000000000000700000000000000068000000000000007b00000000",
            INIT_79 => X"000000ae00000000000000760000000000000057000000000000007400000000",
            INIT_7A => X"0000008d00000000000000a400000000000000ae00000000000000b500000000",
            INIT_7B => X"0000004600000000000000390000000000000045000000000000006300000000",
            INIT_7C => X"0000006000000000000000580000000000000051000000000000005700000000",
            INIT_7D => X"00000070000000000000006b000000000000005e000000000000005d00000000",
            INIT_7E => X"0000005d0000000000000061000000000000006c000000000000006b00000000",
            INIT_7F => X"00000076000000000000007b0000000000000076000000000000006500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE53;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE54 : if BRAM_NAME = "sampleifmap_layersamples_instance54" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000c700000000000000cd00000000000000d200000000000000d900000000",
            INIT_01 => X"000000bd00000000000000cf00000000000000d600000000000000da00000000",
            INIT_02 => X"000000a900000000000000a600000000000000ae00000000000000bb00000000",
            INIT_03 => X"0000008f000000000000008c000000000000009a000000000000009600000000",
            INIT_04 => X"000000df00000000000000db00000000000000bf00000000000000a700000000",
            INIT_05 => X"000000e100000000000000e200000000000000d700000000000000db00000000",
            INIT_06 => X"000000bb00000000000000af00000000000000be00000000000000db00000000",
            INIT_07 => X"000000a200000000000000a100000000000000aa00000000000000c800000000",
            INIT_08 => X"000000d700000000000000dc00000000000000dd00000000000000de00000000",
            INIT_09 => X"000000b300000000000000d300000000000000e100000000000000d800000000",
            INIT_0A => X"000000bc00000000000000be00000000000000c000000000000000b400000000",
            INIT_0B => X"000000db00000000000000d100000000000000ce00000000000000c700000000",
            INIT_0C => X"000000ec00000000000000ec00000000000000eb00000000000000e500000000",
            INIT_0D => X"000000e500000000000000e100000000000000e200000000000000e900000000",
            INIT_0E => X"000000cd00000000000000d000000000000000d400000000000000e700000000",
            INIT_0F => X"000000c800000000000000ba00000000000000b700000000000000d800000000",
            INIT_10 => X"000000e800000000000000e700000000000000e900000000000000ea00000000",
            INIT_11 => X"000000ad00000000000000d900000000000000ef00000000000000e900000000",
            INIT_12 => X"000000b700000000000000ad00000000000000b400000000000000a400000000",
            INIT_13 => X"000000e000000000000000d400000000000000bc00000000000000be00000000",
            INIT_14 => X"000000e100000000000000e300000000000000eb00000000000000da00000000",
            INIT_15 => X"000000e100000000000000d600000000000000df00000000000000e500000000",
            INIT_16 => X"000000d800000000000000e600000000000000e800000000000000ea00000000",
            INIT_17 => X"000000d300000000000000d000000000000000ca00000000000000d100000000",
            INIT_18 => X"000000f200000000000000f400000000000000f400000000000000f500000000",
            INIT_19 => X"0000009e00000000000000e400000000000000f300000000000000f400000000",
            INIT_1A => X"0000009f0000000000000083000000000000009d000000000000009200000000",
            INIT_1B => X"0000009f00000000000000a20000000000000088000000000000009100000000",
            INIT_1C => X"000000d300000000000000c300000000000000cb00000000000000a900000000",
            INIT_1D => X"000000e200000000000000d000000000000000cb00000000000000d100000000",
            INIT_1E => X"000000d500000000000000e400000000000000e900000000000000e600000000",
            INIT_1F => X"000000d400000000000000e000000000000000db00000000000000c700000000",
            INIT_20 => X"000000f400000000000000f400000000000000f300000000000000f500000000",
            INIT_21 => X"0000007500000000000000cf00000000000000f100000000000000f500000000",
            INIT_22 => X"0000006b0000000000000059000000000000006c000000000000006300000000",
            INIT_23 => X"0000005c0000000000000064000000000000005b000000000000006400000000",
            INIT_24 => X"00000095000000000000007c000000000000007c000000000000006600000000",
            INIT_25 => X"000000e900000000000000ca00000000000000b900000000000000b600000000",
            INIT_26 => X"000000cd00000000000000e300000000000000e200000000000000e100000000",
            INIT_27 => X"000000de00000000000000e200000000000000d500000000000000c200000000",
            INIT_28 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_29 => X"0000007e00000000000000d800000000000000ed00000000000000f500000000",
            INIT_2A => X"00000066000000000000005b000000000000005a000000000000004800000000",
            INIT_2B => X"00000063000000000000006b0000000000000067000000000000006500000000",
            INIT_2C => X"0000005d000000000000005b0000000000000059000000000000005900000000",
            INIT_2D => X"000000eb00000000000000d800000000000000be000000000000007e00000000",
            INIT_2E => X"000000c400000000000000d800000000000000df00000000000000e700000000",
            INIT_2F => X"000000ec00000000000000d900000000000000bd00000000000000ae00000000",
            INIT_30 => X"000000f400000000000000f300000000000000f300000000000000f500000000",
            INIT_31 => X"0000009e00000000000000d900000000000000db00000000000000f100000000",
            INIT_32 => X"0000009700000000000000840000000000000072000000000000005000000000",
            INIT_33 => X"0000008a000000000000008f0000000000000084000000000000008c00000000",
            INIT_34 => X"000000780000000000000072000000000000007a000000000000008200000000",
            INIT_35 => X"000000e900000000000000dd000000000000009b000000000000006e00000000",
            INIT_36 => X"000000c000000000000000c600000000000000e000000000000000eb00000000",
            INIT_37 => X"000000eb00000000000000cc00000000000000ab00000000000000a700000000",
            INIT_38 => X"000000f600000000000000f300000000000000f300000000000000f400000000",
            INIT_39 => X"0000009900000000000000d700000000000000c700000000000000e300000000",
            INIT_3A => X"000000ca00000000000000bb0000000000000092000000000000005100000000",
            INIT_3B => X"000000830000000000000083000000000000009e00000000000000cf00000000",
            INIT_3C => X"000000840000000000000083000000000000008d000000000000008100000000",
            INIT_3D => X"000000d7000000000000009f0000000000000084000000000000009f00000000",
            INIT_3E => X"000000d100000000000000d400000000000000d700000000000000e500000000",
            INIT_3F => X"000000dd00000000000000b200000000000000ab00000000000000c500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f500000000000000f400000000000000f300000000000000f400000000",
            INIT_41 => X"0000008200000000000000da00000000000000ce00000000000000e300000000",
            INIT_42 => X"0000008100000000000000800000000000000082000000000000005100000000",
            INIT_43 => X"0000007d0000000000000074000000000000009100000000000000b800000000",
            INIT_44 => X"0000007d000000000000008e0000000000000089000000000000007c00000000",
            INIT_45 => X"000000c600000000000000900000000000000093000000000000009900000000",
            INIT_46 => X"000000dc00000000000000e900000000000000db00000000000000d600000000",
            INIT_47 => X"000000c900000000000000a900000000000000a400000000000000b800000000",
            INIT_48 => X"000000f200000000000000f400000000000000f300000000000000f300000000",
            INIT_49 => X"0000006e00000000000000a800000000000000be00000000000000e400000000",
            INIT_4A => X"0000006e00000000000000770000000000000086000000000000005300000000",
            INIT_4B => X"0000007800000000000000730000000000000080000000000000008f00000000",
            INIT_4C => X"0000007d00000000000000920000000000000083000000000000007d00000000",
            INIT_4D => X"000000c4000000000000008c000000000000009b000000000000009500000000",
            INIT_4E => X"000000e900000000000000f000000000000000f000000000000000e900000000",
            INIT_4F => X"000000dc00000000000000d700000000000000c800000000000000c800000000",
            INIT_50 => X"000000f500000000000000f400000000000000f100000000000000ef00000000",
            INIT_51 => X"0000005f0000000000000082000000000000008500000000000000dc00000000",
            INIT_52 => X"0000006c00000000000000740000000000000074000000000000004e00000000",
            INIT_53 => X"0000006c000000000000006d000000000000006b000000000000006d00000000",
            INIT_54 => X"0000007300000000000000780000000000000078000000000000007300000000",
            INIT_55 => X"000000a7000000000000008f0000000000000096000000000000008800000000",
            INIT_56 => X"000000f300000000000000f500000000000000e400000000000000d000000000",
            INIT_57 => X"000000f400000000000000f500000000000000f500000000000000f400000000",
            INIT_58 => X"000000f400000000000000f200000000000000e900000000000000de00000000",
            INIT_59 => X"0000005900000000000000a500000000000000a900000000000000d800000000",
            INIT_5A => X"00000064000000000000005b0000000000000043000000000000003d00000000",
            INIT_5B => X"000000600000000000000062000000000000005f000000000000005f00000000",
            INIT_5C => X"00000061000000000000005a000000000000005f000000000000006000000000",
            INIT_5D => X"0000007e00000000000000810000000000000079000000000000006900000000",
            INIT_5E => X"000000f300000000000000f800000000000000d8000000000000009b00000000",
            INIT_5F => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_60 => X"000000e300000000000000ec00000000000000df00000000000000d000000000",
            INIT_61 => X"0000006400000000000000b500000000000000b700000000000000bf00000000",
            INIT_62 => X"0000006500000000000000580000000000000038000000000000003700000000",
            INIT_63 => X"0000005400000000000000560000000000000063000000000000006f00000000",
            INIT_64 => X"00000071000000000000005d0000000000000054000000000000005200000000",
            INIT_65 => X"0000008100000000000000700000000000000062000000000000006d00000000",
            INIT_66 => X"000000f400000000000000f500000000000000e200000000000000ae00000000",
            INIT_67 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_68 => X"000000c300000000000000db00000000000000cc00000000000000c800000000",
            INIT_69 => X"00000066000000000000009c000000000000009a00000000000000aa00000000",
            INIT_6A => X"00000066000000000000006c0000000000000063000000000000006800000000",
            INIT_6B => X"00000055000000000000005e0000000000000075000000000000007300000000",
            INIT_6C => X"0000008c000000000000007a000000000000006a000000000000005a00000000",
            INIT_6D => X"0000007c000000000000006c0000000000000068000000000000008000000000",
            INIT_6E => X"000000d400000000000000c300000000000000b3000000000000009600000000",
            INIT_6F => X"000000f400000000000000f400000000000000f500000000000000ef00000000",
            INIT_70 => X"000000a900000000000000cf00000000000000d200000000000000c800000000",
            INIT_71 => X"0000008a0000000000000093000000000000009400000000000000a400000000",
            INIT_72 => X"0000005d000000000000006a000000000000005c000000000000008100000000",
            INIT_73 => X"0000004d0000000000000054000000000000005d000000000000005900000000",
            INIT_74 => X"0000005100000000000000510000000000000051000000000000004c00000000",
            INIT_75 => X"00000052000000000000004b000000000000004a000000000000004f00000000",
            INIT_76 => X"0000008f000000000000008c000000000000007b000000000000006500000000",
            INIT_77 => X"000000f400000000000000f400000000000000f400000000000000bf00000000",
            INIT_78 => X"0000007700000000000000c400000000000000e200000000000000d200000000",
            INIT_79 => X"000000c000000000000000ba0000000000000096000000000000007000000000",
            INIT_7A => X"00000037000000000000004d000000000000004d000000000000006c00000000",
            INIT_7B => X"0000003f000000000000003c000000000000002f000000000000002d00000000",
            INIT_7C => X"00000036000000000000003b000000000000003f000000000000003b00000000",
            INIT_7D => X"00000040000000000000003d0000000000000032000000000000003100000000",
            INIT_7E => X"00000067000000000000005b000000000000004b000000000000004700000000",
            INIT_7F => X"000000f400000000000000f600000000000000e1000000000000008700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE54;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE55 : if BRAM_NAME = "sampleifmap_layersamples_instance55" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000006000000000000000b400000000000000c100000000000000c700000000",
            INIT_01 => X"000000a100000000000000c00000000000000091000000000000005d00000000",
            INIT_02 => X"00000062000000000000005c0000000000000049000000000000005600000000",
            INIT_03 => X"00000047000000000000004f000000000000004f000000000000006800000000",
            INIT_04 => X"0000001b000000000000001e000000000000001c000000000000002500000000",
            INIT_05 => X"0000001c00000000000000160000000000000032000000000000003400000000",
            INIT_06 => X"00000068000000000000005b0000000000000035000000000000001800000000",
            INIT_07 => X"000000f300000000000000f700000000000000ce000000000000008000000000",
            INIT_08 => X"0000007100000000000000c200000000000000c700000000000000d300000000",
            INIT_09 => X"00000047000000000000009f000000000000009d000000000000007800000000",
            INIT_0A => X"0000007c0000000000000074000000000000005a000000000000004400000000",
            INIT_0B => X"0000006600000000000000800000000000000079000000000000009500000000",
            INIT_0C => X"0000006400000000000000700000000000000062000000000000004e00000000",
            INIT_0D => X"00000063000000000000005c0000000000000093000000000000009400000000",
            INIT_0E => X"0000008e0000000000000087000000000000006c000000000000005e00000000",
            INIT_0F => X"000000f500000000000000f200000000000000b7000000000000009c00000000",
            INIT_10 => X"0000006600000000000000b700000000000000ca00000000000000dc00000000",
            INIT_11 => X"0000001e000000000000008400000000000000a5000000000000006e00000000",
            INIT_12 => X"00000053000000000000006b0000000000000062000000000000003900000000",
            INIT_13 => X"0000006400000000000000810000000000000065000000000000005200000000",
            INIT_14 => X"0000009f000000000000009e00000000000000ae000000000000009900000000",
            INIT_15 => X"000000a300000000000000a200000000000000a800000000000000ac00000000",
            INIT_16 => X"00000077000000000000009c00000000000000af00000000000000a000000000",
            INIT_17 => X"000000f700000000000000e40000000000000087000000000000007200000000",
            INIT_18 => X"0000006200000000000000bc00000000000000cf00000000000000db00000000",
            INIT_19 => X"0000002a000000000000006f000000000000008d000000000000005300000000",
            INIT_1A => X"0000003e000000000000004c0000000000000048000000000000003a00000000",
            INIT_1B => X"0000005d00000000000000400000000000000038000000000000003500000000",
            INIT_1C => X"00000065000000000000005b000000000000007c00000000000000a000000000",
            INIT_1D => X"000000670000000000000067000000000000006b000000000000007400000000",
            INIT_1E => X"00000043000000000000007e000000000000009b000000000000006300000000",
            INIT_1F => X"000000f800000000000000d90000000000000076000000000000005100000000",
            INIT_20 => X"0000006500000000000000c700000000000000d200000000000000d900000000",
            INIT_21 => X"0000003c000000000000005d0000000000000058000000000000003800000000",
            INIT_22 => X"00000046000000000000003f000000000000002e000000000000003800000000",
            INIT_23 => X"0000004100000000000000400000000000000036000000000000003c00000000",
            INIT_24 => X"0000006700000000000000690000000000000072000000000000006300000000",
            INIT_25 => X"00000061000000000000005d0000000000000060000000000000006400000000",
            INIT_26 => X"000000490000000000000064000000000000006f000000000000006600000000",
            INIT_27 => X"000000f900000000000000d40000000000000072000000000000005200000000",
            INIT_28 => X"0000007500000000000000ca00000000000000cd00000000000000d100000000",
            INIT_29 => X"0000004400000000000000510000000000000046000000000000005300000000",
            INIT_2A => X"00000033000000000000002b0000000000000023000000000000003200000000",
            INIT_2B => X"0000003f0000000000000057000000000000004d000000000000004400000000",
            INIT_2C => X"0000004800000000000000520000000000000047000000000000003400000000",
            INIT_2D => X"0000005d000000000000003e0000000000000043000000000000004000000000",
            INIT_2E => X"0000006c0000000000000053000000000000003c000000000000005800000000",
            INIT_2F => X"000000fa00000000000000cc000000000000006c000000000000007000000000",
            INIT_30 => X"0000006800000000000000c500000000000000ca00000000000000cd00000000",
            INIT_31 => X"000000490000000000000047000000000000006f000000000000005d00000000",
            INIT_32 => X"0000002200000000000000260000000000000029000000000000003f00000000",
            INIT_33 => X"0000004f000000000000008e0000000000000063000000000000004b00000000",
            INIT_34 => X"0000007600000000000000930000000000000056000000000000001e00000000",
            INIT_35 => X"0000009900000000000000660000000000000072000000000000006300000000",
            INIT_36 => X"0000008d000000000000004a000000000000003f00000000000000b200000000",
            INIT_37 => X"000000f600000000000000c3000000000000005a000000000000007700000000",
            INIT_38 => X"0000005700000000000000b900000000000000c200000000000000c600000000",
            INIT_39 => X"000000630000000000000061000000000000006c000000000000003100000000",
            INIT_3A => X"0000002400000000000000270000000000000033000000000000005f00000000",
            INIT_3B => X"0000003700000000000000570000000000000032000000000000002800000000",
            INIT_3C => X"0000007f0000000000000097000000000000004f000000000000002000000000",
            INIT_3D => X"0000009c00000000000000740000000000000088000000000000007a00000000",
            INIT_3E => X"0000004a00000000000000350000000000000037000000000000009f00000000",
            INIT_3F => X"000000f000000000000000c2000000000000004e000000000000003e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004d00000000000000a900000000000000b400000000000000b600000000",
            INIT_41 => X"00000090000000000000006c000000000000003b000000000000002500000000",
            INIT_42 => X"00000020000000000000002b000000000000003c000000000000006a00000000",
            INIT_43 => X"00000021000000000000001e000000000000001c000000000000001d00000000",
            INIT_44 => X"00000058000000000000003a000000000000002a000000000000002700000000",
            INIT_45 => X"00000075000000000000007a0000000000000079000000000000006a00000000",
            INIT_46 => X"000000320000000000000033000000000000002f000000000000004300000000",
            INIT_47 => X"000000e100000000000000ba0000000000000050000000000000003300000000",
            INIT_48 => X"0000007d00000000000000a400000000000000a500000000000000a800000000",
            INIT_49 => X"0000008d000000000000006f0000000000000060000000000000005b00000000",
            INIT_4A => X"000000240000000000000037000000000000004a000000000000006000000000",
            INIT_4B => X"0000001f000000000000001d000000000000001e000000000000001e00000000",
            INIT_4C => X"000000ae00000000000000400000000000000018000000000000002300000000",
            INIT_4D => X"000000b500000000000000b300000000000000cb00000000000000cd00000000",
            INIT_4E => X"00000030000000000000002b0000000000000026000000000000005700000000",
            INIT_4F => X"000000d300000000000000ae000000000000005b000000000000004200000000",
            INIT_50 => X"000000b400000000000000af00000000000000a300000000000000a200000000",
            INIT_51 => X"0000008d000000000000006c0000000000000076000000000000009800000000",
            INIT_52 => X"00000030000000000000004e0000000000000053000000000000005b00000000",
            INIT_53 => X"0000001d00000000000000190000000000000018000000000000001900000000",
            INIT_54 => X"000000a400000000000000470000000000000026000000000000002700000000",
            INIT_55 => X"000000a600000000000000a900000000000000b100000000000000b800000000",
            INIT_56 => X"00000031000000000000001e000000000000001e000000000000005100000000",
            INIT_57 => X"000000ce00000000000000a9000000000000005f000000000000004e00000000",
            INIT_58 => X"000000a600000000000000b300000000000000ac000000000000009a00000000",
            INIT_59 => X"0000009200000000000000670000000000000075000000000000009200000000",
            INIT_5A => X"0000003600000000000000520000000000000055000000000000005700000000",
            INIT_5B => X"000000250000000000000021000000000000001e000000000000002000000000",
            INIT_5C => X"000000650000000000000056000000000000004d000000000000003600000000",
            INIT_5D => X"00000089000000000000008e0000000000000079000000000000006b00000000",
            INIT_5E => X"000000360000000000000021000000000000001e000000000000003c00000000",
            INIT_5F => X"000000c700000000000000a5000000000000005b000000000000004e00000000",
            INIT_60 => X"00000094000000000000009e00000000000000a900000000000000a600000000",
            INIT_61 => X"0000007100000000000000670000000000000085000000000000008f00000000",
            INIT_62 => X"0000003c000000000000004b0000000000000051000000000000004f00000000",
            INIT_63 => X"0000002c000000000000002a0000000000000027000000000000002a00000000",
            INIT_64 => X"0000004d00000000000000410000000000000036000000000000003000000000",
            INIT_65 => X"0000008b0000000000000083000000000000006e000000000000005a00000000",
            INIT_66 => X"000000360000000000000026000000000000001d000000000000003500000000",
            INIT_67 => X"000000c400000000000000a9000000000000005b000000000000004600000000",
            INIT_68 => X"0000008d0000000000000093000000000000009700000000000000a200000000",
            INIT_69 => X"0000004e000000000000006b0000000000000085000000000000008900000000",
            INIT_6A => X"0000003c0000000000000046000000000000004e000000000000004800000000",
            INIT_6B => X"00000030000000000000002e000000000000002a000000000000003200000000",
            INIT_6C => X"00000042000000000000003b0000000000000033000000000000003100000000",
            INIT_6D => X"0000007100000000000000650000000000000059000000000000004c00000000",
            INIT_6E => X"000000340000000000000023000000000000001d000000000000004500000000",
            INIT_6F => X"000000ba00000000000000ae0000000000000062000000000000003f00000000",
            INIT_70 => X"0000008c000000000000008e000000000000008d000000000000009400000000",
            INIT_71 => X"0000003c000000000000006a000000000000008c000000000000008f00000000",
            INIT_72 => X"000000370000000000000042000000000000004a000000000000004200000000",
            INIT_73 => X"0000003a00000000000000360000000000000034000000000000003900000000",
            INIT_74 => X"000000460000000000000041000000000000003a000000000000003a00000000",
            INIT_75 => X"0000005d00000000000000570000000000000050000000000000004900000000",
            INIT_76 => X"0000003700000000000000260000000000000025000000000000004d00000000",
            INIT_77 => X"000000b400000000000000b30000000000000083000000000000004a00000000",
            INIT_78 => X"000000a200000000000000a00000000000000095000000000000009000000000",
            INIT_79 => X"0000003d000000000000007e0000000000000092000000000000009e00000000",
            INIT_7A => X"00000043000000000000003a0000000000000039000000000000003900000000",
            INIT_7B => X"0000004800000000000000490000000000000045000000000000004600000000",
            INIT_7C => X"0000006200000000000000590000000000000049000000000000004400000000",
            INIT_7D => X"0000006100000000000000630000000000000061000000000000005e00000000",
            INIT_7E => X"0000004700000000000000400000000000000045000000000000005200000000",
            INIT_7F => X"000000ba00000000000000b600000000000000a4000000000000007700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE55;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE56 : if BRAM_NAME = "sampleifmap_layersamples_instance56" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ca00000000000000d000000000000000d000000000000000d700000000",
            INIT_01 => X"000000b900000000000000ca00000000000000d100000000000000d700000000",
            INIT_02 => X"000000a0000000000000009800000000000000a800000000000000b800000000",
            INIT_03 => X"0000009d000000000000009a00000000000000a7000000000000009d00000000",
            INIT_04 => X"000000e100000000000000e100000000000000cb00000000000000b500000000",
            INIT_05 => X"000000e400000000000000e500000000000000db00000000000000de00000000",
            INIT_06 => X"000000c400000000000000b800000000000000c500000000000000dd00000000",
            INIT_07 => X"000000a500000000000000b000000000000000b800000000000000d000000000",
            INIT_08 => X"000000d900000000000000e100000000000000e000000000000000e200000000",
            INIT_09 => X"000000ab00000000000000cc00000000000000dd00000000000000d500000000",
            INIT_0A => X"000000b100000000000000b200000000000000bd00000000000000b400000000",
            INIT_0B => X"000000e000000000000000d000000000000000cd00000000000000c400000000",
            INIT_0C => X"000000f300000000000000f200000000000000f000000000000000ec00000000",
            INIT_0D => X"000000e700000000000000e400000000000000e500000000000000ee00000000",
            INIT_0E => X"000000d200000000000000d400000000000000d600000000000000e700000000",
            INIT_0F => X"000000c500000000000000bf00000000000000be00000000000000de00000000",
            INIT_10 => X"000000eb00000000000000ea00000000000000ea00000000000000eb00000000",
            INIT_11 => X"000000a600000000000000d600000000000000ef00000000000000ea00000000",
            INIT_12 => X"000000b100000000000000a800000000000000b100000000000000a600000000",
            INIT_13 => X"000000df00000000000000ce00000000000000b700000000000000b800000000",
            INIT_14 => X"000000e800000000000000e300000000000000ec00000000000000dc00000000",
            INIT_15 => X"000000e000000000000000d900000000000000e400000000000000eb00000000",
            INIT_16 => X"000000dd00000000000000e600000000000000e900000000000000e900000000",
            INIT_17 => X"000000d200000000000000d100000000000000ce00000000000000d900000000",
            INIT_18 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_19 => X"0000009900000000000000e300000000000000f400000000000000f400000000",
            INIT_1A => X"0000009f0000000000000082000000000000009b000000000000009200000000",
            INIT_1B => X"000000a000000000000000a2000000000000008a000000000000009000000000",
            INIT_1C => X"000000dc00000000000000c200000000000000cd00000000000000ac00000000",
            INIT_1D => X"000000e000000000000000d300000000000000d300000000000000de00000000",
            INIT_1E => X"000000db00000000000000e500000000000000e900000000000000e600000000",
            INIT_1F => X"000000d400000000000000e200000000000000df00000000000000cf00000000",
            INIT_20 => X"000000f400000000000000f400000000000000f400000000000000f500000000",
            INIT_21 => X"0000007000000000000000cd00000000000000f000000000000000f500000000",
            INIT_22 => X"0000006d000000000000005b000000000000006d000000000000006200000000",
            INIT_23 => X"0000005c0000000000000064000000000000005c000000000000006500000000",
            INIT_24 => X"0000009a000000000000007c000000000000007d000000000000006800000000",
            INIT_25 => X"000000e300000000000000c900000000000000c200000000000000c200000000",
            INIT_26 => X"000000d300000000000000e300000000000000de00000000000000dc00000000",
            INIT_27 => X"000000e100000000000000e800000000000000dc00000000000000cb00000000",
            INIT_28 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_29 => X"0000007b00000000000000d400000000000000eb00000000000000f600000000",
            INIT_2A => X"00000069000000000000005f000000000000005d000000000000004700000000",
            INIT_2B => X"00000066000000000000006e000000000000006a000000000000006700000000",
            INIT_2C => X"0000005d000000000000005b0000000000000059000000000000005b00000000",
            INIT_2D => X"000000e600000000000000d900000000000000c5000000000000008100000000",
            INIT_2E => X"000000c600000000000000d600000000000000da00000000000000dd00000000",
            INIT_2F => X"000000ed00000000000000e200000000000000c500000000000000b400000000",
            INIT_30 => X"000000f400000000000000f300000000000000f300000000000000f500000000",
            INIT_31 => X"0000009c00000000000000d500000000000000d600000000000000f000000000",
            INIT_32 => X"0000009a00000000000000890000000000000077000000000000004f00000000",
            INIT_33 => X"00000096000000000000009b000000000000008b000000000000009000000000",
            INIT_34 => X"0000007e00000000000000790000000000000080000000000000008e00000000",
            INIT_35 => X"000000e900000000000000e100000000000000a0000000000000007200000000",
            INIT_36 => X"000000ba00000000000000c000000000000000da00000000000000e900000000",
            INIT_37 => X"000000ec00000000000000d400000000000000b000000000000000a500000000",
            INIT_38 => X"000000f700000000000000f300000000000000f300000000000000f400000000",
            INIT_39 => X"0000009600000000000000d300000000000000c100000000000000e200000000",
            INIT_3A => X"000000c800000000000000bc0000000000000098000000000000005100000000",
            INIT_3B => X"00000090000000000000008d00000000000000a500000000000000cd00000000",
            INIT_3C => X"0000008f000000000000008d0000000000000096000000000000008e00000000",
            INIT_3D => X"000000d600000000000000a3000000000000008c00000000000000a700000000",
            INIT_3E => X"000000d200000000000000d300000000000000d100000000000000e000000000",
            INIT_3F => X"000000dc00000000000000af00000000000000ae00000000000000c700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f500000000000000f400000000000000f300000000000000f400000000",
            INIT_41 => X"0000007f00000000000000d800000000000000ca00000000000000e100000000",
            INIT_42 => X"0000008700000000000000840000000000000086000000000000005100000000",
            INIT_43 => X"00000087000000000000007c000000000000009700000000000000b900000000",
            INIT_44 => X"0000008800000000000000960000000000000091000000000000008600000000",
            INIT_45 => X"000000c0000000000000008e000000000000009e00000000000000a400000000",
            INIT_46 => X"000000d700000000000000e700000000000000d800000000000000cf00000000",
            INIT_47 => X"000000c4000000000000009c000000000000009e00000000000000b100000000",
            INIT_48 => X"000000f200000000000000f400000000000000f200000000000000f200000000",
            INIT_49 => X"0000006e00000000000000a800000000000000bd00000000000000e300000000",
            INIT_4A => X"000000760000000000000080000000000000008c000000000000005300000000",
            INIT_4B => X"00000081000000000000007c0000000000000087000000000000009300000000",
            INIT_4C => X"000000860000000000000097000000000000008b000000000000008500000000",
            INIT_4D => X"000000c1000000000000009100000000000000a4000000000000009e00000000",
            INIT_4E => X"000000e600000000000000ef00000000000000ef00000000000000e500000000",
            INIT_4F => X"000000d700000000000000cc00000000000000be00000000000000c100000000",
            INIT_50 => X"000000f400000000000000f300000000000000ef00000000000000e800000000",
            INIT_51 => X"0000005e0000000000000080000000000000008100000000000000da00000000",
            INIT_52 => X"00000070000000000000007a000000000000007a000000000000004f00000000",
            INIT_53 => X"0000007300000000000000730000000000000070000000000000007100000000",
            INIT_54 => X"0000007e000000000000007f0000000000000080000000000000007c00000000",
            INIT_55 => X"000000aa0000000000000099000000000000009e000000000000009000000000",
            INIT_56 => X"000000f400000000000000f600000000000000e300000000000000ce00000000",
            INIT_57 => X"000000f400000000000000f500000000000000f300000000000000f300000000",
            INIT_58 => X"000000f200000000000000f200000000000000e300000000000000cd00000000",
            INIT_59 => X"00000058000000000000009f00000000000000a100000000000000d300000000",
            INIT_5A => X"00000066000000000000005e0000000000000045000000000000003c00000000",
            INIT_5B => X"0000006600000000000000670000000000000061000000000000006200000000",
            INIT_5C => X"00000067000000000000005f0000000000000064000000000000006800000000",
            INIT_5D => X"000000800000000000000089000000000000007f000000000000007100000000",
            INIT_5E => X"000000f300000000000000f800000000000000d7000000000000009900000000",
            INIT_5F => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_60 => X"000000dc00000000000000e400000000000000d500000000000000bc00000000",
            INIT_61 => X"0000006300000000000000ad00000000000000aa00000000000000b400000000",
            INIT_62 => X"00000066000000000000005a0000000000000039000000000000003700000000",
            INIT_63 => X"0000005500000000000000580000000000000067000000000000007200000000",
            INIT_64 => X"00000073000000000000005d0000000000000055000000000000005500000000",
            INIT_65 => X"0000008600000000000000760000000000000065000000000000007000000000",
            INIT_66 => X"000000f400000000000000f500000000000000e100000000000000b000000000",
            INIT_67 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_68 => X"000000b500000000000000ca00000000000000bc00000000000000b800000000",
            INIT_69 => X"00000063000000000000008d0000000000000086000000000000009800000000",
            INIT_6A => X"00000067000000000000006f0000000000000066000000000000006700000000",
            INIT_6B => X"0000005600000000000000600000000000000078000000000000007600000000",
            INIT_6C => X"00000092000000000000007d000000000000006b000000000000005c00000000",
            INIT_6D => X"0000007f000000000000006e000000000000006a000000000000008400000000",
            INIT_6E => X"000000d200000000000000c300000000000000b3000000000000009800000000",
            INIT_6F => X"000000f400000000000000f400000000000000f500000000000000ee00000000",
            INIT_70 => X"0000009800000000000000bd00000000000000c200000000000000b600000000",
            INIT_71 => X"0000007e000000000000007f000000000000007b000000000000009200000000",
            INIT_72 => X"0000005e0000000000000069000000000000005d000000000000007c00000000",
            INIT_73 => X"0000004f0000000000000055000000000000005d000000000000005a00000000",
            INIT_74 => X"0000005500000000000000540000000000000053000000000000004e00000000",
            INIT_75 => X"00000053000000000000004c000000000000004b000000000000005100000000",
            INIT_76 => X"0000008a000000000000008a000000000000007a000000000000006500000000",
            INIT_77 => X"000000f400000000000000f400000000000000f400000000000000bc00000000",
            INIT_78 => X"0000006500000000000000a700000000000000cc00000000000000bd00000000",
            INIT_79 => X"000000ae00000000000000a9000000000000007d000000000000006500000000",
            INIT_7A => X"00000036000000000000004f000000000000004d000000000000006700000000",
            INIT_7B => X"0000003e000000000000003b000000000000002f000000000000002b00000000",
            INIT_7C => X"000000340000000000000039000000000000003e000000000000003b00000000",
            INIT_7D => X"00000040000000000000003d0000000000000030000000000000002f00000000",
            INIT_7E => X"00000061000000000000005a000000000000004a000000000000004600000000",
            INIT_7F => X"000000f400000000000000f600000000000000df000000000000008000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE56;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE57 : if BRAM_NAME = "sampleifmap_layersamples_instance57" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000054000000000000009700000000000000a400000000000000ae00000000",
            INIT_01 => X"0000009200000000000000ac000000000000007c000000000000005200000000",
            INIT_02 => X"0000005a00000000000000570000000000000049000000000000005300000000",
            INIT_03 => X"00000044000000000000004c000000000000004b000000000000006400000000",
            INIT_04 => X"00000017000000000000001a0000000000000017000000000000002100000000",
            INIT_05 => X"000000190000000000000014000000000000002f000000000000003000000000",
            INIT_06 => X"0000006400000000000000560000000000000032000000000000001500000000",
            INIT_07 => X"000000f300000000000000f700000000000000ca000000000000007800000000",
            INIT_08 => X"0000006800000000000000b300000000000000b400000000000000c000000000",
            INIT_09 => X"00000040000000000000008e0000000000000087000000000000006800000000",
            INIT_0A => X"00000078000000000000006c0000000000000057000000000000004100000000",
            INIT_0B => X"00000062000000000000007d0000000000000076000000000000009500000000",
            INIT_0C => X"00000060000000000000006a0000000000000059000000000000004600000000",
            INIT_0D => X"0000006000000000000000590000000000000090000000000000009000000000",
            INIT_0E => X"0000008b00000000000000820000000000000067000000000000005a00000000",
            INIT_0F => X"000000f400000000000000f100000000000000b2000000000000009700000000",
            INIT_10 => X"0000005e00000000000000ab00000000000000bd00000000000000d100000000",
            INIT_11 => X"0000001c00000000000000760000000000000092000000000000006200000000",
            INIT_12 => X"0000004f0000000000000067000000000000005f000000000000003600000000",
            INIT_13 => X"0000005f00000000000000800000000000000064000000000000005300000000",
            INIT_14 => X"0000009e000000000000009b00000000000000aa000000000000009200000000",
            INIT_15 => X"000000a100000000000000a000000000000000a800000000000000ab00000000",
            INIT_16 => X"00000077000000000000009b00000000000000ac000000000000009e00000000",
            INIT_17 => X"000000f700000000000000e20000000000000080000000000000006f00000000",
            INIT_18 => X"0000005b00000000000000b000000000000000c100000000000000d000000000",
            INIT_19 => X"000000280000000000000064000000000000007f000000000000004c00000000",
            INIT_1A => X"0000003900000000000000490000000000000044000000000000003500000000",
            INIT_1B => X"00000059000000000000003d0000000000000035000000000000003200000000",
            INIT_1C => X"0000006200000000000000570000000000000077000000000000009c00000000",
            INIT_1D => X"0000006400000000000000630000000000000068000000000000007100000000",
            INIT_1E => X"0000003f000000000000007a0000000000000098000000000000006000000000",
            INIT_1F => X"000000f800000000000000d60000000000000070000000000000004d00000000",
            INIT_20 => X"0000005f00000000000000be00000000000000c300000000000000ca00000000",
            INIT_21 => X"000000380000000000000053000000000000004e000000000000003300000000",
            INIT_22 => X"00000044000000000000003c0000000000000027000000000000003300000000",
            INIT_23 => X"0000003d000000000000003b0000000000000033000000000000003900000000",
            INIT_24 => X"000000650000000000000066000000000000006e000000000000005f00000000",
            INIT_25 => X"00000060000000000000005c000000000000005f000000000000006300000000",
            INIT_26 => X"000000460000000000000060000000000000006c000000000000006400000000",
            INIT_27 => X"000000f900000000000000d0000000000000006c000000000000004f00000000",
            INIT_28 => X"0000006e00000000000000c000000000000000c000000000000000c200000000",
            INIT_29 => X"0000003f0000000000000049000000000000003e000000000000004c00000000",
            INIT_2A => X"000000300000000000000028000000000000001d000000000000002e00000000",
            INIT_2B => X"0000003b00000000000000530000000000000048000000000000004100000000",
            INIT_2C => X"00000043000000000000004d0000000000000043000000000000003000000000",
            INIT_2D => X"00000058000000000000003b0000000000000040000000000000003c00000000",
            INIT_2E => X"00000069000000000000004e0000000000000036000000000000005200000000",
            INIT_2F => X"000000f900000000000000c90000000000000065000000000000006b00000000",
            INIT_30 => X"0000006100000000000000bb00000000000000be00000000000000c300000000",
            INIT_31 => X"0000004300000000000000410000000000000063000000000000005500000000",
            INIT_32 => X"0000002000000000000000230000000000000026000000000000003a00000000",
            INIT_33 => X"0000004c000000000000008d0000000000000060000000000000004800000000",
            INIT_34 => X"00000071000000000000008c000000000000004f000000000000001900000000",
            INIT_35 => X"000000920000000000000061000000000000006d000000000000005e00000000",
            INIT_36 => X"0000008a0000000000000045000000000000003a00000000000000ab00000000",
            INIT_37 => X"000000f400000000000000c00000000000000053000000000000007400000000",
            INIT_38 => X"0000005200000000000000b000000000000000b700000000000000bd00000000",
            INIT_39 => X"0000005e00000000000000590000000000000063000000000000002c00000000",
            INIT_3A => X"0000002100000000000000240000000000000030000000000000005a00000000",
            INIT_3B => X"000000340000000000000055000000000000002f000000000000002600000000",
            INIT_3C => X"0000007b0000000000000091000000000000004a000000000000001c00000000",
            INIT_3D => X"0000009700000000000000710000000000000086000000000000007700000000",
            INIT_3E => X"0000004700000000000000320000000000000033000000000000009c00000000",
            INIT_3F => X"000000ee00000000000000c00000000000000047000000000000003b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004800000000000000a300000000000000ad00000000000000ae00000000",
            INIT_41 => X"0000008b00000000000000650000000000000036000000000000002200000000",
            INIT_42 => X"0000001e0000000000000028000000000000003a000000000000006600000000",
            INIT_43 => X"0000001e000000000000001a0000000000000019000000000000001a00000000",
            INIT_44 => X"0000005600000000000000350000000000000026000000000000002500000000",
            INIT_45 => X"0000007200000000000000760000000000000075000000000000006800000000",
            INIT_46 => X"0000002e0000000000000030000000000000002b000000000000003e00000000",
            INIT_47 => X"000000df00000000000000b8000000000000004b000000000000002f00000000",
            INIT_48 => X"00000078000000000000009e00000000000000a000000000000000a200000000",
            INIT_49 => X"0000008800000000000000670000000000000059000000000000005700000000",
            INIT_4A => X"0000002200000000000000340000000000000048000000000000005c00000000",
            INIT_4B => X"0000001d000000000000001b000000000000001b000000000000001c00000000",
            INIT_4C => X"000000af000000000000003d0000000000000015000000000000002000000000",
            INIT_4D => X"000000b400000000000000b100000000000000ca00000000000000cf00000000",
            INIT_4E => X"0000002c00000000000000280000000000000022000000000000005400000000",
            INIT_4F => X"000000d100000000000000ab0000000000000057000000000000003e00000000",
            INIT_50 => X"000000b000000000000000a8000000000000009c000000000000009c00000000",
            INIT_51 => X"0000008800000000000000660000000000000070000000000000009300000000",
            INIT_52 => X"0000002d000000000000004b0000000000000051000000000000005600000000",
            INIT_53 => X"0000001a00000000000000170000000000000016000000000000001600000000",
            INIT_54 => X"000000a400000000000000450000000000000022000000000000002300000000",
            INIT_55 => X"000000a500000000000000a900000000000000b100000000000000b900000000",
            INIT_56 => X"0000002d000000000000001a0000000000000019000000000000004e00000000",
            INIT_57 => X"000000cc00000000000000a7000000000000005c000000000000004b00000000",
            INIT_58 => X"000000a100000000000000ad00000000000000a7000000000000009500000000",
            INIT_59 => X"0000008e00000000000000630000000000000071000000000000008d00000000",
            INIT_5A => X"00000033000000000000004f0000000000000053000000000000005300000000",
            INIT_5B => X"00000022000000000000001f000000000000001c000000000000001d00000000",
            INIT_5C => X"0000006100000000000000510000000000000048000000000000003200000000",
            INIT_5D => X"00000085000000000000008a0000000000000074000000000000006600000000",
            INIT_5E => X"00000032000000000000001d000000000000001b000000000000003700000000",
            INIT_5F => X"000000c600000000000000a40000000000000059000000000000004c00000000",
            INIT_60 => X"00000090000000000000009b00000000000000a600000000000000a400000000",
            INIT_61 => X"0000006c00000000000000630000000000000082000000000000008b00000000",
            INIT_62 => X"0000003800000000000000480000000000000050000000000000004c00000000",
            INIT_63 => X"0000002900000000000000270000000000000024000000000000002600000000",
            INIT_64 => X"00000048000000000000003d0000000000000033000000000000002d00000000",
            INIT_65 => X"00000083000000000000007c0000000000000067000000000000005400000000",
            INIT_66 => X"000000320000000000000021000000000000001a000000000000003100000000",
            INIT_67 => X"000000c300000000000000a90000000000000059000000000000004500000000",
            INIT_68 => X"0000008d0000000000000092000000000000009400000000000000a000000000",
            INIT_69 => X"0000004900000000000000660000000000000082000000000000008700000000",
            INIT_6A => X"000000380000000000000042000000000000004d000000000000004500000000",
            INIT_6B => X"0000002d000000000000002b0000000000000028000000000000002f00000000",
            INIT_6C => X"0000003d00000000000000360000000000000030000000000000002e00000000",
            INIT_6D => X"0000006a000000000000005e0000000000000054000000000000004600000000",
            INIT_6E => X"00000030000000000000001f000000000000001a000000000000004000000000",
            INIT_6F => X"000000ba00000000000000af0000000000000062000000000000003d00000000",
            INIT_70 => X"0000008c000000000000008e000000000000008d000000000000009300000000",
            INIT_71 => X"000000390000000000000068000000000000008b000000000000008f00000000",
            INIT_72 => X"00000034000000000000003f000000000000004a000000000000004000000000",
            INIT_73 => X"0000003600000000000000330000000000000031000000000000003700000000",
            INIT_74 => X"00000042000000000000003d0000000000000036000000000000003600000000",
            INIT_75 => X"000000570000000000000051000000000000004a000000000000004400000000",
            INIT_76 => X"0000003400000000000000230000000000000021000000000000004800000000",
            INIT_77 => X"000000b500000000000000b60000000000000084000000000000004800000000",
            INIT_78 => X"000000a300000000000000a10000000000000096000000000000009200000000",
            INIT_79 => X"0000003a000000000000007c0000000000000091000000000000009d00000000",
            INIT_7A => X"0000004100000000000000390000000000000038000000000000003700000000",
            INIT_7B => X"0000004500000000000000460000000000000042000000000000004300000000",
            INIT_7C => X"0000005f00000000000000570000000000000048000000000000004300000000",
            INIT_7D => X"0000005e0000000000000060000000000000005f000000000000005c00000000",
            INIT_7E => X"00000046000000000000003e0000000000000044000000000000005100000000",
            INIT_7F => X"000000b900000000000000b600000000000000a3000000000000007600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE57;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE58 : if BRAM_NAME = "sampleifmap_layersamples_instance58" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b600000000000000bf00000000000000ca00000000000000d100000000",
            INIT_01 => X"000000af00000000000000c600000000000000d100000000000000d100000000",
            INIT_02 => X"000000a0000000000000009d00000000000000a500000000000000ab00000000",
            INIT_03 => X"0000008f000000000000008d000000000000009a000000000000009500000000",
            INIT_04 => X"000000db00000000000000d600000000000000bc00000000000000a400000000",
            INIT_05 => X"000000d600000000000000d900000000000000ca00000000000000d100000000",
            INIT_06 => X"000000ad00000000000000a100000000000000b100000000000000d000000000",
            INIT_07 => X"000000950000000000000095000000000000009d00000000000000b700000000",
            INIT_08 => X"000000cd00000000000000d200000000000000d400000000000000d400000000",
            INIT_09 => X"000000a300000000000000c800000000000000db00000000000000cf00000000",
            INIT_0A => X"000000b600000000000000b800000000000000b600000000000000a500000000",
            INIT_0B => X"000000d700000000000000cd00000000000000c900000000000000c200000000",
            INIT_0C => X"000000e400000000000000e300000000000000e300000000000000df00000000",
            INIT_0D => X"000000d700000000000000d300000000000000d400000000000000dd00000000",
            INIT_0E => X"000000bb00000000000000c300000000000000cd00000000000000df00000000",
            INIT_0F => X"000000ba00000000000000ad00000000000000aa00000000000000c600000000",
            INIT_10 => X"000000e200000000000000e300000000000000e500000000000000e600000000",
            INIT_11 => X"000000a400000000000000d300000000000000ec00000000000000e300000000",
            INIT_12 => X"000000b800000000000000b700000000000000ad000000000000009f00000000",
            INIT_13 => X"000000e000000000000000cf00000000000000bf00000000000000bc00000000",
            INIT_14 => X"000000d600000000000000e000000000000000e500000000000000db00000000",
            INIT_15 => X"000000d300000000000000c800000000000000d000000000000000d600000000",
            INIT_16 => X"000000c500000000000000db00000000000000e000000000000000de00000000",
            INIT_17 => X"000000c600000000000000c500000000000000bc00000000000000b900000000",
            INIT_18 => X"000000f100000000000000f400000000000000f400000000000000f500000000",
            INIT_19 => X"000000af00000000000000e300000000000000f100000000000000f200000000",
            INIT_1A => X"000000bb00000000000000a100000000000000b000000000000000a800000000",
            INIT_1B => X"000000b600000000000000b800000000000000a000000000000000ae00000000",
            INIT_1C => X"000000ca00000000000000d000000000000000d500000000000000b900000000",
            INIT_1D => X"000000d400000000000000c400000000000000ba00000000000000b900000000",
            INIT_1E => X"000000bb00000000000000d500000000000000dc00000000000000d700000000",
            INIT_1F => X"000000c800000000000000d400000000000000c500000000000000a900000000",
            INIT_20 => X"000000f400000000000000f400000000000000f300000000000000f500000000",
            INIT_21 => X"0000008400000000000000cd00000000000000f100000000000000f500000000",
            INIT_22 => X"000000a7000000000000008a00000000000000a1000000000000008b00000000",
            INIT_23 => X"0000008d000000000000009b000000000000008b000000000000009f00000000",
            INIT_24 => X"000000a4000000000000009900000000000000a6000000000000008e00000000",
            INIT_25 => X"000000e000000000000000c400000000000000a900000000000000a900000000",
            INIT_26 => X"000000b100000000000000d400000000000000d100000000000000d100000000",
            INIT_27 => X"000000d200000000000000cc00000000000000b800000000000000a000000000",
            INIT_28 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_29 => X"0000008100000000000000d700000000000000ee00000000000000f600000000",
            INIT_2A => X"000000aa00000000000000a0000000000000009c000000000000007100000000",
            INIT_2B => X"000000a700000000000000b100000000000000aa00000000000000aa00000000",
            INIT_2C => X"0000008f0000000000000098000000000000009d000000000000009d00000000",
            INIT_2D => X"000000e400000000000000cd00000000000000b3000000000000009400000000",
            INIT_2E => X"000000aa00000000000000c100000000000000ce00000000000000da00000000",
            INIT_2F => X"000000df00000000000000c000000000000000a0000000000000009300000000",
            INIT_30 => X"000000f400000000000000f300000000000000f300000000000000f500000000",
            INIT_31 => X"000000b400000000000000dd00000000000000dd00000000000000f100000000",
            INIT_32 => X"000000cf00000000000000c400000000000000b4000000000000008300000000",
            INIT_33 => X"000000d300000000000000d900000000000000cb00000000000000c800000000",
            INIT_34 => X"000000bf00000000000000c000000000000000c300000000000000cc00000000",
            INIT_35 => X"000000e100000000000000cd00000000000000a600000000000000a300000000",
            INIT_36 => X"000000a900000000000000b100000000000000d500000000000000e300000000",
            INIT_37 => X"000000da00000000000000b20000000000000092000000000000009100000000",
            INIT_38 => X"000000f700000000000000f200000000000000f200000000000000f400000000",
            INIT_39 => X"000000c000000000000000d900000000000000ca00000000000000e600000000",
            INIT_3A => X"000000e800000000000000e000000000000000c2000000000000008600000000",
            INIT_3B => X"000000d100000000000000ce00000000000000d700000000000000ea00000000",
            INIT_3C => X"000000cf00000000000000ca00000000000000d000000000000000cf00000000",
            INIT_3D => X"000000cc000000000000009a00000000000000b400000000000000e000000000",
            INIT_3E => X"000000bc00000000000000c400000000000000c900000000000000dc00000000",
            INIT_3F => X"000000c7000000000000009a000000000000009200000000000000ab00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f500000000000000f300000000000000f300000000000000f500000000",
            INIT_41 => X"000000ae00000000000000df00000000000000d100000000000000e300000000",
            INIT_42 => X"000000c100000000000000c100000000000000ba000000000000008700000000",
            INIT_43 => X"000000c900000000000000c100000000000000cc00000000000000dd00000000",
            INIT_44 => X"000000c600000000000000cd00000000000000cd00000000000000ca00000000",
            INIT_45 => X"000000bc00000000000000a300000000000000d000000000000000dc00000000",
            INIT_46 => X"000000cb00000000000000df00000000000000d100000000000000cb00000000",
            INIT_47 => X"000000b20000000000000094000000000000008b00000000000000a100000000",
            INIT_48 => X"000000f200000000000000f300000000000000f100000000000000f200000000",
            INIT_49 => X"000000a400000000000000c200000000000000cd00000000000000e500000000",
            INIT_4A => X"000000b800000000000000bd00000000000000c1000000000000008c00000000",
            INIT_4B => X"000000c400000000000000c000000000000000c400000000000000ca00000000",
            INIT_4C => X"000000c600000000000000d000000000000000ca00000000000000c700000000",
            INIT_4D => X"000000c800000000000000bc00000000000000e000000000000000d700000000",
            INIT_4E => X"000000e300000000000000ed00000000000000ee00000000000000e600000000",
            INIT_4F => X"000000d300000000000000ca00000000000000ba00000000000000bc00000000",
            INIT_50 => X"000000f400000000000000f300000000000000ee00000000000000ea00000000",
            INIT_51 => X"0000009c00000000000000a900000000000000a000000000000000df00000000",
            INIT_52 => X"000000ac00000000000000b300000000000000b1000000000000008600000000",
            INIT_53 => X"000000b700000000000000b400000000000000ae00000000000000ae00000000",
            INIT_54 => X"000000be00000000000000bc00000000000000be00000000000000bb00000000",
            INIT_55 => X"000000c400000000000000d000000000000000dc00000000000000cd00000000",
            INIT_56 => X"000000f400000000000000f600000000000000e600000000000000d900000000",
            INIT_57 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_58 => X"000000f200000000000000f200000000000000e600000000000000d300000000",
            INIT_59 => X"0000009700000000000000be00000000000000b600000000000000d800000000",
            INIT_5A => X"000000a00000000000000093000000000000006e000000000000006a00000000",
            INIT_5B => X"000000aa00000000000000a6000000000000009f000000000000009e00000000",
            INIT_5C => X"000000a6000000000000009e00000000000000a300000000000000a900000000",
            INIT_5D => X"000000af00000000000000c600000000000000bd00000000000000ad00000000",
            INIT_5E => X"000000f300000000000000f800000000000000e000000000000000b700000000",
            INIT_5F => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_60 => X"000000e100000000000000e900000000000000da00000000000000c400000000",
            INIT_61 => X"0000009f00000000000000c300000000000000b400000000000000bd00000000",
            INIT_62 => X"000000a0000000000000008d000000000000005c000000000000005d00000000",
            INIT_63 => X"0000008c000000000000008f00000000000000a800000000000000ba00000000",
            INIT_64 => X"000000a700000000000000920000000000000089000000000000008b00000000",
            INIT_65 => X"00000096000000000000008f0000000000000083000000000000009800000000",
            INIT_66 => X"000000f400000000000000f300000000000000e300000000000000bc00000000",
            INIT_67 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_68 => X"000000c100000000000000d300000000000000c700000000000000c300000000",
            INIT_69 => X"0000008900000000000000a2000000000000009500000000000000a400000000",
            INIT_6A => X"000000a600000000000000b200000000000000aa000000000000009600000000",
            INIT_6B => X"0000009200000000000000a600000000000000cd00000000000000bd00000000",
            INIT_6C => X"000000d300000000000000c000000000000000ac000000000000009900000000",
            INIT_6D => X"0000008a0000000000000080000000000000008000000000000000af00000000",
            INIT_6E => X"000000d300000000000000bf00000000000000b100000000000000a000000000",
            INIT_6F => X"000000f300000000000000f300000000000000f500000000000000ef00000000",
            INIT_70 => X"000000a200000000000000c800000000000000cf00000000000000c200000000",
            INIT_71 => X"00000089000000000000008e0000000000000088000000000000009c00000000",
            INIT_72 => X"0000009f00000000000000b100000000000000b200000000000000a200000000",
            INIT_73 => X"0000008b000000000000009500000000000000a3000000000000009600000000",
            INIT_74 => X"0000009300000000000000920000000000000092000000000000008d00000000",
            INIT_75 => X"00000085000000000000007f000000000000007c000000000000008600000000",
            INIT_76 => X"000000a600000000000000ad00000000000000a3000000000000009500000000",
            INIT_77 => X"000000f400000000000000f300000000000000f500000000000000cc00000000",
            INIT_78 => X"0000006e00000000000000ad00000000000000d000000000000000c300000000",
            INIT_79 => X"000000b900000000000000b4000000000000008b000000000000007100000000",
            INIT_7A => X"00000057000000000000007f000000000000009a000000000000008500000000",
            INIT_7B => X"0000005f0000000000000059000000000000004c000000000000004900000000",
            INIT_7C => X"00000058000000000000005e0000000000000060000000000000005c00000000",
            INIT_7D => X"0000006700000000000000630000000000000056000000000000005600000000",
            INIT_7E => X"0000009b000000000000008f0000000000000074000000000000006d00000000",
            INIT_7F => X"000000f500000000000000f500000000000000e800000000000000af00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE58;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE59 : if BRAM_NAME = "sampleifmap_layersamples_instance59" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000006500000000000000a100000000000000aa00000000000000b700000000",
            INIT_01 => X"000000a100000000000000b50000000000000088000000000000006000000000",
            INIT_02 => X"0000008700000000000000810000000000000084000000000000008000000000",
            INIT_03 => X"0000006a000000000000007d000000000000007d000000000000008c00000000",
            INIT_04 => X"00000027000000000000002c000000000000002b000000000000003500000000",
            INIT_05 => X"0000002800000000000000230000000000000047000000000000004d00000000",
            INIT_06 => X"0000009700000000000000910000000000000050000000000000002000000000",
            INIT_07 => X"000000f300000000000000f600000000000000db00000000000000a700000000",
            INIT_08 => X"0000007c00000000000000c200000000000000c100000000000000ca00000000",
            INIT_09 => X"0000004900000000000000990000000000000092000000000000007800000000",
            INIT_0A => X"0000009400000000000000830000000000000087000000000000006900000000",
            INIT_0B => X"0000008300000000000000a9000000000000009f00000000000000b800000000",
            INIT_0C => X"0000007a00000000000000840000000000000076000000000000006600000000",
            INIT_0D => X"00000073000000000000006f00000000000000aa00000000000000af00000000",
            INIT_0E => X"000000b500000000000000b20000000000000091000000000000006f00000000",
            INIT_0F => X"000000f400000000000000f200000000000000c500000000000000bb00000000",
            INIT_10 => X"0000007200000000000000b800000000000000c800000000000000d800000000",
            INIT_11 => X"000000240000000000000082000000000000009d000000000000007300000000",
            INIT_12 => X"0000006300000000000000810000000000000095000000000000004f00000000",
            INIT_13 => X"00000084000000000000009d0000000000000081000000000000006f00000000",
            INIT_14 => X"000000b900000000000000b700000000000000c100000000000000b100000000",
            INIT_15 => X"000000bd00000000000000ba00000000000000c100000000000000c800000000",
            INIT_16 => X"0000009700000000000000b600000000000000c700000000000000b500000000",
            INIT_17 => X"000000f600000000000000e800000000000000a2000000000000009400000000",
            INIT_18 => X"0000007100000000000000bb00000000000000cc00000000000000d900000000",
            INIT_19 => X"0000003d0000000000000071000000000000008b000000000000006000000000",
            INIT_1A => X"0000005d00000000000000730000000000000070000000000000004e00000000",
            INIT_1B => X"0000007d000000000000005e0000000000000053000000000000005500000000",
            INIT_1C => X"0000008a000000000000007f000000000000009f00000000000000bf00000000",
            INIT_1D => X"0000008f000000000000008c000000000000009500000000000000a000000000",
            INIT_1E => X"00000063000000000000009f00000000000000bd000000000000008a00000000",
            INIT_1F => X"000000f700000000000000e2000000000000009a000000000000007300000000",
            INIT_20 => X"0000007500000000000000c700000000000000d000000000000000d500000000",
            INIT_21 => X"000000540000000000000063000000000000005c000000000000004900000000",
            INIT_22 => X"0000006900000000000000610000000000000041000000000000004b00000000",
            INIT_23 => X"0000005f00000000000000670000000000000057000000000000005f00000000",
            INIT_24 => X"00000097000000000000009900000000000000a2000000000000008600000000",
            INIT_25 => X"0000008f00000000000000890000000000000090000000000000009600000000",
            INIT_26 => X"0000006f000000000000008f0000000000000099000000000000009300000000",
            INIT_27 => X"000000f700000000000000de0000000000000092000000000000007300000000",
            INIT_28 => X"0000008300000000000000cc00000000000000ce00000000000000cc00000000",
            INIT_29 => X"0000005a000000000000005c0000000000000051000000000000006500000000",
            INIT_2A => X"000000450000000000000039000000000000002d000000000000004600000000",
            INIT_2B => X"00000057000000000000007d000000000000006f000000000000006200000000",
            INIT_2C => X"0000006700000000000000700000000000000066000000000000004a00000000",
            INIT_2D => X"0000007d000000000000005e0000000000000065000000000000006200000000",
            INIT_2E => X"0000009500000000000000710000000000000052000000000000007300000000",
            INIT_2F => X"000000f800000000000000d40000000000000089000000000000009a00000000",
            INIT_30 => X"0000007500000000000000ce00000000000000d000000000000000d100000000",
            INIT_31 => X"0000005e0000000000000056000000000000007a000000000000006900000000",
            INIT_32 => X"0000002f00000000000000330000000000000036000000000000005600000000",
            INIT_33 => X"0000006300000000000000ad0000000000000083000000000000006600000000",
            INIT_34 => X"00000082000000000000009e0000000000000064000000000000002d00000000",
            INIT_35 => X"000000ab000000000000007c000000000000008a000000000000007900000000",
            INIT_36 => X"000000ab000000000000005f000000000000004b00000000000000bb00000000",
            INIT_37 => X"000000fa00000000000000cf0000000000000075000000000000009800000000",
            INIT_38 => X"0000006800000000000000cc00000000000000d600000000000000dd00000000",
            INIT_39 => X"0000008000000000000000720000000000000074000000000000003b00000000",
            INIT_3A => X"0000003000000000000000340000000000000041000000000000007c00000000",
            INIT_3B => X"0000004b000000000000006c0000000000000046000000000000003800000000",
            INIT_3C => X"0000008f00000000000000a6000000000000005f000000000000003000000000",
            INIT_3D => X"000000af000000000000008f00000000000000a7000000000000009100000000",
            INIT_3E => X"000000620000000000000048000000000000004a00000000000000af00000000",
            INIT_3F => X"000000fb00000000000000d60000000000000068000000000000005400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006300000000000000c900000000000000d400000000000000d700000000",
            INIT_41 => X"000000b000000000000000800000000000000044000000000000002f00000000",
            INIT_42 => X"0000002d00000000000000380000000000000050000000000000008700000000",
            INIT_43 => X"0000002f000000000000002b0000000000000027000000000000002800000000",
            INIT_44 => X"0000006e0000000000000050000000000000003c000000000000003700000000",
            INIT_45 => X"0000008b00000000000000900000000000000093000000000000007d00000000",
            INIT_46 => X"0000004300000000000000460000000000000043000000000000005c00000000",
            INIT_47 => X"000000fb00000000000000d9000000000000006d000000000000004500000000",
            INIT_48 => X"0000009d00000000000000cb00000000000000cf00000000000000cf00000000",
            INIT_49 => X"000000aa00000000000000850000000000000075000000000000007300000000",
            INIT_4A => X"0000003000000000000000480000000000000065000000000000007e00000000",
            INIT_4B => X"0000002d00000000000000290000000000000029000000000000002800000000",
            INIT_4C => X"000000c000000000000000530000000000000027000000000000003200000000",
            INIT_4D => X"000000c900000000000000c700000000000000dc00000000000000da00000000",
            INIT_4E => X"0000003f00000000000000380000000000000034000000000000006b00000000",
            INIT_4F => X"000000f700000000000000d2000000000000007e000000000000005a00000000",
            INIT_50 => X"000000d800000000000000ce00000000000000c000000000000000bc00000000",
            INIT_51 => X"000000a10000000000000086000000000000009a00000000000000bf00000000",
            INIT_52 => X"0000003e00000000000000680000000000000073000000000000007900000000",
            INIT_53 => X"0000002900000000000000230000000000000022000000000000002100000000",
            INIT_54 => X"000000b300000000000000550000000000000031000000000000003300000000",
            INIT_55 => X"000000bb00000000000000be00000000000000c000000000000000c700000000",
            INIT_56 => X"0000004200000000000000260000000000000027000000000000006000000000",
            INIT_57 => X"000000f500000000000000d10000000000000085000000000000006f00000000",
            INIT_58 => X"000000c600000000000000cd00000000000000c600000000000000bf00000000",
            INIT_59 => X"000000a00000000000000084000000000000009e00000000000000b500000000",
            INIT_5A => X"00000046000000000000006f0000000000000076000000000000007200000000",
            INIT_5B => X"00000031000000000000002c0000000000000026000000000000002700000000",
            INIT_5C => X"0000007e0000000000000069000000000000005d000000000000004400000000",
            INIT_5D => X"000000a600000000000000ad0000000000000096000000000000008700000000",
            INIT_5E => X"00000047000000000000002a0000000000000028000000000000004800000000",
            INIT_5F => X"000000f200000000000000cf0000000000000082000000000000007100000000",
            INIT_60 => X"000000b800000000000000c600000000000000d100000000000000ce00000000",
            INIT_61 => X"00000085000000000000008200000000000000a300000000000000ab00000000",
            INIT_62 => X"0000004d0000000000000068000000000000006f000000000000006b00000000",
            INIT_63 => X"000000390000000000000035000000000000002f000000000000003200000000",
            INIT_64 => X"0000006800000000000000570000000000000048000000000000003f00000000",
            INIT_65 => X"000000b000000000000000a80000000000000091000000000000007800000000",
            INIT_66 => X"0000004700000000000000300000000000000028000000000000004500000000",
            INIT_67 => X"000000ee00000000000000d4000000000000007e000000000000006600000000",
            INIT_68 => X"000000bd00000000000000c200000000000000c200000000000000c700000000",
            INIT_69 => X"00000065000000000000008600000000000000a600000000000000b200000000",
            INIT_6A => X"0000004f00000000000000600000000000000069000000000000006300000000",
            INIT_6B => X"0000003e000000000000003b0000000000000036000000000000003e00000000",
            INIT_6C => X"00000057000000000000004e0000000000000045000000000000004100000000",
            INIT_6D => X"0000008f00000000000000810000000000000074000000000000006400000000",
            INIT_6E => X"00000047000000000000002c0000000000000027000000000000005700000000",
            INIT_6F => X"000000e800000000000000df0000000000000085000000000000005900000000",
            INIT_70 => X"000000bc00000000000000be00000000000000bc00000000000000c100000000",
            INIT_71 => X"00000050000000000000009000000000000000bc00000000000000bd00000000",
            INIT_72 => X"0000004600000000000000580000000000000063000000000000005a00000000",
            INIT_73 => X"0000004e000000000000004a0000000000000045000000000000004900000000",
            INIT_74 => X"0000005d0000000000000056000000000000004e000000000000004e00000000",
            INIT_75 => X"00000072000000000000006d0000000000000066000000000000006100000000",
            INIT_76 => X"0000004a00000000000000300000000000000030000000000000005e00000000",
            INIT_77 => X"000000e700000000000000e800000000000000ad000000000000006400000000",
            INIT_78 => X"000000cd00000000000000d000000000000000c700000000000000c400000000",
            INIT_79 => X"0000005500000000000000a500000000000000bb00000000000000c800000000",
            INIT_7A => X"00000054000000000000004e000000000000004c000000000000004c00000000",
            INIT_7B => X"0000006300000000000000620000000000000059000000000000005400000000",
            INIT_7C => X"0000007c00000000000000720000000000000063000000000000005e00000000",
            INIT_7D => X"0000007f00000000000000800000000000000081000000000000007d00000000",
            INIT_7E => X"000000600000000000000054000000000000005b000000000000007000000000",
            INIT_7F => X"000000df00000000000000e100000000000000cc000000000000009400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE59;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE0 : if BRAM_NAME = "samplegold_layersamples_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000200000000000000000000000000000000000000000000000500000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000005400000000",
            INIT_06 => X"0000000200000000000000000000000000000002000000000000001b00000000",
            INIT_07 => X"0000000400000000000000000000000000000000000000000000000500000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000004a00000000000000070000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000750000000000000000000000000000001c00000000",
            INIT_0C => X"0000000d000000000000000c0000000000000001000000000000000900000000",
            INIT_0D => X"0000000000000000000000310000000000000000000000000000000000000000",
            INIT_0E => X"0000003600000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000002800000000000000000000000000000054000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000003400000000",
            INIT_11 => X"0000000000000000000000000000000000000058000000000000000000000000",
            INIT_12 => X"0000000000000000000000060000000000000000000000000000000a00000000",
            INIT_13 => X"0000004200000000000000000000000000000000000000000000001f00000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"000000070000000000000000000000000000000000000000000000d900000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000004d00000000000000440000000000000000000000000000000000000000",
            INIT_18 => X"000000a800000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000001b00000000000000040000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000510000000000000016000000000000000000000000",
            INIT_1C => X"0000000000000000000000620000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_1E => X"0000003800000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000120000000000000000000000000000001700000000",
            INIT_21 => X"000000000000000000000012000000000000001d000000000000000600000000",
            INIT_22 => X"0000000000000000000000470000000000000000000000000000000000000000",
            INIT_23 => X"00000000000000000000000e000000000000001a000000000000000000000000",
            INIT_24 => X"0000003400000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000610000000000000000000000000000003700000000",
            INIT_26 => X"00000000000000000000000000000000000000cb000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_28 => X"0000000500000000000000100000000000000024000000000000001700000000",
            INIT_29 => X"00000000000000000000000e000000000000001d000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000009200000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_2D => X"000000000000000000000038000000000000001f000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000d00000000000000090000000000000004000000000000000000000000",
            INIT_30 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_31 => X"000000000000000000000000000000000000004f000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000002900000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000500000000000000080000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000380000000000000000000000000000000000000000",
            INIT_38 => X"000000ab00000000000000ab00000000000000a4000000000000000000000000",
            INIT_39 => X"000000ae00000000000000ac00000000000000a800000000000000ac00000000",
            INIT_3A => X"00000083000000000000009500000000000000a300000000000000ab00000000",
            INIT_3B => X"0000007a000000000000008a0000000000000093000000000000008b00000000",
            INIT_3C => X"000000af00000000000000b000000000000000ab00000000000000a400000000",
            INIT_3D => X"0000009e00000000000000b3000000000000011100000000000000b700000000",
            INIT_3E => X"0000007400000000000000940000000000000095000000000000007000000000",
            INIT_3F => X"0000007800000000000000860000000000000084000000000000006f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ae00000000000000ac00000000000000ad000000000000009a00000000",
            INIT_41 => X"00000054000000000000005e000000000000008e00000000000000ee00000000",
            INIT_42 => X"0000007400000000000000ae00000000000000cd00000000000000e400000000",
            INIT_43 => X"000000aa000000000000006b0000000000000093000000000000005300000000",
            INIT_44 => X"000000b500000000000000ae00000000000000b900000000000000b400000000",
            INIT_45 => X"000000df000000000000007c000000000000007a00000000000000cc00000000",
            INIT_46 => X"000000280000000000000067000000000000009200000000000000d100000000",
            INIT_47 => X"000000bf000000000000013100000000000000e0000000000000008500000000",
            INIT_48 => X"000000f20000000000000123000000000000017d00000000000000fc00000000",
            INIT_49 => X"0000010800000000000000bf000000000000005c000000000000008800000000",
            INIT_4A => X"00000039000000000000004c0000000000000089000000000000008f00000000",
            INIT_4B => X"0000009500000000000000d0000000000000015f00000000000000f400000000",
            INIT_4C => X"000000bc000000000000012e000000000000011f000000000000015c00000000",
            INIT_4D => X"0000008c000000000000011d000000000000012b000000000000006600000000",
            INIT_4E => X"0000010000000000000000480000000000000080000000000000009b00000000",
            INIT_4F => X"000000ee000000000000008000000000000000bb000000000000014400000000",
            INIT_50 => X"0000009100000000000000f70000000000000167000000000000014100000000",
            INIT_51 => X"0000008c00000000000000920000000000000100000000000000015600000000",
            INIT_52 => X"000001610000000000000134000000000000008500000000000000ae00000000",
            INIT_53 => X"0000018300000000000000cd00000000000000be00000000000000c400000000",
            INIT_54 => X"00000123000000000000009200000000000000d8000000000000010f00000000",
            INIT_55 => X"000000ad0000000000000096000000000000009000000000000000f800000000",
            INIT_56 => X"000000c1000000000000018a000000000000016d000000000000009300000000",
            INIT_57 => X"000000bf00000000000000d200000000000000b4000000000000010b00000000",
            INIT_58 => X"000000ad00000000000000c700000000000000c900000000000000b800000000",
            INIT_59 => X"000000ad000000000000009e0000000000000059000000000000005600000000",
            INIT_5A => X"0000012800000000000000ef0000000000000184000000000000018200000000",
            INIT_5B => X"0000012b00000000000000f9000000000000009100000000000000cf00000000",
            INIT_5C => X"000000290000000000000057000000000000009c00000000000000b100000000",
            INIT_5D => X"0000018f00000000000000b300000000000000ce000000000000007d00000000",
            INIT_5E => X"0000019500000000000001b000000000000000fa000000000000017a00000000",
            INIT_5F => X"000000ba000000000000014c000000000000014700000000000000fd00000000",
            INIT_60 => X"000000a7000000000000007e0000000000000061000000000000007000000000",
            INIT_61 => X"00000175000000000000012500000000000000a900000000000000cd00000000",
            INIT_62 => X"000000ae00000000000001770000000000000225000000000000014800000000",
            INIT_63 => X"0000008b000000000000008d00000000000000a900000000000000b200000000",
            INIT_64 => X"000000c900000000000000bb00000000000000ab000000000000009c00000000",
            INIT_65 => X"0000017900000000000000fc00000000000000b600000000000000b900000000",
            INIT_66 => X"0000009b00000000000000a600000000000000ba00000000000001e100000000",
            INIT_67 => X"000000b5000000000000009a0000000000000093000000000000009600000000",
            INIT_68 => X"000000f600000000000000cd00000000000000ce00000000000000c900000000",
            INIT_69 => X"0000016b000000000000013400000000000000ad00000000000000b900000000",
            INIT_6A => X"0000009700000000000000a800000000000000b900000000000000a500000000",
            INIT_6B => X"000000c100000000000000b900000000000000af000000000000009d00000000",
            INIT_6C => X"000000bd00000000000000d200000000000000e000000000000000b900000000",
            INIT_6D => X"0000008100000000000000ce00000000000000b200000000000000b100000000",
            INIT_6E => X"000000bc00000000000000a800000000000000a3000000000000009200000000",
            INIT_6F => X"0000010300000000000000b200000000000000b000000000000000cf00000000",
            INIT_70 => X"000000000000000000000000000000000000009c000000000000010e00000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000033000000000000000000000000",
            INIT_7A => X"00000000000000000000000a0000000000000023000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000090000000000000000000000000000004700000000",
            INIT_7F => X"0000001e00000000000000000000000000000013000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE0;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE1 : if BRAM_NAME = "samplegold_layersamples_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000050000000000000012000000000000000000000000",
            INIT_01 => X"0000002700000000000000000000000000000000000000000000000600000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_03 => X"0000000000000000000000470000000000000011000000000000000000000000",
            INIT_04 => X"0000000a000000000000003a000000000000009c000000000000000400000000",
            INIT_05 => X"0000001200000000000000620000000000000000000000000000000000000000",
            INIT_06 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_07 => X"00000000000000000000000c000000000000002c000000000000000800000000",
            INIT_08 => X"00000000000000000000003f0000000000000038000000000000004800000000",
            INIT_09 => X"0000000000000000000000050000000000000073000000000000000000000000",
            INIT_0A => X"0000001f00000000000000000000000000000004000000000000000000000000",
            INIT_0B => X"0000001000000000000000000000000000000000000000000000002a00000000",
            INIT_0C => X"0000000000000000000000260000000000000018000000000000007a00000000",
            INIT_0D => X"000000110000000000000000000000000000000f000000000000005700000000",
            INIT_0E => X"0000005900000000000000300000000000000000000000000000001700000000",
            INIT_0F => X"000000390000000000000000000000000000002b000000000000000000000000",
            INIT_10 => X"00000000000000000000000e0000000000000000000000000000000700000000",
            INIT_11 => X"00000004000000000000000c0000000000000000000000000000003400000000",
            INIT_12 => X"0000000000000000000000560000000000000052000000000000000000000000",
            INIT_13 => X"0000001c00000000000000000000000000000009000000000000004200000000",
            INIT_14 => X"0000000000000000000000190000000000000008000000000000000600000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"000000800000000000000000000000000000004d000000000000007500000000",
            INIT_17 => X"0000004e00000000000000500000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000008d0000000000000001000000000000001a000000000000000900000000",
            INIT_1A => X"0000005000000000000000940000000000000022000000000000007200000000",
            INIT_1B => X"000000150000000000000038000000000000003b000000000000002900000000",
            INIT_1C => X"0000001e000000000000001d0000000000000013000000000000001000000000",
            INIT_1D => X"00000073000000000000000e000000000000001a000000000000002000000000",
            INIT_1E => X"000000140000000000000009000000000000007a000000000000006d00000000",
            INIT_1F => X"0000000e000000000000000b0000000000000010000000000000001200000000",
            INIT_20 => X"000000290000000000000026000000000000001e000000000000001600000000",
            INIT_21 => X"0000009e000000000000001b0000000000000014000000000000002800000000",
            INIT_22 => X"00000009000000000000001c0000000000000007000000000000004d00000000",
            INIT_23 => X"00000022000000000000001c0000000000000017000000000000001200000000",
            INIT_24 => X"0000003b0000000000000034000000000000001c000000000000002f00000000",
            INIT_25 => X"0000004300000000000000270000000000000023000000000000001100000000",
            INIT_26 => X"0000001500000000000000280000000000000029000000000000000d00000000",
            INIT_27 => X"0000001b00000000000000150000000000000018000000000000001800000000",
            INIT_28 => X"0000000000000000000000000000000000000025000000000000003000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000d00000000000000060000000000000009000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000004000000000000001700000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000300000000000000060000000000000003000000000000000b00000000",
            INIT_37 => X"000000240000000000000000000000000000000a000000000000001100000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"00000008000000000000000e0000000000000005000000000000000000000000",
            INIT_3A => X"0000000a000000000000000a0000000000000006000000000000001500000000",
            INIT_3B => X"00000005000000000000002d0000000000000000000000000000000f00000000",
            INIT_3C => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000400000000000000060000000000000008000000000000000000000000",
            INIT_3E => X"00000014000000000000000b0000000000000017000000000000000600000000",
            INIT_3F => X"000000000000000000000000000000000000003a000000000000001500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"000000140000000000000000000000000000000b000000000000000e00000000",
            INIT_42 => X"000000080000000000000011000000000000000f000000000000001300000000",
            INIT_43 => X"000000000000000000000011000000000000001c000000000000002d00000000",
            INIT_44 => X"00000004000000000000000c0000000000000000000000000000000000000000",
            INIT_45 => X"0000001000000000000000060000000000000000000000000000000d00000000",
            INIT_46 => X"0000002600000000000000000000000000000003000000000000001100000000",
            INIT_47 => X"0000000000000000000000090000000000000025000000000000001d00000000",
            INIT_48 => X"0000000e00000000000000000000000000000008000000000000000700000000",
            INIT_49 => X"0000000b00000000000000110000000000000000000000000000000000000000",
            INIT_4A => X"0000001800000000000000150000000000000000000000000000000000000000",
            INIT_4B => X"0000001100000000000000140000000000000018000000000000001f00000000",
            INIT_4C => X"0000000100000000000000080000000000000005000000000000001800000000",
            INIT_4D => X"000000000000000000000005000000000000001c000000000000000d00000000",
            INIT_4E => X"0000001c00000000000000180000000000000013000000000000000000000000",
            INIT_4F => X"00000010000000000000001b000000000000001e000000000000001d00000000",
            INIT_50 => X"0000003300000000000000230000000000000028000000000000001f00000000",
            INIT_51 => X"0000002600000000000000240000000000000030000000000000003500000000",
            INIT_52 => X"00000000000000000000002a0000000000000031000000000000003400000000",
            INIT_53 => X"00000043000000000000003f000000000000004d000000000000000b00000000",
            INIT_54 => X"0000004d00000000000000490000000000000045000000000000004800000000",
            INIT_55 => X"000000570000000000000053000000000000004e000000000000005300000000",
            INIT_56 => X"000000500000000000000000000000000000003b000000000000003900000000",
            INIT_57 => X"0000004900000000000000480000000000000049000000000000004c00000000",
            INIT_58 => X"0000004f00000000000000540000000000000053000000000000004d00000000",
            INIT_59 => X"0000005800000000000000640000000000000060000000000000005700000000",
            INIT_5A => X"0000004b0000000000000046000000000000001d000000000000003800000000",
            INIT_5B => X"00000051000000000000004e000000000000004a000000000000004c00000000",
            INIT_5C => X"0000005f000000000000005d0000000000000057000000000000005400000000",
            INIT_5D => X"0000004b000000000000005e0000000000000061000000000000005000000000",
            INIT_5E => X"0000004a00000000000000480000000000000044000000000000003e00000000",
            INIT_5F => X"00000051000000000000004f000000000000004a000000000000004e00000000",
            INIT_60 => X"000000610000000000000055000000000000005a000000000000005800000000",
            INIT_61 => X"0000008600000000000000850000000000000086000000000000008100000000",
            INIT_62 => X"00000092000000000000008b0000000000000080000000000000008400000000",
            INIT_63 => X"0000006900000000000000640000000000000072000000000000008600000000",
            INIT_64 => X"0000008000000000000000720000000000000075000000000000006c00000000",
            INIT_65 => X"000000880000000000000088000000000000008d000000000000008b00000000",
            INIT_66 => X"0000005900000000000000780000000000000078000000000000007800000000",
            INIT_67 => X"00000046000000000000002c000000000000001c000000000000003600000000",
            INIT_68 => X"000000710000000000000062000000000000006e000000000000005f00000000",
            INIT_69 => X"00000094000000000000008c000000000000008a000000000000008800000000",
            INIT_6A => X"0000003600000000000000270000000000000035000000000000004100000000",
            INIT_6B => X"000000390000000000000019000000000000001e000000000000002000000000",
            INIT_6C => X"0000007c00000000000000490000000000000015000000000000006100000000",
            INIT_6D => X"0000003900000000000000570000000000000072000000000000008c00000000",
            INIT_6E => X"0000002000000000000000480000000000000018000000000000001f00000000",
            INIT_6F => X"0000005c0000000000000011000000000000000e000000000000002900000000",
            INIT_70 => X"000000850000000000000066000000000000003f000000000000000000000000",
            INIT_71 => X"0000001a000000000000002f0000000000000049000000000000005100000000",
            INIT_72 => X"00000019000000000000002e0000000000000033000000000000001900000000",
            INIT_73 => X"000000030000000000000039000000000000000f000000000000002100000000",
            INIT_74 => X"0000005400000000000000630000000000000059000000000000002d00000000",
            INIT_75 => X"000000100000000000000028000000000000002a000000000000003c00000000",
            INIT_76 => X"0000002900000000000000100000000000000027000000000000005100000000",
            INIT_77 => X"0000001f00000000000000000000000000000010000000000000001700000000",
            INIT_78 => X"0000004000000000000000670000000000000065000000000000004800000000",
            INIT_79 => X"0000005500000000000000170000000000000020000000000000004100000000",
            INIT_7A => X"0000001b0000000000000019000000000000000f000000000000001100000000",
            INIT_7B => X"0000002000000000000000180000000000000006000000000000001e00000000",
            INIT_7C => X"0000002e00000000000000610000000000000055000000000000004000000000",
            INIT_7D => X"0000001b0000000000000062000000000000001a000000000000003000000000",
            INIT_7E => X"00000041000000000000002e0000000000000023000000000000001100000000",
            INIT_7F => X"000000280000000000000000000000000000001f000000000000000b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE1;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE2 : if BRAM_NAME = "samplegold_layersamples_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002100000000000000220000000000000037000000000000002b00000000",
            INIT_01 => X"0000001a0000000000000035000000000000003e000000000000002e00000000",
            INIT_02 => X"00000020000000000000006c0000000000000041000000000000002200000000",
            INIT_03 => X"0000001900000000000000240000000000000000000000000000002100000000",
            INIT_04 => X"0000002700000000000000200000000000000031000000000000003000000000",
            INIT_05 => X"00000029000000000000000f0000000000000018000000000000003600000000",
            INIT_06 => X"000000220000000000000022000000000000006b000000000000006900000000",
            INIT_07 => X"0000000e00000000000000000000000000000044000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000020000000000000002d00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"00000010000000000000000f0000000000000009000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000005900000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000003000000000000000160000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"000000250000000000000024000000000000002a000000000000000000000000",
            INIT_1A => X"0000002a00000000000000230000000000000027000000000000002500000000",
            INIT_1B => X"0000002000000000000000210000000000000023000000000000002a00000000",
            INIT_1C => X"000000210000000000000025000000000000001f000000000000002600000000",
            INIT_1D => X"0000002500000000000000260000000000000027000000000000002a00000000",
            INIT_1E => X"00000022000000000000001b0000000000000020000000000000002300000000",
            INIT_1F => X"00000021000000000000000a000000000000000f000000000000000900000000",
            INIT_20 => X"000000270000000000000026000000000000002b000000000000003100000000",
            INIT_21 => X"0000002c0000000000000025000000000000002c000000000000003100000000",
            INIT_22 => X"0000001200000000000000110000000000000001000000000000003a00000000",
            INIT_23 => X"0000000e0000000000000007000000000000000b000000000000002100000000",
            INIT_24 => X"000000570000000000000000000000000000002d000000000000003600000000",
            INIT_25 => X"0000001000000000000000200000000000000027000000000000003000000000",
            INIT_26 => X"0000003500000000000000150000000000000006000000000000000a00000000",
            INIT_27 => X"0000001e00000000000000020000000000000016000000000000000000000000",
            INIT_28 => X"0000001b000000000000003d0000000000000000000000000000004300000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_2A => X"000000040000000000000028000000000000001a000000000000000100000000",
            INIT_2B => X"0000004300000000000000070000000000000018000000000000000000000000",
            INIT_2C => X"0000001900000000000000100000000000000027000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_2E => X"000000000000000000000000000000000000004f000000000000000900000000",
            INIT_2F => X"00000000000000000000000e0000000000000005000000000000001f00000000",
            INIT_30 => X"0000003b00000000000000020000000000000023000000000000001900000000",
            INIT_31 => X"0000000000000000000000000000000000000004000000000000001200000000",
            INIT_32 => X"0000001c00000000000000020000000000000000000000000000005100000000",
            INIT_33 => X"0000000000000000000000000000000000000015000000000000001300000000",
            INIT_34 => X"0000002c000000000000001c000000000000000c000000000000000e00000000",
            INIT_35 => X"0000004a00000000000000010000000000000011000000000000000000000000",
            INIT_36 => X"00000024000000000000001e0000000000000004000000000000000000000000",
            INIT_37 => X"0000000000000000000000020000000000000000000000000000001c00000000",
            INIT_38 => X"000000070000000000000013000000000000000f000000000000001b00000000",
            INIT_39 => X"00000029000000000000001c0000000000000020000000000000001300000000",
            INIT_3A => X"0000002b00000000000000270000000000000028000000000000000200000000",
            INIT_3B => X"0000002100000000000000000000000000000006000000000000000000000000",
            INIT_3C => X"00000000000000000000000c0000000000000013000000000000000000000000",
            INIT_3D => X"0000000e0000000000000000000000000000000e000000000000002800000000",
            INIT_3E => X"000000230000000000000021000000000000003f000000000000003100000000",
            INIT_3F => X"0000000000000000000000370000000000000000000000000000000400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000019000000000000000000000000",
            INIT_41 => X"0000001d00000000000000090000000000000011000000000000000000000000",
            INIT_42 => X"0000000c00000000000000480000000000000006000000000000001d00000000",
            INIT_43 => X"0000000000000000000000000000000000000039000000000000000000000000",
            INIT_44 => X"0000000900000000000000040000000000000011000000000000001700000000",
            INIT_45 => X"00000013000000000000000a000000000000000f000000000000000f00000000",
            INIT_46 => X"0000001300000000000000440000000000000011000000000000000800000000",
            INIT_47 => X"0000000900000000000000080000000000000000000000000000001700000000",
            INIT_48 => X"0000000e0000000000000010000000000000000f000000000000000e00000000",
            INIT_49 => X"0000000900000000000000040000000000000010000000000000001100000000",
            INIT_4A => X"0000000000000000000000520000000000000013000000000000000200000000",
            INIT_4B => X"0000000f00000000000000050000000000000010000000000000000000000000",
            INIT_4C => X"00000011000000000000000f000000000000000d000000000000000a00000000",
            INIT_4D => X"0000000000000000000000160000000000000015000000000000000500000000",
            INIT_4E => X"0000001100000000000000200000000000000019000000000000000c00000000",
            INIT_4F => X"0000000900000000000000080000000000000011000000000000001d00000000",
            INIT_50 => X"0000000d000000000000000d000000000000000a000000000000000900000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000001200000000000000020000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000005000000000000001200000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"000000010000000000000000000000000000000c000000000000000000000000",
            INIT_5B => X"0000002e000000000000003f000000000000003b000000000000000500000000",
            INIT_5C => X"000000060000000000000000000000000000000b000000000000001c00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_5E => X"0000002600000000000000140000000000000010000000000000000000000000",
            INIT_5F => X"000000210000000000000029000000000000002b000000000000004200000000",
            INIT_60 => X"0000004400000000000000210000000000000004000000000000001300000000",
            INIT_61 => X"0000001200000000000000140000000000000000000000000000000000000000",
            INIT_62 => X"00000029000000000000002b000000000000001e000000000000002c00000000",
            INIT_63 => X"0000001300000000000000270000000000000015000000000000003100000000",
            INIT_64 => X"0000000000000000000000680000000000000046000000000000000f00000000",
            INIT_65 => X"000000310000000000000026000000000000006e000000000000000000000000",
            INIT_66 => X"00000041000000000000004e0000000000000020000000000000001f00000000",
            INIT_67 => X"0000000d00000000000000220000000000000031000000000000002100000000",
            INIT_68 => X"000000000000000000000002000000000000006f000000000000003900000000",
            INIT_69 => X"0000002a00000000000000510000000000000033000000000000003300000000",
            INIT_6A => X"00000028000000000000003b000000000000006c000000000000002300000000",
            INIT_6B => X"00000048000000000000001f0000000000000031000000000000002f00000000",
            INIT_6C => X"0000000b0000000000000000000000000000001e000000000000006200000000",
            INIT_6D => X"0000002000000000000000440000000000000048000000000000006100000000",
            INIT_6E => X"0000003500000000000000300000000000000038000000000000005600000000",
            INIT_6F => X"0000007c00000000000000630000000000000004000000000000003600000000",
            INIT_70 => X"0000003d00000000000000150000000000000042000000000000003b00000000",
            INIT_71 => X"0000002000000000000000290000000000000031000000000000002900000000",
            INIT_72 => X"00000015000000000000002a0000000000000022000000000000003900000000",
            INIT_73 => X"00000048000000000000007a000000000000006f000000000000000000000000",
            INIT_74 => X"0000002d000000000000001b0000000000000036000000000000006300000000",
            INIT_75 => X"0000001f0000000000000026000000000000003a000000000000004000000000",
            INIT_76 => X"000000000000000000000000000000000000001e000000000000001600000000",
            INIT_77 => X"0000007a000000000000004f000000000000006b000000000000008900000000",
            INIT_78 => X"0000007200000000000000680000000000000038000000000000004000000000",
            INIT_79 => X"00000045000000000000003c000000000000002b000000000000003a00000000",
            INIT_7A => X"000000c5000000000000004e0000000000000063000000000000005e00000000",
            INIT_7B => X"000000930000000000000099000000000000004e000000000000008f00000000",
            INIT_7C => X"000000770000000000000087000000000000008b000000000000007c00000000",
            INIT_7D => X"00000096000000000000008e0000000000000085000000000000007600000000",
            INIT_7E => X"000000b100000000000000a70000000000000096000000000000009d00000000",
            INIT_7F => X"00000080000000000000006c00000000000000a5000000000000007700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE2;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE3 : if BRAM_NAME = "samplegold_layersamples_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000087000000000000007f000000000000007f000000000000007f00000000",
            INIT_01 => X"0000009d00000000000000a0000000000000009c000000000000009300000000",
            INIT_02 => X"000000b1000000000000009c00000000000000ac00000000000000a900000000",
            INIT_03 => X"00000082000000000000008a000000000000006e00000000000000a600000000",
            INIT_04 => X"000000a100000000000000910000000000000084000000000000008200000000",
            INIT_05 => X"000000c200000000000000b700000000000000a300000000000000ac00000000",
            INIT_06 => X"000000a5000000000000009b00000000000000a700000000000000aa00000000",
            INIT_07 => X"00000083000000000000008f0000000000000091000000000000008200000000",
            INIT_08 => X"0000009900000000000000970000000000000095000000000000008600000000",
            INIT_09 => X"00000078000000000000009900000000000000bd00000000000000a400000000",
            INIT_0A => X"0000007e000000000000007f000000000000007b000000000000007b00000000",
            INIT_0B => X"00000082000000000000008b000000000000007c000000000000007600000000",
            INIT_0C => X"0000006100000000000000560000000000000053000000000000006500000000",
            INIT_0D => X"00000081000000000000007a0000000000000073000000000000006e00000000",
            INIT_0E => X"00000061000000000000007f0000000000000081000000000000007e00000000",
            INIT_0F => X"0000003200000000000000500000000000000063000000000000006f00000000",
            INIT_10 => X"00000050000000000000002f0000000000000020000000000000001d00000000",
            INIT_11 => X"0000008100000000000000500000000000000047000000000000006900000000",
            INIT_12 => X"0000004e00000000000000670000000000000083000000000000008500000000",
            INIT_13 => X"0000001d0000000000000013000000000000002a000000000000003900000000",
            INIT_14 => X"0000004d0000000000000029000000000000001d000000000000001e00000000",
            INIT_15 => X"0000007f00000000000000730000000000000021000000000000003100000000",
            INIT_16 => X"0000002900000000000000320000000000000053000000000000006700000000",
            INIT_17 => X"000000230000000000000029000000000000001a000000000000001a00000000",
            INIT_18 => X"000000280000000000000031000000000000001f000000000000002200000000",
            INIT_19 => X"0000002b00000000000000690000000000000067000000000000000c00000000",
            INIT_1A => X"0000001800000000000000250000000000000029000000000000003100000000",
            INIT_1B => X"0000001c000000000000002a0000000000000028000000000000001d00000000",
            INIT_1C => X"0000000600000000000000220000000000000022000000000000002000000000",
            INIT_1D => X"0000003600000000000000150000000000000068000000000000006600000000",
            INIT_1E => X"00000004000000000000001e000000000000002f000000000000002700000000",
            INIT_1F => X"0000001e00000000000000190000000000000029000000000000002400000000",
            INIT_20 => X"0000003e0000000000000000000000000000002b000000000000001d00000000",
            INIT_21 => X"0000001c00000000000000270000000000000028000000000000006d00000000",
            INIT_22 => X"0000002700000000000000000000000000000025000000000000002800000000",
            INIT_23 => X"00000026000000000000001a0000000000000019000000000000002200000000",
            INIT_24 => X"0000003b0000000000000022000000000000000c000000000000001d00000000",
            INIT_25 => X"0000001e0000000000000026000000000000000e000000000000004300000000",
            INIT_26 => X"00000026000000000000002b0000000000000022000000000000002d00000000",
            INIT_27 => X"00000012000000000000004f000000000000001e000000000000001600000000",
            INIT_28 => X"00000031000000000000000c000000000000001c000000000000000000000000",
            INIT_29 => X"0000001d000000000000001f0000000000000032000000000000002900000000",
            INIT_2A => X"0000001c00000000000000280000000000000029000000000000003400000000",
            INIT_2B => X"0000000c0000000000000016000000000000005c000000000000003b00000000",
            INIT_2C => X"0000002300000000000000180000000000000000000000000000001600000000",
            INIT_2D => X"00000025000000000000001d0000000000000018000000000000002100000000",
            INIT_2E => X"00000040000000000000000c0000000000000014000000000000001b00000000",
            INIT_2F => X"00000016000000000000000f0000000000000000000000000000005e00000000",
            INIT_30 => X"00000000000000000000000a0000000000000014000000000000000000000000",
            INIT_31 => X"0000000000000000000000040000000000000001000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000040000000000000000000000000000000500000000",
            INIT_43 => X"0000000000000000000000030000000000000001000000000000000000000000",
            INIT_44 => X"0000001100000000000000020000000000000000000000000000000000000000",
            INIT_45 => X"0000000200000000000000000000000000000000000000000000000400000000",
            INIT_46 => X"0000000800000000000000000000000000000005000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000001600000000000000000000000000000000000000000000001500000000",
            INIT_49 => X"0000004400000000000000000000000000000000000000000000001c00000000",
            INIT_4A => X"0000001c00000000000000080000000000000000000000000000000400000000",
            INIT_4B => X"0000003d00000000000000090000000000000000000000000000000000000000",
            INIT_4C => X"0000002400000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"00000000000000000000005f0000000000000000000000000000002200000000",
            INIT_4E => X"0000000000000000000000160000000000000000000000000000000800000000",
            INIT_4F => X"00000000000000000000006d0000000000000000000000000000000000000000",
            INIT_50 => X"0000005f00000000000000000000000000000000000000000000000200000000",
            INIT_51 => X"000000520000000000000000000000000000001c000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000086000000000000000000000000",
            INIT_54 => X"0000000000000000000000330000000000000000000000000000000000000000",
            INIT_55 => X"0000007600000000000000190000000000000000000000000000001800000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_57 => X"000000130000000000000000000000000000000000000000000000d200000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"00000040000000000000005f0000000000000000000000000000000f00000000",
            INIT_5A => X"000000b100000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"00000010000000000000000b0000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"000000000000000000000054000000000000003d000000000000000000000000",
            INIT_5E => X"0000000000000000000000740000000000000000000000000000000500000000",
            INIT_5F => X"00000000000000000000000f0000000000000025000000000000000000000000",
            INIT_60 => X"0000003100000000000000000000000000000007000000000000000000000000",
            INIT_61 => X"000000000000000000000000000000000000002e000000000000000000000000",
            INIT_62 => X"0000000000000000000000200000000000000000000000000000002700000000",
            INIT_63 => X"00000000000000000000000b0000000000000025000000000000002b00000000",
            INIT_64 => X"0000000000000000000000550000000000000000000000000000000d00000000",
            INIT_65 => X"0000000000000000000000000000000000000034000000000000000c00000000",
            INIT_66 => X"0000002f00000000000000040000000000000000000000000000000300000000",
            INIT_67 => X"00000005000000000000005a0000000000000000000000000000002900000000",
            INIT_68 => X"00000000000000000000000000000000000000aa000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000003e00000000",
            INIT_6A => X"0000001f00000000000000160000000000000006000000000000000000000000",
            INIT_6B => X"00000000000000000000004c0000000000000075000000000000000000000000",
            INIT_6C => X"0000001f00000000000000000000000000000000000000000000007a00000000",
            INIT_6D => X"0000000c00000000000000080000000000000000000000000000001a00000000",
            INIT_6E => X"00000000000000000000000d000000000000000c000000000000001000000000",
            INIT_6F => X"0000000000000000000000840000000000000071000000000000000000000000",
            INIT_70 => X"0000000600000000000000000000000000000002000000000000000000000000",
            INIT_71 => X"00000008000000000000000d0000000000000009000000000000000200000000",
            INIT_72 => X"00000000000000000000000e000000000000000f000000000000000600000000",
            INIT_73 => X"00000000000000000000000000000000000000bd000000000000001100000000",
            INIT_74 => X"0000000e00000000000000010000000000000000000000000000000c00000000",
            INIT_75 => X"000000040000000000000010000000000000000b000000000000000b00000000",
            INIT_76 => X"0000000c00000000000000000000000000000000000000000000002000000000",
            INIT_77 => X"0000002500000000000000000000000000000007000000000000002300000000",
            INIT_78 => X"00000000000000000000000b0000000000000006000000000000001800000000",
            INIT_79 => X"00000000000000000000002d000000000000000f000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000002500000000000000160000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000004000000000000001c00000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000e00000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE3;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE4 : if BRAM_NAME = "samplegold_layersamples_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000000000000c000000000000004500000000",
            INIT_01 => X"0000002700000000000000000000000000000018000000000000001d00000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_03 => X"00000001000000000000002b0000000000000025000000000000004e00000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000006000000000000001e00000000",
            INIT_06 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"00000000000000000000000a0000000000000010000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_0B => X"0000000000000000000000070000000000000009000000000000000000000000",
            INIT_0C => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000002900000000000000000000000000000000000000000000000a00000000",
            INIT_0E => X"0000000000000000000000000000000000000022000000000000006400000000",
            INIT_0F => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_11 => X"000000280000000000000000000000000000001a000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000600000000000000050000000000000000000000000000000000000000",
            INIT_16 => X"000000050000000000000000000000000000002b000000000000002000000000",
            INIT_17 => X"00000007000000000000000b0000000000000000000000000000000100000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000600000000000000540000000000000000000000000000000000000000",
            INIT_1A => X"0000003100000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"000000000000000000000000000000000000001f000000000000003a00000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_1D => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_1E => X"0000001a0000000000000037000000000000003f000000000000000000000000",
            INIT_1F => X"0000001000000000000000050000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"00000008000000000000002f0000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"000000320000000000000065000000000000002b000000000000002700000000",
            INIT_24 => X"0000006800000000000000500000000000000000000000000000000000000000",
            INIT_25 => X"00000013000000000000001e0000000000000043000000000000004600000000",
            INIT_26 => X"0000000000000000000000000000000000000009000000000000000500000000",
            INIT_27 => X"0000001900000000000000490000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000056000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_2B => X"0000004100000000000000510000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_2D => X"0000001300000000000000060000000000000000000000000000000200000000",
            INIT_2E => X"0000000000000000000000260000000000000000000000000000000800000000",
            INIT_2F => X"0000001f000000000000004e000000000000000b000000000000000000000000",
            INIT_30 => X"0000000000000000000000010000000000000024000000000000002400000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"000000a600000000000000a80000000000000000000000000000000000000000",
            INIT_33 => X"000000a400000000000000ad00000000000000ad00000000000000af00000000",
            INIT_34 => X"0000009100000000000000aa00000000000000b700000000000000b800000000",
            INIT_35 => X"00000096000000000000008f0000000000000086000000000000007b00000000",
            INIT_36 => X"000000b500000000000000b300000000000000ab000000000000008a00000000",
            INIT_37 => X"000000b300000000000000c400000000000000b400000000000000b200000000",
            INIT_38 => X"0000004f0000000000000057000000000000006400000000000000a000000000",
            INIT_39 => X"000000920000000000000080000000000000005d000000000000005200000000",
            INIT_3A => X"000000b100000000000000b6000000000000008d000000000000007200000000",
            INIT_3B => X"000000350000000000000054000000000000008b00000000000000b600000000",
            INIT_3C => X"0000003b00000000000000460000000000000065000000000000004100000000",
            INIT_3D => X"0000002a00000000000000850000000000000051000000000000003500000000",
            INIT_3E => X"000000a200000000000000b700000000000000b9000000000000009400000000",
            INIT_3F => X"00000034000000000000003f0000000000000071000000000000007f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000014000000000000003d0000000000000043000000000000006900000000",
            INIT_41 => X"000000a3000000000000002f0000000000000076000000000000001e00000000",
            INIT_42 => X"000000ac00000000000000c600000000000000bf00000000000000ad00000000",
            INIT_43 => X"00000063000000000000001c0000000000000036000000000000005a00000000",
            INIT_44 => X"0000001f000000000000003b0000000000000040000000000000006900000000",
            INIT_45 => X"000000a400000000000000770000000000000039000000000000004f00000000",
            INIT_46 => X"0000006800000000000000670000000000000057000000000000008400000000",
            INIT_47 => X"0000006200000000000000ac0000000000000021000000000000004900000000",
            INIT_48 => X"0000002f000000000000002c000000000000003e000000000000001f00000000",
            INIT_49 => X"00000077000000000000007c000000000000005a000000000000004400000000",
            INIT_4A => X"0000005d000000000000007b0000000000000095000000000000006e00000000",
            INIT_4B => X"0000002e000000000000003d000000000000009e000000000000002400000000",
            INIT_4C => X"0000005c00000000000000420000000000000043000000000000003500000000",
            INIT_4D => X"00000080000000000000007c0000000000000069000000000000005400000000",
            INIT_4E => X"0000002a0000000000000041000000000000004700000000000000ae00000000",
            INIT_4F => X"000000380000000000000022000000000000003e000000000000008f00000000",
            INIT_50 => X"0000006d000000000000005a0000000000000058000000000000004b00000000",
            INIT_51 => X"0000003600000000000000740000000000000065000000000000002b00000000",
            INIT_52 => X"00000064000000000000005f0000000000000048000000000000003b00000000",
            INIT_53 => X"0000005e00000000000000220000000000000004000000000000004400000000",
            INIT_54 => X"000000220000000000000069000000000000005a00000000000000a300000000",
            INIT_55 => X"000000630000000000000053000000000000004b000000000000005e00000000",
            INIT_56 => X"0000000800000000000000400000000000000059000000000000006a00000000",
            INIT_57 => X"0000009400000000000000a7000000000000004c000000000000000800000000",
            INIT_58 => X"000000b3000000000000001f0000000000000074000000000000006d00000000",
            INIT_59 => X"0000004d00000000000000850000000000000077000000000000007c00000000",
            INIT_5A => X"0000002000000000000000110000000000000015000000000000001f00000000",
            INIT_5B => X"00000024000000000000002d000000000000003c000000000000002900000000",
            INIT_5C => X"0000002200000000000000de0000000000000059000000000000004f00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"000000000000000000000000000000000000008d000000000000006f00000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000005a00000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000c00000000000000000000000000000000000000000000000900000000",
            INIT_6B => X"0000000e0000000000000011000000000000000b000000000000001100000000",
            INIT_6C => X"0000000d0000000000000011000000000000000d000000000000000900000000",
            INIT_6D => X"000000090000000000000003000000000000000e000000000000000d00000000",
            INIT_6E => X"0000000900000000000000060000000000000013000000000000000f00000000",
            INIT_6F => X"0000000000000000000000070000000000000014000000000000000800000000",
            INIT_70 => X"0000000000000000000000270000000000000009000000000000002100000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_72 => X"0000000900000000000000000000000000000013000000000000000b00000000",
            INIT_73 => X"0000003a000000000000000e0000000000000007000000000000001200000000",
            INIT_74 => X"0000003100000000000000000000000000000000000000000000001000000000",
            INIT_75 => X"000000000000000000000000000000000000002e000000000000002600000000",
            INIT_76 => X"00000001000000000000000a0000000000000000000000000000005e00000000",
            INIT_77 => X"0000002700000000000000140000000000000000000000000000000f00000000",
            INIT_78 => X"0000001a00000000000000540000000000000000000000000000001500000000",
            INIT_79 => X"0000007d00000000000000000000000000000013000000000000003500000000",
            INIT_7A => X"0000001800000000000000000000000000000037000000000000000000000000",
            INIT_7B => X"0000002200000000000000390000000000000052000000000000002800000000",
            INIT_7C => X"0000000700000000000000490000000000000023000000000000000000000000",
            INIT_7D => X"00000009000000000000006c0000000000000000000000000000002d00000000",
            INIT_7E => X"0000004c0000000000000000000000000000001b000000000000004e00000000",
            INIT_7F => X"000000000000000000000040000000000000003b000000000000005100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE4;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE5 : if BRAM_NAME = "samplegold_layersamples_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000270000000000000000000000000000005f000000000000006b00000000",
            INIT_01 => X"00000013000000000000003f0000000000000068000000000000001400000000",
            INIT_02 => X"0000004100000000000000000000000000000000000000000000004700000000",
            INIT_03 => X"0000007900000000000000000000000000000059000000000000004a00000000",
            INIT_04 => X"0000002800000000000000000000000000000002000000000000003900000000",
            INIT_05 => X"000000210000000000000023000000000000004e000000000000005700000000",
            INIT_06 => X"0000003200000000000000900000000000000000000000000000000000000000",
            INIT_07 => X"00000045000000000000005a0000000000000000000000000000004200000000",
            INIT_08 => X"00000065000000000000002c0000000000000013000000000000000000000000",
            INIT_09 => X"0000001d0000000000000000000000000000007d000000000000002400000000",
            INIT_0A => X"00000000000000000000000f0000000000000031000000000000002600000000",
            INIT_0B => X"00000000000000000000005b0000000000000000000000000000002800000000",
            INIT_0C => X"0000003000000000000000460000000000000000000000000000000000000000",
            INIT_0D => X"0000001500000000000000440000000000000000000000000000008f00000000",
            INIT_0E => X"0000002d0000000000000015000000000000002f000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000007000000000000005400000000",
            INIT_10 => X"00000089000000000000002c0000000000000000000000000000001700000000",
            INIT_11 => X"000000000000000000000023000000000000008d000000000000000000000000",
            INIT_12 => X"0000000000000000000000280000000000000069000000000000004e00000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"000000000000000000000054000000000000000c000000000000000000000000",
            INIT_15 => X"000000110000000000000010000000000000006400000000000000c200000000",
            INIT_16 => X"0000000800000000000000080000000000000009000000000000001c00000000",
            INIT_17 => X"00000021000000000000001b000000000000000f000000000000000c00000000",
            INIT_18 => X"000000b600000000000000410000000000000000000000000000000000000000",
            INIT_19 => X"000000110000000000000011000000000000001a000000000000001400000000",
            INIT_1A => X"0000001500000000000000030000000000000004000000000000000800000000",
            INIT_1B => X"0000000600000000000000310000000000000003000000000000001700000000",
            INIT_1C => X"0000000b00000000000000410000000000000091000000000000000000000000",
            INIT_1D => X"0000000c000000000000000e0000000000000010000000000000002000000000",
            INIT_1E => X"00000000000000000000001f0000000000000014000000000000001200000000",
            INIT_1F => X"0000000700000000000000110000000000000040000000000000003700000000",
            INIT_20 => X"000000150000000000000000000000000000001f000000000000001d00000000",
            INIT_21 => X"000000220000000000000011000000000000000b000000000000001a00000000",
            INIT_22 => X"00000050000000000000002f0000000000000000000000000000001000000000",
            INIT_23 => X"00000053000000000000004b0000000000000053000000000000004d00000000",
            INIT_24 => X"000000550000000000000054000000000000004a000000000000004f00000000",
            INIT_25 => X"000000400000000000000047000000000000004a000000000000004e00000000",
            INIT_26 => X"0000004a0000000000000049000000000000004b000000000000004800000000",
            INIT_27 => X"000000490000000000000058000000000000004a000000000000004f00000000",
            INIT_28 => X"00000054000000000000004f0000000000000068000000000000004c00000000",
            INIT_29 => X"0000002600000000000000340000000000000041000000000000002c00000000",
            INIT_2A => X"00000032000000000000004f0000000000000048000000000000003a00000000",
            INIT_2B => X"00000049000000000000004b0000000000000057000000000000005200000000",
            INIT_2C => X"00000009000000000000001f0000000000000040000000000000007c00000000",
            INIT_2D => X"0000001700000000000000530000000000000050000000000000006200000000",
            INIT_2E => X"0000005b0000000000000000000000000000008e000000000000003600000000",
            INIT_2F => X"00000056000000000000002f0000000000000059000000000000004700000000",
            INIT_30 => X"0000008e0000000000000000000000000000003a000000000000004500000000",
            INIT_31 => X"000000000000000000000036000000000000005c000000000000004300000000",
            INIT_32 => X"000000040000000000000082000000000000002500000000000000b200000000",
            INIT_33 => X"00000065000000000000008f0000000000000053000000000000007a00000000",
            INIT_34 => X"00000075000000000000006a0000000000000000000000000000004500000000",
            INIT_35 => X"0000009400000000000000000000000000000050000000000000003200000000",
            INIT_36 => X"00000044000000000000003b00000000000000a1000000000000006800000000",
            INIT_37 => X"0000006c000000000000006d00000000000000aa000000000000008900000000",
            INIT_38 => X"00000029000000000000008b00000000000000a9000000000000000000000000",
            INIT_39 => X"0000009500000000000000950000000000000036000000000000004a00000000",
            INIT_3A => X"0000003800000000000000000000000000000086000000000000006f00000000",
            INIT_3B => X"00000000000000000000008a0000000000000089000000000000009700000000",
            INIT_3C => X"0000002f000000000000002b000000000000006b00000000000000be00000000",
            INIT_3D => X"0000005600000000000000a40000000000000095000000000000005600000000",
            INIT_3E => X"000000be000000000000002a0000000000000009000000000000007700000000",
            INIT_3F => X"000000990000000000000000000000000000007b000000000000006700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005a0000000000000041000000000000001c000000000000007700000000",
            INIT_41 => X"0000004200000000000000b2000000000000007900000000000000ad00000000",
            INIT_42 => X"0000004d00000000000000740000000000000050000000000000005600000000",
            INIT_43 => X"00000077000000000000003e000000000000005c000000000000002900000000",
            INIT_44 => X"00000097000000000000003b0000000000000032000000000000001600000000",
            INIT_45 => X"0000008d000000000000000e00000000000000d6000000000000007a00000000",
            INIT_46 => X"0000003f0000000000000080000000000000002b000000000000002c00000000",
            INIT_47 => X"000000030000000000000021000000000000006d000000000000005d00000000",
            INIT_48 => X"0000007f0000000000000042000000000000005f000000000000002600000000",
            INIT_49 => X"0000006000000000000000ec000000000000000000000000000000ce00000000",
            INIT_4A => X"0000004a000000000000009d0000000000000092000000000000002300000000",
            INIT_4B => X"00000028000000000000000f000000000000000d000000000000001500000000",
            INIT_4C => X"0000009d00000000000000600000000000000006000000000000004300000000",
            INIT_4D => X"0000003f000000000000009e0000000000000111000000000000001600000000",
            INIT_4E => X"00000029000000000000002a000000000000004a000000000000004300000000",
            INIT_4F => X"0000004000000000000000300000000000000030000000000000002700000000",
            INIT_50 => X"000000ac00000000000000270000000000000001000000000000004300000000",
            INIT_51 => X"0000002f0000000000000036000000000000003600000000000000e100000000",
            INIT_52 => X"0000002800000000000000230000000000000025000000000000002e00000000",
            INIT_53 => X"0000005400000000000000300000000000000036000000000000003700000000",
            INIT_54 => X"0000006600000000000000f30000000000000000000000000000002a00000000",
            INIT_55 => X"00000028000000000000002f0000000000000042000000000000002b00000000",
            INIT_56 => X"0000003e0000000000000037000000000000002d000000000000002900000000",
            INIT_57 => X"0000002f000000000000005e0000000000000057000000000000001800000000",
            INIT_58 => X"0000001e000000000000003a0000000000000055000000000000002b00000000",
            INIT_59 => X"0000003600000000000000290000000000000038000000000000003200000000",
            INIT_5A => X"000000570000000000000014000000000000002b000000000000004100000000",
            INIT_5B => X"0000003b0000000000000034000000000000003a000000000000006f00000000",
            INIT_5C => X"0000004200000000000000340000000000000039000000000000003800000000",
            INIT_5D => X"0000002f000000000000002f0000000000000039000000000000004600000000",
            INIT_5E => X"0000002c00000000000000320000000000000032000000000000003400000000",
            INIT_5F => X"0000003b000000000000003a000000000000003b000000000000004000000000",
            INIT_60 => X"000000370000000000000039000000000000001f000000000000003700000000",
            INIT_61 => X"000000080000000000000000000000000000000c000000000000002700000000",
            INIT_62 => X"0000002400000000000000300000000000000037000000000000002300000000",
            INIT_63 => X"0000003c00000000000000400000000000000041000000000000004f00000000",
            INIT_64 => X"0000000100000000000000130000000000000025000000000000001100000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000001c0000000000000000000000000000002e000000000000001a00000000",
            INIT_67 => X"0000001f000000000000002e000000000000003d000000000000004400000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000003800000000000000000000000000000000000000000000002500000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"00000002000000000000003d0000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"00000000000000000000001c0000000000000047000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000022000000000000000400000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000001a00000000000000030000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE5;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE6 : if BRAM_NAME = "samplegold_layersamples_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000031000000000000001b000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000002400000000000000240000000000000000000000000000000000000000",
            INIT_14 => X"0000001c000000000000001f000000000000001e000000000000002000000000",
            INIT_15 => X"0000002400000000000000200000000000000029000000000000002700000000",
            INIT_16 => X"00000021000000000000001e0000000000000029000000000000002d00000000",
            INIT_17 => X"00000021000000000000001d000000000000001f000000000000001e00000000",
            INIT_18 => X"0000001d00000000000000000000000000000017000000000000002100000000",
            INIT_19 => X"000000000000000000000000000000000000003d000000000000002800000000",
            INIT_1A => X"00000019000000000000001d0000000000000023000000000000000700000000",
            INIT_1B => X"00000023000000000000001f0000000000000031000000000000003b00000000",
            INIT_1C => X"0000002200000000000000330000000000000042000000000000002400000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"000000000000000000000014000000000000001e000000000000000000000000",
            INIT_1F => X"0000001b000000000000001a0000000000000019000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000d0000000000000015000000000000000a000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000014000000000000001100000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_24 => X"0000000000000000000000180000000000000006000000000000000900000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000001e00000000000000000000000000000008000000000000002200000000",
            INIT_27 => X"00000000000000000000001f000000000000002b000000000000004400000000",
            INIT_28 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_2A => X"00000020000000000000002b0000000000000002000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_2C => X"00000000000000000000000c0000000000000000000000000000000100000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000a00000000000000250000000000000032000000000000000000000000",
            INIT_30 => X"00000000000000000000000d000000000000000d000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000013000000000000001000000000",
            INIT_32 => X"0000003800000000000000080000000000000000000000000000000c00000000",
            INIT_33 => X"0000001e00000000000000000000000000000000000000000000000d00000000",
            INIT_34 => X"000000000000000000000018000000000000003d000000000000001500000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_36 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_37 => X"000000330000000000000028000000000000000e000000000000000000000000",
            INIT_38 => X"0000001e00000000000000000000000000000000000000000000000700000000",
            INIT_39 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_3A => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_3C => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000004700000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"00000000000000000000000d0000000000000012000000000000002e00000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000100000000000000120000000000000017000000000000000700000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"00000000000000000000001c000000000000000e000000000000000000000000",
            INIT_52 => X"0000000c000000000000000d0000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000290000000000000022000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"00000004000000000000000e0000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_5A => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_5F => X"0000000900000000000000150000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_62 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"000000060000000000000014000000000000001d000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_6A => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"00000000000000000000000c0000000000000005000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000001400000000000000040000000000000000000000000000000000000000",
            INIT_6F => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000070000000000000000000000000000001600000000",
            INIT_71 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_72 => X"0000002f00000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000023000000000000002e00000000",
            INIT_74 => X"0000001b00000000000000190000000000000005000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000021000000000000002d00000000",
            INIT_76 => X"000000000000000000000000000000000000000e000000000000001500000000",
            INIT_77 => X"0000000000000000000000010000000000000002000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"00000003000000000000000b000000000000000b000000000000001c00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"000000000000000000000003000000000000001f000000000000003100000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE6;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE7 : if BRAM_NAME = "samplegold_layersamples_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_01 => X"0000000a00000000000000030000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000070000000000000005000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000003d00000000",
            INIT_13 => X"0000000000000000000000330000000000000000000000000000000000000000",
            INIT_14 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000c00000000000000000000000000000008000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000002000000000000002700000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000006800000000",
            INIT_1B => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_1C => X"000000000000000000000070000000000000005c000000000000001600000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"000000000000000000000073000000000000001b000000000000000000000000",
            INIT_1F => X"00000042000000000000000b0000000000000001000000000000003c00000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"00000020000000000000002e0000000000000022000000000000001100000000",
            INIT_22 => X"0000001a00000000000000170000000000000000000000000000010400000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000001400000000000000120000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000260000000000000000000000000000001100000000",
            INIT_2E => X"0000008e00000000000000080000000000000000000000000000000000000000",
            INIT_2F => X"00000044000000000000002e0000000000000023000000000000001600000000",
            INIT_30 => X"0000002700000000000000000000000000000000000000000000003a00000000",
            INIT_31 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_32 => X"00000000000000000000007a0000000000000001000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"000000000000000000000032000000000000001a000000000000001d00000000",
            INIT_35 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_36 => X"00000000000000000000000c000000000000003b000000000000000200000000",
            INIT_37 => X"00000001000000000000002e0000000000000036000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000021000000000000001a00000000",
            INIT_39 => X"0000000c000000000000000a0000000000000005000000000000000700000000",
            INIT_3A => X"0000004300000000000000330000000000000016000000000000001e00000000",
            INIT_3B => X"0000001500000000000000100000000000000000000000000000000900000000",
            INIT_3C => X"0000020f000000000000020f000000000000020f000000000000002000000000",
            INIT_3D => X"0000021100000000000002110000000000000210000000000000020f00000000",
            INIT_3E => X"00000210000000000000020e000000000000020f000000000000020f00000000",
            INIT_3F => X"00000212000000000000020f0000000000000210000000000000021000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000021100000000000002120000000000000212000000000000021100000000",
            INIT_41 => X"0000021200000000000002110000000000000210000000000000021000000000",
            INIT_42 => X"0000020a00000000000001e000000000000001cb000000000000020800000000",
            INIT_43 => X"0000020c00000000000002140000000000000211000000000000021100000000",
            INIT_44 => X"0000021400000000000002130000000000000214000000000000020e00000000",
            INIT_45 => X"000001b600000000000001ee000000000000020f000000000000021000000000",
            INIT_46 => X"000002130000000000000201000000000000019d000000000000018500000000",
            INIT_47 => X"00000211000000000000020d0000000000000217000000000000021400000000",
            INIT_48 => X"000001f100000000000002170000000000000217000000000000021700000000",
            INIT_49 => X"000001b900000000000001c400000000000001e300000000000001fb00000000",
            INIT_4A => X"00000219000000000000021900000000000001ff00000000000001b200000000",
            INIT_4B => X"0000020100000000000001700000000000000145000000000000021c00000000",
            INIT_4C => X"0000020b00000000000002030000000000000212000000000000020d00000000",
            INIT_4D => X"000001c300000000000001f5000000000000020b000000000000020900000000",
            INIT_4E => X"0000021e00000000000001d10000000000000178000000000000019900000000",
            INIT_4F => X"000001b900000000000001f900000000000001c300000000000001a000000000",
            INIT_50 => X"000001a7000000000000018a000000000000017b00000000000001d700000000",
            INIT_51 => X"000001bb00000000000001cb00000000000001f900000000000001e300000000",
            INIT_52 => X"000000fe000000000000021b00000000000001d8000000000000018b00000000",
            INIT_53 => X"000001c000000000000001ba000000000000017e000000000000013400000000",
            INIT_54 => X"000001be000000000000014500000000000000da00000000000000c000000000",
            INIT_55 => X"0000018a000000000000018b00000000000001bc00000000000001eb00000000",
            INIT_56 => X"00000132000000000000009500000000000001b4000000000000018c00000000",
            INIT_57 => X"0000019d00000000000001c30000000000000180000000000000010f00000000",
            INIT_58 => X"00000159000000000000017700000000000001a600000000000001ca00000000",
            INIT_59 => X"0000017400000000000001470000000000000128000000000000012d00000000",
            INIT_5A => X"000001a300000000000001cf0000000000000112000000000000019000000000",
            INIT_5B => X"000001de00000000000001e800000000000001f200000000000001ce00000000",
            INIT_5C => X"0000017f000000000000016e0000000000000186000000000000019200000000",
            INIT_5D => X"0000014100000000000001480000000000000147000000000000015b00000000",
            INIT_5E => X"0000013e000000000000013a0000000000000128000000000000012c00000000",
            INIT_5F => X"0000012800000000000001480000000000000154000000000000014900000000",
            INIT_60 => X"000000ce00000000000000f400000000000000f3000000000000012a00000000",
            INIT_61 => X"0000000a000000000000010d00000000000000dc00000000000000cd00000000",
            INIT_62 => X"0000002f00000000000000200000000000000027000000000000003700000000",
            INIT_63 => X"00000087000000000000007d000000000000006f000000000000004f00000000",
            INIT_64 => X"000000b80000000000000080000000000000006c000000000000007200000000",
            INIT_65 => X"0000001a0000000000000000000000000000010400000000000000d700000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000002c00000000",
            INIT_67 => X"00000071000000000000006a0000000000000079000000000000008e00000000",
            INIT_68 => X"000000e800000000000000d100000000000000c4000000000000009e00000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000012400000000",
            INIT_6A => X"0000009100000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000008800000000000000a200000000000000ba00000000000000ca00000000",
            INIT_6C => X"00000164000000000000010900000000000000be000000000000009d00000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000003a00000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"000000cb000000000000007c0000000000000033000000000000000700000000",
            INIT_70 => X"000000140000000000000181000000000000012300000000000000f400000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000004000000000000000250000000000000000000000000000000000000000",
            INIT_73 => X"0000010e00000000000000eb00000000000000df00000000000000ae00000000",
            INIT_74 => X"0000007a00000000000000780000000000000193000000000000014500000000",
            INIT_75 => X"0000007b000000000000007b000000000000007a000000000000007a00000000",
            INIT_76 => X"0000007a000000000000007a000000000000007b000000000000007b00000000",
            INIT_77 => X"0000007a000000000000007a000000000000007a000000000000007d00000000",
            INIT_78 => X"0000007c000000000000007c000000000000007a000000000000007c00000000",
            INIT_79 => X"0000007c000000000000007b000000000000007c000000000000007b00000000",
            INIT_7A => X"0000008d000000000000006e0000000000000078000000000000007a00000000",
            INIT_7B => X"0000007d000000000000007b000000000000007b000000000000008700000000",
            INIT_7C => X"0000007b000000000000007d000000000000007e000000000000007d00000000",
            INIT_7D => X"00000073000000000000007f000000000000007b000000000000007d00000000",
            INIT_7E => X"000000950000000000000081000000000000005b000000000000007900000000",
            INIT_7F => X"0000007e000000000000007e000000000000007d000000000000007c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE7;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE8 : if BRAM_NAME = "samplegold_layersamples_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007f000000000000007d000000000000007f000000000000007900000000",
            INIT_01 => X"0000004b000000000000005a000000000000008a000000000000006d00000000",
            INIT_02 => X"0000007c000000000000007f0000000000000037000000000000003a00000000",
            INIT_03 => X"0000009a0000000000000088000000000000007e000000000000007d00000000",
            INIT_04 => X"00000065000000000000007f0000000000000080000000000000009e00000000",
            INIT_05 => X"0000007400000000000000740000000000000070000000000000007700000000",
            INIT_06 => X"000000a400000000000000880000000000000080000000000000007a00000000",
            INIT_07 => X"0000007100000000000000340000000000000024000000000000008400000000",
            INIT_08 => X"000000a000000000000000850000000000000088000000000000007b00000000",
            INIT_09 => X"0000003f00000000000000670000000000000098000000000000009e00000000",
            INIT_0A => X"00000083000000000000006e0000000000000014000000000000002f00000000",
            INIT_0B => X"00000061000000000000008d000000000000009b000000000000007e00000000",
            INIT_0C => X"00000033000000000000001d0000000000000000000000000000004900000000",
            INIT_0D => X"0000008500000000000000860000000000000080000000000000007200000000",
            INIT_0E => X"0000002e000000000000009c0000000000000082000000000000008800000000",
            INIT_0F => X"000000670000000000000085000000000000002d000000000000002500000000",
            INIT_10 => X"00000072000000000000004f0000000000000032000000000000001600000000",
            INIT_11 => X"0000002b00000000000000260000000000000030000000000000005900000000",
            INIT_12 => X"0000005400000000000000550000000000000051000000000000003100000000",
            INIT_13 => X"00000078000000000000007a0000000000000054000000000000002a00000000",
            INIT_14 => X"00000058000000000000004b0000000000000052000000000000008c00000000",
            INIT_15 => X"00000071000000000000006b000000000000005b000000000000006200000000",
            INIT_16 => X"0000008a0000000000000081000000000000007b000000000000006100000000",
            INIT_17 => X"0000006100000000000000780000000000000086000000000000008b00000000",
            INIT_18 => X"0000004a0000000000000036000000000000005b000000000000004f00000000",
            INIT_19 => X"000000420000000000000030000000000000002d000000000000003100000000",
            INIT_1A => X"0000003b000000000000002a0000000000000028000000000000000d00000000",
            INIT_1B => X"000000610000000000000066000000000000005d000000000000004c00000000",
            INIT_1C => X"0000002b0000000000000031000000000000003f000000000000005000000000",
            INIT_1D => X"000000000000000000000035000000000000001f000000000000002a00000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000002600000000000000080000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000031000000000000002700000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000002b000000000000002e000000000000004a000000000000008100000000",
            INIT_24 => X"000000240000000000000014000000000000002d000000000000003300000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000004500000000",
            INIT_26 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"00000000000000000000000b0000000000000024000000000000003e00000000",
            INIT_28 => X"0000005500000000000000320000000000000018000000000000000900000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"00000015000000000000000f0000000000000000000000000000000000000000",
            INIT_2C => X"0000001400000000000000530000000000000034000000000000002300000000",
            INIT_2D => X"0000001400000000000000140000000000000014000000000000001400000000",
            INIT_2E => X"0000001200000000000000130000000000000014000000000000001300000000",
            INIT_2F => X"0000001300000000000000130000000000000016000000000000001400000000",
            INIT_30 => X"0000001400000000000000140000000000000013000000000000001400000000",
            INIT_31 => X"0000001400000000000000140000000000000013000000000000001400000000",
            INIT_32 => X"0000001000000000000000120000000000000013000000000000001400000000",
            INIT_33 => X"0000001400000000000000140000000000000017000000000000001a00000000",
            INIT_34 => X"0000001300000000000000140000000000000014000000000000001400000000",
            INIT_35 => X"0000001600000000000000120000000000000014000000000000001300000000",
            INIT_36 => X"000000180000000000000029000000000000001d000000000000000f00000000",
            INIT_37 => X"0000001400000000000000130000000000000014000000000000001a00000000",
            INIT_38 => X"0000001300000000000000130000000000000018000000000000001b00000000",
            INIT_39 => X"0000001c0000000000000015000000000000000b000000000000001400000000",
            INIT_3A => X"000000160000000000000029000000000000002a000000000000002700000000",
            INIT_3B => X"0000002600000000000000140000000000000014000000000000001600000000",
            INIT_3C => X"0000001300000000000000130000000000000017000000000000002800000000",
            INIT_3D => X"000000180000000000000017000000000000000d000000000000001700000000",
            INIT_3E => X"0000001d000000000000001c0000000000000018000000000000001b00000000",
            INIT_3F => X"00000023000000000000002b0000000000000015000000000000002500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001200000000000000100000000000000012000000000000000800000000",
            INIT_41 => X"0000001f000000000000001f0000000000000019000000000000001800000000",
            INIT_42 => X"0000001300000000000000240000000000000028000000000000002b00000000",
            INIT_43 => X"00000026000000000000002e000000000000002d000000000000001600000000",
            INIT_44 => X"00000035000000000000003d0000000000000010000000000000002800000000",
            INIT_45 => X"000000150000000000000013000000000000001e000000000000003400000000",
            INIT_46 => X"000000210000000000000014000000000000001d000000000000001900000000",
            INIT_47 => X"0000000e00000000000000200000000000000015000000000000003f00000000",
            INIT_48 => X"00000009000000000000001a000000000000002d000000000000002500000000",
            INIT_49 => X"000000300000000000000031000000000000002c000000000000001d00000000",
            INIT_4A => X"00000031000000000000001b000000000000002a000000000000002a00000000",
            INIT_4B => X"0000001800000000000000160000000000000025000000000000001900000000",
            INIT_4C => X"0000002b000000000000002f0000000000000018000000000000001800000000",
            INIT_4D => X"000000270000000000000026000000000000002d000000000000002800000000",
            INIT_4E => X"0000003b00000000000000110000000000000030000000000000002700000000",
            INIT_4F => X"0000004400000000000000440000000000000043000000000000003d00000000",
            INIT_50 => X"00000046000000000000003c0000000000000046000000000000004500000000",
            INIT_51 => X"00000033000000000000003b0000000000000045000000000000003b00000000",
            INIT_52 => X"00000033000000000000002e000000000000002a000000000000002b00000000",
            INIT_53 => X"0000004500000000000000370000000000000030000000000000003400000000",
            INIT_54 => X"0000004500000000000000480000000000000046000000000000004700000000",
            INIT_55 => X"0000001e00000000000000300000000000000042000000000000004200000000",
            INIT_56 => X"0000001c0000000000000021000000000000001a000000000000001c00000000",
            INIT_57 => X"0000003f00000000000000390000000000000022000000000000001b00000000",
            INIT_58 => X"0000002d000000000000003f0000000000000044000000000000004200000000",
            INIT_59 => X"0000000f0000000000000014000000000000001d000000000000001700000000",
            INIT_5A => X"0000001900000000000000180000000000000014000000000000001000000000",
            INIT_5B => X"0000001600000000000000220000000000000011000000000000001500000000",
            INIT_5C => X"0000001300000000000000140000000000000004000000000000000800000000",
            INIT_5D => X"000000120000000000000012000000000000000d000000000000000c00000000",
            INIT_5E => X"0000001400000000000000150000000000000016000000000000001300000000",
            INIT_5F => X"0000000b00000000000000000000000000000000000000000000001100000000",
            INIT_60 => X"0000000c00000000000000070000000000000000000000000000000c00000000",
            INIT_61 => X"0000000b00000000000000090000000000000014000000000000000d00000000",
            INIT_62 => X"0000000a00000000000000120000000000000011000000000000001000000000",
            INIT_63 => X"0000000000000000000000000000000000000010000000000000000a00000000",
            INIT_64 => X"0000000e000000000000000c0000000000000009000000000000000700000000",
            INIT_65 => X"0000002c000000000000002c000000000000002c000000000000002a00000000",
            INIT_66 => X"0000002c000000000000002c000000000000002c000000000000002c00000000",
            INIT_67 => X"0000002b0000000000000029000000000000002a000000000000002e00000000",
            INIT_68 => X"0000002a000000000000002c000000000000002c000000000000002c00000000",
            INIT_69 => X"0000002b000000000000002b000000000000002b000000000000002b00000000",
            INIT_6A => X"0000002a000000000000002b000000000000002c000000000000002b00000000",
            INIT_6B => X"0000002b000000000000002a0000000000000022000000000000001900000000",
            INIT_6C => X"0000002d000000000000002c000000000000002b000000000000002b00000000",
            INIT_6D => X"0000002c000000000000002c000000000000002b000000000000002c00000000",
            INIT_6E => X"0000000800000000000000170000000000000021000000000000002b00000000",
            INIT_6F => X"0000002c000000000000002b000000000000002f000000000000002900000000",
            INIT_70 => X"0000002900000000000000220000000000000020000000000000002b00000000",
            INIT_71 => X"0000002d0000000000000021000000000000002d000000000000002e00000000",
            INIT_72 => X"000000020000000000000004000000000000000b000000000000001900000000",
            INIT_73 => X"0000002900000000000000260000000000000023000000000000002800000000",
            INIT_74 => X"0000002f00000000000000280000000000000014000000000000000400000000",
            INIT_75 => X"0000002500000000000000300000000000000023000000000000002d00000000",
            INIT_76 => X"000000120000000000000017000000000000001c000000000000002500000000",
            INIT_77 => X"0000001100000000000000260000000000000027000000000000001400000000",
            INIT_78 => X"0000002c000000000000002c0000000000000034000000000000001800000000",
            INIT_79 => X"00000028000000000000002c000000000000002b000000000000002800000000",
            INIT_7A => X"00000001000000000000000b0000000000000003000000000000000f00000000",
            INIT_7B => X"0000001200000000000000010000000000000027000000000000002600000000",
            INIT_7C => X"000000000000000000000013000000000000001b000000000000001700000000",
            INIT_7D => X"0000002b000000000000001f0000000000000000000000000000000000000000",
            INIT_7E => X"0000002700000000000000280000000000000024000000000000002700000000",
            INIT_7F => X"00000013000000000000000a0000000000000009000000000000002500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE8;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE9 : if BRAM_NAME = "samplegold_layersamples_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001f00000000000000000000000000000016000000000000003200000000",
            INIT_01 => X"0000000000000000000000000000000000000014000000000000002000000000",
            INIT_02 => X"0000001600000000000000050000000000000001000000000000000000000000",
            INIT_03 => X"0000002e0000000000000015000000000000002a000000000000002d00000000",
            INIT_04 => X"00000005000000000000001e000000000000001b000000000000002a00000000",
            INIT_05 => X"0000000e000000000000000f0000000000000013000000000000001400000000",
            INIT_06 => X"000000300000000000000000000000000000000b000000000000000e00000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_0B => X"0000000200000000000000020000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000d00000000000000240000000000000004000000000000001a00000000",
            INIT_0F => X"00000000000000000000000f0000000000000009000000000000000900000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000002200000000000000210000000000000027000000000000001200000000",
            INIT_12 => X"00000010000000000000001f0000000000000010000000000000000800000000",
            INIT_13 => X"0000005a0000000000000065000000000000000e000000000000000b00000000",
            INIT_14 => X"00000033000000000000004c0000000000000060000000000000006500000000",
            INIT_15 => X"000000000000000000000027000000000000002a000000000000002400000000",
            INIT_16 => X"0000001000000000000000100000000000000016000000000000001000000000",
            INIT_17 => X"0000008d00000000000000a70000000000000051000000000000001100000000",
            INIT_18 => X"0000002800000000000000370000000000000037000000000000005000000000",
            INIT_19 => X"0000001300000000000000000000000000000027000000000000002500000000",
            INIT_1A => X"0000000e0000000000000010000000000000000e000000000000001000000000",
            INIT_1B => X"000000460000000000000036000000000000004e000000000000002700000000",
            INIT_1C => X"0000002500000000000000260000000000000023000000000000003600000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000002500000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"000000000000000000000007000000000000001c000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_2B => X"0000000000000000000000000000000000000020000000000000000000000000",
            INIT_2C => X"00000015000000000000001f000000000000001d000000000000000000000000",
            INIT_2D => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000100000000000000120000000000000011000000000000000900000000",
            INIT_30 => X"0000000100000000000000170000000000000000000000000000000000000000",
            INIT_31 => X"00000008000000000000000e0000000000000003000000000000000800000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000001900000000000000030000000000000021000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000011000000000000001700000000",
            INIT_35 => X"00000025000000000000001c0000000000000014000000000000000000000000",
            INIT_36 => X"0000000200000000000000010000000000000000000000000000000500000000",
            INIT_37 => X"00000024000000000000000d000000000000000d000000000000000a00000000",
            INIT_38 => X"000000000000000000000000000000000000002a000000000000001500000000",
            INIT_39 => X"0000000000000000000000090000000000000008000000000000000000000000",
            INIT_3A => X"00000004000000000000000c0000000000000004000000000000000000000000",
            INIT_3B => X"0000000000000000000000030000000000000047000000000000001600000000",
            INIT_3C => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000800000000000000100000000000000007000000000000000000000000",
            INIT_3F => X"0000000000000000000000070000000000000000000000000000003000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"00000000000000000000000b0000000000000000000000000000000500000000",
            INIT_42 => X"000000230000000000000010000000000000000d000000000000000900000000",
            INIT_43 => X"000000250000000000000020000000000000001c000000000000002200000000",
            INIT_44 => X"0000000b000000000000000c0000000000000010000000000000001c00000000",
            INIT_45 => X"0000000c000000000000000a0000000000000008000000000000000500000000",
            INIT_46 => X"0000003200000000000000100000000000000015000000000000000f00000000",
            INIT_47 => X"0000001f0000000000000019000000000000000c000000000000000300000000",
            INIT_48 => X"0000000400000000000000060000000000000000000000000000000400000000",
            INIT_49 => X"000000070000000000000007000000000000000c000000000000000700000000",
            INIT_4A => X"00000025000000000000002e0000000000000015000000000000001300000000",
            INIT_4B => X"000000630000000000000021000000000000001b000000000000001200000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000001c0000000000000015000000000000000a000000000000000100000000",
            INIT_4E => X"0000001c00000000000000220000000000000022000000000000000000000000",
            INIT_4F => X"00000000000000000000003b0000000000000022000000000000002100000000",
            INIT_50 => X"0000001d00000000000000050000000000000000000000000000000000000000",
            INIT_51 => X"00000000000000000000001b000000000000001b000000000000001500000000",
            INIT_52 => X"0000002200000000000000240000000000000024000000000000002100000000",
            INIT_53 => X"000000010000000000000005000000000000002e000000000000002100000000",
            INIT_54 => X"0000001a00000000000000160000000000000018000000000000002400000000",
            INIT_55 => X"00000090000000000000008f0000000000000019000000000000001900000000",
            INIT_56 => X"0000009100000000000000910000000000000090000000000000009000000000",
            INIT_57 => X"00000092000000000000008e0000000000000090000000000000009100000000",
            INIT_58 => X"0000009000000000000000900000000000000091000000000000009400000000",
            INIT_59 => X"0000009200000000000000920000000000000091000000000000009100000000",
            INIT_5A => X"0000009200000000000000920000000000000092000000000000009200000000",
            INIT_5B => X"0000009d00000000000000960000000000000092000000000000009000000000",
            INIT_5C => X"0000009300000000000000920000000000000091000000000000009700000000",
            INIT_5D => X"0000009200000000000000920000000000000090000000000000009100000000",
            INIT_5E => X"0000009700000000000000940000000000000092000000000000009100000000",
            INIT_5F => X"0000009c00000000000000980000000000000090000000000000009b00000000",
            INIT_60 => X"0000009b00000000000000940000000000000093000000000000009300000000",
            INIT_61 => X"0000009100000000000000920000000000000098000000000000009800000000",
            INIT_62 => X"00000085000000000000008b0000000000000095000000000000009200000000",
            INIT_63 => X"0000009d00000000000000a30000000000000083000000000000008700000000",
            INIT_64 => X"000000a900000000000000ad0000000000000099000000000000009900000000",
            INIT_65 => X"0000008c0000000000000092000000000000009000000000000000a800000000",
            INIT_66 => X"0000009d0000000000000095000000000000008e000000000000009100000000",
            INIT_67 => X"000000a300000000000000a500000000000000a800000000000000a400000000",
            INIT_68 => X"0000009b0000000000000071000000000000006a00000000000000a000000000",
            INIT_69 => X"0000009f00000000000000920000000000000099000000000000008800000000",
            INIT_6A => X"00000088000000000000009e000000000000009e000000000000009e00000000",
            INIT_6B => X"000000a10000000000000090000000000000006c000000000000007900000000",
            INIT_6C => X"0000007c000000000000009a000000000000009e000000000000009f00000000",
            INIT_6D => X"0000007d000000000000006f0000000000000056000000000000009000000000",
            INIT_6E => X"00000095000000000000009a000000000000009d000000000000009100000000",
            INIT_6F => X"0000004d000000000000009e000000000000009a000000000000009000000000",
            INIT_70 => X"00000090000000000000008b000000000000006c000000000000007000000000",
            INIT_71 => X"00000096000000000000008f0000000000000071000000000000006100000000",
            INIT_72 => X"00000071000000000000006d0000000000000079000000000000008900000000",
            INIT_73 => X"0000008b00000000000000590000000000000088000000000000007400000000",
            INIT_74 => X"0000009f00000000000000940000000000000075000000000000006000000000",
            INIT_75 => X"000000890000000000000082000000000000008300000000000000aa00000000",
            INIT_76 => X"0000009e00000000000000940000000000000091000000000000009200000000",
            INIT_77 => X"000000b000000000000000a00000000000000095000000000000009400000000",
            INIT_78 => X"000000a600000000000000ac00000000000000af00000000000000b000000000",
            INIT_79 => X"0000009100000000000000810000000000000099000000000000009600000000",
            INIT_7A => X"0000007500000000000000700000000000000074000000000000007d00000000",
            INIT_7B => X"000000680000000000000063000000000000005d000000000000004e00000000",
            INIT_7C => X"00000088000000000000008b0000000000000079000000000000006e00000000",
            INIT_7D => X"00000069000000000000006e0000000000000077000000000000008500000000",
            INIT_7E => X"0000000900000000000000610000000000000061000000000000006b00000000",
            INIT_7F => X"0000000300000000000000060000000000000014000000000000002500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE9;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE10 : if BRAM_NAME = "samplegold_layersamples_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000049000000000000003d0000000000000035000000000000000e00000000",
            INIT_01 => X"0000004600000000000000450000000000000042000000000000004500000000",
            INIT_02 => X"0000000b00000000000000000000000000000053000000000000004c00000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_04 => X"0000000000000000000000000000000000000008000000000000004c00000000",
            INIT_05 => X"00000048000000000000002a0000000000000027000000000000001400000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000006a00000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000007b00000000000000590000000000000044000000000000002700000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000004300000000000000310000000000000011000000000000000000000000",
            INIT_0D => X"0000000c000000000000007e0000000000000061000000000000004f00000000",
            INIT_0E => X"0000000b000000000000000b000000000000000b000000000000000b00000000",
            INIT_0F => X"0000000e000000000000000c000000000000000b000000000000000b00000000",
            INIT_10 => X"0000000c000000000000000a0000000000000007000000000000000a00000000",
            INIT_11 => X"0000000b000000000000000c000000000000000b000000000000000b00000000",
            INIT_12 => X"0000000b000000000000000b000000000000000b000000000000000b00000000",
            INIT_13 => X"00000002000000000000000a000000000000000c000000000000000b00000000",
            INIT_14 => X"0000000b000000000000000b0000000000000007000000000000000000000000",
            INIT_15 => X"0000000c000000000000000c000000000000000c000000000000000b00000000",
            INIT_16 => X"00000009000000000000000b000000000000000c000000000000000d00000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_18 => X"0000000b000000000000000c000000000000000b000000000000000000000000",
            INIT_19 => X"0000000d00000000000000080000000000000001000000000000000000000000",
            INIT_1A => X"00000010000000000000000a0000000000000009000000000000000b00000000",
            INIT_1B => X"0000000000000000000000000000000000000002000000000000000600000000",
            INIT_1C => X"0000000000000000000000090000000000000006000000000000000400000000",
            INIT_1D => X"0000000b000000000000000e0000000000000000000000000000000000000000",
            INIT_1E => X"00000004000000000000000b0000000000000006000000000000000d00000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_21 => X"000000020000000000000001000000000000000d000000000000000000000000",
            INIT_22 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000030000000000000005000000000000000800000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_25 => X"0000000000000000000000120000000000000000000000000000000300000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"00000006000000000000000f0000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000011000000000000000c00000000",
            INIT_2A => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"000000140000000000000014000000000000000e000000000000001900000000",
            INIT_38 => X"000000000000000000000000000000000000000f000000000000001500000000",
            INIT_39 => X"0000000400000000000000050000000000000000000000000000000000000000",
            INIT_3A => X"00000024000000000000000d000000000000000c000000000000000500000000",
            INIT_3B => X"0000001b000000000000001d0000000000000019000000000000001500000000",
            INIT_3C => X"000000440000000000000049000000000000000d000000000000001800000000",
            INIT_3D => X"0000001b00000000000000200000000000000021000000000000003700000000",
            INIT_3E => X"0000001b00000000000000280000000000000009000000000000001100000000",
            INIT_3F => X"00000019000000000000001a0000000000000018000000000000001700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002000000000000000310000000000000039000000000000001900000000",
            INIT_41 => X"0000001300000000000000190000000000000019000000000000002200000000",
            INIT_42 => X"000000210000000000000028000000000000002f000000000000000900000000",
            INIT_43 => X"00000013000000000000001d000000000000001f000000000000001f00000000",
            INIT_44 => X"00000021000000000000002a0000000000000028000000000000001c00000000",
            INIT_45 => X"0000000900000000000000120000000000000019000000000000001d00000000",
            INIT_46 => X"0000000200000000000000020000000000000002000000000000000000000000",
            INIT_47 => X"0000000000000000000000030000000000000003000000000000000300000000",
            INIT_48 => X"0000000300000000000000040000000000000000000000000000000300000000",
            INIT_49 => X"0000000000000000000000040000000000000002000000000000000200000000",
            INIT_4A => X"0000000400000000000000020000000000000003000000000000000300000000",
            INIT_4B => X"0000000000000000000000010000000000000005000000000000000200000000",
            INIT_4C => X"00000001000000000000001f000000000000003b000000000000000000000000",
            INIT_4D => X"0000000700000000000000050000000000000004000000000000000300000000",
            INIT_4E => X"0000000000000000000000050000000000000001000000000000000500000000",
            INIT_4F => X"0000000000000000000000010000000000000000000000000000000b00000000",
            INIT_50 => X"000000040000000000000001000000000000004a000000000000003f00000000",
            INIT_51 => X"000000070000000000000000000000000000000f000000000000000400000000",
            INIT_52 => X"0000003300000000000000000000000000000003000000000000000500000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000500000000000000030000000000000003000000000000003900000000",
            INIT_55 => X"0000000c0000000000000056000000000000005f000000000000003f00000000",
            INIT_56 => X"0000000000000000000000160000000000000000000000000000000500000000",
            INIT_57 => X"0000001600000000000000000000000000000000000000000000000500000000",
            INIT_58 => X"0000000000000000000000130000000000000073000000000000002500000000",
            INIT_59 => X"00000019000000000000000d000000000000000a000000000000000000000000",
            INIT_5A => X"0000004400000000000000400000000000000044000000000000000400000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"00000075000000000000003f0000000000000017000000000000004f00000000",
            INIT_5D => X"0000000000000000000000000000000000000025000000000000003d00000000",
            INIT_5E => X"00000004000000000000004e0000000000000038000000000000002800000000",
            INIT_5F => X"0000001c00000000000000250000000000000011000000000000000700000000",
            INIT_60 => X"00000002000000000000001c0000000000000069000000000000005b00000000",
            INIT_61 => X"000000000000000000000000000000000000000b000000000000006c00000000",
            INIT_62 => X"0000000000000000000000050000000000000019000000000000000000000000",
            INIT_63 => X"000000160000000000000000000000000000000b000000000000000000000000",
            INIT_64 => X"000000060000000000000000000000000000000000000000000000d600000000",
            INIT_65 => X"0000000000000000000000160000000000000000000000000000001600000000",
            INIT_66 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_67 => X"00000070000000000000001d000000000000002b000000000000002200000000",
            INIT_68 => X"000000350000000000000039000000000000003f000000000000003300000000",
            INIT_69 => X"00000015000000000000000e0000000000000007000000000000002600000000",
            INIT_6A => X"0000001100000000000000000000000000000014000000000000000000000000",
            INIT_6B => X"0000004100000000000000140000000000000028000000000000001a00000000",
            INIT_6C => X"0000005800000000000000490000000000000037000000000000001d00000000",
            INIT_6D => X"00000020000000000000002f0000000000000040000000000000004600000000",
            INIT_6E => X"0000000a000000000000002c0000000000000024000000000000001f00000000",
            INIT_6F => X"00000000000000000000004a0000000000000000000000000000002300000000",
            INIT_70 => X"0000004c000000000000001a0000000000000000000000000000000000000000",
            INIT_71 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"00000028000000000000000c000000000000000e000000000000000000000000",
            INIT_73 => X"0000000000000000000000240000000000000026000000000000000000000000",
            INIT_74 => X"0000001700000000000000e90000000000000009000000000000000000000000",
            INIT_75 => X"0000001e000000000000000f0000000000000000000000000000000600000000",
            INIT_76 => X"000000000000000000000033000000000000001d000000000000000d00000000",
            INIT_77 => X"000000030000000000000000000000000000000a000000000000000000000000",
            INIT_78 => X"000000000000000000000022000000000000007d000000000000000400000000",
            INIT_79 => X"0000000b00000000000000170000000000000009000000000000000e00000000",
            INIT_7A => X"0000000000000000000000000000000000000034000000000000002700000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"000000280000000000000004000000000000001b000000000000002b00000000",
            INIT_7D => X"0000001e00000000000000170000000000000007000000000000000700000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000002c00000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE10;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE11 : if BRAM_NAME = "samplegold_layersamples_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000260000000000000012000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000003a00000000000000020000000000000000000000000000000000000000",
            INIT_08 => X"00000000000000000000001d0000000000000028000000000000002000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000001c0000000000000084000000000000008a000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"00000000000000000000005b0000000000000073000000000000005e00000000",
            INIT_11 => X"0000002c00000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"00000081000000000000009a000000000000007c000000000000002a00000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000005300000000",
            INIT_14 => X"0000009c00000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"000000000000000000000000000000000000005300000000000000a500000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000006200000000000000670000000000000041000000000000000300000000",
            INIT_18 => X"00000000000000000000002c000000000000005f000000000000005f00000000",
            INIT_19 => X"0000000000000000000000000000000000000024000000000000000600000000",
            INIT_1A => X"00000032000000000000004e0000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000003000000000000000150000000000000000000000000000000000000000",
            INIT_1E => X"0000001500000000000000140000000000000000000000000000001900000000",
            INIT_1F => X"0000004800000000000000690000000000000054000000000000002800000000",
            INIT_20 => X"0000007a00000000000000810000000000000085000000000000003f00000000",
            INIT_21 => X"0000001a00000000000000330000000000000051000000000000006a00000000",
            INIT_22 => X"00000023000000000000002b0000000000000014000000000000002000000000",
            INIT_23 => X"00000052000000000000000a000000000000000d000000000000000a00000000",
            INIT_24 => X"00000096000000000000007f000000000000005c000000000000005400000000",
            INIT_25 => X"000000780000000000000093000000000000009c00000000000000a800000000",
            INIT_26 => X"000000030000000000000030000000000000004e000000000000006700000000",
            INIT_27 => X"0000002000000000000000110000000000000000000000000000000000000000",
            INIT_28 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000003b000000000000001b0000000000000000000000000000000000000000",
            INIT_2C => X"000000580000000000000008000000000000000d000000000000002700000000",
            INIT_2D => X"0000004600000000000000000000000000000000000000000000000d00000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000004100000000",
            INIT_2F => X"0000000c000000000000000c0000000000000002000000000000000000000000",
            INIT_30 => X"00000018000000000000000f0000000000000005000000000000000600000000",
            INIT_31 => X"0000000000000000000000000000000000000037000000000000005a00000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"00000000000000000000001b0000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000009900000000000000980000000000000000000000000000000000000000",
            INIT_37 => X"00000099000000000000009a0000000000000099000000000000009900000000",
            INIT_38 => X"00000097000000000000009a0000000000000099000000000000009900000000",
            INIT_39 => X"000000990000000000000099000000000000009b000000000000009500000000",
            INIT_3A => X"0000009900000000000000990000000000000098000000000000009a00000000",
            INIT_3B => X"0000009800000000000000980000000000000098000000000000009800000000",
            INIT_3C => X"0000007100000000000000690000000000000095000000000000009900000000",
            INIT_3D => X"0000009900000000000000980000000000000099000000000000009400000000",
            INIT_3E => X"0000009900000000000000990000000000000097000000000000009500000000",
            INIT_3F => X"0000008200000000000000950000000000000098000000000000009b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008b0000000000000072000000000000003e000000000000005600000000",
            INIT_41 => X"00000092000000000000009a0000000000000099000000000000009900000000",
            INIT_42 => X"0000009b000000000000009c000000000000009a000000000000009500000000",
            INIT_43 => X"000000760000000000000076000000000000008f000000000000008100000000",
            INIT_44 => X"0000009600000000000000a9000000000000007b000000000000007000000000",
            INIT_45 => X"0000002f0000000000000010000000000000009a000000000000009800000000",
            INIT_46 => X"0000008600000000000000970000000000000097000000000000008400000000",
            INIT_47 => X"000000840000000000000099000000000000009200000000000000a900000000",
            INIT_48 => X"0000006600000000000000350000000000000041000000000000006200000000",
            INIT_49 => X"000000a400000000000000a60000000000000091000000000000009800000000",
            INIT_4A => X"00000046000000000000004c0000000000000077000000000000007600000000",
            INIT_4B => X"00000076000000000000006f000000000000006c000000000000005500000000",
            INIT_4C => X"0000009800000000000000b00000000000000072000000000000008a00000000",
            INIT_4D => X"0000007a0000000000000043000000000000000f000000000000000000000000",
            INIT_4E => X"0000005000000000000000190000000000000000000000000000007100000000",
            INIT_4F => X"0000004a0000000000000066000000000000008900000000000000a100000000",
            INIT_50 => X"00000008000000000000005b000000000000004b000000000000004c00000000",
            INIT_51 => X"0000005f000000000000006c000000000000003c000000000000007300000000",
            INIT_52 => X"00000038000000000000007a00000000000000b4000000000000007d00000000",
            INIT_53 => X"00000058000000000000003c0000000000000026000000000000002400000000",
            INIT_54 => X"0000008600000000000000970000000000000086000000000000006b00000000",
            INIT_55 => X"00000078000000000000009700000000000000ad000000000000009800000000",
            INIT_56 => X"0000005a000000000000006d000000000000004e000000000000007000000000",
            INIT_57 => X"0000002300000000000000330000000000000045000000000000005400000000",
            INIT_58 => X"0000000800000000000000070000000000000056000000000000001d00000000",
            INIT_59 => X"0000000d0000000000000013000000000000000b000000000000000700000000",
            INIT_5A => X"0000000800000000000000070000000000000019000000000000001400000000",
            INIT_5B => X"0000003700000000000000230000000000000010000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"00000000000000000000004b0000000000000032000000000000000700000000",
            INIT_60 => X"000000000000000000000000000000000000000f000000000000001500000000",
            INIT_61 => X"00000007000000000000001c0000000000000018000000000000000000000000",
            INIT_62 => X"0000004c00000000000000530000000000000030000000000000000e00000000",
            INIT_63 => X"0000000000000000000000000000000000000064000000000000003800000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000005400000000000000650000000000000052000000000000005a00000000",
            INIT_66 => X"00000064000000000000004a0000000000000018000000000000002b00000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000007d00000000",
            INIT_68 => X"0000004900000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"000000580000000000000027000000000000003b000000000000007700000000",
            INIT_6A => X"0000007800000000000000660000000000000058000000000000007300000000",
            INIT_6B => X"000000000000000000000004000000000000000b000000000000000000000000",
            INIT_6C => X"0000003800000000000000250000000000000001000000000000000100000000",
            INIT_6D => X"000000520000000000000066000000000000007f000000000000004f00000000",
            INIT_6E => X"0000004700000000000000800000000000000070000000000000006200000000",
            INIT_6F => X"0000004200000000000000430000000000000043000000000000004300000000",
            INIT_70 => X"0000004300000000000000450000000000000043000000000000004300000000",
            INIT_71 => X"0000004300000000000000420000000000000041000000000000004300000000",
            INIT_72 => X"0000004300000000000000470000000000000041000000000000004300000000",
            INIT_73 => X"0000004300000000000000420000000000000043000000000000004300000000",
            INIT_74 => X"0000006700000000000000430000000000000044000000000000004100000000",
            INIT_75 => X"000000420000000000000044000000000000002a000000000000002300000000",
            INIT_76 => X"0000004200000000000000440000000000000048000000000000004100000000",
            INIT_77 => X"0000004000000000000000460000000000000041000000000000004400000000",
            INIT_78 => X"0000001000000000000000580000000000000052000000000000005900000000",
            INIT_79 => X"0000004200000000000000430000000000000044000000000000001a00000000",
            INIT_7A => X"00000043000000000000003c000000000000003d000000000000002e00000000",
            INIT_7B => X"0000006500000000000000200000000000000063000000000000004400000000",
            INIT_7C => X"000000000000000000000021000000000000003f000000000000003a00000000",
            INIT_7D => X"0000002f0000000000000040000000000000003f000000000000004000000000",
            INIT_7E => X"0000004200000000000000430000000000000008000000000000001600000000",
            INIT_7F => X"0000003700000000000000490000000000000020000000000000005800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE11;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE12 : if BRAM_NAME = "samplegold_layersamples_instance12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004900000000000000590000000000000060000000000000004f00000000",
            INIT_01 => X"0000001a000000000000002d0000000000000038000000000000000900000000",
            INIT_02 => X"0000006d00000000000000390000000000000049000000000000002500000000",
            INIT_03 => X"00000058000000000000003c0000000000000047000000000000004800000000",
            INIT_04 => X"00000000000000000000004b000000000000002e000000000000003c00000000",
            INIT_05 => X"0000001e00000000000000150000000000000035000000000000003200000000",
            INIT_06 => X"0000000000000000000000840000000000000057000000000000002000000000",
            INIT_07 => X"0000005f00000000000000460000000000000000000000000000000000000000",
            INIT_08 => X"0000001d0000000000000054000000000000004e000000000000006500000000",
            INIT_09 => X"0000000000000000000000310000000000000000000000000000000000000000",
            INIT_0A => X"0000005700000000000000060000000000000040000000000000003200000000",
            INIT_0B => X"0000000c000000000000002f000000000000003d000000000000004300000000",
            INIT_0C => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_0D => X"0000002b00000000000000150000000000000021000000000000003200000000",
            INIT_0E => X"00000036000000000000006f000000000000003b000000000000005000000000",
            INIT_0F => X"000000430000000000000053000000000000003c000000000000004700000000",
            INIT_10 => X"000000450000000000000000000000000000003a000000000000004100000000",
            INIT_11 => X"0000003300000000000000360000000000000038000000000000003400000000",
            INIT_12 => X"0000003c0000000000000021000000000000002a000000000000003f00000000",
            INIT_13 => X"0000001500000000000000130000000000000036000000000000002500000000",
            INIT_14 => X"0000001d00000000000000000000000000000019000000000000000e00000000",
            INIT_15 => X"00000028000000000000001c000000000000001a000000000000001c00000000",
            INIT_16 => X"0000002100000000000000320000000000000030000000000000002a00000000",
            INIT_17 => X"0000000600000000000000090000000000000000000000000000001200000000",
            INIT_18 => X"0000002000000000000000280000000000000000000000000000001f00000000",
            INIT_19 => X"0000000c00000000000000000000000000000000000000000000000700000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000002200000000000000000000000000000022000000000000002700000000",
            INIT_1C => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_1D => X"00000063000000000000006c0000000000000000000000000000000000000000",
            INIT_1E => X"000000000000000000000022000000000000004f000000000000005f00000000",
            INIT_1F => X"0000000000000000000000630000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"000000010000000000000037000000000000000f000000000000000000000000",
            INIT_22 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_23 => X"000000000000000000000000000000000000005f000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000300000000000000040000000000000005000000000000001200000000",
            INIT_27 => X"000000ac00000000000000ac00000000000000ac00000000000000b100000000",
            INIT_28 => X"000000af00000000000000ad00000000000000ad00000000000000ab00000000",
            INIT_29 => X"000000ad00000000000000ab00000000000000ad00000000000000ab00000000",
            INIT_2A => X"000000b100000000000000ac00000000000000ac00000000000000ad00000000",
            INIT_2B => X"000000ad00000000000000ae00000000000000ad00000000000000ad00000000",
            INIT_2C => X"000000af00000000000000af00000000000000ac00000000000000ad00000000",
            INIT_2D => X"000000ae0000000000000099000000000000008900000000000000ca00000000",
            INIT_2E => X"000000ac00000000000000af00000000000000ad00000000000000ad00000000",
            INIT_2F => X"000000b100000000000000ab00000000000000af00000000000000ad00000000",
            INIT_30 => X"000000b100000000000000ad00000000000000bf00000000000000a800000000",
            INIT_31 => X"000000ad00000000000000b1000000000000007c000000000000005c00000000",
            INIT_32 => X"000000ab00000000000000ab000000000000009e00000000000000ae00000000",
            INIT_33 => X"0000008800000000000000d000000000000000af00000000000000ae00000000",
            INIT_34 => X"0000007b0000000000000095000000000000009200000000000000ca00000000",
            INIT_35 => X"000000ae00000000000000ad00000000000000b0000000000000005000000000",
            INIT_36 => X"000000ac000000000000007d0000000000000068000000000000007d00000000",
            INIT_37 => X"000000b5000000000000008700000000000000c600000000000000ad00000000",
            INIT_38 => X"000000a600000000000000b300000000000000b3000000000000009b00000000",
            INIT_39 => X"0000007400000000000000a80000000000000063000000000000009800000000",
            INIT_3A => X"0000009d00000000000000a2000000000000007f000000000000006300000000",
            INIT_3B => X"0000008f0000000000000092000000000000008e00000000000000b000000000",
            INIT_3C => X"0000009c000000000000008700000000000000a000000000000000c100000000",
            INIT_3D => X"000000530000000000000070000000000000009c000000000000002c00000000",
            INIT_3E => X"000000b500000000000000b5000000000000007a000000000000007c00000000",
            INIT_3F => X"000000a2000000000000002a0000000000000020000000000000002a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000096000000000000009800000000000000ac00000000000000ae00000000",
            INIT_41 => X"0000006400000000000000210000000000000000000000000000006f00000000",
            INIT_42 => X"00000057000000000000009c0000000000000096000000000000002f00000000",
            INIT_43 => X"0000008300000000000000950000000000000091000000000000009b00000000",
            INIT_44 => X"0000004e000000000000005b000000000000004a000000000000006000000000",
            INIT_45 => X"0000006800000000000000770000000000000085000000000000000000000000",
            INIT_46 => X"000000c4000000000000009d00000000000000b0000000000000008000000000",
            INIT_47 => X"0000008a000000000000007c000000000000007b000000000000007400000000",
            INIT_48 => X"0000000000000000000000810000000000000079000000000000007700000000",
            INIT_49 => X"000000750000000000000076000000000000006a000000000000007800000000",
            INIT_4A => X"00000064000000000000006c0000000000000084000000000000007b00000000",
            INIT_4B => X"0000003f00000000000000640000000000000054000000000000007300000000",
            INIT_4C => X"0000001000000000000000280000000000000041000000000000004200000000",
            INIT_4D => X"0000002300000000000000230000000000000026000000000000002f00000000",
            INIT_4E => X"000000480000000000000048000000000000003e000000000000003600000000",
            INIT_4F => X"0000003a0000000000000023000000000000002d000000000000003900000000",
            INIT_50 => X"0000003400000000000000000000000000000025000000000000003700000000",
            INIT_51 => X"0000000000000000000000000000000000000003000000000000002000000000",
            INIT_52 => X"0000000a000000000000000e0000000000000011000000000000002800000000",
            INIT_53 => X"00000036000000000000004f000000000000003d000000000000001800000000",
            INIT_54 => X"0000001b00000000000000030000000000000000000000000000002900000000",
            INIT_55 => X"0000007e00000000000000000000000000000000000000000000000100000000",
            INIT_56 => X"0000004c000000000000005a0000000000000061000000000000005f00000000",
            INIT_57 => X"0000007f00000000000000390000000000000031000000000000003800000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000004d000000000000003a0000000000000000000000000000000000000000",
            INIT_5A => X"0000004500000000000000170000000000000010000000000000002700000000",
            INIT_5B => X"000000050000000000000081000000000000004a000000000000003b00000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000010000000000000004000000000000000000000000",
            INIT_5E => X"000000470000000000000044000000000000004d000000000000003b00000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000005300000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE12;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE13 : if BRAM_NAME = "samplegold_layersamples_instance13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000003b00000000000000130000000000000000000000000000000000000000",
            INIT_12 => X"000000000000000000000000000000000000001f000000000000003100000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000400000000000000160000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000002a00000000000000410000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000370000000000000027000000000000000700000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000003f00000000000000400000000000000003000000000000000e00000000",
            INIT_2C => X"0000000000000000000000000000000000000004000000000000002c00000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000100000000000000046000000000000005700000000",
            INIT_2F => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_30 => X"00000036000000000000001a0000000000000000000000000000000000000000",
            INIT_31 => X"00000000000000000000000f0000000000000030000000000000002000000000",
            INIT_32 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_33 => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000002c000000000000001a0000000000000002000000000000000000000000",
            INIT_39 => X"00000036000000000000003c000000000000000f000000000000001300000000",
            INIT_3A => X"0000000800000000000000140000000000000027000000000000003200000000",
            INIT_3B => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_3D => X"0000005e000000000000004a0000000000000034000000000000004400000000",
            INIT_3E => X"00000053000000000000005b0000000000000065000000000000006700000000",
            INIT_3F => X"000000110000000000000027000000000000003e000000000000004300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000001100000000000000040000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_43 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000002000000000000000080000000000000000000000000000000600000000",
            INIT_45 => X"000000130000000000000017000000000000002e000000000000003800000000",
            INIT_46 => X"0000005b00000000000000510000000000000056000000000000003100000000",
            INIT_47 => X"0000000000000000000000000000000000000040000000000000007400000000",
            INIT_48 => X"00000015000000000000000e0000000000000009000000000000000000000000",
            INIT_49 => X"00000039000000000000000f0000000000000010000000000000001600000000",
            INIT_4A => X"00000000000000000000004800000000000000ad000000000000009700000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_4D => X"00000027000000000000000c0000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"000000170000000000000004000000000000000b000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000002000000000000000c00000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000001d000000000000001e000000000000001d000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_63 => X"000000430000000000000012000000000000000d000000000000000000000000",
            INIT_64 => X"000000000000000000000024000000000000004b000000000000005800000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"00000013000000000000001d000000000000002b000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000002b00000000000000070000000000000000000000000000000000000000",
            INIT_69 => X"0000001a000000000000002a0000000000000036000000000000003800000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000001300000000000000090000000000000000000000000000000000000000",
            INIT_6F => X"0000001a0000000000000024000000000000001c000000000000001100000000",
            INIT_70 => X"0000003c00000000000000370000000000000031000000000000002f00000000",
            INIT_71 => X"0000003300000000000000370000000000000000000000000000002200000000",
            INIT_72 => X"0000000b000000000000001a0000000000000026000000000000002600000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"000000300000000000000024000000000000001d000000000000001000000000",
            INIT_77 => X"00000015000000000000001f0000000000000029000000000000003600000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_79 => X"0000000000000000000000000000000000000007000000000000000400000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_7D => X"0000000000000000000000000000000000000005000000000000000200000000",
            INIT_7E => X"0000000000000000000000030000000000000017000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000021000000000000001000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE13;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE14 : if BRAM_NAME = "samplegold_layersamples_instance14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"000000110000000000000045000000000000003b000000000000001e00000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000004100000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000024000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000002700000000000000000000000000000000000000000000000100000000",
            INIT_1B => X"00000022000000000000000a0000000000000000000000000000000700000000",
            INIT_1C => X"0000000000000000000000000000000000000005000000000000000500000000",
            INIT_1D => X"00000000000000000000003a0000000000000031000000000000000000000000",
            INIT_1E => X"00000000000000000000000b0000000000000000000000000000003700000000",
            INIT_1F => X"0000000000000000000000160000000000000024000000000000000000000000",
            INIT_20 => X"00000017000000000000001b0000000000000002000000000000000a00000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000003700000000",
            INIT_22 => X"0000002800000000000000120000000000000003000000000000000000000000",
            INIT_23 => X"000000000000000000000000000000000000000e000000000000002300000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000004b00000000000000000000000000000000000000000000000700000000",
            INIT_26 => X"0000000800000000000000140000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000290000000000000000000000000000000400000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000003000000000000003800000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"00000000000000000000001f0000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000035000000000000000000000000",
            INIT_32 => X"00000000000000000000002e000000000000000a000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000200000000000000060000000000000006000000000000000400000000",
            INIT_3E => X"00000000000000000000001f0000000000000000000000000000000000000000",
            INIT_3F => X"0000000300000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000001ef000000000000018d00000000000001a2000000000000000000000000",
            INIT_41 => X"0000021700000000000001ff000000000000020900000000000001f400000000",
            INIT_42 => X"0000020f00000000000002250000000000000216000000000000021100000000",
            INIT_43 => X"0000021d00000000000002280000000000000216000000000000022800000000",
            INIT_44 => X"000001e800000000000001f2000000000000018c00000000000001aa00000000",
            INIT_45 => X"0000020f00000000000001fc00000000000001ec000000000000020900000000",
            INIT_46 => X"0000022500000000000001c400000000000001d6000000000000020e00000000",
            INIT_47 => X"000001a7000000000000021b0000000000000224000000000000021200000000",
            INIT_48 => X"000001fb00000000000001df00000000000001e1000000000000017700000000",
            INIT_49 => X"000001da00000000000001bf00000000000001d700000000000001dc00000000",
            INIT_4A => X"000001f500000000000001f90000000000000180000000000000017300000000",
            INIT_4B => X"0000014e000000000000017f000000000000020a000000000000020200000000",
            INIT_4C => X"000001c300000000000001c700000000000001b8000000000000019f00000000",
            INIT_4D => X"000000dd0000000000000123000000000000018200000000000001ba00000000",
            INIT_4E => X"000001ad000000000000016900000000000000d400000000000000da00000000",
            INIT_4F => X"000000e600000000000000ca00000000000000d800000000000001ab00000000",
            INIT_50 => X"0000013000000000000001220000000000000112000000000000010000000000",
            INIT_51 => X"000000c300000000000000cb00000000000000da000000000000012100000000",
            INIT_52 => X"000000e90000000000000135000000000000011700000000000000d300000000",
            INIT_53 => X"000000cd00000000000000ca00000000000000bd00000000000000b300000000",
            INIT_54 => X"000000e8000000000000010b00000000000000f5000000000000010600000000",
            INIT_55 => X"0000017e000000000000010b00000000000000db00000000000000d900000000",
            INIT_56 => X"000000d000000000000000b10000000000000155000000000000011a00000000",
            INIT_57 => X"0000012a00000000000000e000000000000000aa00000000000000b200000000",
            INIT_58 => X"0000012900000000000001240000000000000136000000000000012d00000000",
            INIT_59 => X"0000015b000000000000018f000000000000015f000000000000012f00000000",
            INIT_5A => X"0000010c00000000000000fd000000000000006a00000000000000ff00000000",
            INIT_5B => X"00000189000000000000017a0000000000000155000000000000012700000000",
            INIT_5C => X"000001230000000000000166000000000000016a000000000000018a00000000",
            INIT_5D => X"000000d700000000000001580000000000000157000000000000012600000000",
            INIT_5E => X"0000012f00000000000000fc00000000000000f900000000000000dc00000000",
            INIT_5F => X"0000015d00000000000001630000000000000170000000000000017300000000",
            INIT_60 => X"00000148000000000000013d0000000000000152000000000000015300000000",
            INIT_61 => X"0000012f0000000000000122000000000000014d000000000000015600000000",
            INIT_62 => X"000001430000000000000148000000000000011100000000000000e900000000",
            INIT_63 => X"0000013b000000000000015d000000000000015a000000000000014b00000000",
            INIT_64 => X"0000013c000000000000015d0000000000000160000000000000012f00000000",
            INIT_65 => X"00000127000000000000009d00000000000000bd000000000000010100000000",
            INIT_66 => X"0000010f000000000000010b000000000000012f000000000000013700000000",
            INIT_67 => X"000000d100000000000000b50000000000000122000000000000014700000000",
            INIT_68 => X"0000008e00000000000000cb00000000000000fe000000000000011f00000000",
            INIT_69 => X"0000011f0000000000000109000000000000004f000000000000006b00000000",
            INIT_6A => X"0000010e00000000000000c800000000000000b700000000000000fb00000000",
            INIT_6B => X"000000b700000000000000b700000000000000af00000000000000ea00000000",
            INIT_6C => X"0000003700000000000000520000000000000079000000000000008c00000000",
            INIT_6D => X"000000b200000000000000cb00000000000000c6000000000000001500000000",
            INIT_6E => X"0000008700000000000000970000000000000097000000000000009300000000",
            INIT_6F => X"0000005000000000000000710000000000000075000000000000008500000000",
            INIT_70 => X"00000014000000000000001c0000000000000032000000000000005000000000",
            INIT_71 => X"0000004400000000000000380000000000000032000000000000003400000000",
            INIT_72 => X"0000004e00000000000000570000000000000051000000000000004f00000000",
            INIT_73 => X"0000002300000000000000360000000000000055000000000000006800000000",
            INIT_74 => X"0000000f0000000000000017000000000000001a000000000000001700000000",
            INIT_75 => X"00000039000000000000002e0000000000000023000000000000001400000000",
            INIT_76 => X"0000005e000000000000002c0000000000000041000000000000003f00000000",
            INIT_77 => X"000000120000000000000010000000000000001c000000000000003300000000",
            INIT_78 => X"0000006300000000000000530000000000000000000000000000001f00000000",
            INIT_79 => X"0000007e0000000000000083000000000000007d000000000000007f00000000",
            INIT_7A => X"0000008b00000000000000860000000000000076000000000000008300000000",
            INIT_7B => X"0000008100000000000000790000000000000085000000000000008000000000",
            INIT_7C => X"0000008400000000000000610000000000000055000000000000008300000000",
            INIT_7D => X"0000008200000000000000750000000000000080000000000000007300000000",
            INIT_7E => X"0000008c00000000000000690000000000000082000000000000008300000000",
            INIT_7F => X"000000870000000000000087000000000000007a000000000000008e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE14;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE15 : if BRAM_NAME = "samplegold_layersamples_instance15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000068000000000000007d000000000000005c000000000000005300000000",
            INIT_01 => X"00000083000000000000006b000000000000006b000000000000007600000000",
            INIT_02 => X"0000009900000000000000900000000000000031000000000000008a00000000",
            INIT_03 => X"00000053000000000000008a0000000000000082000000000000007600000000",
            INIT_04 => X"0000006e000000000000007a0000000000000077000000000000005300000000",
            INIT_05 => X"000000490000000000000046000000000000005d000000000000006d00000000",
            INIT_06 => X"000000a6000000000000006a000000000000003e000000000000003b00000000",
            INIT_07 => X"0000004300000000000000540000000000000084000000000000007d00000000",
            INIT_08 => X"0000006e0000000000000068000000000000006b000000000000005200000000",
            INIT_09 => X"0000001b0000000000000024000000000000004b000000000000006500000000",
            INIT_0A => X"0000003400000000000000350000000000000012000000000000002200000000",
            INIT_0B => X"0000000800000000000000100000000000000013000000000000004900000000",
            INIT_0C => X"00000031000000000000001a0000000000000017000000000000001400000000",
            INIT_0D => X"000000230000000000000011000000000000001d000000000000002400000000",
            INIT_0E => X"00000000000000000000004c0000000000000000000000000000002b00000000",
            INIT_0F => X"0000003000000000000000160000000000000013000000000000002600000000",
            INIT_10 => X"00000016000000000000002f000000000000002a000000000000004900000000",
            INIT_11 => X"000000610000000000000048000000000000001c000000000000000f00000000",
            INIT_12 => X"0000001f0000000000000000000000000000003e000000000000002d00000000",
            INIT_13 => X"000000490000000000000032000000000000001d000000000000001200000000",
            INIT_14 => X"0000005c000000000000004d0000000000000051000000000000004f00000000",
            INIT_15 => X"0000004400000000000000570000000000000059000000000000003900000000",
            INIT_16 => X"0000004800000000000000450000000000000000000000000000000000000000",
            INIT_17 => X"0000006400000000000000650000000000000069000000000000006400000000",
            INIT_18 => X"0000001600000000000000450000000000000041000000000000005800000000",
            INIT_19 => X"000000310000000000000042000000000000003e000000000000002e00000000",
            INIT_1A => X"0000004600000000000000330000000000000019000000000000004a00000000",
            INIT_1B => X"000000450000000000000040000000000000004a000000000000005200000000",
            INIT_1C => X"0000004b000000000000004e0000000000000050000000000000004b00000000",
            INIT_1D => X"00000024000000000000002a000000000000003d000000000000004500000000",
            INIT_1E => X"0000004100000000000000480000000000000043000000000000004c00000000",
            INIT_1F => X"000000180000000000000030000000000000005f000000000000005c00000000",
            INIT_20 => X"0000002e00000000000000460000000000000054000000000000003700000000",
            INIT_21 => X"0000005400000000000000000000000000000000000000000000000f00000000",
            INIT_22 => X"00000019000000000000001c0000000000000027000000000000004400000000",
            INIT_23 => X"0000001b00000000000000110000000000000034000000000000005100000000",
            INIT_24 => X"000000000000000000000001000000000000000f000000000000001e00000000",
            INIT_25 => X"0000003f00000000000000420000000000000000000000000000000000000000",
            INIT_26 => X"0000002600000000000000240000000000000021000000000000003300000000",
            INIT_27 => X"00000009000000000000000d000000000000000a000000000000001200000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000060000000000000006000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_30 => X"0000003900000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000002a00000000000000300000000000000031000000000000003c00000000",
            INIT_32 => X"000000180000000000000019000000000000001d000000000000002700000000",
            INIT_33 => X"0000001c00000000000000160000000000000019000000000000001800000000",
            INIT_34 => X"00000031000000000000002d000000000000001c000000000000001500000000",
            INIT_35 => X"0000001a00000000000000180000000000000022000000000000002300000000",
            INIT_36 => X"0000000b00000000000000170000000000000015000000000000001400000000",
            INIT_37 => X"0000001000000000000000180000000000000014000000000000002700000000",
            INIT_38 => X"00000018000000000000002a0000000000000022000000000000001900000000",
            INIT_39 => X"0000000a00000000000000120000000000000007000000000000001600000000",
            INIT_3A => X"0000001a00000000000000150000000000000016000000000000000f00000000",
            INIT_3B => X"0000000f00000000000000090000000000000011000000000000001500000000",
            INIT_3C => X"0000000e000000000000000a0000000000000026000000000000001900000000",
            INIT_3D => X"00000008000000000000000b000000000000000a000000000000000200000000",
            INIT_3E => X"0000001f00000000000000240000000000000036000000000000001600000000",
            INIT_3F => X"0000002000000000000000080000000000000003000000000000001700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000110000000000000010000000000000001a000000000000001e00000000",
            INIT_41 => X"000000360000000000000022000000000000001d000000000000000f00000000",
            INIT_42 => X"0000000d00000000000000320000000000000030000000000000002d00000000",
            INIT_43 => X"0000002e000000000000002e000000000000000b000000000000000200000000",
            INIT_44 => X"0000002d0000000000000025000000000000002f000000000000002100000000",
            INIT_45 => X"0000002c000000000000002f0000000000000039000000000000003000000000",
            INIT_46 => X"0000000200000000000000060000000000000015000000000000003400000000",
            INIT_47 => X"000000350000000000000031000000000000002d000000000000001900000000",
            INIT_48 => X"0000003e000000000000003d0000000000000037000000000000003200000000",
            INIT_49 => X"0000001b000000000000002e0000000000000037000000000000004300000000",
            INIT_4A => X"0000002600000000000000030000000000000016000000000000000c00000000",
            INIT_4B => X"00000039000000000000003c000000000000003b000000000000004000000000",
            INIT_4C => X"0000003300000000000000390000000000000039000000000000003b00000000",
            INIT_4D => X"00000011000000000000001a000000000000001f000000000000003000000000",
            INIT_4E => X"0000003e000000000000001b0000000000000028000000000000001500000000",
            INIT_4F => X"0000003b000000000000003f0000000000000040000000000000003900000000",
            INIT_50 => X"0000002a00000000000000330000000000000035000000000000003900000000",
            INIT_51 => X"0000001d00000000000000160000000000000017000000000000002800000000",
            INIT_52 => X"0000003f000000000000004d000000000000000c000000000000001b00000000",
            INIT_53 => X"0000003600000000000000410000000000000038000000000000003600000000",
            INIT_54 => X"00000023000000000000002a0000000000000021000000000000002a00000000",
            INIT_55 => X"0000001b0000000000000017000000000000001a000000000000002100000000",
            INIT_56 => X"0000003b00000000000000400000000000000044000000000000001e00000000",
            INIT_57 => X"000000280000000000000034000000000000002d000000000000003700000000",
            INIT_58 => X"0000001e0000000000000019000000000000002d000000000000003500000000",
            INIT_59 => X"0000001600000000000000240000000000000021000000000000002400000000",
            INIT_5A => X"0000003f0000000000000034000000000000003c000000000000003100000000",
            INIT_5B => X"0000002c000000000000002c0000000000000026000000000000003900000000",
            INIT_5C => X"00000026000000000000001f0000000000000024000000000000002400000000",
            INIT_5D => X"0000002d00000000000000240000000000000021000000000000002400000000",
            INIT_5E => X"00000028000000000000002f0000000000000032000000000000002f00000000",
            INIT_5F => X"000000210000000000000024000000000000002e000000000000002900000000",
            INIT_60 => X"0000002400000000000000220000000000000027000000000000002500000000",
            INIT_61 => X"0000002a00000000000000260000000000000025000000000000002500000000",
            INIT_62 => X"0000002000000000000000200000000000000026000000000000002700000000",
            INIT_63 => X"0000001e000000000000002b0000000000000024000000000000002400000000",
            INIT_64 => X"0000002300000000000000260000000000000022000000000000002600000000",
            INIT_65 => X"0000001f000000000000001e000000000000001e000000000000002000000000",
            INIT_66 => X"0000002000000000000000210000000000000023000000000000002100000000",
            INIT_67 => X"00000021000000000000002b000000000000001d000000000000001f00000000",
            INIT_68 => X"0000001700000000000000230000000000000023000000000000002500000000",
            INIT_69 => X"0000000a00000000000000070000000000000000000000000000000000000000",
            INIT_6A => X"0000001f00000000000000220000000000000019000000000000001200000000",
            INIT_6B => X"0000002b00000000000000270000000000000027000000000000002700000000",
            INIT_6C => X"0000000000000000000000290000000000000026000000000000002300000000",
            INIT_6D => X"000000240000000000000017000000000000001b000000000000000a00000000",
            INIT_6E => X"0000002a00000000000000280000000000000028000000000000002200000000",
            INIT_6F => X"0000002700000000000000310000000000000027000000000000001500000000",
            INIT_70 => X"00000017000000000000000b000000000000002e000000000000002e00000000",
            INIT_71 => X"0000002800000000000000330000000000000025000000000000002a00000000",
            INIT_72 => X"0000000000000000000000320000000000000033000000000000002800000000",
            INIT_73 => X"0000003500000000000000280000000000000037000000000000002e00000000",
            INIT_74 => X"0000003a0000000000000022000000000000001c000000000000003600000000",
            INIT_75 => X"0000003300000000000000390000000000000040000000000000003d00000000",
            INIT_76 => X"0000000000000000000000000000000000000006000000000000001e00000000",
            INIT_77 => X"00000049000000000000003e0000000000000032000000000000000c00000000",
            INIT_78 => X"0000002a0000000000000019000000000000000f000000000000001400000000",
            INIT_79 => X"00000009000000000000001e000000000000002e000000000000002c00000000",
            INIT_7A => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000240000000000000024000000000000003400000000",
            INIT_7C => X"0000000000000000000000060000000000000001000000000000000400000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000d0000000000000022000000000000000c000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000010000000000000003900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE15;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE16 : if BRAM_NAME = "samplegold_layersamples_instance16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000004300000000000000210000000000000032000000000000001b00000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000002000000000000000020000000000000002000000000000000000000000",
            INIT_06 => X"0000000700000000000000000000000000000025000000000000002c00000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000002100000000000000200000000000000002000000000000000900000000",
            INIT_0A => X"0000000000000000000000360000000000000017000000000000001800000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000c000000000000000a0000000000000001000000000000000000000000",
            INIT_0D => X"0000001300000000000000150000000000000015000000000000001000000000",
            INIT_0E => X"0000000000000000000000000000000000000010000000000000000d00000000",
            INIT_0F => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_10 => X"0000001300000000000000050000000000000000000000000000000000000000",
            INIT_11 => X"0000000200000000000000000000000000000003000000000000000c00000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_13 => X"00000001000000000000000a0000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000300000000000000030000000000000002000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_20 => X"0000000100000000000000000000000000000000000000000000000100000000",
            INIT_21 => X"0000000300000000000000020000000000000000000000000000000300000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000090000000000000003000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_27 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"000000080000000000000000000000000000000b000000000000000200000000",
            INIT_2A => X"00000008000000000000000b0000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000070000000000000029000000000000000000000000",
            INIT_2C => X"0000000300000000000000000000000000000000000000000000000200000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_2E => X"0000000200000000000000040000000000000000000000000000000000000000",
            INIT_2F => X"0000000d00000000000000240000000000000036000000000000002600000000",
            INIT_30 => X"0000001a000000000000000e0000000000000011000000000000000b00000000",
            INIT_31 => X"0000000800000000000000140000000000000016000000000000002300000000",
            INIT_32 => X"0000000b00000000000000070000000000000000000000000000000100000000",
            INIT_33 => X"000000190000000000000016000000000000001e000000000000000d00000000",
            INIT_34 => X"0000000f00000000000000080000000000000011000000000000001800000000",
            INIT_35 => X"000000010000000000000005000000000000000a000000000000000700000000",
            INIT_36 => X"000000060000000000000016000000000000000b000000000000000d00000000",
            INIT_37 => X"0000001900000000000000000000000000000013000000000000000000000000",
            INIT_38 => X"000000130000000000000015000000000000000a000000000000000b00000000",
            INIT_39 => X"0000000500000000000000000000000000000002000000000000000000000000",
            INIT_3A => X"0000000000000000000000110000000000000020000000000000000d00000000",
            INIT_3B => X"0000000000000000000000020000000000000000000000000000001f00000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000700000000000000030000000000000001000000000000000000000000",
            INIT_3E => X"000000000000000000000000000000000000000d000000000000001d00000000",
            INIT_3F => X"0000001500000000000000060000000000000008000000000000000800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000a00000000000000010000000000000000000000000000000100000000",
            INIT_41 => X"000000130000000000000000000000000000000f000000000000000700000000",
            INIT_42 => X"0000001400000000000000000000000000000002000000000000000700000000",
            INIT_43 => X"0000000800000000000000050000000000000009000000000000000000000000",
            INIT_44 => X"0000000c000000000000000b0000000000000009000000000000000300000000",
            INIT_45 => X"000000020000000000000007000000000000000a000000000000000500000000",
            INIT_46 => X"000000080000000000000015000000000000000b000000000000000700000000",
            INIT_47 => X"0000001600000000000000010000000000000009000000000000000500000000",
            INIT_48 => X"0000002600000000000000050000000000000003000000000000000e00000000",
            INIT_49 => X"0000000f000000000000000d000000000000000b000000000000001900000000",
            INIT_4A => X"000000080000000000000028000000000000001a000000000000001200000000",
            INIT_4B => X"0000002b000000000000000d000000000000000a000000000000000300000000",
            INIT_4C => X"0000001800000000000000170000000000000001000000000000000000000000",
            INIT_4D => X"0000001900000000000000180000000000000015000000000000001500000000",
            INIT_4E => X"0000000b00000000000000100000000000000022000000000000001600000000",
            INIT_4F => X"0000000f000000000000001e000000000000001b000000000000000e00000000",
            INIT_50 => X"00000017000000000000001a0000000000000019000000000000001900000000",
            INIT_51 => X"00000017000000000000001a000000000000000f000000000000002000000000",
            INIT_52 => X"00000020000000000000001d000000000000001e000000000000002100000000",
            INIT_53 => X"00000020000000000000001d000000000000001f000000000000002000000000",
            INIT_54 => X"0000001800000000000000190000000000000018000000000000001700000000",
            INIT_55 => X"0000001b000000000000001e000000000000001c000000000000001700000000",
            INIT_56 => X"0000001e00000000000000210000000000000021000000000000001f00000000",
            INIT_57 => X"0000002700000000000000200000000000000020000000000000001e00000000",
            INIT_58 => X"0000001d0000000000000016000000000000001b000000000000000800000000",
            INIT_59 => X"0000009c00000000000000ab000000000000001a000000000000001d00000000",
            INIT_5A => X"000000a200000000000000b100000000000000b200000000000000b900000000",
            INIT_5B => X"000000a300000000000000a1000000000000009e00000000000000a200000000",
            INIT_5C => X"000000a00000000000000096000000000000009b000000000000009600000000",
            INIT_5D => X"000000aa000000000000008d00000000000000a3000000000000009500000000",
            INIT_5E => X"0000009a000000000000009300000000000000a3000000000000009c00000000",
            INIT_5F => X"0000008d000000000000009d0000000000000099000000000000009d00000000",
            INIT_60 => X"00000093000000000000009d0000000000000091000000000000009800000000",
            INIT_61 => X"000000870000000000000095000000000000007a000000000000009200000000",
            INIT_62 => X"00000090000000000000008e0000000000000084000000000000009100000000",
            INIT_63 => X"0000009a000000000000008c0000000000000084000000000000009100000000",
            INIT_64 => X"0000007a000000000000008e0000000000000091000000000000008e00000000",
            INIT_65 => X"0000007100000000000000710000000000000079000000000000006200000000",
            INIT_66 => X"0000007f00000000000000710000000000000076000000000000007300000000",
            INIT_67 => X"0000008a0000000000000087000000000000007e000000000000007b00000000",
            INIT_68 => X"0000005d000000000000006d0000000000000071000000000000007f00000000",
            INIT_69 => X"0000006c000000000000006b0000000000000070000000000000006d00000000",
            INIT_6A => X"0000006b0000000000000067000000000000007d000000000000007300000000",
            INIT_6B => X"000000670000000000000054000000000000004b000000000000006800000000",
            INIT_6C => X"0000005b0000000000000051000000000000005c000000000000005700000000",
            INIT_6D => X"0000007900000000000000630000000000000060000000000000005500000000",
            INIT_6E => X"0000005c0000000000000066000000000000006c000000000000007a00000000",
            INIT_6F => X"00000034000000000000005a0000000000000048000000000000005c00000000",
            INIT_70 => X"0000006f0000000000000062000000000000005f000000000000007300000000",
            INIT_71 => X"0000007a000000000000008c0000000000000081000000000000008b00000000",
            INIT_72 => X"0000007700000000000000750000000000000079000000000000007800000000",
            INIT_73 => X"0000007500000000000000260000000000000051000000000000005300000000",
            INIT_74 => X"0000009300000000000000810000000000000068000000000000006b00000000",
            INIT_75 => X"00000098000000000000009c00000000000000a1000000000000009c00000000",
            INIT_76 => X"0000005d00000000000000630000000000000072000000000000008300000000",
            INIT_77 => X"0000008c000000000000008e0000000000000032000000000000002d00000000",
            INIT_78 => X"000000ab00000000000000ab00000000000000a6000000000000009b00000000",
            INIT_79 => X"000000640000000000000081000000000000009200000000000000a800000000",
            INIT_7A => X"0000005a000000000000006c0000000000000066000000000000005e00000000",
            INIT_7B => X"00000093000000000000007e000000000000007f000000000000006400000000",
            INIT_7C => X"0000008e0000000000000093000000000000009a000000000000009f00000000",
            INIT_7D => X"0000007a0000000000000083000000000000007b000000000000008900000000",
            INIT_7E => X"00000050000000000000005c000000000000006a000000000000007300000000",
            INIT_7F => X"0000008a000000000000009a000000000000009c000000000000009a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE16;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE17 : if BRAM_NAME = "samplegold_layersamples_instance17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000006a000000000000008c0000000000000098000000000000009500000000",
            INIT_01 => X"0000006c00000000000000780000000000000081000000000000006c00000000",
            INIT_02 => X"00000097000000000000003d0000000000000044000000000000005300000000",
            INIT_03 => X"0000006f0000000000000075000000000000008f000000000000009500000000",
            INIT_04 => X"0000006100000000000000580000000000000076000000000000008b00000000",
            INIT_05 => X"0000004400000000000000540000000000000059000000000000006500000000",
            INIT_06 => X"00000080000000000000007d0000000000000029000000000000003a00000000",
            INIT_07 => X"0000006d000000000000006e0000000000000067000000000000007800000000",
            INIT_08 => X"0000005600000000000000560000000000000055000000000000005700000000",
            INIT_09 => X"0000002f00000000000000370000000000000042000000000000004400000000",
            INIT_0A => X"00000047000000000000004b000000000000004f000000000000002800000000",
            INIT_0B => X"0000004e00000000000000480000000000000047000000000000004700000000",
            INIT_0C => X"000000390000000000000043000000000000003e000000000000004a00000000",
            INIT_0D => X"0000002c000000000000002d000000000000002d000000000000003000000000",
            INIT_0E => X"0000003400000000000000310000000000000027000000000000002500000000",
            INIT_0F => X"00000038000000000000003f0000000000000039000000000000003700000000",
            INIT_10 => X"00000028000000000000002e0000000000000037000000000000004200000000",
            INIT_11 => X"00000000000000000000001f000000000000002d000000000000002c00000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000100000000000000020000000000000000000000000000000000000000",
            INIT_14 => X"0000000b000000000000000b000000000000000b000000000000000200000000",
            INIT_15 => X"000000000000000000000000000000000000000a000000000000000300000000",
            INIT_16 => X"0000000a00000000000000000000000000000002000000000000000000000000",
            INIT_17 => X"0000000000000000000000070000000000000003000000000000000400000000",
            INIT_18 => X"00000007000000000000000f0000000000000007000000000000000c00000000",
            INIT_19 => X"00000006000000000000000a0000000000000000000000000000000c00000000",
            INIT_1A => X"000000090000000000000012000000000000000e000000000000001300000000",
            INIT_1B => X"00000000000000000000000c000000000000000b000000000000000b00000000",
            INIT_1C => X"0000001000000000000000120000000000000010000000000000000200000000",
            INIT_1D => X"00000016000000000000000b0000000000000013000000000000000900000000",
            INIT_1E => X"0000000b0000000000000019000000000000001d000000000000001b00000000",
            INIT_1F => X"0000000600000000000000000000000000000002000000000000000000000000",
            INIT_20 => X"000000000000000000000022000000000000000e000000000000000500000000",
            INIT_21 => X"0000000900000000000000010000000000000001000000000000000200000000",
            INIT_22 => X"0000000000000000000000000000000000000004000000000000000800000000",
            INIT_23 => X"0000000a00000000000000070000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000010000000000000001000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000001300000000000000180000000000000006000000000000000100000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"000000240000000000000016000000000000001e000000000000001000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000001200000000000000070000000000000000000000000000000000000000",
            INIT_2F => X"000000000000000000000018000000000000001f000000000000001200000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000700000000000000060000000000000000000000000000000300000000",
            INIT_33 => X"000000000000000000000000000000000000000d000000000000000f00000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000900000000000000030000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_3A => X"0000000700000000000000080000000000000005000000000000000200000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"00000000000000000000000d0000000000000005000000000000000600000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000600000000000000040000000000000008000000000000000000000000",
            INIT_42 => X"0000000500000000000000020000000000000005000000000000000600000000",
            INIT_43 => X"0000000100000000000000000000000000000001000000000000000200000000",
            INIT_44 => X"0000000000000000000000070000000000000004000000000000000100000000",
            INIT_45 => X"0000000600000000000000070000000000000006000000000000000600000000",
            INIT_46 => X"00000008000000000000000a000000000000000b000000000000000700000000",
            INIT_47 => X"0000000100000000000000040000000000000006000000000000000800000000",
            INIT_48 => X"00000005000000000000000c0000000000000004000000000000000800000000",
            INIT_49 => X"0000000f00000000000000050000000000000005000000000000000700000000",
            INIT_4A => X"0000000a000000000000001f0000000000000029000000000000000000000000",
            INIT_4B => X"00000000000000000000000c000000000000000a000000000000000a00000000",
            INIT_4C => X"0000000f00000000000000040000000000000008000000000000001800000000",
            INIT_4D => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_4E => X"0000000d00000000000000000000000000000029000000000000002a00000000",
            INIT_4F => X"00000014000000000000000b000000000000000a000000000000000400000000",
            INIT_50 => X"0000000000000000000000210000000000000052000000000000000000000000",
            INIT_51 => X"000000280000000000000000000000000000001a000000000000000100000000",
            INIT_52 => X"0000000000000000000000090000000000000000000000000000002e00000000",
            INIT_53 => X"0000000000000000000000300000000000000020000000000000000000000000",
            INIT_54 => X"0000000d00000000000000000000000000000041000000000000008400000000",
            INIT_55 => X"00000025000000000000002a0000000000000000000000000000002200000000",
            INIT_56 => X"0000000000000000000000120000000000000006000000000000002600000000",
            INIT_57 => X"0000003800000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000003c0000000000000020000000000000008c000000000000005000000000",
            INIT_59 => X"0000004800000000000000230000000000000030000000000000002500000000",
            INIT_5A => X"00000000000000000000002b0000000000000039000000000000003200000000",
            INIT_5B => X"0000000c00000000000000150000000000000000000000000000000000000000",
            INIT_5C => X"0000001e000000000000002d0000000000000000000000000000003000000000",
            INIT_5D => X"00000000000000000000001e0000000000000000000000000000001600000000",
            INIT_5E => X"0000000400000000000000000000000000000009000000000000000000000000",
            INIT_5F => X"00000000000000000000000c0000000000000034000000000000000000000000",
            INIT_60 => X"0000000700000000000000180000000000000000000000000000002500000000",
            INIT_61 => X"0000000000000000000000250000000000000040000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"000000000000000000000000000000000000001d000000000000003900000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000007000000000000000600000000",
            INIT_66 => X"000000450000000000000000000000000000000e000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000002a00000000",
            INIT_68 => X"000000230000000000000041000000000000001a000000000000000900000000",
            INIT_69 => X"00000000000000000000000f000000000000000d000000000000000400000000",
            INIT_6A => X"0000000300000000000000170000000000000000000000000000000e00000000",
            INIT_6B => X"00000000000000000000000c0000000000000000000000000000000100000000",
            INIT_6C => X"0000000e00000000000000090000000000000013000000000000001c00000000",
            INIT_6D => X"0000002800000000000000000000000000000000000000000000000400000000",
            INIT_6E => X"000000000000000000000000000000000000000a000000000000001100000000",
            INIT_6F => X"00000006000000000000002f000000000000001a000000000000000000000000",
            INIT_70 => X"0000003900000000000000290000000000000000000000000000000500000000",
            INIT_71 => X"0000002100000000000000460000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_73 => X"0000000000000000000000110000000000000053000000000000000000000000",
            INIT_74 => X"00000000000000000000003d000000000000000b000000000000000100000000",
            INIT_75 => X"0000000000000000000000050000000000000019000000000000000000000000",
            INIT_76 => X"0000000000000000000000030000000000000000000000000000000400000000",
            INIT_77 => X"0000001200000000000000000000000000000016000000000000003d00000000",
            INIT_78 => X"0000000500000000000000060000000000000019000000000000001c00000000",
            INIT_79 => X"000000140000000000000000000000000000000c000000000000000b00000000",
            INIT_7A => X"0000001800000000000000000000000000000003000000000000000000000000",
            INIT_7B => X"0000000f0000000000000016000000000000000e000000000000001800000000",
            INIT_7C => X"0000001e00000000000000030000000000000012000000000000001300000000",
            INIT_7D => X"0000000000000000000000020000000000000005000000000000000000000000",
            INIT_7E => X"0000000b00000000000000010000000000000000000000000000000600000000",
            INIT_7F => X"000000040000000000000006000000000000000b000000000000000900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE17;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE18 : if BRAM_NAME = "samplegold_layersamples_instance18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000480000000000000000000000000000000500000000",
            INIT_01 => X"0000000d00000000000000060000000000000001000000000000000900000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"000000000000000000000033000000000000000a000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_0B => X"00000025000000000000002c0000000000000000000000000000000000000000",
            INIT_0C => X"0000000500000000000000310000000000000030000000000000000e00000000",
            INIT_0D => X"0000000f00000000000000100000000000000001000000000000000400000000",
            INIT_0E => X"0000000700000000000000100000000000000020000000000000001900000000",
            INIT_0F => X"0000005900000000000000530000000000000000000000000000000200000000",
            INIT_10 => X"0000003600000000000000810000000000000082000000000000003900000000",
            INIT_11 => X"0000005e000000000000005c000000000000006d000000000000004400000000",
            INIT_12 => X"0000006500000000000000750000000000000072000000000000006f00000000",
            INIT_13 => X"0000000d00000000000000000000000000000017000000000000004700000000",
            INIT_14 => X"0000004900000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000040000000000000012000000000000000500000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000037000000000000002200000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"00000015000000000000000c0000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000020000000000000014000000000000003800000000",
            INIT_20 => X"00000023000000000000003b000000000000000d000000000000000000000000",
            INIT_21 => X"0000001d0000000000000026000000000000000b000000000000000500000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000002800000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000900000000000000000000000000000003000000000000003a00000000",
            INIT_27 => X"0000000d00000000000000410000000000000046000000000000003800000000",
            INIT_28 => X"0000003e000000000000001a0000000000000000000000000000000000000000",
            INIT_29 => X"0000001200000000000000220000000000000006000000000000003100000000",
            INIT_2A => X"0000002b00000000000000410000000000000047000000000000002a00000000",
            INIT_2B => X"0000000c0000000000000010000000000000001c000000000000002200000000",
            INIT_2C => X"000000010000000000000000000000000000000e000000000000000100000000",
            INIT_2D => X"0000001a00000000000000140000000000000015000000000000002c00000000",
            INIT_2E => X"0000001400000000000000090000000000000026000000000000002700000000",
            INIT_2F => X"00000046000000000000003f0000000000000028000000000000001000000000",
            INIT_30 => X"0000001900000000000000390000000000000039000000000000003100000000",
            INIT_31 => X"0000000d000000000000002b000000000000002a000000000000000a00000000",
            INIT_32 => X"00000003000000000000000b0000000000000016000000000000001200000000",
            INIT_33 => X"0000001700000000000000210000000000000034000000000000003000000000",
            INIT_34 => X"0000001300000000000000230000000000000026000000000000001900000000",
            INIT_35 => X"0000000c00000000000000130000000000000000000000000000000000000000",
            INIT_36 => X"0000000800000000000000000000000000000000000000000000000a00000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_38 => X"0000002400000000000000100000000000000006000000000000000000000000",
            INIT_39 => X"0000000600000000000000080000000000000008000000000000000900000000",
            INIT_3A => X"000000560000000000000042000000000000000d000000000000000300000000",
            INIT_3B => X"00000082000000000000007b000000000000006f000000000000006b00000000",
            INIT_3C => X"0000009700000000000000950000000000000087000000000000009000000000",
            INIT_3D => X"000000980000000000000094000000000000009c000000000000008d00000000",
            INIT_3E => X"0000007c0000000000000061000000000000004d000000000000009c00000000",
            INIT_3F => X"0000008900000000000000840000000000000088000000000000007a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007600000000000000670000000000000095000000000000008900000000",
            INIT_41 => X"0000009f0000000000000097000000000000009500000000000000a200000000",
            INIT_42 => X"0000008700000000000000890000000000000066000000000000005a00000000",
            INIT_43 => X"00000074000000000000007f0000000000000086000000000000009600000000",
            INIT_44 => X"0000008b0000000000000078000000000000002c000000000000008200000000",
            INIT_45 => X"00000057000000000000009b0000000000000091000000000000008800000000",
            INIT_46 => X"0000008d00000000000000840000000000000082000000000000006800000000",
            INIT_47 => X"00000023000000000000006f000000000000007b000000000000008900000000",
            INIT_48 => X"0000004c00000000000000120000000000000013000000000000000000000000",
            INIT_49 => X"0000001b000000000000000d0000000000000084000000000000007c00000000",
            INIT_4A => X"0000003d00000000000000360000000000000036000000000000001d00000000",
            INIT_4B => X"000000190000000000000011000000000000001f000000000000003500000000",
            INIT_4C => X"0000005400000000000000730000000000000045000000000000001500000000",
            INIT_4D => X"00000029000000000000003a0000000000000021000000000000004000000000",
            INIT_4E => X"0000003400000000000000410000000000000044000000000000002f00000000",
            INIT_4F => X"0000005800000000000000210000000000000021000000000000001600000000",
            INIT_50 => X"0000002b00000000000000680000000000000067000000000000009400000000",
            INIT_51 => X"0000002800000000000000060000000000000018000000000000002200000000",
            INIT_52 => X"0000002e000000000000002e0000000000000029000000000000003000000000",
            INIT_53 => X"0000007d0000000000000080000000000000004b000000000000004400000000",
            INIT_54 => X"0000002d00000000000000000000000000000069000000000000005400000000",
            INIT_55 => X"00000056000000000000005e000000000000004e000000000000003e00000000",
            INIT_56 => X"0000003d0000000000000043000000000000004b000000000000005100000000",
            INIT_57 => X"0000006500000000000000670000000000000042000000000000002b00000000",
            INIT_58 => X"000000090000000000000017000000000000005a000000000000002600000000",
            INIT_59 => X"0000002500000000000000320000000000000035000000000000002300000000",
            INIT_5A => X"000000480000000000000051000000000000002e000000000000002300000000",
            INIT_5B => X"000000530000000000000058000000000000006e000000000000007e00000000",
            INIT_5C => X"00000040000000000000003c0000000000000005000000000000005600000000",
            INIT_5D => X"0000004e00000000000000430000000000000022000000000000002700000000",
            INIT_5E => X"0000005a000000000000004e0000000000000035000000000000004000000000",
            INIT_5F => X"000000150000000000000010000000000000002d000000000000004a00000000",
            INIT_60 => X"0000001700000000000000270000000000000025000000000000001a00000000",
            INIT_61 => X"00000000000000000000001b0000000000000027000000000000001d00000000",
            INIT_62 => X"00000007000000000000001e000000000000003a000000000000003000000000",
            INIT_63 => X"0000002400000000000000090000000000000003000000000000000800000000",
            INIT_64 => X"0000000f00000000000000000000000000000002000000000000001800000000",
            INIT_65 => X"0000001c00000000000000130000000000000011000000000000004000000000",
            INIT_66 => X"0000000000000000000000000000000000000008000000000000001300000000",
            INIT_67 => X"00000008000000000000001b0000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000040000000000000012000000000000000000000000",
            INIT_6A => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_6D => X"00000000000000000000000c0000000000000011000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"000000000000000000000005000000000000000a000000000000000400000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_72 => X"0000005200000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000003d000000000000003e0000000000000024000000000000001a00000000",
            INIT_74 => X"000000310000000000000053000000000000003f000000000000004200000000",
            INIT_75 => X"0000004f000000000000003f0000000000000054000000000000004100000000",
            INIT_76 => X"0000001e0000000000000053000000000000003d000000000000004500000000",
            INIT_77 => X"00000048000000000000003a0000000000000049000000000000002200000000",
            INIT_78 => X"0000007300000000000000380000000000000040000000000000003f00000000",
            INIT_79 => X"000000470000000000000054000000000000002e000000000000001100000000",
            INIT_7A => X"000000200000000000000026000000000000005a000000000000003900000000",
            INIT_7B => X"0000004d00000000000000450000000000000039000000000000004b00000000",
            INIT_7C => X"0000000000000000000000ab000000000000002b000000000000003700000000",
            INIT_7D => X"000000320000000000000042000000000000005a000000000000002d00000000",
            INIT_7E => X"0000003b00000000000000310000000000000025000000000000005e00000000",
            INIT_7F => X"000000490000000000000054000000000000003d000000000000004b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE18;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE19 : if BRAM_NAME = "samplegold_layersamples_instance19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000400000000000000000000000000000047000000000000005900000000",
            INIT_01 => X"0000002b0000000000000038000000000000003c000000000000000000000000",
            INIT_02 => X"000000250000000000000009000000000000001c000000000000002100000000",
            INIT_03 => X"00000039000000000000004c000000000000002b000000000000002300000000",
            INIT_04 => X"000000000000000000000000000000000000001a000000000000002b00000000",
            INIT_05 => X"000000000000000000000000000000000000000d000000000000003500000000",
            INIT_06 => X"0000000700000000000000000000000000000000000000000000002d00000000",
            INIT_07 => X"0000001b000000000000001d0000000000000036000000000000001100000000",
            INIT_08 => X"0000000300000000000000590000000000000004000000000000000000000000",
            INIT_09 => X"00000022000000000000001c0000000000000003000000000000005e00000000",
            INIT_0A => X"0000001900000000000000270000000000000000000000000000000000000000",
            INIT_0B => X"00000000000000000000000e000000000000000c000000000000002000000000",
            INIT_0C => X"0000008000000000000000280000000000000066000000000000002700000000",
            INIT_0D => X"0000000800000000000000080000000000000012000000000000001300000000",
            INIT_0E => X"0000003d00000000000000300000000000000027000000000000001a00000000",
            INIT_0F => X"00000013000000000000000d000000000000005e000000000000003600000000",
            INIT_10 => X"0000002400000000000000000000000000000073000000000000003200000000",
            INIT_11 => X"0000003a000000000000001c0000000000000000000000000000003400000000",
            INIT_12 => X"0000001600000000000000300000000000000038000000000000004000000000",
            INIT_13 => X"0000002d000000000000001f0000000000000000000000000000004500000000",
            INIT_14 => X"000000000000000000000026000000000000002f000000000000003800000000",
            INIT_15 => X"0000001c00000000000000230000000000000030000000000000001900000000",
            INIT_16 => X"000000240000000000000030000000000000003e000000000000002800000000",
            INIT_17 => X"0000004600000000000000480000000000000040000000000000002500000000",
            INIT_18 => X"000000260000000000000023000000000000000c000000000000001a00000000",
            INIT_19 => X"00000050000000000000001a0000000000000025000000000000004000000000",
            INIT_1A => X"00000041000000000000001b0000000000000000000000000000003e00000000",
            INIT_1B => X"0000001d0000000000000021000000000000002e000000000000003f00000000",
            INIT_1C => X"0000002000000000000000470000000000000024000000000000000000000000",
            INIT_1D => X"0000003700000000000000550000000000000000000000000000000600000000",
            INIT_1E => X"000000220000000000000028000000000000001a000000000000001200000000",
            INIT_1F => X"0000000000000000000000150000000000000011000000000000001500000000",
            INIT_20 => X"0000002200000000000000290000000000000043000000000000003100000000",
            INIT_21 => X"0000001d00000000000000100000000000000017000000000000001900000000",
            INIT_22 => X"0000002600000000000000040000000000000016000000000000001900000000",
            INIT_23 => X"0000000d000000000000000f0000000000000003000000000000000400000000",
            INIT_24 => X"0000000d000000000000000a0000000000000001000000000000000b00000000",
            INIT_25 => X"000000230000000000000000000000000000000f000000000000000900000000",
            INIT_26 => X"000000000000000000000009000000000000000a000000000000000d00000000",
            INIT_27 => X"0000000000000000000000000000000000000004000000000000000100000000",
            INIT_28 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"00000002000000000000003e0000000000000000000000000000001300000000",
            INIT_2A => X"0000002300000000000000000000000000000000000000000000000600000000",
            INIT_2B => X"00000098000000000000007d000000000000005800000000000000a500000000",
            INIT_2C => X"000000be00000000000000a600000000000000a0000000000000009f00000000",
            INIT_2D => X"000000aa00000000000000b700000000000000ae000000000000009700000000",
            INIT_2E => X"000000ab00000000000000a500000000000000b300000000000000b600000000",
            INIT_2F => X"000000a200000000000000a6000000000000007e000000000000006200000000",
            INIT_30 => X"0000009c00000000000000ac00000000000000a700000000000000a700000000",
            INIT_31 => X"000000bd000000000000009c000000000000006e00000000000000da00000000",
            INIT_32 => X"0000006200000000000000b1000000000000009f00000000000000b700000000",
            INIT_33 => X"000000a600000000000000a100000000000000aa000000000000007a00000000",
            INIT_34 => X"000001020000000000000085000000000000008d00000000000000b500000000",
            INIT_35 => X"000000ae00000000000000c10000000000000088000000000000001f00000000",
            INIT_36 => X"00000083000000000000005e00000000000000ac000000000000009600000000",
            INIT_37 => X"000000b0000000000000009500000000000000a9000000000000009300000000",
            INIT_38 => X"0000003400000000000000910000000000000094000000000000009f00000000",
            INIT_39 => X"0000008200000000000000970000000000000049000000000000004300000000",
            INIT_3A => X"0000004a000000000000005f0000000000000052000000000000006500000000",
            INIT_3B => X"0000009500000000000000700000000000000068000000000000006e00000000",
            INIT_3C => X"00000036000000000000003f0000000000000054000000000000006c00000000",
            INIT_3D => X"00000018000000000000004c0000000000000089000000000000002600000000",
            INIT_3E => X"0000004200000000000000260000000000000059000000000000002300000000",
            INIT_3F => X"0000004900000000000000680000000000000047000000000000003f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009f00000000000000500000000000000015000000000000004f00000000",
            INIT_41 => X"00000047000000000000002a0000000000000079000000000000005d00000000",
            INIT_42 => X"0000006900000000000000400000000000000014000000000000004a00000000",
            INIT_43 => X"00000053000000000000004f000000000000005e000000000000005a00000000",
            INIT_44 => X"0000005500000000000000be0000000000000076000000000000003200000000",
            INIT_45 => X"00000040000000000000004b0000000000000043000000000000009b00000000",
            INIT_46 => X"0000007a000000000000006d000000000000005b000000000000003c00000000",
            INIT_47 => X"0000004e000000000000009d0000000000000078000000000000008000000000",
            INIT_48 => X"0000004200000000000000b0000000000000007f000000000000006500000000",
            INIT_49 => X"000000610000000000000035000000000000005c000000000000005600000000",
            INIT_4A => X"0000007c000000000000007c000000000000007f000000000000007c00000000",
            INIT_4B => X"00000065000000000000003b0000000000000090000000000000005d00000000",
            INIT_4C => X"0000005b000000000000006b000000000000007c000000000000007600000000",
            INIT_4D => X"000000660000000000000068000000000000004b000000000000002900000000",
            INIT_4E => X"000000640000000000000079000000000000006c000000000000006400000000",
            INIT_4F => X"0000007f0000000000000087000000000000006e000000000000006f00000000",
            INIT_50 => X"0000005b00000000000000400000000000000047000000000000007a00000000",
            INIT_51 => X"0000005700000000000000500000000000000073000000000000006200000000",
            INIT_52 => X"0000005a0000000000000011000000000000006f000000000000009500000000",
            INIT_53 => X"00000042000000000000005a0000000000000075000000000000007600000000",
            INIT_54 => X"00000082000000000000005a000000000000000e000000000000003900000000",
            INIT_55 => X"00000085000000000000001d0000000000000038000000000000004e00000000",
            INIT_56 => X"0000004e000000000000004c0000000000000037000000000000005700000000",
            INIT_57 => X"0000002b00000000000000270000000000000038000000000000004200000000",
            INIT_58 => X"0000004100000000000000640000000000000052000000000000001800000000",
            INIT_59 => X"0000003200000000000000400000000000000041000000000000003f00000000",
            INIT_5A => X"0000001800000000000000360000000000000039000000000000003600000000",
            INIT_5B => X"0000002000000000000000140000000000000016000000000000003b00000000",
            INIT_5C => X"0000001f00000000000000150000000000000020000000000000002100000000",
            INIT_5D => X"0000000b000000000000002e0000000000000023000000000000002300000000",
            INIT_5E => X"0000001a000000000000001c0000000000000022000000000000003b00000000",
            INIT_5F => X"0000000700000000000000130000000000000012000000000000000d00000000",
            INIT_60 => X"000000140000000000000011000000000000000d000000000000000b00000000",
            INIT_61 => X"000000580000000000000000000000000000002a000000000000001800000000",
            INIT_62 => X"00000009000000000000000c0000000000000015000000000000001200000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000003100000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE19;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE20 : if BRAM_NAME = "samplegold_layersamples_instance20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_26 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"00000008000000000000000d000000000000000f000000000000000000000000",
            INIT_28 => X"0000003a00000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000001e0000000000000050000000000000001a000000000000002700000000",
            INIT_2A => X"00000032000000000000003b000000000000001e000000000000001700000000",
            INIT_2B => X"0000003e0000000000000043000000000000003c000000000000003400000000",
            INIT_2C => X"0000000000000000000000000000000000000019000000000000002b00000000",
            INIT_2D => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000003000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000350000000000000025000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000013000000000000001500000000",
            INIT_39 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000004000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000023000000000000002f0000000000000021000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000001000000000000000000000000000000000000000000000000e00000000",
            INIT_43 => X"0000002000000000000000220000000000000002000000000000000000000000",
            INIT_44 => X"0000000000000000000000150000000000000009000000000000001000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_47 => X"0000000000000000000000090000000000000009000000000000000000000000",
            INIT_48 => X"000000150000000000000000000000000000000c000000000000000a00000000",
            INIT_49 => X"0000001700000000000000190000000000000010000000000000001900000000",
            INIT_4A => X"0000000f000000000000000e0000000000000000000000000000000000000000",
            INIT_4B => X"00000001000000000000000f0000000000000001000000000000000000000000",
            INIT_4C => X"0000000a000000000000001a0000000000000020000000000000000000000000",
            INIT_4D => X"00000006000000000000000a0000000000000004000000000000000000000000",
            INIT_4E => X"0000000500000000000000000000000000000000000000000000000200000000",
            INIT_4F => X"0000000000000000000000000000000000000001000000000000000600000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_51 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"000000040000000000000004000000000000000a000000000000000000000000",
            INIT_53 => X"00000000000000000000001c0000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000001200000000000000000000000000000007000000000000000200000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_5F => X"0000000e00000000000000150000000000000008000000000000000500000000",
            INIT_60 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_62 => X"0000001d0000000000000016000000000000001d000000000000002000000000",
            INIT_63 => X"000000230000000000000020000000000000000f000000000000001b00000000",
            INIT_64 => X"000000050000000000000011000000000000001b000000000000002600000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_66 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000003000000000000000100000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000001400000000000000140000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000008000000000000000500000000",
            INIT_71 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000700000000000000000000000000000000000000000000001000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000009000000000000000200000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_77 => X"0000000000000000000000140000000000000015000000000000000000000000",
            INIT_78 => X"000000100000000000000017000000000000000a000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000001000000000000000900000000",
            INIT_7A => X"000000000000000000000005000000000000001b000000000000001100000000",
            INIT_7B => X"0000001800000000000000120000000000000000000000000000000000000000",
            INIT_7C => X"0000000b0000000000000002000000000000000a000000000000000600000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000001300000000000000180000000000000000000000000000000000000000",
            INIT_7F => X"00000000000000000000000a0000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE20;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE21 : if BRAM_NAME = "samplegold_layersamples_instance21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"000000060000000000000019000000000000001a000000000000002000000000",
            INIT_02 => X"0000000d00000000000000030000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000600000000000000060000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000001000000000000002300000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000001d00000000000000000000000000000003000000000000000a00000000",
            INIT_10 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_14 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000020000000000000014000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_19 => X"0000000b00000000000000000000000000000000000000000000000800000000",
            INIT_1A => X"0000000000000000000000000000000000000025000000000000000500000000",
            INIT_1B => X"0000000000000000000000000000000000000002000000000000000800000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_27 => X"0000000000000000000000130000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_2B => X"000000000000000000000001000000000000000c000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"000000000000000000000003000000000000000b000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"00000000000000000000001e0000000000000000000000000000000000000000",
            INIT_32 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000290000000000000088000000000000003d00000000",
            INIT_34 => X"0000001f0000000000000088000000000000001f000000000000004600000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000044000000000000000000000000",
            INIT_41 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"000000070000000000000001000000000000000d000000000000000300000000",
            INIT_43 => X"0000004000000000000000160000000000000000000000000000000000000000",
            INIT_44 => X"0000018500000000000001b70000000000000189000000000000000000000000",
            INIT_45 => X"00000194000000000000019b0000000000000187000000000000016e00000000",
            INIT_46 => X"0000019b00000000000001970000000000000193000000000000019000000000",
            INIT_47 => X"000001d100000000000001c800000000000001aa000000000000019600000000",
            INIT_48 => X"0000014300000000000001b400000000000001bd000000000000018a00000000",
            INIT_49 => X"0000014d0000000000000144000000000000014c000000000000013b00000000",
            INIT_4A => X"00000170000000000000015d000000000000015a000000000000015300000000",
            INIT_4B => X"0000018500000000000001d700000000000001d100000000000001c400000000",
            INIT_4C => X"00000147000000000000013600000000000001a800000000000001b000000000",
            INIT_4D => X"0000015800000000000001430000000000000126000000000000013b00000000",
            INIT_4E => X"000001b60000000000000162000000000000015a000000000000015a00000000",
            INIT_4F => X"000001ac000000000000018200000000000001dd00000000000001d400000000",
            INIT_50 => X"00000156000000000000014b000000000000012d000000000000019000000000",
            INIT_51 => X"000001510000000000000159000000000000014f000000000000014900000000",
            INIT_52 => X"000001c900000000000001810000000000000168000000000000015600000000",
            INIT_53 => X"000001ac00000000000001aa000000000000019500000000000001d200000000",
            INIT_54 => X"0000016a00000000000001630000000000000166000000000000018300000000",
            INIT_55 => X"00000172000000000000016e0000000000000175000000000000017800000000",
            INIT_56 => X"000001cc00000000000001c900000000000001b800000000000001a500000000",
            INIT_57 => X"000001af000000000000017e000000000000019f00000000000001b600000000",
            INIT_58 => X"000001b700000000000001b100000000000001a500000000000001ab00000000",
            INIT_59 => X"000001bb00000000000001b000000000000001ab00000000000001ab00000000",
            INIT_5A => X"000001c700000000000001d100000000000001cb00000000000001c700000000",
            INIT_5B => X"0000015600000000000000fd000000000000012a000000000000019900000000",
            INIT_5C => X"000001d000000000000001d300000000000001cd00000000000001b800000000",
            INIT_5D => X"000001c500000000000001c300000000000001c400000000000001c500000000",
            INIT_5E => X"000001de00000000000001d700000000000001cd00000000000001c700000000",
            INIT_5F => X"0000011000000000000000b0000000000000014500000000000001c300000000",
            INIT_60 => X"000001c100000000000001ce00000000000001d4000000000000019600000000",
            INIT_61 => X"000001c300000000000001c500000000000001c200000000000001c200000000",
            INIT_62 => X"000001e700000000000001ea00000000000001de00000000000001c600000000",
            INIT_63 => X"000000b8000000000000008600000000000000b200000000000001d400000000",
            INIT_64 => X"000001ba000000000000018d0000000000000150000000000000010100000000",
            INIT_65 => X"000001c500000000000001c200000000000001c500000000000001c900000000",
            INIT_66 => X"000001b900000000000001e500000000000001e200000000000001de00000000",
            INIT_67 => X"0000007e00000000000000640000000000000040000000000000009900000000",
            INIT_68 => X"0000010900000000000000b4000000000000008e000000000000009200000000",
            INIT_69 => X"000001d400000000000001c300000000000001a2000000000000015c00000000",
            INIT_6A => X"0000014700000000000001b500000000000001df00000000000001db00000000",
            INIT_6B => X"00000145000000000000011300000000000000b000000000000000d200000000",
            INIT_6C => X"0000014600000000000000d600000000000000f500000000000000e400000000",
            INIT_6D => X"00000156000000000000015600000000000001ae000000000000019300000000",
            INIT_6E => X"000001130000000000000138000000000000013d000000000000014700000000",
            INIT_6F => X"0000012e0000000000000149000000000000013f000000000000010b00000000",
            INIT_70 => X"0000015300000000000001550000000000000141000000000000014700000000",
            INIT_71 => X"000000c600000000000000d400000000000000cd000000000000015800000000",
            INIT_72 => X"000000a300000000000000a500000000000000af00000000000000b900000000",
            INIT_73 => X"000000a200000000000000a500000000000000ae00000000000000b700000000",
            INIT_74 => X"0000009a00000000000000a400000000000000aa00000000000000a300000000",
            INIT_75 => X"000000620000000000000065000000000000006e000000000000006600000000",
            INIT_76 => X"0000005500000000000000500000000000000050000000000000005a00000000",
            INIT_77 => X"0000004400000000000000440000000000000046000000000000005500000000",
            INIT_78 => X"00000043000000000000009b0000000000000050000000000000004400000000",
            INIT_79 => X"00000046000000000000004a0000000000000049000000000000004900000000",
            INIT_7A => X"00000060000000000000005f0000000000000057000000000000005800000000",
            INIT_7B => X"0000006e00000000000000460000000000000049000000000000005800000000",
            INIT_7C => X"0000006d0000000000000067000000000000009e00000000000000af00000000",
            INIT_7D => X"0000005b000000000000005f0000000000000050000000000000004400000000",
            INIT_7E => X"0000005700000000000000510000000000000057000000000000005300000000",
            INIT_7F => X"0000006900000000000000600000000000000057000000000000005800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE21;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE22 : if BRAM_NAME = "samplegold_layersamples_instance22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000600000000000000078000000000000006d000000000000006c00000000",
            INIT_01 => X"0000006b00000000000000790000000000000070000000000000003c00000000",
            INIT_02 => X"0000007700000000000000740000000000000073000000000000007900000000",
            INIT_03 => X"0000007400000000000000750000000000000077000000000000007600000000",
            INIT_04 => X"0000005200000000000000720000000000000072000000000000006b00000000",
            INIT_05 => X"00000054000000000000003e000000000000004a000000000000004000000000",
            INIT_06 => X"00000059000000000000004d0000000000000049000000000000004a00000000",
            INIT_07 => X"0000006200000000000000780000000000000072000000000000007b00000000",
            INIT_08 => X"00000051000000000000003e000000000000004d000000000000007000000000",
            INIT_09 => X"0000005700000000000000520000000000000042000000000000005400000000",
            INIT_0A => X"0000007400000000000000530000000000000059000000000000005100000000",
            INIT_0B => X"0000006f000000000000005d0000000000000079000000000000007400000000",
            INIT_0C => X"0000005c00000000000000590000000000000054000000000000006500000000",
            INIT_0D => X"0000005800000000000000610000000000000061000000000000005900000000",
            INIT_0E => X"0000006f00000000000000690000000000000073000000000000005c00000000",
            INIT_0F => X"0000006e000000000000006b0000000000000065000000000000007300000000",
            INIT_10 => X"00000058000000000000004f000000000000004e000000000000006500000000",
            INIT_11 => X"0000005500000000000000510000000000000053000000000000005b00000000",
            INIT_12 => X"00000071000000000000006e0000000000000070000000000000006900000000",
            INIT_13 => X"0000007a0000000000000014000000000000003d000000000000006d00000000",
            INIT_14 => X"000000750000000000000075000000000000007e000000000000009e00000000",
            INIT_15 => X"0000006f0000000000000071000000000000006a000000000000006f00000000",
            INIT_16 => X"0000007b000000000000007a0000000000000075000000000000007200000000",
            INIT_17 => X"0000000f00000000000000000000000000000048000000000000007400000000",
            INIT_18 => X"00000073000000000000007b000000000000009c000000000000009400000000",
            INIT_19 => X"0000006d000000000000006c000000000000006e000000000000006d00000000",
            INIT_1A => X"0000007a000000000000007e0000000000000071000000000000006b00000000",
            INIT_1B => X"0000000f00000000000000000000000000000060000000000000007200000000",
            INIT_1C => X"00000082000000000000009a0000000000000095000000000000004c00000000",
            INIT_1D => X"00000070000000000000006f000000000000006e000000000000007c00000000",
            INIT_1E => X"000000760000000000000078000000000000007c000000000000007200000000",
            INIT_1F => X"0000000900000000000000010000000000000000000000000000006e00000000",
            INIT_20 => X"0000008a000000000000003c0000000000000011000000000000000300000000",
            INIT_21 => X"00000075000000000000007f0000000000000096000000000000009e00000000",
            INIT_22 => X"0000004100000000000000780000000000000077000000000000008100000000",
            INIT_23 => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000008f0000000000000072000000000000004b000000000000003500000000",
            INIT_26 => X"00000091000000000000008d000000000000008a000000000000008d00000000",
            INIT_27 => X"00000080000000000000007a000000000000005b000000000000006900000000",
            INIT_28 => X"0000006f00000000000000620000000000000070000000000000006300000000",
            INIT_29 => X"00000025000000000000001f000000000000007f000000000000007f00000000",
            INIT_2A => X"0000001100000000000000140000000000000017000000000000001c00000000",
            INIT_2B => X"0000003c00000000000000360000000000000036000000000000001800000000",
            INIT_2C => X"00000049000000000000004e0000000000000048000000000000003e00000000",
            INIT_2D => X"00000014000000000000001b0000000000000009000000000000004900000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000002000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000002700000000000000280000000000000030000000000000003100000000",
            INIT_36 => X"0000002500000000000000260000000000000023000000000000002700000000",
            INIT_37 => X"0000002700000000000000250000000000000024000000000000002500000000",
            INIT_38 => X"0000003100000000000000240000000000000021000000000000002000000000",
            INIT_39 => X"0000001a00000000000000130000000000000026000000000000003400000000",
            INIT_3A => X"00000019000000000000001a0000000000000019000000000000001500000000",
            INIT_3B => X"0000002800000000000000230000000000000024000000000000001800000000",
            INIT_3C => X"00000036000000000000002f0000000000000025000000000000002500000000",
            INIT_3D => X"0000001e0000000000000019000000000000001c000000000000003500000000",
            INIT_3E => X"00000020000000000000001e0000000000000023000000000000001d00000000",
            INIT_3F => X"000000270000000000000022000000000000001f000000000000001f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001a000000000000002b0000000000000033000000000000002600000000",
            INIT_41 => X"00000018000000000000001b000000000000001a000000000000001800000000",
            INIT_42 => X"0000001400000000000000100000000000000016000000000000001700000000",
            INIT_43 => X"00000024000000000000002a0000000000000025000000000000001b00000000",
            INIT_44 => X"0000002b000000000000002b0000000000000038000000000000003000000000",
            INIT_45 => X"0000002a000000000000002d000000000000002f000000000000002b00000000",
            INIT_46 => X"0000002b000000000000002e0000000000000025000000000000002b00000000",
            INIT_47 => X"00000027000000000000001f000000000000002d000000000000002d00000000",
            INIT_48 => X"00000032000000000000002f0000000000000037000000000000002f00000000",
            INIT_49 => X"0000002d00000000000000300000000000000030000000000000003000000000",
            INIT_4A => X"0000002c000000000000002e0000000000000028000000000000002c00000000",
            INIT_4B => X"000000220000000000000031000000000000001c000000000000002d00000000",
            INIT_4C => X"0000002f0000000000000030000000000000002a000000000000001600000000",
            INIT_4D => X"0000002b000000000000002b000000000000002e000000000000002f00000000",
            INIT_4E => X"0000002c000000000000002a000000000000002b000000000000002b00000000",
            INIT_4F => X"0000001f000000000000002d0000000000000029000000000000001900000000",
            INIT_50 => X"000000280000000000000025000000000000001b000000000000001200000000",
            INIT_51 => X"0000002b0000000000000029000000000000002b000000000000002a00000000",
            INIT_52 => X"00000014000000000000002f000000000000002d000000000000002c00000000",
            INIT_53 => X"0000002400000000000000250000000000000023000000000000002100000000",
            INIT_54 => X"0000001e00000000000000130000000000000009000000000000000f00000000",
            INIT_55 => X"0000002b000000000000002e000000000000002f000000000000002300000000",
            INIT_56 => X"0000001f0000000000000011000000000000002f000000000000002b00000000",
            INIT_57 => X"00000014000000000000002b0000000000000019000000000000002300000000",
            INIT_58 => X"00000010000000000000000a0000000000000012000000000000001400000000",
            INIT_59 => X"00000027000000000000001e0000000000000018000000000000001b00000000",
            INIT_5A => X"0000002300000000000000260000000000000016000000000000002d00000000",
            INIT_5B => X"00000021000000000000001d0000000000000036000000000000002700000000",
            INIT_5C => X"0000001d000000000000002b0000000000000018000000000000002600000000",
            INIT_5D => X"00000025000000000000001f000000000000001a000000000000001f00000000",
            INIT_5E => X"0000001b000000000000001c000000000000001f000000000000001000000000",
            INIT_5F => X"0000002200000000000000220000000000000028000000000000001c00000000",
            INIT_60 => X"0000003800000000000000300000000000000038000000000000003000000000",
            INIT_61 => X"000000190000000000000039000000000000003d000000000000003300000000",
            INIT_62 => X"0000001900000000000000200000000000000026000000000000002a00000000",
            INIT_63 => X"0000002300000000000000200000000000000021000000000000001d00000000",
            INIT_64 => X"0000002200000000000000210000000000000022000000000000002200000000",
            INIT_65 => X"0000001800000000000000120000000000000020000000000000002200000000",
            INIT_66 => X"00000012000000000000000e0000000000000014000000000000001700000000",
            INIT_67 => X"0000000d000000000000000d0000000000000011000000000000001400000000",
            INIT_68 => X"0000000d000000000000000e000000000000000d000000000000000d00000000",
            INIT_69 => X"000000110000000000000012000000000000000d000000000000001100000000",
            INIT_6A => X"000000100000000000000013000000000000000f000000000000000e00000000",
            INIT_6B => X"0000000b000000000000000f000000000000000d000000000000000e00000000",
            INIT_6C => X"000000000000000000000009000000000000000b000000000000000800000000",
            INIT_6D => X"000000130000000000000000000000000000000d000000000000001e00000000",
            INIT_6E => X"0000001500000000000000110000000000000010000000000000001c00000000",
            INIT_6F => X"0000001400000000000000130000000000000014000000000000001400000000",
            INIT_70 => X"0000001500000000000000200000000000000020000000000000001a00000000",
            INIT_71 => X"00000042000000000000002f0000000000000005000000000000000800000000",
            INIT_72 => X"0000004900000000000000490000000000000046000000000000004900000000",
            INIT_73 => X"0000002200000000000000460000000000000046000000000000004600000000",
            INIT_74 => X"000000050000000000000013000000000000001c000000000000001c00000000",
            INIT_75 => X"0000004f000000000000004c0000000000000040000000000000000800000000",
            INIT_76 => X"0000004a000000000000004c000000000000005b000000000000005400000000",
            INIT_77 => X"0000001b000000000000003d0000000000000045000000000000004900000000",
            INIT_78 => X"000000130000000000000004000000000000000f000000000000001900000000",
            INIT_79 => X"00000035000000000000003a0000000000000039000000000000003700000000",
            INIT_7A => X"0000004100000000000000360000000000000034000000000000003f00000000",
            INIT_7B => X"0000001400000000000000140000000000000039000000000000003000000000",
            INIT_7C => X"0000000f00000000000000060000000000000006000000000000000d00000000",
            INIT_7D => X"00000017000000000000000d000000000000000f000000000000001100000000",
            INIT_7E => X"0000002200000000000000190000000000000014000000000000001400000000",
            INIT_7F => X"0000001600000000000000110000000000000012000000000000001700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE22;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE23 : if BRAM_NAME = "samplegold_layersamples_instance23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000c000000000000000c0000000000000010000000000000000e00000000",
            INIT_01 => X"0000001000000000000000140000000000000012000000000000000b00000000",
            INIT_02 => X"0000001000000000000000140000000000000014000000000000000f00000000",
            INIT_03 => X"00000000000000000000001c0000000000000011000000000000001100000000",
            INIT_04 => X"000000170000000000000028000000000000002b000000000000000000000000",
            INIT_05 => X"0000001200000000000000120000000000000012000000000000001300000000",
            INIT_06 => X"0000001400000000000000130000000000000013000000000000001600000000",
            INIT_07 => X"0000001000000000000000110000000000000020000000000000001400000000",
            INIT_08 => X"0000002f00000000000000380000000000000018000000000000000000000000",
            INIT_09 => X"0000001600000000000000130000000000000016000000000000001d00000000",
            INIT_0A => X"0000000e00000000000000100000000000000012000000000000001300000000",
            INIT_0B => X"0000001d000000000000001b000000000000001d000000000000002700000000",
            INIT_0C => X"00000037000000000000002d0000000000000020000000000000000000000000",
            INIT_0D => X"00000012000000000000001b0000000000000027000000000000003500000000",
            INIT_0E => X"0000002b000000000000000f0000000000000011000000000000001300000000",
            INIT_0F => X"00000000000000000000001c000000000000001c000000000000002100000000",
            INIT_10 => X"0000002000000000000000220000000000000021000000000000001c00000000",
            INIT_11 => X"0000003300000000000000330000000000000029000000000000001900000000",
            INIT_12 => X"0000001c000000000000002b0000000000000017000000000000002400000000",
            INIT_13 => X"000000000000000000000000000000000000000a000000000000001d00000000",
            INIT_14 => X"00000006000000000000000e0000000000000023000000000000000200000000",
            INIT_15 => X"0000001f00000000000000230000000000000001000000000000000100000000",
            INIT_16 => X"0000002800000000000000290000000000000038000000000000001c00000000",
            INIT_17 => X"00000026000000000000001e000000000000002b000000000000002a00000000",
            INIT_18 => X"0000001800000000000000060000000000000016000000000000002700000000",
            INIT_19 => X"0000000a00000000000000090000000000000011000000000000000c00000000",
            INIT_1A => X"0000001700000000000000120000000000000012000000000000001a00000000",
            INIT_1B => X"00000020000000000000001a0000000000000019000000000000001a00000000",
            INIT_1C => X"0000001b0000000000000019000000000000001a000000000000001600000000",
            INIT_1D => X"00000018000000000000001b0000000000000019000000000000001c00000000",
            INIT_1E => X"0000001800000000000000180000000000000014000000000000001800000000",
            INIT_1F => X"0000001900000000000000190000000000000016000000000000001700000000",
            INIT_20 => X"0000001900000000000000190000000000000019000000000000001800000000",
            INIT_21 => X"00000018000000000000001a0000000000000010000000000000001600000000",
            INIT_22 => X"000000180000000000000018000000000000001a000000000000001700000000",
            INIT_23 => X"000000160000000000000017000000000000001b000000000000001700000000",
            INIT_24 => X"0000000d0000000000000016000000000000001e000000000000001800000000",
            INIT_25 => X"0000000000000000000000000000000000000003000000000000000f00000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"00000007000000000000002f0000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000060000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002f00000000000000130000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_44 => X"00000033000000000000001f0000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000009000000000000002d00000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_48 => X"00000011000000000000001c000000000000001c000000000000000000000000",
            INIT_49 => X"0000002100000000000000350000000000000029000000000000001c00000000",
            INIT_4A => X"0000000600000000000000000000000000000000000000000000000800000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"000000000000000000000016000000000000000e000000000000000000000000",
            INIT_4D => X"0000002000000000000000060000000000000000000000000000000000000000",
            INIT_4E => X"00000004000000000000000f0000000000000000000000000000000600000000",
            INIT_4F => X"0000000000000000000000090000000000000008000000000000000600000000",
            INIT_50 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_53 => X"0000000500000000000000030000000000000006000000000000000100000000",
            INIT_54 => X"0000000b000000000000000c0000000000000005000000000000000e00000000",
            INIT_55 => X"0000000e000000000000000a000000000000000e000000000000000f00000000",
            INIT_56 => X"0000001e000000000000001b000000000000001d000000000000001400000000",
            INIT_57 => X"00000020000000000000001e000000000000001e000000000000001f00000000",
            INIT_58 => X"0000001e0000000000000021000000000000001e000000000000001f00000000",
            INIT_59 => X"0000000a0000000000000026000000000000001b000000000000001d00000000",
            INIT_5A => X"00000019000000000000001e0000000000000019000000000000001800000000",
            INIT_5B => X"00000019000000000000001c0000000000000018000000000000001a00000000",
            INIT_5C => X"0000001c0000000000000022000000000000001c000000000000001b00000000",
            INIT_5D => X"0000009a00000000000000850000000000000032000000000000003400000000",
            INIT_5E => X"00000083000000000000007c0000000000000078000000000000008600000000",
            INIT_5F => X"0000007f000000000000007c000000000000007b000000000000007e00000000",
            INIT_60 => X"00000084000000000000007f000000000000007e000000000000008000000000",
            INIT_61 => X"0000009800000000000000ab0000000000000092000000000000008900000000",
            INIT_62 => X"0000004c00000000000000500000000000000046000000000000004c00000000",
            INIT_63 => X"000000560000000000000050000000000000004e000000000000005000000000",
            INIT_64 => X"00000090000000000000008e0000000000000083000000000000005a00000000",
            INIT_65 => X"0000002e000000000000009e00000000000000a9000000000000009200000000",
            INIT_66 => X"000000180000000000000019000000000000001d000000000000002e00000000",
            INIT_67 => X"0000003b000000000000002e000000000000002e000000000000002600000000",
            INIT_68 => X"0000008f00000000000000950000000000000094000000000000007b00000000",
            INIT_69 => X"0000003a000000000000001b000000000000008300000000000000a500000000",
            INIT_6A => X"00000044000000000000003c0000000000000034000000000000004800000000",
            INIT_6B => X"0000005d00000000000000470000000000000040000000000000004200000000",
            INIT_6C => X"000000a30000000000000090000000000000009a000000000000009700000000",
            INIT_6D => X"0000007e000000000000007d0000000000000085000000000000009900000000",
            INIT_6E => X"0000007e00000000000000800000000000000080000000000000008100000000",
            INIT_6F => X"0000009900000000000000850000000000000087000000000000007c00000000",
            INIT_70 => X"00000096000000000000009c0000000000000093000000000000009a00000000",
            INIT_71 => X"0000008500000000000000830000000000000087000000000000009100000000",
            INIT_72 => X"0000008600000000000000860000000000000082000000000000008500000000",
            INIT_73 => X"0000009a0000000000000096000000000000009a000000000000009000000000",
            INIT_74 => X"00000086000000000000006f000000000000008a000000000000009300000000",
            INIT_75 => X"0000009900000000000000990000000000000098000000000000008e00000000",
            INIT_76 => X"0000009500000000000000950000000000000093000000000000009600000000",
            INIT_77 => X"00000099000000000000009a000000000000009a000000000000009900000000",
            INIT_78 => X"00000046000000000000003a000000000000008000000000000000a000000000",
            INIT_79 => X"0000009500000000000000960000000000000090000000000000008500000000",
            INIT_7A => X"0000009600000000000000920000000000000091000000000000009000000000",
            INIT_7B => X"0000009a000000000000009a000000000000009b000000000000009500000000",
            INIT_7C => X"00000036000000000000002b0000000000000088000000000000009600000000",
            INIT_7D => X"0000008900000000000000840000000000000083000000000000005c00000000",
            INIT_7E => X"0000009800000000000000960000000000000093000000000000009100000000",
            INIT_7F => X"0000009400000000000000930000000000000094000000000000009b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE23;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE24 : if BRAM_NAME = "samplegold_layersamples_instance24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002800000000000000270000000000000035000000000000009300000000",
            INIT_01 => X"0000007e000000000000005f0000000000000039000000000000002300000000",
            INIT_02 => X"00000094000000000000008b0000000000000087000000000000008800000000",
            INIT_03 => X"0000007f00000000000000950000000000000093000000000000009300000000",
            INIT_04 => X"00000036000000000000002d0000000000000017000000000000003400000000",
            INIT_05 => X"0000002f00000000000000270000000000000027000000000000003400000000",
            INIT_06 => X"00000088000000000000008d0000000000000074000000000000005700000000",
            INIT_07 => X"0000008c000000000000008b000000000000008b000000000000008e00000000",
            INIT_08 => X"000000910000000000000080000000000000006a000000000000007700000000",
            INIT_09 => X"0000008d000000000000007b0000000000000088000000000000007900000000",
            INIT_0A => X"0000004e00000000000000450000000000000093000000000000009600000000",
            INIT_0B => X"0000004000000000000000420000000000000045000000000000004a00000000",
            INIT_0C => X"0000005b00000000000000590000000000000056000000000000004200000000",
            INIT_0D => X"0000006300000000000000660000000000000062000000000000005d00000000",
            INIT_0E => X"0000003b000000000000003f0000000000000031000000000000006200000000",
            INIT_0F => X"0000002b000000000000002c000000000000002d000000000000003400000000",
            INIT_10 => X"0000002100000000000000210000000000000028000000000000002a00000000",
            INIT_11 => X"0000003600000000000000200000000000000020000000000000002000000000",
            INIT_12 => X"0000001e000000000000001f000000000000001f000000000000001100000000",
            INIT_13 => X"0000001b000000000000001b000000000000001e000000000000001a00000000",
            INIT_14 => X"0000001a0000000000000019000000000000001b000000000000001d00000000",
            INIT_15 => X"00000000000000000000005b0000000000000048000000000000002100000000",
            INIT_16 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"00000022000000000000001d0000000000000023000000000000000000000000",
            INIT_1B => X"000000200000000000000029000000000000002a000000000000002600000000",
            INIT_1C => X"0000000000000000000000000000000000000029000000000000002400000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"00000021000000000000000a000000000000000c000000000000002400000000",
            INIT_1F => X"0000000a000000000000000b000000000000000c000000000000001500000000",
            INIT_20 => X"0000000000000000000000000000000000000004000000000000000b00000000",
            INIT_21 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"000000070000000000000006000000000000000a000000000000000600000000",
            INIT_23 => X"000000010000000000000008000000000000000b000000000000000400000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000001f00000000000000020000000000000000000000000000000000000000",
            INIT_35 => X"000000030000000000000009000000000000000f000000000000001000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000001500000000000000230000000000000000000000000000000000000000",
            INIT_39 => X"0000001100000000000000140000000000000018000000000000001400000000",
            INIT_3A => X"0000000000000000000000000000000000000003000000000000000600000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000001000000000000000120000000000000017000000000000000500000000",
            INIT_3D => X"0000000d000000000000001c000000000000000a000000000000000e00000000",
            INIT_3E => X"0000000000000000000000000000000000000002000000000000001400000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000600000000000000020000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000002000000000000000800000000",
            INIT_45 => X"0000000100000000000000010000000000000001000000000000000100000000",
            INIT_46 => X"0000001700000000000000260000000000000005000000000000000100000000",
            INIT_47 => X"0000001e0000000000000020000000000000001c000000000000001800000000",
            INIT_48 => X"0000001e000000000000001c000000000000001d000000000000001a00000000",
            INIT_49 => X"00000018000000000000001b000000000000001b000000000000001e00000000",
            INIT_4A => X"000000180000000000000019000000000000002b000000000000001000000000",
            INIT_4B => X"0000001e000000000000001e000000000000001f000000000000001a00000000",
            INIT_4C => X"0000002200000000000000220000000000000023000000000000002100000000",
            INIT_4D => X"00000018000000000000000a0000000000000018000000000000002000000000",
            INIT_4E => X"000000050000000000000000000000000000000f000000000000003000000000",
            INIT_4F => X"0000000600000000000000000000000000000004000000000000001b00000000",
            INIT_50 => X"0000000100000000000000010000000000000003000000000000000000000000",
            INIT_51 => X"0000002d00000000000000050000000000000009000000000000001200000000",
            INIT_52 => X"0000002600000000000000000000000000000000000000000000001d00000000",
            INIT_53 => X"0000001d000000000000002d0000000000000012000000000000002b00000000",
            INIT_54 => X"0000001a0000000000000033000000000000001d000000000000002100000000",
            INIT_55 => X"00000015000000000000002e000000000000000a000000000000000900000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_57 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_58 => X"00000007000000000000002c000000000000000e000000000000000000000000",
            INIT_59 => X"000000000000000000000016000000000000001e000000000000000c00000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000800000000000000000000000000000000000000000000000700000000",
            INIT_5C => X"0000000f000000000000000b000000000000002c000000000000000000000000",
            INIT_5D => X"0000000000000000000000010000000000000013000000000000000300000000",
            INIT_5E => X"0000000e000000000000000e000000000000000e000000000000000a00000000",
            INIT_5F => X"0000002d000000000000000e0000000000000000000000000000000800000000",
            INIT_60 => X"00000007000000000000000a000000000000000a000000000000000100000000",
            INIT_61 => X"0000000000000000000000120000000000000010000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"00000008000000000000000b0000000000000000000000000000000000000000",
            INIT_64 => X"000000000000000000000015000000000000000b000000000000000500000000",
            INIT_65 => X"0000002d000000000000006d0000000000000038000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000003000000000000000c00000000",
            INIT_67 => X"0000000a00000000000000080000000000000002000000000000000700000000",
            INIT_68 => X"0000000000000000000000000000000000000023000000000000001000000000",
            INIT_69 => X"00000065000000000000007d0000000000000000000000000000000000000000",
            INIT_6A => X"0000000500000000000000000000000000000000000000000000001500000000",
            INIT_6B => X"0000000900000000000000010000000000000003000000000000000100000000",
            INIT_6C => X"0000000000000000000000000000000000000009000000000000002300000000",
            INIT_6D => X"0000006b0000000000000053000000000000001f000000000000000000000000",
            INIT_6E => X"000000010000000000000028000000000000002d000000000000005900000000",
            INIT_6F => X"00000023000000000000000a0000000000000005000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000005000000000000000a00000000",
            INIT_71 => X"0000001c00000000000000120000000000000022000000000000001600000000",
            INIT_72 => X"0000005a0000000000000066000000000000007a000000000000002600000000",
            INIT_73 => X"00000009000000000000002b0000000000000012000000000000003400000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_75 => X"0000000000000000000000000000000000000032000000000000000000000000",
            INIT_76 => X"0000001200000000000000440000000000000000000000000000000000000000",
            INIT_77 => X"0000002d000000000000002c0000000000000045000000000000001400000000",
            INIT_78 => X"000000220000000000000003000000000000003b000000000000003200000000",
            INIT_79 => X"0000002500000000000000170000000000000022000000000000004e00000000",
            INIT_7A => X"0000002900000000000000290000000000000026000000000000001600000000",
            INIT_7B => X"0000000000000000000000000000000000000002000000000000000600000000",
            INIT_7C => X"0000001e00000000000000060000000000000000000000000000000000000000",
            INIT_7D => X"0000002400000000000000190000000000000018000000000000000800000000",
            INIT_7E => X"000000020000000000000025000000000000001a000000000000002400000000",
            INIT_7F => X"0000000800000000000000150000000000000010000000000000001b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE24;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE25 : if BRAM_NAME = "samplegold_layersamples_instance25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000300000000000000110000000000000010000000000000000d00000000",
            INIT_01 => X"0000000700000000000000050000000000000008000000000000000000000000",
            INIT_02 => X"0000000200000000000000000000000000000016000000000000000900000000",
            INIT_03 => X"0000000800000000000000000000000000000008000000000000000200000000",
            INIT_04 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_05 => X"0000000800000000000000130000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000002100000000000000260000000000000026000000000000000900000000",
            INIT_0C => X"0000002500000000000000240000000000000023000000000000001f00000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000100000000000000080000000000000003000000000000000000000000",
            INIT_17 => X"0000000000000000000000030000000000000005000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"00000000000000000000002b0000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000007d000000000000005f0000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000007400000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000001000000000000005700000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000004f00000000000000090000000000000000000000000000000000000000",
            INIT_26 => X"0000000e000000000000003f0000000000000087000000000000009800000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000200000000000000180000000000000025000000000000001800000000",
            INIT_2A => X"000000b300000000000000ad0000000000000060000000000000001900000000",
            INIT_2B => X"0000000000000000000000000000000000000032000000000000008500000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000007c00000000000000780000000000000000000000000000000000000000",
            INIT_30 => X"0000007f000000000000009f0000000000000095000000000000008b00000000",
            INIT_31 => X"000000440000000000000069000000000000005b000000000000005300000000",
            INIT_32 => X"0000004f000000000000003a0000000000000033000000000000004500000000",
            INIT_33 => X"0000000000000000000000000000000000000005000000000000004d00000000",
            INIT_34 => X"0000000500000000000000010000000000000000000000000000000000000000",
            INIT_35 => X"00000044000000000000003c0000000000000031000000000000001f00000000",
            INIT_36 => X"0000005c00000000000000540000000000000054000000000000004e00000000",
            INIT_37 => X"0000002900000000000000320000000000000037000000000000003400000000",
            INIT_38 => X"00000019000000000000001b0000000000000022000000000000002200000000",
            INIT_39 => X"00000009000000000000000c000000000000000d000000000000001000000000",
            INIT_3A => X"0000000700000000000000000000000000000003000000000000000a00000000",
            INIT_3B => X"0000000200000000000000010000000000000001000000000000000300000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000006800000000000000620000000000000024000000000000000000000000",
            INIT_3F => X"0000006800000000000000650000000000000062000000000000005500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006b000000000000006c0000000000000069000000000000006600000000",
            INIT_41 => X"00000088000000000000007a000000000000006a000000000000006b00000000",
            INIT_42 => X"0000005c000000000000005b0000000000000058000000000000008300000000",
            INIT_43 => X"00000058000000000000005a0000000000000063000000000000006500000000",
            INIT_44 => X"0000006100000000000000610000000000000064000000000000006300000000",
            INIT_45 => X"0000007b00000000000000740000000000000071000000000000006c00000000",
            INIT_46 => X"0000007900000000000000590000000000000055000000000000005400000000",
            INIT_47 => X"00000098000000000000008c000000000000008e000000000000007e00000000",
            INIT_48 => X"0000009b00000000000000960000000000000097000000000000009600000000",
            INIT_49 => X"0000005500000000000000770000000000000076000000000000007900000000",
            INIT_4A => X"0000006a000000000000007c0000000000000057000000000000005300000000",
            INIT_4B => X"0000006800000000000000750000000000000073000000000000006c00000000",
            INIT_4C => X"0000008000000000000000650000000000000069000000000000006100000000",
            INIT_4D => X"000000550000000000000056000000000000006d000000000000006700000000",
            INIT_4E => X"0000004f00000000000000510000000000000058000000000000005d00000000",
            INIT_4F => X"000000520000000000000054000000000000005d000000000000004e00000000",
            INIT_50 => X"0000006e0000000000000075000000000000006f000000000000005d00000000",
            INIT_51 => X"00000048000000000000005a0000000000000062000000000000006900000000",
            INIT_52 => X"0000007900000000000000720000000000000073000000000000005a00000000",
            INIT_53 => X"0000007800000000000000720000000000000072000000000000007700000000",
            INIT_54 => X"0000006f000000000000006c0000000000000067000000000000007500000000",
            INIT_55 => X"0000002e000000000000003e0000000000000047000000000000006e00000000",
            INIT_56 => X"0000006d000000000000006b0000000000000059000000000000002f00000000",
            INIT_57 => X"00000069000000000000006c000000000000006b000000000000006e00000000",
            INIT_58 => X"0000007500000000000000690000000000000069000000000000006900000000",
            INIT_59 => X"00000042000000000000006c0000000000000075000000000000006d00000000",
            INIT_5A => X"0000006d000000000000006c0000000000000053000000000000003a00000000",
            INIT_5B => X"0000006b000000000000006a000000000000006d000000000000006800000000",
            INIT_5C => X"0000007b000000000000007c0000000000000067000000000000006900000000",
            INIT_5D => X"00000031000000000000001b0000000000000076000000000000007d00000000",
            INIT_5E => X"0000004f00000000000000390000000000000027000000000000002f00000000",
            INIT_5F => X"00000067000000000000006a000000000000006e000000000000006200000000",
            INIT_60 => X"0000007b000000000000007f000000000000007e000000000000006500000000",
            INIT_61 => X"0000002600000000000000130000000000000000000000000000007100000000",
            INIT_62 => X"000000030000000000000004000000000000002e000000000000003300000000",
            INIT_63 => X"000000680000000000000059000000000000003a000000000000001a00000000",
            INIT_64 => X"000000550000000000000079000000000000007b000000000000007700000000",
            INIT_65 => X"00000087000000000000004a000000000000005d000000000000006f00000000",
            INIT_66 => X"0000005c000000000000006f0000000000000060000000000000008a00000000",
            INIT_67 => X"00000041000000000000006e0000000000000083000000000000008e00000000",
            INIT_68 => X"00000028000000000000002c0000000000000031000000000000003a00000000",
            INIT_69 => X"0000002700000000000000470000000000000039000000000000001600000000",
            INIT_6A => X"0000003e0000000000000039000000000000003c000000000000002d00000000",
            INIT_6B => X"0000003400000000000000340000000000000031000000000000002a00000000",
            INIT_6C => X"0000002d00000000000000370000000000000035000000000000003400000000",
            INIT_6D => X"0000000e0000000000000012000000000000002a000000000000002d00000000",
            INIT_6E => X"0000000000000000000000030000000000000007000000000000000800000000",
            INIT_6F => X"0000000400000000000000090000000000000007000000000000000000000000",
            INIT_70 => X"00000010000000000000000d0000000000000014000000000000000f00000000",
            INIT_71 => X"0000001a00000000000000180000000000000018000000000000001500000000",
            INIT_72 => X"00000045000000000000001f000000000000001d000000000000001c00000000",
            INIT_73 => X"00000024000000000000001e000000000000001f000000000000001900000000",
            INIT_74 => X"00000033000000000000002b0000000000000028000000000000002000000000",
            INIT_75 => X"00000029000000000000002a000000000000002e000000000000002d00000000",
            INIT_76 => X"0000000100000000000000260000000000000052000000000000002b00000000",
            INIT_77 => X"0000001e000000000000002f000000000000004a000000000000002700000000",
            INIT_78 => X"0000002b00000000000000250000000000000031000000000000002a00000000",
            INIT_79 => X"0000001b000000000000002b000000000000002a000000000000002800000000",
            INIT_7A => X"0000002500000000000000080000000000000036000000000000002800000000",
            INIT_7B => X"0000004e000000000000002b0000000000000074000000000000004400000000",
            INIT_7C => X"00000053000000000000005b0000000000000048000000000000005d00000000",
            INIT_7D => X"0000003a000000000000002b0000000000000046000000000000005800000000",
            INIT_7E => X"0000004100000000000000290000000000000009000000000000003900000000",
            INIT_7F => X"0000003d000000000000001a0000000000000041000000000000006700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE25;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE26 : if BRAM_NAME = "samplegold_layersamples_instance26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000029000000000000002f000000000000002d000000000000001b00000000",
            INIT_01 => X"0000003800000000000000380000000000000033000000000000002700000000",
            INIT_02 => X"0000002700000000000000510000000000000028000000000000001100000000",
            INIT_03 => X"0000001d000000000000002b0000000000000025000000000000001f00000000",
            INIT_04 => X"00000026000000000000001b0000000000000039000000000000002500000000",
            INIT_05 => X"0000002600000000000000350000000000000035000000000000000000000000",
            INIT_06 => X"0000002c000000000000004c0000000000000033000000000000002700000000",
            INIT_07 => X"000000330000000000000027000000000000002b000000000000002f00000000",
            INIT_08 => X"00000038000000000000000c0000000000000026000000000000003700000000",
            INIT_09 => X"0000003f000000000000002b000000000000003a000000000000003700000000",
            INIT_0A => X"0000002f00000000000000310000000000000031000000000000004b00000000",
            INIT_0B => X"00000034000000000000003b0000000000000034000000000000002b00000000",
            INIT_0C => X"000000380000000000000039000000000000002e000000000000002d00000000",
            INIT_0D => X"0000004800000000000000590000000000000021000000000000003500000000",
            INIT_0E => X"000000360000000000000033000000000000001d000000000000001100000000",
            INIT_0F => X"0000003b00000000000000450000000000000040000000000000003d00000000",
            INIT_10 => X"00000039000000000000003c000000000000003c000000000000004000000000",
            INIT_11 => X"00000070000000000000004b000000000000003f000000000000001600000000",
            INIT_12 => X"0000003d000000000000001e0000000000000000000000000000002b00000000",
            INIT_13 => X"0000003d00000000000000380000000000000043000000000000004200000000",
            INIT_14 => X"000000180000000000000036000000000000003b000000000000003a00000000",
            INIT_15 => X"000000c1000000000000004e0000000000000043000000000000003c00000000",
            INIT_16 => X"0000003300000000000000080000000000000000000000000000000000000000",
            INIT_17 => X"0000003e000000000000003d0000000000000032000000000000004500000000",
            INIT_18 => X"0000003a0000000000000019000000000000003b000000000000003d00000000",
            INIT_19 => X"0000000500000000000000dc0000000000000055000000000000003e00000000",
            INIT_1A => X"0000001500000000000000080000000000000009000000000000000000000000",
            INIT_1B => X"0000003b00000000000000340000000000000026000000000000000000000000",
            INIT_1C => X"0000003d000000000000003c0000000000000013000000000000003a00000000",
            INIT_1D => X"00000000000000000000004a0000000000000031000000000000006f00000000",
            INIT_1E => X"000000000000000000000023000000000000001a000000000000000000000000",
            INIT_1F => X"00000021000000000000000a0000000000000000000000000000000000000000",
            INIT_20 => X"0000005200000000000000550000000000000054000000000000002c00000000",
            INIT_21 => X"00000024000000000000003f0000000000000068000000000000004e00000000",
            INIT_22 => X"0000003d00000000000000330000000000000045000000000000004500000000",
            INIT_23 => X"0000001d00000000000000370000000000000035000000000000003300000000",
            INIT_24 => X"0000002200000000000000260000000000000026000000000000002300000000",
            INIT_25 => X"0000003a000000000000001a0000000000000021000000000000002800000000",
            INIT_26 => X"0000003500000000000000300000000000000036000000000000003100000000",
            INIT_27 => X"0000001500000000000000240000000000000038000000000000004100000000",
            INIT_28 => X"0000000d0000000000000014000000000000000f000000000000001900000000",
            INIT_29 => X"0000000d000000000000000c0000000000000009000000000000000a00000000",
            INIT_2A => X"0000000000000000000000040000000000000005000000000000000300000000",
            INIT_2B => X"0000000500000000000000080000000000000021000000000000000000000000",
            INIT_2C => X"0000000500000000000000000000000000000008000000000000000000000000",
            INIT_2D => X"0000000700000000000000010000000000000007000000000000000000000000",
            INIT_2E => X"0000003300000000000000000000000000000000000000000000000400000000",
            INIT_2F => X"0000007d000000000000009e000000000000007f000000000000004600000000",
            INIT_30 => X"0000007c000000000000008a0000000000000087000000000000006700000000",
            INIT_31 => X"000000840000000000000085000000000000007f000000000000008100000000",
            INIT_32 => X"0000004a000000000000008d0000000000000085000000000000007600000000",
            INIT_33 => X"0000006e00000000000000b8000000000000009e000000000000007600000000",
            INIT_34 => X"0000008b000000000000007b000000000000008f000000000000007d00000000",
            INIT_35 => X"0000007a00000000000000730000000000000089000000000000008400000000",
            INIT_36 => X"00000077000000000000004d0000000000000094000000000000009500000000",
            INIT_37 => X"000000590000000000000080000000000000009c000000000000009a00000000",
            INIT_38 => X"000000710000000000000069000000000000004f000000000000007300000000",
            INIT_39 => X"000000950000000000000068000000000000005f000000000000006200000000",
            INIT_3A => X"000000b400000000000000730000000000000054000000000000009400000000",
            INIT_3B => X"0000008400000000000000770000000000000077000000000000008800000000",
            INIT_3C => X"0000007c000000000000009d000000000000007e000000000000007100000000",
            INIT_3D => X"0000008e0000000000000093000000000000004f000000000000008900000000",
            INIT_3E => X"0000009c000000000000008c0000000000000074000000000000006f00000000",
            INIT_3F => X"0000007300000000000000750000000000000077000000000000007500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005f00000000000000720000000000000085000000000000007d00000000",
            INIT_41 => X"0000007a000000000000008d000000000000008d000000000000008600000000",
            INIT_42 => X"000000800000000000000082000000000000008a000000000000008a00000000",
            INIT_43 => X"0000008b0000000000000087000000000000007b000000000000007f00000000",
            INIT_44 => X"0000008f000000000000007b000000000000007f000000000000008400000000",
            INIT_45 => X"000000ad0000000000000077000000000000008b000000000000009100000000",
            INIT_46 => X"0000007e00000000000000550000000000000047000000000000009d00000000",
            INIT_47 => X"0000009a00000000000000980000000000000095000000000000008c00000000",
            INIT_48 => X"0000009300000000000000910000000000000094000000000000008f00000000",
            INIT_49 => X"000000b000000000000000980000000000000070000000000000008f00000000",
            INIT_4A => X"0000005f000000000000001a000000000000004900000000000000c200000000",
            INIT_4B => X"00000090000000000000009c000000000000009a000000000000009200000000",
            INIT_4C => X"0000008a00000000000000920000000000000090000000000000009400000000",
            INIT_4D => X"000000af00000000000000a10000000000000097000000000000007100000000",
            INIT_4E => X"0000003e0000000000000016000000000000002300000000000000fc00000000",
            INIT_4F => X"00000095000000000000007e0000000000000084000000000000006b00000000",
            INIT_50 => X"00000072000000000000008d0000000000000093000000000000009400000000",
            INIT_51 => X"0000010f00000000000000b6000000000000009d000000000000009700000000",
            INIT_52 => X"0000002a000000000000002d000000000000001c000000000000001d00000000",
            INIT_53 => X"0000006a000000000000005c0000000000000020000000000000003e00000000",
            INIT_54 => X"0000009900000000000000690000000000000088000000000000007e00000000",
            INIT_55 => X"00000084000000000000009000000000000000cf000000000000009900000000",
            INIT_56 => X"0000005b00000000000000660000000000000000000000000000001f00000000",
            INIT_57 => X"000000550000000000000000000000000000003d000000000000003a00000000",
            INIT_58 => X"0000008d000000000000008d000000000000005d000000000000007600000000",
            INIT_59 => X"00000064000000000000009f0000000000000082000000000000008900000000",
            INIT_5A => X"0000006900000000000000830000000000000081000000000000004e00000000",
            INIT_5B => X"0000007900000000000000760000000000000067000000000000007800000000",
            INIT_5C => X"0000004d00000000000000500000000000000051000000000000004000000000",
            INIT_5D => X"00000033000000000000003c0000000000000046000000000000004700000000",
            INIT_5E => X"00000048000000000000004e000000000000004a000000000000005800000000",
            INIT_5F => X"0000003d000000000000004d000000000000005a000000000000004e00000000",
            INIT_60 => X"000000370000000000000031000000000000003e000000000000003800000000",
            INIT_61 => X"0000003000000000000000280000000000000029000000000000002b00000000",
            INIT_62 => X"0000002000000000000000240000000000000021000000000000002b00000000",
            INIT_63 => X"0000002500000000000000370000000000000000000000000000001f00000000",
            INIT_64 => X"000000180000000000000026000000000000001d000000000000002400000000",
            INIT_65 => X"000000230000000000000028000000000000001c000000000000002500000000",
            INIT_66 => X"0000000e00000000000000100000000000000022000000000000002400000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000004c00000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE26;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE27 : if BRAM_NAME = "samplegold_layersamples_instance27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000004d000000000000004d0000000000000034000000000000002a00000000",
            INIT_25 => X"0000003b00000000000000440000000000000047000000000000003c00000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_27 => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000500000000000000100000000000000000000000000000000f00000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000a00000000000000170000000000000000000000000000000000000000",
            INIT_2C => X"00000016000000000000000d0000000000000007000000000000000400000000",
            INIT_2D => X"00000000000000000000000a0000000000000013000000000000001f00000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000004000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000010000000000000003200000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000c000000000000000d0000000000000000000000000000000000000000",
            INIT_3F => X"00000015000000000000003b0000000000000052000000000000003900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000f00000000000000200000000000000043000000000000000000000000",
            INIT_43 => X"00000065000000000000004d000000000000001d000000000000000700000000",
            INIT_44 => X"0000000000000000000000030000000000000035000000000000005f00000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000003000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"000000580000000000000053000000000000004f000000000000004700000000",
            INIT_4A => X"0000003500000000000000290000000000000023000000000000003f00000000",
            INIT_4B => X"000000180000000000000009000000000000001a000000000000001700000000",
            INIT_4C => X"000000000000000000000000000000000000001f000000000000002500000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000002a00000000000000240000000000000014000000000000000000000000",
            INIT_4F => X"00000042000000000000003a0000000000000034000000000000003100000000",
            INIT_50 => X"0000002b0000000000000030000000000000002d000000000000004300000000",
            INIT_51 => X"00000019000000000000001c000000000000001f000000000000002200000000",
            INIT_52 => X"00000008000000000000000d000000000000000f000000000000001500000000",
            INIT_53 => X"0000000000000000000000000000000000000008000000000000000700000000",
            INIT_54 => X"0000000300000000000000040000000000000007000000000000000c00000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000b0000000000000012000000000000000a000000000000000500000000",
            INIT_61 => X"0000001300000000000000100000000000000011000000000000000e00000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_63 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000060000000000000029000000000000000200000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000230000000000000023000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000003c00000000000000260000000000000002000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_7C => X"00000018000000000000003f0000000000000045000000000000002000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE27;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE28 : if BRAM_NAME = "samplegold_layersamples_instance28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000004d000000000000004a0000000000000047000000000000003c00000000",
            INIT_02 => X"0000003e000000000000004a0000000000000046000000000000004f00000000",
            INIT_03 => X"0000002c000000000000002c0000000000000033000000000000002b00000000",
            INIT_04 => X"000000000000000000000022000000000000001d000000000000002300000000",
            INIT_05 => X"0000000d000000000000000a0000000000000003000000000000000000000000",
            INIT_06 => X"0000001900000000000000180000000000000013000000000000000e00000000",
            INIT_07 => X"00000020000000000000001e000000000000001c000000000000001b00000000",
            INIT_08 => X"0000000000000000000000000000000000000017000000000000002000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"00000007000000000000002f0000000000000000000000000000000c00000000",
            INIT_11 => X"000000040000000000000000000000000000004b000000000000000000000000",
            INIT_12 => X"0000004200000000000000000000000000000000000000000000000100000000",
            INIT_13 => X"0000000000000000000000100000000000000025000000000000000000000000",
            INIT_14 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_15 => X"00000000000000000000002c0000000000000000000000000000002500000000",
            INIT_16 => X"0000000000000000000000640000000000000000000000000000000d00000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000004700000000",
            INIT_18 => X"0000004900000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000020000000000000000000000000000002b00000000",
            INIT_1A => X"000000050000000000000000000000000000004c000000000000003f00000000",
            INIT_1B => X"0000000000000000000000720000000000000000000000000000000e00000000",
            INIT_1C => X"00000000000000000000004e0000000000000000000000000000000000000000",
            INIT_1D => X"0000005200000000000000000000000000000064000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000003a00000000",
            INIT_1F => X"0000000000000000000000000000000000000078000000000000000000000000",
            INIT_20 => X"0000005600000000000000000000000000000007000000000000004100000000",
            INIT_21 => X"000000000000000000000004000000000000002a000000000000000b00000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000004a00000000000000000000000000000000000000000000006b00000000",
            INIT_24 => X"00000000000000000000002f0000000000000000000000000000000600000000",
            INIT_25 => X"00000000000000000000003f0000000000000000000000000000000000000000",
            INIT_26 => X"0000004600000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_28 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_29 => X"0000001200000000000000000000000000000010000000000000000000000000",
            INIT_2A => X"00000017000000000000002d0000000000000000000000000000000000000000",
            INIT_2B => X"0000002300000000000000000000000000000013000000000000000000000000",
            INIT_2C => X"00000000000000000000000e0000000000000000000000000000000900000000",
            INIT_2D => X"0000000000000000000000010000000000000000000000000000000e00000000",
            INIT_2E => X"0000000000000000000000000000000000000015000000000000000a00000000",
            INIT_2F => X"0000000000000000000000030000000000000000000000000000000300000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000270000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000130000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000003900000000000000000000000000000031000000000000000200000000",
            INIT_36 => X"00000000000000000000000c0000000000000024000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000005600000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"00000000000000000000004c0000000000000025000000000000001800000000",
            INIT_3A => X"00000024000000000000001d0000000000000000000000000000001600000000",
            INIT_3B => X"0000001c00000000000000000000000000000000000000000000000100000000",
            INIT_3C => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_3D => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_3E => X"000000000000000000000000000000000000001b000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"000000000000000000000009000000000000003c000000000000000000000000",
            INIT_42 => X"0000002e00000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_44 => X"0000000500000000000000000000000000000012000000000000004c00000000",
            INIT_45 => X"0000000000000000000000000000000000000036000000000000004000000000",
            INIT_46 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_47 => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"00000065000000000000002f000000000000007c000000000000008300000000",
            INIT_49 => X"0000006200000000000000330000000000000012000000000000007100000000",
            INIT_4A => X"0000008100000000000000a2000000000000009c000000000000006600000000",
            INIT_4B => X"0000006a0000000000000057000000000000008600000000000000b800000000",
            INIT_4C => X"000000850000000000000087000000000000007700000000000000b500000000",
            INIT_4D => X"0000006900000000000000450000000000000021000000000000000400000000",
            INIT_4E => X"000000d400000000000000810000000000000095000000000000009b00000000",
            INIT_4F => X"0000007e00000000000000ad000000000000009b00000000000000c700000000",
            INIT_50 => X"00000000000000000000006b0000000000000084000000000000007500000000",
            INIT_51 => X"000000970000000000000079000000000000008c000000000000004900000000",
            INIT_52 => X"0000012500000000000000f90000000000000094000000000000004c00000000",
            INIT_53 => X"000000b4000000000000005200000000000000de00000000000000df00000000",
            INIT_54 => X"000000c000000000000000290000000000000057000000000000009300000000",
            INIT_55 => X"000000630000000000000080000000000000002500000000000000a800000000",
            INIT_56 => X"0000010b000000000000013f000000000000010d00000000000000d400000000",
            INIT_57 => X"000000dc000000000000010f000000000000006400000000000000b700000000",
            INIT_58 => X"0000007400000000000000eb0000000000000098000000000000005800000000",
            INIT_59 => X"000000f300000000000000df00000000000000d2000000000000006b00000000",
            INIT_5A => X"0000006d0000000000000119000000000000013100000000000000fb00000000",
            INIT_5B => X"000000ae000000000000013100000000000000f4000000000000004c00000000",
            INIT_5C => X"000000ff000000000000009e00000000000000db00000000000000db00000000",
            INIT_5D => X"000000fc00000000000000d700000000000000f000000000000000f900000000",
            INIT_5E => X"0000006a000000000000005e0000000000000118000000000000011e00000000",
            INIT_5F => X"000000e00000000000000127000000000000011700000000000000d400000000",
            INIT_60 => X"000000d000000000000000e700000000000000cb00000000000000dc00000000",
            INIT_61 => X"00000100000000000000010a00000000000000e600000000000000db00000000",
            INIT_62 => X"000000d7000000000000008c0000000000000086000000000000011b00000000",
            INIT_63 => X"000000a20000000000000120000000000000012300000000000000fd00000000",
            INIT_64 => X"000001060000000000000107000000000000010100000000000000f400000000",
            INIT_65 => X"000001050000000000000106000000000000012b00000000000000f300000000",
            INIT_66 => X"000000e400000000000000f700000000000000cb000000000000005500000000",
            INIT_67 => X"0000010400000000000000fc000000000000011c00000000000000fa00000000",
            INIT_68 => X"0000010e00000000000001260000000000000122000000000000011800000000",
            INIT_69 => X"0000006f00000000000000be00000000000000f8000000000000011300000000",
            INIT_6A => X"000000c3000000000000008c00000000000000cb00000000000000e800000000",
            INIT_6B => X"0000013e000000000000011e00000000000000ff00000000000000dc00000000",
            INIT_6C => X"0000010a000000000000010d000000000000013c000000000000013b00000000",
            INIT_6D => X"000000a700000000000000ca000000000000008600000000000000bf00000000",
            INIT_6E => X"000000d700000000000000d8000000000000009900000000000000bb00000000",
            INIT_6F => X"000001450000000000000164000000000000014400000000000000cc00000000",
            INIT_70 => X"000000d10000000000000102000000000000010d000000000000011a00000000",
            INIT_71 => X"00000165000000000000010b000000000000010800000000000000cc00000000",
            INIT_72 => X"000000fb00000000000000e000000000000000e600000000000000fa00000000",
            INIT_73 => X"0000010f00000000000001430000000000000152000000000000014000000000",
            INIT_74 => X"000000da00000000000000d20000000000000104000000000000012b00000000",
            INIT_75 => X"00000179000000000000016400000000000000f1000000000000010900000000",
            INIT_76 => X"0000012d000000000000010300000000000000eb000000000000012d00000000",
            INIT_77 => X"00000138000000000000012e00000000000000fb00000000000000de00000000",
            INIT_78 => X"000000e4000000000000009b00000000000000b400000000000000fc00000000",
            INIT_79 => X"0000017e000000000000013c0000000000000069000000000000008300000000",
            INIT_7A => X"000000d700000000000001020000000000000107000000000000014600000000",
            INIT_7B => X"000000e90000000000000128000000000000012700000000000000e800000000",
            INIT_7C => X"0000007900000000000000fa000000000000007b000000000000006200000000",
            INIT_7D => X"0000019000000000000001570000000000000087000000000000003100000000",
            INIT_7E => X"000000ca00000000000001230000000000000136000000000000017100000000",
            INIT_7F => X"0000008e00000000000000cd00000000000000df00000000000000e500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE28;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE29 : if BRAM_NAME = "samplegold_layersamples_instance29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000000000014200000000000000c100000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000001600000000000000100000000000000000000000000000000000000000",
            INIT_0F => X"0000002c00000000000000000000000000000000000000000000000200000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"00000013000000000000000b000000000000000d000000000000000000000000",
            INIT_13 => X"00000012000000000000003b0000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"00000000000000000000001b0000000000000000000000000000000400000000",
            INIT_17 => X"00000006000000000000002a0000000000000010000000000000000000000000",
            INIT_18 => X"0000000a0000000000000000000000000000000c000000000000000000000000",
            INIT_19 => X"0000000c00000000000000080000000000000018000000000000001000000000",
            INIT_1A => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_1B => X"00000007000000000000001b000000000000000c000000000000000b00000000",
            INIT_1C => X"00000004000000000000001d0000000000000021000000000000000000000000",
            INIT_1D => X"0000000000000000000000390000000000000012000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_1F => X"00000000000000000000004b0000000000000013000000000000001000000000",
            INIT_20 => X"0000002f000000000000001d0000000000000022000000000000002800000000",
            INIT_21 => X"0000000c000000000000002e0000000000000027000000000000001f00000000",
            INIT_22 => X"0000000000000000000000050000000000000009000000000000000000000000",
            INIT_23 => X"0000001d000000000000005e0000000000000004000000000000001000000000",
            INIT_24 => X"0000001f00000000000000260000000000000034000000000000002900000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_26 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_27 => X"0000003800000000000000570000000000000000000000000000000000000000",
            INIT_28 => X"0000001a00000000000000260000000000000031000000000000002d00000000",
            INIT_29 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000003900000000000000430000000000000038000000000000001900000000",
            INIT_2C => X"00000000000000000000001f0000000000000026000000000000001700000000",
            INIT_2D => X"00000068000000000000003b0000000000000000000000000000000e00000000",
            INIT_2E => X"0000002300000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"000000280000000000000053000000000000002e000000000000003200000000",
            INIT_30 => X"000000020000000000000000000000000000000c000000000000003b00000000",
            INIT_31 => X"0000005c00000000000000200000000000000000000000000000000000000000",
            INIT_32 => X"0000000300000000000000000000000000000000000000000000001200000000",
            INIT_33 => X"0000002c000000000000003e000000000000000f000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_35 => X"0000005500000000000000240000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_37 => X"00000007000000000000003c0000000000000038000000000000000700000000",
            INIT_38 => X"00000000000000000000002a0000000000000000000000000000000000000000",
            INIT_39 => X"0000000a00000000000000020000000000000000000000000000000b00000000",
            INIT_3A => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000100000000000000070000000000000005000000000000000000000000",
            INIT_3D => X"0000000000000000000000100000000000000003000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000016000000000000000800000000",
            INIT_42 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000700000000000000000000000000000000000000000000000100000000",
            INIT_45 => X"0000000800000000000000000000000000000000000000000000001100000000",
            INIT_46 => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_47 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"00000000000000000000000a0000000000000002000000000000000000000000",
            INIT_4C => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"00000003000000000000000a0000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_5F => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000003000000000000000100000000",
            INIT_71 => X"000000050000000000000016000000000000000c000000000000001300000000",
            INIT_72 => X"0000001b0000000000000015000000000000001f000000000000000000000000",
            INIT_73 => X"000000290000000000000009000000000000001d000000000000002300000000",
            INIT_74 => X"00000017000000000000000e0000000000000022000000000000000a00000000",
            INIT_75 => X"0000000000000000000000060000000000000011000000000000000f00000000",
            INIT_76 => X"00000015000000000000001a0000000000000010000000000000001f00000000",
            INIT_77 => X"0000000b0000000000000032000000000000000f000000000000001a00000000",
            INIT_78 => X"0000000d00000000000000130000000000000011000000000000002500000000",
            INIT_79 => X"0000001c0000000000000000000000000000000d000000000000000800000000",
            INIT_7A => X"0000000500000000000000120000000000000016000000000000001900000000",
            INIT_7B => X"00000014000000000000001a0000000000000039000000000000001900000000",
            INIT_7C => X"00000014000000000000001d0000000000000001000000000000001600000000",
            INIT_7D => X"000000130000000000000026000000000000000e000000000000000500000000",
            INIT_7E => X"0000003500000000000000000000000000000026000000000000000300000000",
            INIT_7F => X"0000000800000000000000190000000000000021000000000000002c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE29;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE30 : if BRAM_NAME = "samplegold_layersamples_instance30" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001d00000000000000000000000000000030000000000000000300000000",
            INIT_01 => X"0000001a00000000000000050000000000000020000000000000002300000000",
            INIT_02 => X"0000002f00000000000000290000000000000029000000000000002700000000",
            INIT_03 => X"0000000500000000000000000000000000000017000000000000002800000000",
            INIT_04 => X"0000002400000000000000000000000000000018000000000000003500000000",
            INIT_05 => X"0000001e00000000000000330000000000000032000000000000003000000000",
            INIT_06 => X"00000025000000000000002e0000000000000023000000000000002600000000",
            INIT_07 => X"0000002a00000000000000000000000000000000000000000000001700000000",
            INIT_08 => X"0000004a00000000000000390000000000000013000000000000002400000000",
            INIT_09 => X"0000004300000000000000390000000000000043000000000000003b00000000",
            INIT_0A => X"0000001d0000000000000022000000000000003a000000000000003d00000000",
            INIT_0B => X"00000014000000000000001e0000000000000006000000000000000000000000",
            INIT_0C => X"00000045000000000000003f000000000000002e000000000000002100000000",
            INIT_0D => X"000000460000000000000045000000000000004a000000000000004d00000000",
            INIT_0E => X"00000000000000000000001e0000000000000025000000000000004700000000",
            INIT_0F => X"0000001e000000000000001d0000000000000020000000000000001500000000",
            INIT_10 => X"0000004800000000000000540000000000000019000000000000004d00000000",
            INIT_11 => X"0000004700000000000000480000000000000045000000000000004700000000",
            INIT_12 => X"000000190000000000000000000000000000002e000000000000004700000000",
            INIT_13 => X"00000015000000000000001a0000000000000003000000000000001800000000",
            INIT_14 => X"0000004c000000000000003f000000000000003d000000000000005800000000",
            INIT_15 => X"000000240000000000000042000000000000003d000000000000004600000000",
            INIT_16 => X"0000001a00000000000000050000000000000023000000000000000c00000000",
            INIT_17 => X"0000000800000000000000240000000000000023000000000000001100000000",
            INIT_18 => X"000000450000000000000039000000000000004a000000000000005400000000",
            INIT_19 => X"0000002400000000000000360000000000000041000000000000004200000000",
            INIT_1A => X"0000001600000000000000340000000000000018000000000000001500000000",
            INIT_1B => X"000000440000000000000033000000000000000b000000000000002300000000",
            INIT_1C => X"0000004900000000000000370000000000000045000000000000004f00000000",
            INIT_1D => X"0000000d000000000000002c000000000000003d000000000000004a00000000",
            INIT_1E => X"0000002300000000000000260000000000000049000000000000003000000000",
            INIT_1F => X"0000004c0000000000000049000000000000002d000000000000001900000000",
            INIT_20 => X"0000003f0000000000000053000000000000003f000000000000004a00000000",
            INIT_21 => X"00000008000000000000000b000000000000002a000000000000003500000000",
            INIT_22 => X"00000026000000000000002c0000000000000043000000000000003500000000",
            INIT_23 => X"0000003d000000000000001b000000000000002e000000000000002100000000",
            INIT_24 => X"000000210000000000000046000000000000003e000000000000004c00000000",
            INIT_25 => X"0000000a00000000000000120000000000000012000000000000001500000000",
            INIT_26 => X"000000200000000000000035000000000000004e000000000000004b00000000",
            INIT_27 => X"0000004c00000000000000300000000000000023000000000000001b00000000",
            INIT_28 => X"0000001b000000000000000d000000000000002d000000000000004c00000000",
            INIT_29 => X"0000003a000000000000001c0000000000000026000000000000004000000000",
            INIT_2A => X"00000033000000000000004a0000000000000021000000000000003900000000",
            INIT_2B => X"0000002a000000000000003b000000000000004a000000000000003800000000",
            INIT_2C => X"0000002800000000000000450000000000000015000000000000004800000000",
            INIT_2D => X"0000003600000000000000300000000000000024000000000000002700000000",
            INIT_2E => X"00000044000000000000002e000000000000004a000000000000001800000000",
            INIT_2F => X"00000054000000000000002a000000000000003f000000000000002c00000000",
            INIT_30 => X"00000036000000000000002a000000000000003d000000000000000000000000",
            INIT_31 => X"00000012000000000000002e0000000000000029000000000000002900000000",
            INIT_32 => X"0000003500000000000000410000000000000040000000000000003e00000000",
            INIT_33 => X"00000016000000000000004e000000000000003e000000000000002f00000000",
            INIT_34 => X"0000004700000000000000250000000000000036000000000000003600000000",
            INIT_35 => X"0000005a000000000000001e000000000000001c000000000000003000000000",
            INIT_36 => X"0000000500000000000000590000000000000021000000000000005100000000",
            INIT_37 => X"0000002d00000000000000230000000000000054000000000000005300000000",
            INIT_38 => X"0000000a00000000000000570000000000000026000000000000002000000000",
            INIT_39 => X"00000019000000000000003e0000000000000037000000000000003100000000",
            INIT_3A => X"0000004f00000000000000460000000000000042000000000000003c00000000",
            INIT_3B => X"0000000a0000000000000029000000000000002c000000000000004900000000",
            INIT_3C => X"00000004000000000000002a000000000000005e000000000000001200000000",
            INIT_3D => X"0000002c00000000000000020000000000000034000000000000005700000000",
            INIT_3E => X"0000004400000000000000270000000000000039000000000000003000000000",
            INIT_3F => X"0000000c0000000000000000000000000000002e000000000000002900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000230000000000000028000000000000003f000000000000004e00000000",
            INIT_41 => X"0000001b00000000000000270000000000000005000000000000001600000000",
            INIT_42 => X"0000001300000000000000250000000000000006000000000000001000000000",
            INIT_43 => X"0000003e00000000000000220000000000000000000000000000003f00000000",
            INIT_44 => X"0000001000000000000000000000000000000031000000000000003600000000",
            INIT_45 => X"0000000b00000000000000000000000000000012000000000000001c00000000",
            INIT_46 => X"0000002700000000000000060000000000000005000000000000001a00000000",
            INIT_47 => X"00000030000000000000003f0000000000000026000000000000000c00000000",
            INIT_48 => X"000000190000000000000000000000000000003e000000000000003300000000",
            INIT_49 => X"00000005000000000000000f000000000000000f000000000000000000000000",
            INIT_4A => X"0000000400000000000000190000000000000012000000000000001400000000",
            INIT_4B => X"000000440000000000000026000000000000002a000000000000003300000000",
            INIT_4C => X"000000050000000000000000000000000000003d000000000000001e00000000",
            INIT_4D => X"0000000a00000000000000070000000000000002000000000000000800000000",
            INIT_4E => X"0000001c000000000000003e0000000000000020000000000000000000000000",
            INIT_4F => X"0000004b000000000000003c0000000000000024000000000000003600000000",
            INIT_50 => X"00000000000000000000000a0000000000000035000000000000001600000000",
            INIT_51 => X"0000000900000000000000060000000000000009000000000000000b00000000",
            INIT_52 => X"00000030000000000000001d000000000000003c000000000000001b00000000",
            INIT_53 => X"000000450000000000000021000000000000004b000000000000001d00000000",
            INIT_54 => X"000000000000000000000000000000000000000e000000000000002a00000000",
            INIT_55 => X"000000210000000000000011000000000000000a000000000000001100000000",
            INIT_56 => X"0000001d0000000000000043000000000000004f000000000000004000000000",
            INIT_57 => X"0000002e00000000000000360000000000000034000000000000003400000000",
            INIT_58 => X"0000000c00000000000000000000000000000017000000000000001200000000",
            INIT_59 => X"0000004f000000000000002e000000000000000a000000000000000000000000",
            INIT_5A => X"0000002b000000000000005d0000000000000066000000000000002d00000000",
            INIT_5B => X"0000000f00000000000000460000000000000040000000000000003400000000",
            INIT_5C => X"0000000900000000000000000000000000000016000000000000003e00000000",
            INIT_5D => X"00000028000000000000003a000000000000004c000000000000000000000000",
            INIT_5E => X"0000002700000000000000610000000000000081000000000000002a00000000",
            INIT_5F => X"0000003300000000000000490000000000000040000000000000003100000000",
            INIT_60 => X"0000000d0000000000000000000000000000001a000000000000002300000000",
            INIT_61 => X"00000010000000000000002c000000000000006f000000000000003e00000000",
            INIT_62 => X"0000002000000000000000280000000000000042000000000000002e00000000",
            INIT_63 => X"0000003f0000000000000044000000000000002a000000000000002d00000000",
            INIT_64 => X"0000002e000000000000002e000000000000003a000000000000003b00000000",
            INIT_65 => X"0000003c000000000000001f000000000000003e000000000000002600000000",
            INIT_66 => X"0000002d00000000000000240000000000000019000000000000004600000000",
            INIT_67 => X"00000038000000000000003a0000000000000036000000000000002e00000000",
            INIT_68 => X"0000003f000000000000002c000000000000002b000000000000004300000000",
            INIT_69 => X"0000003f000000000000003b0000000000000032000000000000004600000000",
            INIT_6A => X"00000040000000000000002f0000000000000019000000000000000f00000000",
            INIT_6B => X"00000048000000000000003b0000000000000036000000000000004300000000",
            INIT_6C => X"0000002f0000000000000052000000000000004d000000000000005100000000",
            INIT_6D => X"0000000a0000000000000027000000000000003c000000000000003b00000000",
            INIT_6E => X"000000400000000000000020000000000000004e000000000000004100000000",
            INIT_6F => X"0000006800000000000000510000000000000043000000000000001600000000",
            INIT_70 => X"0000006600000000000000320000000000000056000000000000005600000000",
            INIT_71 => X"000000490000000000000022000000000000002c000000000000004300000000",
            INIT_72 => X"0000003d00000000000000400000000000000018000000000000002a00000000",
            INIT_73 => X"00000062000000000000005b000000000000004b000000000000005300000000",
            INIT_74 => X"0000006800000000000000690000000000000022000000000000004100000000",
            INIT_75 => X"0000000b000000000000003b000000000000004a000000000000002700000000",
            INIT_76 => X"000000350000000000000043000000000000003d000000000000003700000000",
            INIT_77 => X"0000002c00000000000000690000000000000056000000000000003500000000",
            INIT_78 => X"0000005c00000000000000680000000000000055000000000000001c00000000",
            INIT_79 => X"0000002b00000000000000050000000000000014000000000000002e00000000",
            INIT_7A => X"0000002d0000000000000015000000000000001d000000000000002700000000",
            INIT_7B => X"00000038000000000000002e0000000000000061000000000000003b00000000",
            INIT_7C => X"0000002500000000000000620000000000000059000000000000005100000000",
            INIT_7D => X"0000000d000000000000001b0000000000000023000000000000000d00000000",
            INIT_7E => X"0000002d000000000000002e0000000000000023000000000000001200000000",
            INIT_7F => X"00000055000000000000003c0000000000000031000000000000005000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE30;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE31 : if BRAM_NAME = "samplegold_layersamples_instance31" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000013000000000000005c000000000000005d000000000000005b00000000",
            INIT_01 => X"0000002e0000000000000027000000000000001f000000000000002500000000",
            INIT_02 => X"00000038000000000000003d000000000000002f000000000000001f00000000",
            INIT_03 => X"0000004000000000000000510000000000000056000000000000002000000000",
            INIT_04 => X"0000002700000000000000550000000000000044000000000000005500000000",
            INIT_05 => X"0000002500000000000000310000000000000030000000000000003000000000",
            INIT_06 => X"00000046000000000000002c000000000000001d000000000000002900000000",
            INIT_07 => X"0000004f0000000000000036000000000000003c000000000000004900000000",
            INIT_08 => X"00000044000000000000004f0000000000000035000000000000005400000000",
            INIT_09 => X"0000002300000000000000290000000000000037000000000000003600000000",
            INIT_0A => X"0000003a000000000000005e0000000000000037000000000000002100000000",
            INIT_0B => X"000000520000000000000057000000000000002d000000000000004000000000",
            INIT_0C => X"0000003a000000000000003d000000000000004b000000000000005700000000",
            INIT_0D => X"000000160000000000000020000000000000002e000000000000002b00000000",
            INIT_0E => X"0000006f000000000000006a000000000000006d000000000000003400000000",
            INIT_0F => X"0000005700000000000000490000000000000043000000000000004c00000000",
            INIT_10 => X"0000002c00000000000000390000000000000031000000000000005000000000",
            INIT_11 => X"0000002e0000000000000014000000000000001d000000000000003500000000",
            INIT_12 => X"0000006b000000000000004a000000000000003c000000000000006b00000000",
            INIT_13 => X"0000005000000000000000480000000000000046000000000000005500000000",
            INIT_14 => X"00000029000000000000003b000000000000003a000000000000002e00000000",
            INIT_15 => X"0000005400000000000000390000000000000010000000000000002400000000",
            INIT_16 => X"00000069000000000000004d000000000000000f000000000000003600000000",
            INIT_17 => X"00000058000000000000004e000000000000004f000000000000005b00000000",
            INIT_18 => X"0000001e00000000000000360000000000000039000000000000003b00000000",
            INIT_19 => X"0000001c000000000000005f000000000000003d000000000000001500000000",
            INIT_1A => X"00000025000000000000001d000000000000001b000000000000002d00000000",
            INIT_1B => X"0000002800000000000000280000000000000026000000000000001c00000000",
            INIT_1C => X"000000370000000000000028000000000000002d000000000000002f00000000",
            INIT_1D => X"000000310000000000000027000000000000002b000000000000002200000000",
            INIT_1E => X"0000001b000000000000002d000000000000001b000000000000002700000000",
            INIT_1F => X"0000002600000000000000250000000000000025000000000000002400000000",
            INIT_20 => X"0000002000000000000000390000000000000022000000000000002b00000000",
            INIT_21 => X"000000270000000000000029000000000000001d000000000000001f00000000",
            INIT_22 => X"0000002b00000000000000210000000000000030000000000000002100000000",
            INIT_23 => X"0000001f000000000000002c0000000000000025000000000000002800000000",
            INIT_24 => X"000000240000000000000028000000000000002b000000000000002900000000",
            INIT_25 => X"0000002700000000000000280000000000000017000000000000002600000000",
            INIT_26 => X"0000004100000000000000380000000000000023000000000000003500000000",
            INIT_27 => X"00000034000000000000001f0000000000000034000000000000001e00000000",
            INIT_28 => X"0000002c00000000000000170000000000000028000000000000002e00000000",
            INIT_29 => X"0000002600000000000000290000000000000025000000000000000c00000000",
            INIT_2A => X"0000002a000000000000002e000000000000003d000000000000003300000000",
            INIT_2B => X"0000003600000000000000410000000000000035000000000000003200000000",
            INIT_2C => X"0000000c00000000000000300000000000000024000000000000001d00000000",
            INIT_2D => X"0000004400000000000000290000000000000035000000000000001f00000000",
            INIT_2E => X"00000045000000000000003a0000000000000023000000000000003d00000000",
            INIT_2F => X"0000001f00000000000000380000000000000039000000000000004200000000",
            INIT_30 => X"0000002400000000000000170000000000000030000000000000003000000000",
            INIT_31 => X"00000044000000000000003b0000000000000041000000000000002800000000",
            INIT_32 => X"000000330000000000000035000000000000003c000000000000003800000000",
            INIT_33 => X"000000360000000000000023000000000000003c000000000000003900000000",
            INIT_34 => X"0000001e0000000000000020000000000000001d000000000000002d00000000",
            INIT_35 => X"0000003b0000000000000030000000000000003f000000000000002f00000000",
            INIT_36 => X"00000029000000000000003b000000000000003e000000000000003b00000000",
            INIT_37 => X"0000002900000000000000380000000000000026000000000000003200000000",
            INIT_38 => X"000000240000000000000025000000000000002a000000000000002400000000",
            INIT_39 => X"0000003200000000000000320000000000000030000000000000002d00000000",
            INIT_3A => X"0000002d0000000000000035000000000000003e000000000000003600000000",
            INIT_3B => X"0000002b000000000000001e000000000000002f000000000000002900000000",
            INIT_3C => X"000000250000000000000021000000000000001a000000000000002b00000000",
            INIT_3D => X"0000002c00000000000000320000000000000027000000000000002a00000000",
            INIT_3E => X"0000002100000000000000300000000000000034000000000000003600000000",
            INIT_3F => X"0000003400000000000000250000000000000029000000000000002500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002200000000000000280000000000000028000000000000001c00000000",
            INIT_41 => X"00000030000000000000002e0000000000000028000000000000002c00000000",
            INIT_42 => X"00000014000000000000002f0000000000000039000000000000003800000000",
            INIT_43 => X"000000350000000000000049000000000000002d000000000000003300000000",
            INIT_44 => X"0000003300000000000000260000000000000022000000000000002a00000000",
            INIT_45 => X"00000035000000000000002b0000000000000030000000000000002d00000000",
            INIT_46 => X"00000020000000000000002b0000000000000032000000000000003d00000000",
            INIT_47 => X"0000004100000000000000520000000000000046000000000000002c00000000",
            INIT_48 => X"0000002a000000000000002c0000000000000026000000000000002700000000",
            INIT_49 => X"000000340000000000000039000000000000002b000000000000003000000000",
            INIT_4A => X"0000002c0000000000000028000000000000002b000000000000003700000000",
            INIT_4B => X"0000004900000000000000510000000000000049000000000000002b00000000",
            INIT_4C => X"0000002b0000000000000028000000000000003a000000000000003b00000000",
            INIT_4D => X"0000001f00000000000000350000000000000039000000000000002f00000000",
            INIT_4E => X"00000026000000000000002b000000000000002c000000000000003900000000",
            INIT_4F => X"00000049000000000000004b0000000000000044000000000000003200000000",
            INIT_50 => X"0000002200000000000000230000000000000042000000000000004600000000",
            INIT_51 => X"00000029000000000000002c0000000000000038000000000000003100000000",
            INIT_52 => X"00000005000000000000000a0000000000000000000000000000000000000000",
            INIT_53 => X"000000230000000000000000000000000000004b000000000000000000000000",
            INIT_54 => X"0000006d00000000000000000000000000000023000000000000000e00000000",
            INIT_55 => X"0000000000000000000000010000000000000045000000000000000000000000",
            INIT_56 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_57 => X"000000000000000000000031000000000000000d000000000000003f00000000",
            INIT_58 => X"0000000000000000000000870000000000000000000000000000001200000000",
            INIT_59 => X"0000001e00000000000000000000000000000000000000000000002100000000",
            INIT_5A => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000310000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000079000000000000002700000000",
            INIT_5D => X"0000000000000000000000470000000000000000000000000000000000000000",
            INIT_5E => X"00000000000000000000002a0000000000000000000000000000000000000000",
            INIT_5F => X"000000250000000000000000000000000000004c000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000004b00000000",
            INIT_61 => X"0000000000000000000000000000000000000073000000000000000000000000",
            INIT_62 => X"0000003000000000000000000000000000000005000000000000004100000000",
            INIT_63 => X"000000480000000000000000000000000000000d000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000002500000000000000000000000000000001000000000000008000000000",
            INIT_66 => X"0000000000000000000000230000000000000000000000000000001900000000",
            INIT_67 => X"0000000000000000000000500000000000000000000000000000000d00000000",
            INIT_68 => X"0000004300000000000000000000000000000000000000000000001100000000",
            INIT_69 => X"0000000b00000000000000000000000000000000000000000000003f00000000",
            INIT_6A => X"0000001000000000000000010000000000000005000000000000000000000000",
            INIT_6B => X"0000001800000000000000000000000000000010000000000000000700000000",
            INIT_6C => X"0000001f00000000000000370000000000000000000000000000000000000000",
            INIT_6D => X"0000002e00000000000000000000000000000000000000000000000300000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"00000000000000000000000c0000000000000000000000000000002f00000000",
            INIT_70 => X"000000120000000000000008000000000000000e000000000000000400000000",
            INIT_71 => X"00000002000000000000001b0000000000000000000000000000003900000000",
            INIT_72 => X"000000110000000000000000000000000000000d000000000000000100000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"00000015000000000000002f0000000000000000000000000000000000000000",
            INIT_75 => X"00000000000000000000000b0000000000000007000000000000004600000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000003700000000000000000000000000000026000000000000000000000000",
            INIT_78 => X"0000000000000000000000040000000000000024000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000005e00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_7C => X"0000003300000000000000250000000000000000000000000000001300000000",
            INIT_7D => X"0000000900000000000000000000000000000000000000000000000f00000000",
            INIT_7E => X"00000000000000000000001d0000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000072000000000000003600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE31;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE32 : if BRAM_NAME = "samplegold_layersamples_instance32" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000018000000000000002c000000000000000000000000",
            INIT_01 => X"0000000000000000000000040000000000000000000000000000005800000000",
            INIT_02 => X"000000000000000000000001000000000000002c000000000000000000000000",
            INIT_03 => X"0000000000000000000000060000000000000098000000000000006000000000",
            INIT_04 => X"0000002f00000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"000000000000000000000000000000000000000b000000000000001b00000000",
            INIT_06 => X"0000000000000000000000000000000000000022000000000000004100000000",
            INIT_07 => X"0000000000000000000000000000000000000088000000000000008000000000",
            INIT_08 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000006c00000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"00000002000000000000002a0000000000000010000000000000000c00000000",
            INIT_0D => X"0000000000000000000000220000000000000000000000000000000800000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"000000000000000000000020000000000000001c000000000000000000000000",
            INIT_10 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"00000005000000000000000f0000000000000003000000000000003300000000",
            INIT_13 => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000006000000000000001600000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000033000000000000000a00000000",
            INIT_18 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000003500000000",
            INIT_1D => X"0000000000000000000000000000000000000023000000000000000c00000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"000000000000000000000000000000000000000c000000000000000500000000",
            INIT_21 => X"000000000000000000000000000000000000001f000000000000000000000000",
            INIT_22 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000a00000000000000000000000000000000000000000000000100000000",
            INIT_24 => X"0000000400000000000000030000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000900000000000000000000000000000006000000000000000000000000",
            INIT_28 => X"0000002400000000000000000000000000000000000000000000001900000000",
            INIT_29 => X"000000000000000000000000000000000000002a000000000000002100000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"00000000000000000000003b0000000000000024000000000000000000000000",
            INIT_2C => X"0000001700000000000000160000000000000030000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000049000000000000001900000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000001000000000000000600000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_36 => X"0000001200000000000000070000000000000000000000000000000000000000",
            INIT_37 => X"000000000000000000000071000000000000004d000000000000000f00000000",
            INIT_38 => X"0000000e000000000000000a0000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000059000000000000004500000000",
            INIT_3A => X"00000013000000000000003f0000000000000000000000000000000000000000",
            INIT_3B => X"00000000000000000000007b0000000000000073000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"000000030000000000000000000000000000000a000000000000000000000000",
            INIT_3E => X"0000000100000000000000000000000000000011000000000000003500000000",
            INIT_3F => X"0000000000000000000000610000000000000047000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000280000000000000050000000000000003300000000",
            INIT_42 => X"0000002000000000000000340000000000000000000000000000000000000000",
            INIT_43 => X"0000003700000000000000000000000000000028000000000000003f00000000",
            INIT_44 => X"00000040000000000000004c000000000000003a000000000000003300000000",
            INIT_45 => X"0000002e00000000000000250000000000000064000000000000002600000000",
            INIT_46 => X"0000003000000000000000480000000000000046000000000000003400000000",
            INIT_47 => X"0000001100000000000000280000000000000000000000000000002f00000000",
            INIT_48 => X"00000027000000000000004e000000000000003e000000000000004600000000",
            INIT_49 => X"0000004400000000000000680000000000000037000000000000007700000000",
            INIT_4A => X"0000002300000000000000280000000000000021000000000000002b00000000",
            INIT_4B => X"0000003e0000000000000057000000000000003f000000000000000000000000",
            INIT_4C => X"0000008500000000000000370000000000000019000000000000002e00000000",
            INIT_4D => X"0000000e00000000000000540000000000000059000000000000006100000000",
            INIT_4E => X"00000025000000000000001b0000000000000042000000000000005e00000000",
            INIT_4F => X"0000005300000000000000000000000000000049000000000000007400000000",
            INIT_50 => X"00000058000000000000008c0000000000000074000000000000001a00000000",
            INIT_51 => X"0000007500000000000000260000000000000021000000000000006200000000",
            INIT_52 => X"0000006800000000000000600000000000000031000000000000003a00000000",
            INIT_53 => X"0000007a00000000000000650000000000000059000000000000001f00000000",
            INIT_54 => X"00000059000000000000006a000000000000006e000000000000006f00000000",
            INIT_55 => X"0000005a00000000000000650000000000000014000000000000000000000000",
            INIT_56 => X"000000510000000000000068000000000000007b000000000000003d00000000",
            INIT_57 => X"00000055000000000000006b0000000000000075000000000000008500000000",
            INIT_58 => X"00000000000000000000004e0000000000000067000000000000009500000000",
            INIT_59 => X"000000650000000000000062000000000000005f000000000000002b00000000",
            INIT_5A => X"00000073000000000000006d0000000000000077000000000000006d00000000",
            INIT_5B => X"000000880000000000000072000000000000006f000000000000005e00000000",
            INIT_5C => X"0000002c0000000000000014000000000000006e000000000000005a00000000",
            INIT_5D => X"0000007f00000000000000610000000000000066000000000000005300000000",
            INIT_5E => X"000000840000000000000086000000000000007a000000000000006400000000",
            INIT_5F => X"00000074000000000000007d0000000000000080000000000000008c00000000",
            INIT_60 => X"0000006e00000000000000520000000000000000000000000000005700000000",
            INIT_61 => X"00000065000000000000007d000000000000004d000000000000004900000000",
            INIT_62 => X"0000007e000000000000008d000000000000007e000000000000008c00000000",
            INIT_63 => X"0000003e00000000000000560000000000000084000000000000007900000000",
            INIT_64 => X"0000002a000000000000003a000000000000005c000000000000001900000000",
            INIT_65 => X"0000007e00000000000000670000000000000042000000000000004b00000000",
            INIT_66 => X"0000007a0000000000000085000000000000008a000000000000008e00000000",
            INIT_67 => X"000000580000000000000033000000000000003f000000000000007600000000",
            INIT_68 => X"00000051000000000000003a0000000000000053000000000000001e00000000",
            INIT_69 => X"000000900000000000000094000000000000004d000000000000006900000000",
            INIT_6A => X"0000006f00000000000000700000000000000070000000000000007e00000000",
            INIT_6B => X"0000006d000000000000006d000000000000004a000000000000005d00000000",
            INIT_6C => X"0000003f0000000000000068000000000000007300000000000000ba00000000",
            INIT_6D => X"00000077000000000000008b000000000000008f000000000000006b00000000",
            INIT_6E => X"00000064000000000000007e0000000000000089000000000000006e00000000",
            INIT_6F => X"000000730000000000000058000000000000004d000000000000005f00000000",
            INIT_70 => X"00000068000000000000005c000000000000008d000000000000009100000000",
            INIT_71 => X"0000007800000000000000570000000000000058000000000000008300000000",
            INIT_72 => X"00000043000000000000005a000000000000006c000000000000008800000000",
            INIT_73 => X"00000072000000000000003e0000000000000029000000000000005000000000",
            INIT_74 => X"0000006c00000000000000770000000000000095000000000000009200000000",
            INIT_75 => X"0000007b000000000000007e000000000000008b000000000000004b00000000",
            INIT_76 => X"0000004c000000000000004b0000000000000013000000000000006b00000000",
            INIT_77 => X"0000008d00000000000000680000000000000026000000000000002400000000",
            INIT_78 => X"00000077000000000000008e00000000000000a4000000000000009500000000",
            INIT_79 => X"000000400000000000000059000000000000005f000000000000005900000000",
            INIT_7A => X"0000000200000000000000b70000000000000052000000000000004500000000",
            INIT_7B => X"0000003e00000000000000000000000000000000000000000000001400000000",
            INIT_7C => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_7D => X"000000780000000000000000000000000000002d000000000000000000000000",
            INIT_7E => X"0000000d000000000000000d0000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000470000000000000000000000000000001000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE32;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE33 : if BRAM_NAME = "samplegold_layersamples_instance33" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000c0000000000000000000000000000000100000000",
            INIT_01 => X"00000000000000000000006e0000000000000000000000000000002e00000000",
            INIT_02 => X"0000000600000000000000100000000000000016000000000000001700000000",
            INIT_03 => X"000000000000000000000000000000000000003e000000000000001300000000",
            INIT_04 => X"0000000000000000000000320000000000000000000000000000000a00000000",
            INIT_05 => X"0000000e00000000000000020000000000000049000000000000000000000000",
            INIT_06 => X"0000002300000000000000150000000000000000000000000000002700000000",
            INIT_07 => X"0000004000000000000000170000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000036000000000000000000000000",
            INIT_09 => X"00000029000000000000005a0000000000000012000000000000003d00000000",
            INIT_0A => X"0000000000000000000000160000000000000050000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000059000000000000000400000000",
            INIT_0C => X"0000002500000000000000000000000000000009000000000000000000000000",
            INIT_0D => X"00000000000000000000004c000000000000008f000000000000001300000000",
            INIT_0E => X"0000000a00000000000000000000000000000051000000000000001400000000",
            INIT_0F => X"00000016000000000000001d0000000000000000000000000000002f00000000",
            INIT_10 => X"0000001000000000000000390000000000000000000000000000002900000000",
            INIT_11 => X"0000000000000000000000000000000000000038000000000000009500000000",
            INIT_12 => X"0000002000000000000000160000000000000035000000000000002800000000",
            INIT_13 => X"000000190000000000000014000000000000001a000000000000000b00000000",
            INIT_14 => X"0000007d00000000000000000000000000000037000000000000000700000000",
            INIT_15 => X"0000001200000000000000000000000000000000000000000000002900000000",
            INIT_16 => X"000000120000000000000000000000000000002b000000000000002300000000",
            INIT_17 => X"0000000a00000000000000100000000000000011000000000000002c00000000",
            INIT_18 => X"00000000000000000000007d000000000000000f000000000000004500000000",
            INIT_19 => X"000000000000000000000014000000000000001f000000000000000000000000",
            INIT_1A => X"0000001900000000000000260000000000000004000000000000004700000000",
            INIT_1B => X"000000410000000000000018000000000000002b000000000000001900000000",
            INIT_1C => X"0000002e0000000000000008000000000000004d000000000000003700000000",
            INIT_1D => X"0000000000000000000000190000000000000000000000000000002800000000",
            INIT_1E => X"0000003400000000000000210000000000000015000000000000002300000000",
            INIT_1F => X"000000070000000000000053000000000000002d000000000000002400000000",
            INIT_20 => X"0000002d00000000000000000000000000000059000000000000000000000000",
            INIT_21 => X"0000000000000000000000200000000000000000000000000000000000000000",
            INIT_22 => X"0000002700000000000000350000000000000036000000000000002f00000000",
            INIT_23 => X"00000000000000000000000d0000000000000035000000000000002b00000000",
            INIT_24 => X"0000000000000000000000440000000000000000000000000000000000000000",
            INIT_25 => X"0000002400000000000000000000000000000000000000000000003100000000",
            INIT_26 => X"0000002a00000000000000100000000000000043000000000000002e00000000",
            INIT_27 => X"0000000300000000000000170000000000000003000000000000003a00000000",
            INIT_28 => X"00000026000000000000002f000000000000003f000000000000000000000000",
            INIT_29 => X"00000003000000000000004b0000000000000013000000000000000000000000",
            INIT_2A => X"0000003b00000000000000420000000000000022000000000000002d00000000",
            INIT_2B => X"000000000000000000000030000000000000000b000000000000000000000000",
            INIT_2C => X"00000016000000000000003a000000000000001b000000000000000000000000",
            INIT_2D => X"0000001700000000000000000000000000000025000000000000000300000000",
            INIT_2E => X"0000000000000000000000710000000000000042000000000000002400000000",
            INIT_2F => X"0000000000000000000000080000000000000043000000000000000000000000",
            INIT_30 => X"0000001f000000000000002d0000000000000025000000000000000000000000",
            INIT_31 => X"00000029000000000000000d0000000000000021000000000000000c00000000",
            INIT_32 => X"0000000000000000000000000000000000000021000000000000003500000000",
            INIT_33 => X"0000001e00000000000000040000000000000030000000000000003300000000",
            INIT_34 => X"00000008000000000000002b0000000000000000000000000000005f00000000",
            INIT_35 => X"000000000000000000000066000000000000002e000000000000002b00000000",
            INIT_36 => X"0000003b0000000000000024000000000000000000000000000000bb00000000",
            INIT_37 => X"0000006200000000000000250000000000000038000000000000003700000000",
            INIT_38 => X"0000004800000000000000000000000000000023000000000000000000000000",
            INIT_39 => X"000000c300000000000000000000000000000065000000000000001b00000000",
            INIT_3A => X"0000003e000000000000004a000000000000004b000000000000000000000000",
            INIT_3B => X"0000000000000000000000530000000000000032000000000000003300000000",
            INIT_3C => X"00000056000000000000001d0000000000000033000000000000000f00000000",
            INIT_3D => X"0000003e00000000000000a80000000000000000000000000000001e00000000",
            INIT_3E => X"0000004900000000000000000000000000000055000000000000005a00000000",
            INIT_3F => X"0000005600000000000000000000000000000011000000000000004a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000630000000000000000000000000000005900000000",
            INIT_41 => X"000000a000000000000000580000000000000097000000000000000c00000000",
            INIT_42 => X"0000003e000000000000009f0000000000000000000000000000004f00000000",
            INIT_43 => X"00000000000000000000008a0000000000000043000000000000000000000000",
            INIT_44 => X"0000002a00000000000000500000000000000024000000000000003500000000",
            INIT_45 => X"0000006900000000000000cc000000000000005c000000000000007400000000",
            INIT_46 => X"0000000500000000000000910000000000000063000000000000000000000000",
            INIT_47 => X"000000570000000000000023000000000000005a000000000000004600000000",
            INIT_48 => X"0000008600000000000000000000000000000066000000000000005200000000",
            INIT_49 => X"00000000000000000000006600000000000000d4000000000000005600000000",
            INIT_4A => X"0000004f0000000000000070000000000000007b000000000000002a00000000",
            INIT_4B => X"0000004d000000000000005a0000000000000046000000000000005900000000",
            INIT_4C => X"0000003c000000000000007a0000000000000044000000000000004f00000000",
            INIT_4D => X"000000360000000000000014000000000000005d00000000000000bb00000000",
            INIT_4E => X"0000003e000000000000004e0000000000000079000000000000006800000000",
            INIT_4F => X"0000004d00000000000000540000000000000069000000000000005b00000000",
            INIT_50 => X"000000a9000000000000004d0000000000000091000000000000004c00000000",
            INIT_51 => X"000000540000000000000051000000000000002e000000000000003600000000",
            INIT_52 => X"00000068000000000000003a0000000000000099000000000000003300000000",
            INIT_53 => X"000000520000000000000077000000000000006a000000000000006100000000",
            INIT_54 => X"0000004500000000000000850000000000000059000000000000008600000000",
            INIT_55 => X"0000005b000000000000002b000000000000005e000000000000005f00000000",
            INIT_56 => X"0000006e00000000000000620000000000000067000000000000002800000000",
            INIT_57 => X"0000008f0000000000000074000000000000006b000000000000007e00000000",
            INIT_58 => X"0000001e000000000000008f000000000000000c000000000000003e00000000",
            INIT_59 => X"000000600000000000000026000000000000001a000000000000006100000000",
            INIT_5A => X"0000007f0000000000000087000000000000007d000000000000001600000000",
            INIT_5B => X"0000003600000000000000710000000000000074000000000000006a00000000",
            INIT_5C => X"0000009200000000000000470000000000000045000000000000004000000000",
            INIT_5D => X"0000004a00000000000000210000000000000074000000000000001f00000000",
            INIT_5E => X"0000005a000000000000008c0000000000000074000000000000007a00000000",
            INIT_5F => X"0000005f00000000000000320000000000000076000000000000007200000000",
            INIT_60 => X"0000008200000000000000ab0000000000000046000000000000004000000000",
            INIT_61 => X"00000087000000000000005a0000000000000035000000000000007000000000",
            INIT_62 => X"0000008300000000000000680000000000000079000000000000003a00000000",
            INIT_63 => X"0000006e00000000000000550000000000000014000000000000007e00000000",
            INIT_64 => X"0000009300000000000000860000000000000020000000000000000000000000",
            INIT_65 => X"000000070000000000000072000000000000005a000000000000006200000000",
            INIT_66 => X"0000009600000000000000820000000000000071000000000000005f00000000",
            INIT_67 => X"0000003200000000000000790000000000000039000000000000000000000000",
            INIT_68 => X"0000008d0000000000000092000000000000001f000000000000000000000000",
            INIT_69 => X"0000004e0000000000000068000000000000005f000000000000007e00000000",
            INIT_6A => X"00000024000000000000005e0000000000000073000000000000005f00000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE33;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE34 : if BRAM_NAME = "samplegold_layersamples_instance34" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000400000000000000010000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000004000000000000001500000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_2D => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"000000000000000000000000000000000000000b000000000000001400000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000007000000000000000b00000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000001c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"000000000000000000000000000000000000001d000000000000000000000000",
            INIT_42 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_43 => X"0000000b00000000000000000000000000000001000000000000000000000000",
            INIT_44 => X"0000001a00000000000000270000000000000005000000000000000200000000",
            INIT_45 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_47 => X"0000000300000000000000030000000000000000000000000000000000000000",
            INIT_48 => X"000000000000000000000000000000000000000c000000000000000800000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000600000000000000120000000000000018000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000900000000000000080000000000000000000000000000000000000000",
            INIT_4F => X"00000014000000000000000e0000000000000000000000000000000500000000",
            INIT_50 => X"00000002000000000000001c0000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000260000000000000049000000000000000000000000",
            INIT_53 => X"0000000000000000000000130000000000000010000000000000000700000000",
            INIT_54 => X"0000000000000000000000370000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"00000002000000000000000d0000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000040000000000000001f00000000",
            INIT_58 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000f000000000000003b000000000000001f000000000000000300000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000040000000000000012000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_7E => X"0000000c00000000000000000000000000000001000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE34;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE35 : if BRAM_NAME = "samplegold_layersamples_instance35" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_0A => X"0000001a0000000000000023000000000000000e000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_0E => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000a00000000000000030000000000000000000000000000000000000000",
            INIT_10 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_12 => X"0000002f000000000000001d0000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000800000000000000000000000000000029000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000016000000000000000d00000000",
            INIT_18 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_1A => X"0000000c00000000000000000000000000000014000000000000000000000000",
            INIT_1B => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000100000000000000140000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_24 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_26 => X"0000005a00000000000000000000000000000000000000000000000e00000000",
            INIT_27 => X"0000000000000000000000000000000000000028000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_29 => X"0000001300000000000000000000000000000000000000000000001900000000",
            INIT_2A => X"000000150000000000000072000000000000000b000000000000000000000000",
            INIT_2B => X"00000007000000000000000a0000000000000000000000000000000000000000",
            INIT_2C => X"0000001900000000000000450000000000000000000000000000000000000000",
            INIT_2D => X"00000010000000000000000d0000000000000000000000000000000000000000",
            INIT_2E => X"00000000000000000000005f0000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000026000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_31 => X"0000000000000000000000350000000000000008000000000000000000000000",
            INIT_32 => X"000000000000000000000000000000000000004a000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000003100000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000049000000000000003a00000000",
            INIT_36 => X"0000003b00000000000000000000000000000000000000000000005500000000",
            INIT_37 => X"00000000000000000000004b0000000000000000000000000000000000000000",
            INIT_38 => X"0000002800000000000000040000000000000000000000000000000000000000",
            INIT_39 => X"0000001f00000000000000000000000000000000000000000000006d00000000",
            INIT_3A => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000019000000000000000000000000",
            INIT_3C => X"00000055000000000000001b0000000000000005000000000000000000000000",
            INIT_3D => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_3E => X"0000001600000000000000180000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000700000000000000050000000000000027000000000000000c00000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_42 => X"0000000000000000000000190000000000000000000000000000000000000000",
            INIT_43 => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000300000000000000000000000000000002300000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_46 => X"000000020000000000000000000000000000001c000000000000001a00000000",
            INIT_47 => X"0000000500000000000000270000000000000004000000000000000000000000",
            INIT_48 => X"0000002000000000000000040000000000000000000000000000001800000000",
            INIT_49 => X"0000000500000000000000000000000000000008000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"000000000000000000000000000000000000000a000000000000000c00000000",
            INIT_4C => X"000000a000000000000000ac000000000000009d000000000000001000000000",
            INIT_4D => X"00000074000000000000008e00000000000000a000000000000000a300000000",
            INIT_4E => X"0000004600000000000000320000000000000050000000000000007700000000",
            INIT_4F => X"0000004000000000000000610000000000000043000000000000003e00000000",
            INIT_50 => X"000000bc00000000000000a900000000000000d300000000000000dc00000000",
            INIT_51 => X"0000008a000000000000008d00000000000000ae00000000000000bb00000000",
            INIT_52 => X"0000004b00000000000000410000000000000013000000000000005b00000000",
            INIT_53 => X"000000d0000000000000004f0000000000000061000000000000006d00000000",
            INIT_54 => X"000000d300000000000000cc00000000000000c600000000000000de00000000",
            INIT_55 => X"0000009f000000000000009a00000000000000ab00000000000000c700000000",
            INIT_56 => X"0000005c00000000000000520000000000000079000000000000006a00000000",
            INIT_57 => X"000000e600000000000000c50000000000000066000000000000005f00000000",
            INIT_58 => X"000000cd00000000000000dc00000000000000db00000000000000d000000000",
            INIT_59 => X"000000b700000000000000ac000000000000009c00000000000000b900000000",
            INIT_5A => X"00000058000000000000004a000000000000005a000000000000009a00000000",
            INIT_5B => X"000000df00000000000000dc00000000000000b5000000000000006c00000000",
            INIT_5C => X"000000c900000000000000d200000000000000e200000000000000dd00000000",
            INIT_5D => X"000000b000000000000000a9000000000000009300000000000000d200000000",
            INIT_5E => X"0000006c000000000000005e0000000000000051000000000000006400000000",
            INIT_5F => X"000000f000000000000000fb00000000000000e5000000000000009500000000",
            INIT_60 => X"000000c50000000000000100000000000000011700000000000000d500000000",
            INIT_61 => X"00000030000000000000009500000000000000af000000000000009800000000",
            INIT_62 => X"0000009500000000000000640000000000000047000000000000004300000000",
            INIT_63 => X"000000f100000000000000fb000000000000011d00000000000000fb00000000",
            INIT_64 => X"000000eb00000000000000d100000000000000f2000000000000012700000000",
            INIT_65 => X"0000002f000000000000001f000000000000008800000000000000ed00000000",
            INIT_66 => X"000000ee00000000000000700000000000000051000000000000004900000000",
            INIT_67 => X"0000013a000000000000014000000000000000f7000000000000010e00000000",
            INIT_68 => X"0000012e00000000000001370000000000000137000000000000010300000000",
            INIT_69 => X"00000097000000000000003c000000000000002200000000000000a800000000",
            INIT_6A => X"0000012000000000000000fc0000000000000087000000000000004100000000",
            INIT_6B => X"000000df0000000000000119000000000000012c00000000000000bc00000000",
            INIT_6C => X"0000004100000000000000ae00000000000000d600000000000000d000000000",
            INIT_6D => X"0000004900000000000000d20000000000000036000000000000000000000000",
            INIT_6E => X"0000006d000000000000013b00000000000000f8000000000000008f00000000",
            INIT_6F => X"000000e800000000000000ab000000000000010000000000000000c000000000",
            INIT_70 => X"0000000b000000000000000f000000000000001b000000000000007f00000000",
            INIT_71 => X"000000a600000000000000900000000000000104000000000000003a00000000",
            INIT_72 => X"0000001d0000000000000049000000000000010d00000000000000d800000000",
            INIT_73 => X"0000002b0000000000000085000000000000003e000000000000003400000000",
            INIT_74 => X"00000038000000000000001c0000000000000000000000000000000000000000",
            INIT_75 => X"000000bb000000000000009f00000000000000ce00000000000000e800000000",
            INIT_76 => X"0000004a000000000000005c00000000000000af00000000000000e100000000",
            INIT_77 => X"0000000000000000000000000000000000000035000000000000005e00000000",
            INIT_78 => X"00000065000000000000002e0000000000000000000000000000000000000000",
            INIT_79 => X"000000b500000000000000c300000000000000a200000000000000d100000000",
            INIT_7A => X"0000008d0000000000000083000000000000009500000000000000e600000000",
            INIT_7B => X"0000000000000000000000060000000000000021000000000000005a00000000",
            INIT_7C => X"0000007a00000000000000210000000000000021000000000000000000000000",
            INIT_7D => X"0000009100000000000000a800000000000000af000000000000009700000000",
            INIT_7E => X"0000008700000000000000b1000000000000008c000000000000008600000000",
            INIT_7F => X"0000006c0000000000000052000000000000005e000000000000007000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE35;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE36 : if BRAM_NAME = "samplegold_layersamples_instance36" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009f0000000000000066000000000000005e000000000000005b00000000",
            INIT_01 => X"000000a600000000000000a900000000000000a400000000000000b900000000",
            INIT_02 => X"00000082000000000000008d000000000000009900000000000000b600000000",
            INIT_03 => X"0000009500000000000000a30000000000000088000000000000006f00000000",
            INIT_04 => X"0000000000000000000000000000000000000071000000000000007b00000000",
            INIT_05 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000003000000000000000200000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000b00000000000000030000000000000013000000000000000000000000",
            INIT_0D => X"0000000300000000000000000000000000000003000000000000000a00000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_10 => X"000000110000000000000012000000000000000c000000000000001500000000",
            INIT_11 => X"000000100000000000000000000000000000000a000000000000000a00000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_13 => X"00000015000000000000000f0000000000000000000000000000000000000000",
            INIT_14 => X"0000000a0000000000000010000000000000000c000000000000000d00000000",
            INIT_15 => X"0000002000000000000000000000000000000000000000000000000700000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_17 => X"0000001900000000000000030000000000000035000000000000000000000000",
            INIT_18 => X"00000004000000000000001d000000000000000b000000000000001100000000",
            INIT_19 => X"0000000500000000000000130000000000000000000000000000003500000000",
            INIT_1A => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000001100000000000000220000000000000038000000000000002a00000000",
            INIT_1C => X"0000000000000000000000170000000000000031000000000000000d00000000",
            INIT_1D => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"000000310000000000000023000000000000001f000000000000004900000000",
            INIT_20 => X"0000002f0000000000000037000000000000000c000000000000001b00000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_22 => X"0000003500000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000003f000000000000004a0000000000000006000000000000002300000000",
            INIT_24 => X"00000039000000000000003c000000000000003e000000000000001a00000000",
            INIT_25 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000003400000000000000480000000000000000000000000000000000000000",
            INIT_27 => X"000000020000000000000038000000000000006b000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_29 => X"00000000000000000000003f0000000000000000000000000000000000000000",
            INIT_2A => X"000000000000000000000034000000000000003c000000000000000800000000",
            INIT_2B => X"0000004800000000000000150000000000000026000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000001200000000000000000000000000000058000000000000000000000000",
            INIT_2E => X"000000000000000000000000000000000000001f000000000000001c00000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000001c000000000000000f0000000000000023000000000000002300000000",
            INIT_32 => X"0000000000000000000000000000000000000038000000000000001100000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000d00000000000000320000000000000011000000000000002400000000",
            INIT_36 => X"0000002200000000000000000000000000000000000000000000000b00000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000c00000000000000090000000000000015000000000000000e00000000",
            INIT_3A => X"0000001400000000000000110000000000000010000000000000000000000000",
            INIT_3B => X"0000000b00000000000000040000000000000001000000000000000300000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000300000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000003000000000000000a00000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"00000007000000000000000f0000000000000002000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000700000000000000010000000000000000000000000000000900000000",
            INIT_64 => X"0000000600000000000000040000000000000001000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_68 => X"00000007000000000000000e0000000000000012000000000000000d00000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"00000000000000000000000e000000000000000e000000000000000c00000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000007600000000000000770000000000000068000000000000005600000000",
            INIT_76 => X"00000068000000000000006d0000000000000078000000000000007700000000",
            INIT_77 => X"0000003e00000000000000480000000000000046000000000000004a00000000",
            INIT_78 => X"00000066000000000000003d0000000000000051000000000000004200000000",
            INIT_79 => X"0000007e000000000000007b0000000000000074000000000000006d00000000",
            INIT_7A => X"0000005d000000000000007a0000000000000080000000000000008000000000",
            INIT_7B => X"000000590000000000000053000000000000004a000000000000003f00000000",
            INIT_7C => X"0000006a000000000000005c000000000000004d000000000000005000000000",
            INIT_7D => X"00000083000000000000007f000000000000007e000000000000007600000000",
            INIT_7E => X"00000048000000000000007b0000000000000089000000000000007c00000000",
            INIT_7F => X"0000005a00000000000000600000000000000059000000000000006000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE36;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE37 : if BRAM_NAME = "samplegold_layersamples_instance37" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007600000000000000730000000000000055000000000000005300000000",
            INIT_01 => X"0000008600000000000000890000000000000082000000000000007f00000000",
            INIT_02 => X"00000070000000000000007c000000000000007e000000000000007b00000000",
            INIT_03 => X"0000005800000000000000580000000000000052000000000000005500000000",
            INIT_04 => X"0000007d00000000000000770000000000000068000000000000005600000000",
            INIT_05 => X"0000006400000000000000680000000000000084000000000000008400000000",
            INIT_06 => X"000000490000000000000071000000000000007e000000000000006500000000",
            INIT_07 => X"0000005800000000000000560000000000000058000000000000005300000000",
            INIT_08 => X"0000007800000000000000780000000000000072000000000000006500000000",
            INIT_09 => X"0000005100000000000000630000000000000049000000000000006b00000000",
            INIT_0A => X"0000004c00000000000000370000000000000059000000000000006600000000",
            INIT_0B => X"0000006d000000000000006a0000000000000057000000000000004f00000000",
            INIT_0C => X"0000006800000000000000620000000000000062000000000000006d00000000",
            INIT_0D => X"00000054000000000000004d0000000000000038000000000000005500000000",
            INIT_0E => X"0000004c00000000000000390000000000000028000000000000003d00000000",
            INIT_0F => X"0000006100000000000000750000000000000055000000000000005300000000",
            INIT_10 => X"0000006e00000000000000630000000000000064000000000000006900000000",
            INIT_11 => X"000000350000000000000051000000000000005a000000000000006a00000000",
            INIT_12 => X"00000043000000000000004f000000000000003c000000000000002c00000000",
            INIT_13 => X"00000055000000000000005f0000000000000074000000000000006600000000",
            INIT_14 => X"00000072000000000000005e0000000000000062000000000000005d00000000",
            INIT_15 => X"000000240000000000000034000000000000005c000000000000006200000000",
            INIT_16 => X"0000006100000000000000210000000000000060000000000000004000000000",
            INIT_17 => X"0000007300000000000000250000000000000054000000000000007500000000",
            INIT_18 => X"0000005b000000000000006c0000000000000050000000000000006800000000",
            INIT_19 => X"0000004a0000000000000034000000000000002b000000000000003300000000",
            INIT_1A => X"0000007300000000000000680000000000000019000000000000006d00000000",
            INIT_1B => X"0000003e00000000000000300000000000000023000000000000005400000000",
            INIT_1C => X"0000003000000000000000440000000000000077000000000000004300000000",
            INIT_1D => X"000000730000000000000048000000000000003b000000000000003000000000",
            INIT_1E => X"00000056000000000000006a000000000000006d000000000000002b00000000",
            INIT_1F => X"0000005d00000000000000470000000000000055000000000000004200000000",
            INIT_20 => X"00000019000000000000001a000000000000001a000000000000004700000000",
            INIT_21 => X"00000051000000000000005c0000000000000043000000000000002a00000000",
            INIT_22 => X"0000006a000000000000005d0000000000000072000000000000006f00000000",
            INIT_23 => X"0000004d00000000000000620000000000000063000000000000005800000000",
            INIT_24 => X"0000002000000000000000190000000000000024000000000000003200000000",
            INIT_25 => X"00000066000000000000005c0000000000000039000000000000003e00000000",
            INIT_26 => X"00000044000000000000005b0000000000000065000000000000007100000000",
            INIT_27 => X"00000053000000000000005d0000000000000074000000000000005c00000000",
            INIT_28 => X"0000004a00000000000000520000000000000049000000000000004900000000",
            INIT_29 => X"0000006f0000000000000066000000000000004f000000000000005500000000",
            INIT_2A => X"00000072000000000000005f000000000000006e000000000000006700000000",
            INIT_2B => X"000000630000000000000067000000000000006e000000000000007500000000",
            INIT_2C => X"0000005c00000000000000660000000000000070000000000000006c00000000",
            INIT_2D => X"00000004000000000000001f0000000000000000000000000000005a00000000",
            INIT_2E => X"0000000000000000000000090000000000000002000000000000000300000000",
            INIT_2F => X"00000009000000000000000d0000000000000000000000000000000a00000000",
            INIT_30 => X"000000000000000000000012000000000000000e000000000000000700000000",
            INIT_31 => X"0000000900000000000000010000000000000007000000000000000600000000",
            INIT_32 => X"0000000000000000000000000000000000000003000000000000000300000000",
            INIT_33 => X"000000090000000000000018000000000000000a000000000000000000000000",
            INIT_34 => X"0000000200000000000000030000000000000000000000000000000500000000",
            INIT_35 => X"0000000300000000000000060000000000000009000000000000001700000000",
            INIT_36 => X"00000000000000000000000b0000000000000000000000000000000300000000",
            INIT_37 => X"000000090000000000000000000000000000000f000000000000000000000000",
            INIT_38 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000090000000000000007000000000000000700000000",
            INIT_3A => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_3B => X"0000000c00000000000000010000000000000000000000000000000000000000",
            INIT_3C => X"0000000a00000000000000110000000000000004000000000000000500000000",
            INIT_3D => X"0000000000000000000000000000000000000009000000000000000900000000",
            INIT_3E => X"00000000000000000000000a0000000000000003000000000000000000000000",
            INIT_3F => X"0000000500000000000000070000000000000013000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000600000000000000150000000000000003000000000000002900000000",
            INIT_41 => X"0000001300000000000000000000000000000003000000000000000800000000",
            INIT_42 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_43 => X"00000050000000000000000e000000000000000c000000000000001e00000000",
            INIT_44 => X"0000000400000000000000000000000000000006000000000000000a00000000",
            INIT_45 => X"0000001200000000000000000000000000000000000000000000001900000000",
            INIT_46 => X"0000001c00000000000000000000000000000000000000000000001200000000",
            INIT_47 => X"000000290000000000000002000000000000000e000000000000001500000000",
            INIT_48 => X"00000000000000000000000f0000000000000005000000000000000000000000",
            INIT_49 => X"0000000000000000000000050000000000000003000000000000000000000000",
            INIT_4A => X"0000000d00000000000000190000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000080000000000000025000000000000000000000000",
            INIT_4D => X"00000000000000000000000e000000000000000b000000000000001600000000",
            INIT_4E => X"000000000000000000000020000000000000002f000000000000000700000000",
            INIT_4F => X"000000000000000000000000000000000000001f000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000013000000000000003c00000000",
            INIT_51 => X"0000000c00000000000000040000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000024000000000000002400000000",
            INIT_53 => X"0000002f00000000000000000000000000000007000000000000000e00000000",
            INIT_54 => X"00000000000000000000002a0000000000000007000000000000002c00000000",
            INIT_55 => X"0000001a000000000000000e000000000000001d000000000000000600000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000002d00000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000001a000000000000000a0000000000000000000000000000000800000000",
            INIT_59 => X"0000002600000000000000230000000000000032000000000000001800000000",
            INIT_5A => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_5C => X"0000001300000000000000070000000000000000000000000000000000000000",
            INIT_5D => X"000000350000000000000009000000000000002b000000000000001f00000000",
            INIT_5E => X"0000000400000000000000000000000000000001000000000000000000000000",
            INIT_5F => X"0000000000000000000000080000000000000007000000000000000000000000",
            INIT_60 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000040000000000000000000000000000000f00000000",
            INIT_7D => X"000000000000000000000006000000000000001c000000000000000000000000",
            INIT_7E => X"000000000000000000000000000000000000000d000000000000000800000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE37;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE38 : if BRAM_NAME = "samplegold_layersamples_instance38" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001200000000000000000000000000000003000000000000000800000000",
            INIT_01 => X"0000002500000000000000140000000000000000000000000000000700000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000001200000000000000330000000000000000000000000000000800000000",
            INIT_05 => X"000000140000000000000011000000000000000d000000000000000000000000",
            INIT_06 => X"0000000e00000000000000000000000000000000000000000000000100000000",
            INIT_07 => X"0000002200000000000000060000000000000000000000000000000000000000",
            INIT_08 => X"000000000000000000000010000000000000002c000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000500000000000000150000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_0C => X"000000070000000000000000000000000000001b000000000000000200000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"000000000000000000000015000000000000001a000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_12 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000006400000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000005d0000000000000052000000000000005b000000000000005300000000",
            INIT_1F => X"0000004d00000000000000580000000000000061000000000000005d00000000",
            INIT_20 => X"0000003b00000000000000390000000000000035000000000000003900000000",
            INIT_21 => X"000000570000000000000053000000000000003a000000000000003500000000",
            INIT_22 => X"00000062000000000000005f000000000000005c000000000000006200000000",
            INIT_23 => X"0000004200000000000000610000000000000061000000000000006600000000",
            INIT_24 => X"0000003c0000000000000039000000000000003a000000000000003000000000",
            INIT_25 => X"0000005d000000000000004d000000000000004f000000000000003e00000000",
            INIT_26 => X"000000670000000000000069000000000000005e000000000000006000000000",
            INIT_27 => X"00000048000000000000005c0000000000000067000000000000006300000000",
            INIT_28 => X"0000003d000000000000003e0000000000000039000000000000004800000000",
            INIT_29 => X"0000005e000000000000005c000000000000004b000000000000005400000000",
            INIT_2A => X"0000006000000000000000640000000000000069000000000000006300000000",
            INIT_2B => X"00000053000000000000005e0000000000000060000000000000005700000000",
            INIT_2C => X"00000047000000000000003c000000000000003c000000000000003e00000000",
            INIT_2D => X"0000006300000000000000610000000000000058000000000000004d00000000",
            INIT_2E => X"0000004e00000000000000440000000000000048000000000000005b00000000",
            INIT_2F => X"0000003800000000000000490000000000000053000000000000004d00000000",
            INIT_30 => X"000000530000000000000037000000000000003a000000000000003a00000000",
            INIT_31 => X"0000004f000000000000005b0000000000000058000000000000005000000000",
            INIT_32 => X"00000038000000000000003e0000000000000032000000000000003700000000",
            INIT_33 => X"0000003a000000000000002b0000000000000041000000000000003e00000000",
            INIT_34 => X"0000004a00000000000000460000000000000023000000000000003900000000",
            INIT_35 => X"0000005500000000000000410000000000000051000000000000004a00000000",
            INIT_36 => X"0000003e0000000000000034000000000000002e000000000000004500000000",
            INIT_37 => X"0000003500000000000000390000000000000029000000000000003600000000",
            INIT_38 => X"0000004a00000000000000470000000000000030000000000000004300000000",
            INIT_39 => X"000000410000000000000056000000000000004c000000000000003f00000000",
            INIT_3A => X"00000031000000000000003c000000000000003b000000000000003a00000000",
            INIT_3B => X"0000004a000000000000003b0000000000000034000000000000002b00000000",
            INIT_3C => X"0000002a00000000000000480000000000000040000000000000003100000000",
            INIT_3D => X"0000003e00000000000000410000000000000047000000000000004c00000000",
            INIT_3E => X"0000002900000000000000310000000000000039000000000000003700000000",
            INIT_3F => X"0000003700000000000000480000000000000039000000000000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000031000000000000001d000000000000003e000000000000003200000000",
            INIT_41 => X"0000003a000000000000004a0000000000000039000000000000004d00000000",
            INIT_42 => X"0000002d000000000000002b000000000000002b000000000000002f00000000",
            INIT_43 => X"00000034000000000000003c0000000000000047000000000000003300000000",
            INIT_44 => X"0000002f00000000000000280000000000000026000000000000004b00000000",
            INIT_45 => X"00000022000000000000002e000000000000003d000000000000002c00000000",
            INIT_46 => X"00000036000000000000002a000000000000002f000000000000002900000000",
            INIT_47 => X"0000004d000000000000003c000000000000003d000000000000004e00000000",
            INIT_48 => X"0000003600000000000000410000000000000047000000000000005300000000",
            INIT_49 => X"00000016000000000000001c0000000000000025000000000000002e00000000",
            INIT_4A => X"0000004900000000000000370000000000000031000000000000002b00000000",
            INIT_4B => X"0000004b00000000000000420000000000000042000000000000004900000000",
            INIT_4C => X"0000003f0000000000000049000000000000003e000000000000003e00000000",
            INIT_4D => X"00000024000000000000002b000000000000002f000000000000003100000000",
            INIT_4E => X"0000003e000000000000003c0000000000000026000000000000003600000000",
            INIT_4F => X"0000004100000000000000430000000000000044000000000000004700000000",
            INIT_50 => X"000000420000000000000045000000000000004b000000000000003f00000000",
            INIT_51 => X"0000004000000000000000460000000000000042000000000000004600000000",
            INIT_52 => X"0000004a0000000000000040000000000000004a000000000000003b00000000",
            INIT_53 => X"0000004800000000000000470000000000000048000000000000004700000000",
            INIT_54 => X"0000004400000000000000480000000000000047000000000000004600000000",
            INIT_55 => X"000000450000000000000047000000000000004b000000000000004800000000",
            INIT_56 => X"0000000100000000000000000000000000000003000000000000000000000000",
            INIT_57 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000090000000000000008000000000000000000000000",
            INIT_59 => X"000000000000000000000000000000000000001a000000000000000400000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"00000011000000000000000d0000000000000024000000000000000000000000",
            INIT_5D => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_60 => X"0000000800000000000000080000000000000000000000000000000600000000",
            INIT_61 => X"00000000000000000000000e0000000000000000000000000000000200000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_63 => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_64 => X"0000000900000000000000130000000000000000000000000000000000000000",
            INIT_65 => X"0000000300000000000000000000000000000011000000000000001200000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000060000000000000028000000000000000000000000",
            INIT_68 => X"0000009b000000000000000c0000000000000009000000000000001b00000000",
            INIT_69 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_6A => X"0000000000000000000000030000000000000000000000000000002200000000",
            INIT_6B => X"0000002500000000000000000000000000000000000000000000002100000000",
            INIT_6C => X"00000046000000000000007a0000000000000017000000000000000a00000000",
            INIT_6D => X"0000000d000000000000000e0000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000d00000000000000180000000000000000000000000000000000000000",
            INIT_70 => X"00000000000000000000007e0000000000000000000000000000000b00000000",
            INIT_71 => X"0000000000000000000000000000000000000029000000000000000600000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_73 => X"000000000000000000000016000000000000002c000000000000000000000000",
            INIT_74 => X"000000000000000000000000000000000000005b000000000000000000000000",
            INIT_75 => X"0000001e00000000000000000000000000000033000000000000003700000000",
            INIT_76 => X"000000000000000000000000000000000000000f000000000000002000000000",
            INIT_77 => X"0000000000000000000000000000000000000047000000000000005400000000",
            INIT_78 => X"0000009600000000000000000000000000000000000000000000006800000000",
            INIT_79 => X"0000000000000000000000230000000000000000000000000000003100000000",
            INIT_7A => X"0000004700000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000004a00000000000000000000000000000000000000000000006d00000000",
            INIT_7C => X"0000003c000000000000002d0000000000000000000000000000000000000000",
            INIT_7D => X"000000000000000000000000000000000000004b000000000000002400000000",
            INIT_7E => X"0000009000000000000000220000000000000017000000000000001200000000",
            INIT_7F => X"00000014000000000000000e0000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE38;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE39 : if BRAM_NAME = "samplegold_layersamples_instance39" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_02 => X"0000001700000000000000490000000000000048000000000000002b00000000",
            INIT_03 => X"0000002d00000000000000020000000000000000000000000000000b00000000",
            INIT_04 => X"00000000000000000000000c0000000000000000000000000000000000000000",
            INIT_05 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000350000000000000015000000000000002a00000000",
            INIT_07 => X"00000000000000000000001d0000000000000000000000000000003a00000000",
            INIT_08 => X"0000000000000000000000000000000000000023000000000000000700000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000001000000000000000000000000000000000000000000000000200000000",
            INIT_0B => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000009000000000000000a00000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000600000000000000090000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000050000000000000000000000000000000700000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000018000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000400000000000000100000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000090000000000000008000000000000000100000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000003100000000",
            INIT_22 => X"0000003300000000000000000000000000000000000000000000000900000000",
            INIT_23 => X"0000002100000000000000050000000000000000000000000000001e00000000",
            INIT_24 => X"0000000000000000000000010000000000000006000000000000000c00000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_26 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000800000000000000000000000000000003000000000000000000000000",
            INIT_29 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"00000000000000000000000a0000000000000005000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000240000000000000019000000000000000b00000000",
            INIT_2E => X"0000007000000000000000640000000000000043000000000000004d00000000",
            INIT_2F => X"0000000000000000000000000000000000000003000000000000002400000000",
            INIT_30 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_31 => X"000000000000000000000018000000000000001e000000000000007500000000",
            INIT_32 => X"0000000000000000000000000000000000000025000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_34 => X"00000000000000000000000b0000000000000017000000000000001500000000",
            INIT_35 => X"00000057000000000000004b000000000000004e000000000000006900000000",
            INIT_36 => X"000000000000000000000016000000000000002e000000000000002100000000",
            INIT_37 => X"00000000000000000000000c0000000000000000000000000000002a00000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_39 => X"0000001500000000000000150000000000000000000000000000000000000000",
            INIT_3A => X"0000002f00000000000000200000000000000024000000000000001000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000002d00000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"00000017000000000000000c0000000000000000000000000000000000000000",
            INIT_3F => X"0000000700000000000000000000000000000019000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"00000000000000000000000c0000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"000000a900000000000000710000000000000000000000000000000000000000",
            INIT_47 => X"0000008c000000000000008d0000000000000094000000000000008c00000000",
            INIT_48 => X"0000004100000000000000460000000000000077000000000000007800000000",
            INIT_49 => X"0000005f00000000000000480000000000000045000000000000004800000000",
            INIT_4A => X"0000009300000000000000930000000000000098000000000000003b00000000",
            INIT_4B => X"0000009600000000000000a0000000000000009e000000000000009900000000",
            INIT_4C => X"0000004800000000000000370000000000000060000000000000008e00000000",
            INIT_4D => X"0000004d00000000000000570000000000000062000000000000004e00000000",
            INIT_4E => X"000000a200000000000000a20000000000000094000000000000008100000000",
            INIT_4F => X"0000009f000000000000009a00000000000000a700000000000000a500000000",
            INIT_50 => X"0000006300000000000000800000000000000065000000000000009200000000",
            INIT_51 => X"0000007000000000000000600000000000000057000000000000006100000000",
            INIT_52 => X"000000a700000000000000a9000000000000009a000000000000009c00000000",
            INIT_53 => X"000000980000000000000093000000000000009c00000000000000ac00000000",
            INIT_54 => X"0000004b000000000000005c0000000000000086000000000000009200000000",
            INIT_55 => X"000000970000000000000071000000000000005f000000000000005f00000000",
            INIT_56 => X"000000a500000000000000af00000000000000a500000000000000a400000000",
            INIT_57 => X"0000009000000000000000810000000000000097000000000000008b00000000",
            INIT_58 => X"000000580000000000000056000000000000004b000000000000008d00000000",
            INIT_59 => X"000000ac00000000000000900000000000000070000000000000005b00000000",
            INIT_5A => X"0000008a00000000000000a9000000000000009c00000000000000a900000000",
            INIT_5B => X"0000006c0000000000000082000000000000005a000000000000006c00000000",
            INIT_5C => X"0000005c000000000000004f000000000000004d000000000000001f00000000",
            INIT_5D => X"0000009100000000000000a00000000000000095000000000000009d00000000",
            INIT_5E => X"00000067000000000000006f00000000000000a8000000000000009d00000000",
            INIT_5F => X"0000001f000000000000004e0000000000000093000000000000009900000000",
            INIT_60 => X"0000005d00000000000000510000000000000054000000000000003d00000000",
            INIT_61 => X"000000b1000000000000008c000000000000009000000000000000a500000000",
            INIT_62 => X"00000091000000000000009c00000000000000af00000000000000a400000000",
            INIT_63 => X"0000003e0000000000000024000000000000005a000000000000008800000000",
            INIT_64 => X"000000a80000000000000073000000000000004a000000000000007300000000",
            INIT_65 => X"00000088000000000000008b000000000000007a000000000000009700000000",
            INIT_66 => X"000000500000000000000065000000000000006f000000000000008400000000",
            INIT_67 => X"00000086000000000000004c0000000000000002000000000000000000000000",
            INIT_68 => X"0000008c00000000000000a40000000000000068000000000000002a00000000",
            INIT_69 => X"0000005100000000000000950000000000000062000000000000003400000000",
            INIT_6A => X"0000002a000000000000001c000000000000006c000000000000009e00000000",
            INIT_6B => X"00000030000000000000009e0000000000000050000000000000003400000000",
            INIT_6C => X"0000000700000000000000700000000000000090000000000000007900000000",
            INIT_6D => X"000000620000000000000026000000000000001c000000000000003d00000000",
            INIT_6E => X"0000002500000000000000130000000000000018000000000000001400000000",
            INIT_6F => X"0000006c00000000000000380000000000000094000000000000005400000000",
            INIT_70 => X"0000005e0000000000000078000000000000006d000000000000008900000000",
            INIT_71 => X"00000004000000000000003b0000000000000078000000000000006000000000",
            INIT_72 => X"0000003900000000000000170000000000000000000000000000000300000000",
            INIT_73 => X"0000007d00000000000000890000000000000052000000000000006300000000",
            INIT_74 => X"0000006b0000000000000081000000000000007b000000000000007e00000000",
            INIT_75 => X"000000280000000000000038000000000000005b000000000000007100000000",
            INIT_76 => X"0000003200000000000000470000000000000021000000000000001600000000",
            INIT_77 => X"0000006e000000000000007f0000000000000071000000000000006300000000",
            INIT_78 => X"0000008800000000000000720000000000000049000000000000007300000000",
            INIT_79 => X"0000005b000000000000005d0000000000000061000000000000006800000000",
            INIT_7A => X"0000004500000000000000710000000000000064000000000000007200000000",
            INIT_7B => X"0000008a00000000000000770000000000000096000000000000006d00000000",
            INIT_7C => X"0000006d0000000000000080000000000000008b000000000000007e00000000",
            INIT_7D => X"00000084000000000000007e0000000000000064000000000000006d00000000",
            INIT_7E => X"0000004f000000000000006f000000000000006a000000000000007b00000000",
            INIT_7F => X"0000002100000000000000100000000000000020000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE39;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE40 : if BRAM_NAME = "samplegold_layersamples_instance40" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003a000000000000000f0000000000000027000000000000001800000000",
            INIT_01 => X"00000000000000000000000f0000000000000008000000000000000a00000000",
            INIT_02 => X"000000310000000000000020000000000000002d000000000000000000000000",
            INIT_03 => X"0000001900000000000000190000000000000019000000000000001d00000000",
            INIT_04 => X"00000013000000000000003d0000000000000019000000000000002700000000",
            INIT_05 => X"0000001f000000000000000a000000000000000b000000000000000000000000",
            INIT_06 => X"0000001700000000000000050000000000000041000000000000001000000000",
            INIT_07 => X"0000002900000000000000240000000000000018000000000000001900000000",
            INIT_08 => X"00000000000000000000003e0000000000000028000000000000000a00000000",
            INIT_09 => X"000000110000000000000013000000000000000b000000000000002400000000",
            INIT_0A => X"00000012000000000000001e000000000000000f000000000000003f00000000",
            INIT_0B => X"00000025000000000000002c0000000000000027000000000000002300000000",
            INIT_0C => X"0000003600000000000000240000000000000025000000000000001000000000",
            INIT_0D => X"00000027000000000000000b0000000000000000000000000000001400000000",
            INIT_0E => X"000000190000000000000019000000000000001b000000000000000800000000",
            INIT_0F => X"00000029000000000000000b000000000000001d000000000000002200000000",
            INIT_10 => X"00000000000000000000005d000000000000001a000000000000000000000000",
            INIT_11 => X"000000290000000000000000000000000000000e000000000000001000000000",
            INIT_12 => X"000000000000000000000028000000000000001d000000000000000000000000",
            INIT_13 => X"0000000000000000000000450000000000000026000000000000004400000000",
            INIT_14 => X"0000000a0000000000000000000000000000004b000000000000002700000000",
            INIT_15 => X"0000003000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000004f00000000000000140000000000000007000000000000003000000000",
            INIT_17 => X"0000005200000000000000020000000000000000000000000000003e00000000",
            INIT_18 => X"0000000600000000000000000000000000000000000000000000003500000000",
            INIT_19 => X"00000023000000000000003b0000000000000000000000000000002800000000",
            INIT_1A => X"000000190000000000000030000000000000003c000000000000000000000000",
            INIT_1B => X"0000003b00000000000000600000000000000037000000000000003100000000",
            INIT_1C => X"0000002a00000000000000300000000000000000000000000000000000000000",
            INIT_1D => X"0000000100000000000000430000000000000028000000000000000000000000",
            INIT_1E => X"0000002d00000000000000270000000000000054000000000000001100000000",
            INIT_1F => X"0000000000000000000000210000000000000077000000000000003e00000000",
            INIT_20 => X"0000000000000000000000390000000000000070000000000000000000000000",
            INIT_21 => X"0000000e0000000000000000000000000000009c000000000000002900000000",
            INIT_22 => X"0000002c00000000000000530000000000000000000000000000007100000000",
            INIT_23 => X"000000000000000000000000000000000000000d000000000000000800000000",
            INIT_24 => X"0000003400000000000000000000000000000039000000000000009100000000",
            INIT_25 => X"000000150000000000000000000000000000000000000000000000a300000000",
            INIT_26 => X"00000001000000000000001c0000000000000059000000000000000000000000",
            INIT_27 => X"0000008700000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"00000034000000000000001d000000000000000d000000000000003b00000000",
            INIT_29 => X"0000003700000000000000040000000000000010000000000000003f00000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_2B => X"0000001600000000000000210000000000000000000000000000000000000000",
            INIT_2C => X"0000004000000000000000130000000000000017000000000000002300000000",
            INIT_2D => X"00000029000000000000003a0000000000000006000000000000003300000000",
            INIT_2E => X"0000000000000000000000000000000000000008000000000000000d00000000",
            INIT_2F => X"0000000000000000000000240000000000000000000000000000000100000000",
            INIT_30 => X"0000000300000000000000440000000000000013000000000000004500000000",
            INIT_31 => X"0000002400000000000000180000000000000042000000000000000000000000",
            INIT_32 => X"0000000000000000000000180000000000000002000000000000001b00000000",
            INIT_33 => X"000000300000000000000005000000000000001b000000000000002d00000000",
            INIT_34 => X"0000001e000000000000001b0000000000000026000000000000001400000000",
            INIT_35 => X"0000000c000000000000001d0000000000000025000000000000002900000000",
            INIT_36 => X"00000003000000000000002c0000000000000024000000000000000f00000000",
            INIT_37 => X"0000004800000000000000510000000000000027000000000000008100000000",
            INIT_38 => X"0000002f00000000000000520000000000000048000000000000005700000000",
            INIT_39 => X"0000002e0000000000000027000000000000001f000000000000005a00000000",
            INIT_3A => X"0000006200000000000000490000000000000015000000000000001f00000000",
            INIT_3B => X"0000005400000000000000520000000000000052000000000000007600000000",
            INIT_3C => X"0000006400000000000000480000000000000058000000000000005500000000",
            INIT_3D => X"0000002a00000000000000280000000000000012000000000000002500000000",
            INIT_3E => X"000000530000000000000081000000000000002e000000000000004000000000",
            INIT_3F => X"0000006300000000000000590000000000000059000000000000005400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000600000000000000059000000000000003d000000000000006600000000",
            INIT_41 => X"00000034000000000000002a000000000000003c000000000000001b00000000",
            INIT_42 => X"0000005f000000000000004e0000000000000077000000000000003300000000",
            INIT_43 => X"0000006600000000000000650000000000000063000000000000005300000000",
            INIT_44 => X"0000004e000000000000005c0000000000000046000000000000005700000000",
            INIT_45 => X"00000030000000000000001c0000000000000036000000000000006100000000",
            INIT_46 => X"00000057000000000000005f000000000000004f000000000000005700000000",
            INIT_47 => X"000000550000000000000062000000000000005f000000000000006500000000",
            INIT_48 => X"0000008a000000000000004d0000000000000038000000000000006000000000",
            INIT_49 => X"0000000000000000000000330000000000000030000000000000001e00000000",
            INIT_4A => X"0000006900000000000000650000000000000050000000000000006600000000",
            INIT_4B => X"0000007a00000000000000590000000000000087000000000000003900000000",
            INIT_4C => X"0000000e000000000000006a000000000000005a000000000000002c00000000",
            INIT_4D => X"0000003e00000000000000000000000000000024000000000000002a00000000",
            INIT_4E => X"0000005a000000000000004b0000000000000079000000000000007900000000",
            INIT_4F => X"0000003f0000000000000030000000000000007b000000000000008f00000000",
            INIT_50 => X"00000020000000000000000d000000000000004d000000000000008000000000",
            INIT_51 => X"0000008400000000000000000000000000000046000000000000002700000000",
            INIT_52 => X"0000006f000000000000008f000000000000004a000000000000005e00000000",
            INIT_53 => X"0000009e000000000000007d0000000000000075000000000000005a00000000",
            INIT_54 => X"0000004b00000000000000220000000000000005000000000000004f00000000",
            INIT_55 => X"0000007200000000000000770000000000000003000000000000005500000000",
            INIT_56 => X"00000059000000000000009f0000000000000058000000000000005900000000",
            INIT_57 => X"000000320000000000000099000000000000006b000000000000006600000000",
            INIT_58 => X"00000065000000000000009d000000000000000d000000000000000000000000",
            INIT_59 => X"0000000000000000000000d30000000000000077000000000000000000000000",
            INIT_5A => X"00000072000000000000003400000000000000ac000000000000004500000000",
            INIT_5B => X"00000000000000000000001f0000000000000022000000000000003d00000000",
            INIT_5C => X"00000019000000000000006a00000000000000d0000000000000000000000000",
            INIT_5D => X"00000017000000000000000000000000000000d1000000000000007500000000",
            INIT_5E => X"0000002900000000000000810000000000000012000000000000004300000000",
            INIT_5F => X"000000000000000000000000000000000000001b000000000000001500000000",
            INIT_60 => X"00000054000000000000003b000000000000006300000000000000cf00000000",
            INIT_61 => X"000000160000000000000025000000000000004e000000000000007a00000000",
            INIT_62 => X"0000000800000000000000060000000000000022000000000000004700000000",
            INIT_63 => X"0000005e00000000000000020000000000000000000000000000000000000000",
            INIT_64 => X"0000004d00000000000000460000000000000053000000000000004500000000",
            INIT_65 => X"0000005900000000000000370000000000000053000000000000007400000000",
            INIT_66 => X"0000000000000000000000100000000000000018000000000000003800000000",
            INIT_67 => X"0000005600000000000000000000000000000019000000000000000000000000",
            INIT_68 => X"0000007800000000000000330000000000000075000000000000002a00000000",
            INIT_69 => X"0000003a0000000000000070000000000000002a000000000000003500000000",
            INIT_6A => X"00000033000000000000001d0000000000000034000000000000003e00000000",
            INIT_6B => X"00000036000000000000004e0000000000000047000000000000001900000000",
            INIT_6C => X"0000004d0000000000000051000000000000003f000000000000006200000000",
            INIT_6D => X"00000044000000000000004a0000000000000055000000000000004a00000000",
            INIT_6E => X"00000056000000000000004e000000000000003c000000000000003800000000",
            INIT_6F => X"0000001b0000000000000005000000000000001b000000000000002600000000",
            INIT_70 => X"0000001e00000000000000210000000000000022000000000000002400000000",
            INIT_71 => X"0000000800000000000000050000000000000003000000000000000f00000000",
            INIT_72 => X"0000000300000000000000000000000000000004000000000000000400000000",
            INIT_73 => X"0000002000000000000000250000000000000022000000000000001e00000000",
            INIT_74 => X"0000002400000000000000270000000000000028000000000000002300000000",
            INIT_75 => X"0000000800000000000000080000000000000001000000000000001000000000",
            INIT_76 => X"0000001200000000000000070000000000000007000000000000000600000000",
            INIT_77 => X"0000002700000000000000290000000000000025000000000000002000000000",
            INIT_78 => X"000000200000000000000030000000000000002b000000000000002b00000000",
            INIT_79 => X"0000000c00000000000000040000000000000000000000000000000000000000",
            INIT_7A => X"00000016000000000000001c0000000000000008000000000000001000000000",
            INIT_7B => X"0000003000000000000000250000000000000027000000000000002300000000",
            INIT_7C => X"00000023000000000000002a0000000000000029000000000000002c00000000",
            INIT_7D => X"0000000e000000000000000f0000000000000011000000000000001e00000000",
            INIT_7E => X"00000024000000000000001a0000000000000017000000000000000c00000000",
            INIT_7F => X"000000260000000000000022000000000000002e000000000000002400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE40;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE41 : if BRAM_NAME = "samplegold_layersamples_instance41" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000023000000000000002a000000000000001d000000000000001b00000000",
            INIT_01 => X"0000000c000000000000000b000000000000000e000000000000000f00000000",
            INIT_02 => X"0000002000000000000000220000000000000015000000000000002d00000000",
            INIT_03 => X"000000060000000000000000000000000000000d000000000000002f00000000",
            INIT_04 => X"0000000e00000000000000130000000000000013000000000000001f00000000",
            INIT_05 => X"00000000000000000000000b000000000000000c000000000000000a00000000",
            INIT_06 => X"0000001b00000000000000160000000000000010000000000000002200000000",
            INIT_07 => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_08 => X"0000000400000000000000000000000000000003000000000000000000000000",
            INIT_09 => X"0000000e00000000000000000000000000000008000000000000000800000000",
            INIT_0A => X"0000001000000000000000080000000000000011000000000000000f00000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_0C => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_0D => X"0000000b0000000000000004000000000000000c000000000000000000000000",
            INIT_0E => X"00000016000000000000001c0000000000000004000000000000000d00000000",
            INIT_0F => X"00000011000000000000000f000000000000000f000000000000001400000000",
            INIT_10 => X"0000000000000000000000000000000000000004000000000000000400000000",
            INIT_11 => X"0000000000000000000000000000000000000004000000000000001300000000",
            INIT_12 => X"00000005000000000000001c000000000000000d000000000000000d00000000",
            INIT_13 => X"0000000000000000000000040000000000000007000000000000000000000000",
            INIT_14 => X"0000000f00000000000000000000000000000000000000000000000200000000",
            INIT_15 => X"0000000000000000000000070000000000000000000000000000000a00000000",
            INIT_16 => X"0000002500000000000000160000000000000023000000000000000e00000000",
            INIT_17 => X"0000000000000000000000080000000000000000000000000000000400000000",
            INIT_18 => X"00000008000000000000001a0000000000000000000000000000000000000000",
            INIT_19 => X"000000000000000000000000000000000000000c000000000000000700000000",
            INIT_1A => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_1B => X"00000009000000000000000d0000000000000000000000000000000000000000",
            INIT_1C => X"00000007000000000000000f000000000000001c000000000000000600000000",
            INIT_1D => X"00000016000000000000000d0000000000000018000000000000001700000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_1F => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_20 => X"0000000f0000000000000011000000000000001d000000000000000f00000000",
            INIT_21 => X"00000013000000000000000b000000000000000d000000000000001200000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_23 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000c000000000000000d0000000000000018000000000000000700000000",
            INIT_25 => X"00000010000000000000001c0000000000000013000000000000000c00000000",
            INIT_26 => X"0000001000000000000000130000000000000014000000000000001600000000",
            INIT_27 => X"00000000000000000000000a000000000000000a000000000000001100000000",
            INIT_28 => X"00000034000000000000002c000000000000002a000000000000002e00000000",
            INIT_29 => X"00000029000000000000002c0000000000000029000000000000003200000000",
            INIT_2A => X"0000001d0000000000000016000000000000001f000000000000002300000000",
            INIT_2B => X"000000260000000000000027000000000000001d000000000000002500000000",
            INIT_2C => X"0000003300000000000000260000000000000028000000000000002700000000",
            INIT_2D => X"0000002600000000000000280000000000000029000000000000003100000000",
            INIT_2E => X"00000023000000000000002d0000000000000025000000000000002e00000000",
            INIT_2F => X"0000002b00000000000000240000000000000014000000000000002900000000",
            INIT_30 => X"00000038000000000000002f000000000000002e000000000000002800000000",
            INIT_31 => X"0000002600000000000000000000000000000000000000000000002100000000",
            INIT_32 => X"0000002300000000000000230000000000000033000000000000003800000000",
            INIT_33 => X"0000003000000000000000250000000000000029000000000000001f00000000",
            INIT_34 => X"00000038000000000000003a000000000000003f000000000000003a00000000",
            INIT_35 => X"00000032000000000000002f000000000000002d000000000000002f00000000",
            INIT_36 => X"00000017000000000000002e000000000000002c000000000000002600000000",
            INIT_37 => X"0000002e0000000000000026000000000000002a000000000000002300000000",
            INIT_38 => X"0000003d0000000000000035000000000000000a000000000000002300000000",
            INIT_39 => X"0000003100000000000000250000000000000039000000000000003100000000",
            INIT_3A => X"0000000c000000000000001e0000000000000013000000000000002c00000000",
            INIT_3B => X"0000000700000000000000000000000000000038000000000000002100000000",
            INIT_3C => X"00000036000000000000001c000000000000003a000000000000004100000000",
            INIT_3D => X"0000002b000000000000002b0000000000000023000000000000003f00000000",
            INIT_3E => X"0000001e000000000000001f0000000000000021000000000000000d00000000",
            INIT_3F => X"0000000000000000000000280000000000000015000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002600000000000000280000000000000000000000000000000000000000",
            INIT_41 => X"0000002e0000000000000030000000000000001c000000000000001900000000",
            INIT_42 => X"0000000000000000000000210000000000000022000000000000001000000000",
            INIT_43 => X"0000000c00000000000000060000000000000016000000000000000500000000",
            INIT_44 => X"00000017000000000000002a0000000000000013000000000000000400000000",
            INIT_45 => X"0000000b000000000000002a0000000000000029000000000000000000000000",
            INIT_46 => X"0000002700000000000000220000000000000034000000000000000d00000000",
            INIT_47 => X"0000006b000000000000004e000000000000005c000000000000004100000000",
            INIT_48 => X"00000002000000000000000f0000000000000034000000000000007400000000",
            INIT_49 => X"0000000b000000000000000d000000000000003e000000000000002800000000",
            INIT_4A => X"00000048000000000000002f0000000000000031000000000000004a00000000",
            INIT_4B => X"0000000d000000000000003b000000000000003b000000000000000000000000",
            INIT_4C => X"0000000f0000000000000000000000000000001a000000000000001200000000",
            INIT_4D => X"0000003e000000000000002f000000000000002e000000000000003900000000",
            INIT_4E => X"000000640000000000000058000000000000005d000000000000002000000000",
            INIT_4F => X"0000002300000000000000390000000000000039000000000000006500000000",
            INIT_50 => X"0000004400000000000000170000000000000018000000000000001900000000",
            INIT_51 => X"000000170000000000000000000000000000001e000000000000002d00000000",
            INIT_52 => X"0000002d000000000000003c000000000000000c000000000000000000000000",
            INIT_53 => X"00000020000000000000002a000000000000001b000000000000001d00000000",
            INIT_54 => X"000000330000000000000034000000000000001d000000000000004800000000",
            INIT_55 => X"00000039000000000000001b000000000000002c000000000000003100000000",
            INIT_56 => X"0000000000000000000000060000000000000018000000000000002100000000",
            INIT_57 => X"0000002800000000000000160000000000000000000000000000000000000000",
            INIT_58 => X"00000040000000000000003b0000000000000043000000000000003300000000",
            INIT_59 => X"0000002d000000000000001b0000000000000037000000000000003b00000000",
            INIT_5A => X"0000000700000000000000120000000000000017000000000000003900000000",
            INIT_5B => X"00000028000000000000000e0000000000000001000000000000000000000000",
            INIT_5C => X"0000002200000000000000330000000000000024000000000000002800000000",
            INIT_5D => X"000000430000000000000041000000000000002a000000000000001a00000000",
            INIT_5E => X"00000028000000000000002c0000000000000038000000000000003d00000000",
            INIT_5F => X"000000000000000000000018000000000000002d000000000000002a00000000",
            INIT_60 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_63 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000020000000000000005000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000200000000000000010000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_6E => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000003000000000000000300000000",
            INIT_71 => X"0000000b00000000000000080000000000000008000000000000000e00000000",
            INIT_72 => X"0000000000000000000000090000000000000000000000000000000700000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"00000005000000000000001c0000000000000025000000000000000000000000",
            INIT_75 => X"00000004000000000000000a0000000000000000000000000000000600000000",
            INIT_76 => X"00000000000000000000000f0000000000000003000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"00000011000000000000000b0000000000000000000000000000000000000000",
            INIT_7F => X"0000001d000000000000001f0000000000000011000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE41;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE42 : if BRAM_NAME = "samplegold_layersamples_instance42" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000000000001d000000000000002f00000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"00000027000000000000002c0000000000000006000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_04 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_05 => X"0000000400000000000000030000000000000000000000000000000000000000",
            INIT_06 => X"0000001b000000000000000b0000000000000000000000000000000000000000",
            INIT_07 => X"0000001100000000000000110000000000000026000000000000001b00000000",
            INIT_08 => X"00000000000000000000000a0000000000000000000000000000000700000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000d00000000000000010000000000000000000000000000000000000000",
            INIT_0C => X"0000000600000000000000000000000000000018000000000000000500000000",
            INIT_0D => X"0000001900000000000000090000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000f00000000000000060000000000000001000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000002f00000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000400000000000000010000000000000000000000000000000000000000",
            INIT_22 => X"0000002800000000000000000000000000000000000000000000002200000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000001000000000000000020000000000000004000000000000000000000000",
            INIT_25 => X"000000000000000000000006000000000000000a000000000000000f00000000",
            INIT_26 => X"000000000000000000000000000000000000000b000000000000000b00000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_28 => X"0000000b00000000000000090000000000000011000000000000000600000000",
            INIT_29 => X"000000030000000000000000000000000000002c000000000000003800000000",
            INIT_2A => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000052000000000000004800000000",
            INIT_2D => X"000000090000000000000000000000000000004b000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000340000000000000008000000000000000000000000",
            INIT_30 => X"0000007300000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000200000000000000000000000000000000000000000000007700000000",
            INIT_32 => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000110000000000000000000000000000000d00000000",
            INIT_34 => X"0000000000000000000000ab00000000000000b5000000000000006300000000",
            INIT_35 => X"0000007900000000000000020000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_37 => X"00000099000000000000003f0000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000b000000000000002b0000000000000075000000000000004800000000",
            INIT_3A => X"00000000000000000000000e000000000000000000000000000000cb00000000",
            INIT_3B => X"0000000000000000000000220000000000000072000000000000001d00000000",
            INIT_3C => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000480000000000000000000000000000000000000000",
            INIT_3E => X"0000005c00000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000006000000000000009800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000000000000000000000000000000000005e000000000000000100000000",
            INIT_41 => X"0000002d00000000000000000000000000000014000000000000000000000000",
            INIT_42 => X"00000082000000000000005b0000000000000025000000000000000000000000",
            INIT_43 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_44 => X"000000000000000000000000000000000000001a000000000000003b00000000",
            INIT_45 => X"0000000000000000000000310000000000000010000000000000000f00000000",
            INIT_46 => X"0000000000000000000000680000000000000053000000000000007c00000000",
            INIT_47 => X"0000000000000000000000000000000000000035000000000000000000000000",
            INIT_48 => X"00000010000000000000000c0000000000000000000000000000004200000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000004000000000",
            INIT_4C => X"0000000000000000000000090000000000000009000000000000000000000000",
            INIT_4D => X"00000013000000000000000b0000000000000014000000000000000f00000000",
            INIT_4E => X"0000002500000000000000000000000000000003000000000000000a00000000",
            INIT_4F => X"0000000700000000000000040000000000000000000000000000000000000000",
            INIT_50 => X"0000005e00000000000000530000000000000064000000000000001500000000",
            INIT_51 => X"00000035000000000000002e0000000000000041000000000000004e00000000",
            INIT_52 => X"0000000c000000000000002d000000000000001a000000000000001b00000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_54 => X"00000015000000000000002f0000000000000045000000000000004e00000000",
            INIT_55 => X"00000004000000000000000f0000000000000008000000000000001000000000",
            INIT_56 => X"0000000000000000000000240000000000000000000000000000000200000000",
            INIT_57 => X"0000002500000000000000000000000000000007000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000002000000000000001200000000",
            INIT_59 => X"0000000a00000000000000070000000000000004000000000000000100000000",
            INIT_5A => X"0000000a00000000000000240000000000000054000000000000001600000000",
            INIT_5B => X"0000000000000000000000000000000000000006000000000000002900000000",
            INIT_5C => X"0000000e00000000000000040000000000000000000000000000000000000000",
            INIT_5D => X"0000003700000000000000320000000000000030000000000000002300000000",
            INIT_5E => X"0000000e000000000000001b0000000000000001000000000000000900000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000005800000000000000300000000000000011000000000000000000000000",
            INIT_61 => X"0000004000000000000000a400000000000000ac000000000000006d00000000",
            INIT_62 => X"0000000000000000000000000000000000000022000000000000002800000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000010400000000000000fa0000000000000093000000000000002300000000",
            INIT_65 => X"0000002f00000000000001720000000000000115000000000000011300000000",
            INIT_66 => X"000000020000000000000000000000000000002b000000000000001d00000000",
            INIT_67 => X"0000005700000000000000130000000000000000000000000000000200000000",
            INIT_68 => X"00000016000000000000001a0000000000000087000000000000008600000000",
            INIT_69 => X"0000000000000000000000d700000000000001ef00000000000000ad00000000",
            INIT_6A => X"0000000600000000000000050000000000000000000000000000001e00000000",
            INIT_6B => X"00000058000000000000005d000000000000005c000000000000003a00000000",
            INIT_6C => X"000001af000000000000011e00000000000000a4000000000000006600000000",
            INIT_6D => X"000000010000000000000010000000000000010500000000000001f800000000",
            INIT_6E => X"00000036000000000000002f0000000000000001000000000000008f00000000",
            INIT_6F => X"000000a0000000000000002c000000000000003b000000000000006500000000",
            INIT_70 => X"000001c2000000000000020500000000000001fa00000000000001e400000000",
            INIT_71 => X"0000014b00000000000000b80000000000000078000000000000005b00000000",
            INIT_72 => X"00000040000000000000006b000000000000011c000000000000002400000000",
            INIT_73 => X"000001ce00000000000000da0000000000000000000000000000000000000000",
            INIT_74 => X"000001570000000000000188000000000000016600000000000001c300000000",
            INIT_75 => X"0000004800000000000001050000000000000154000000000000015200000000",
            INIT_76 => X"00000000000000000000001f000000000000009600000000000000fe00000000",
            INIT_77 => X"0000013d00000000000001b30000000000000109000000000000003800000000",
            INIT_78 => X"0000015a00000000000001440000000000000046000000000000003d00000000",
            INIT_79 => X"0000003d0000000000000018000000000000003500000000000000fe00000000",
            INIT_7A => X"000000930000000000000000000000000000000800000000000000c500000000",
            INIT_7B => X"0000002400000000000000be00000000000001bf000000000000015d00000000",
            INIT_7C => X"00000063000000000000011c0000000000000071000000000000000600000000",
            INIT_7D => X"000000d200000000000000550000000000000000000000000000000000000000",
            INIT_7E => X"00000193000000000000011c00000000000000aa000000000000003200000000",
            INIT_7F => X"00000049000000000000006c000000000000009d00000000000001aa00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE42;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE43 : if BRAM_NAME = "samplegold_layersamples_instance43" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000000000000000000b7000000000000000000000000",
            INIT_01 => X"00000017000000000000006a0000000000000035000000000000000000000000",
            INIT_02 => X"00000099000000000000009a0000000000000089000000000000005b00000000",
            INIT_03 => X"00000000000000000000004b0000000000000063000000000000002c00000000",
            INIT_04 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"00000000000000000000000d0000000000000029000000000000001900000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_07 => X"0000000000000000000000000000000000000011000000000000001900000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000001000000000000000300000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000001a00000000000000010000000000000000000000000000000000000000",
            INIT_1D => X"0000000a0000000000000056000000000000005b000000000000002900000000",
            INIT_1E => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000f00000000000000310000000000000031000000000000001200000000",
            INIT_21 => X"0000000000000000000000950000000000000035000000000000000600000000",
            INIT_22 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"00000000000000000000001e0000000000000072000000000000003000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_28 => X"000000880000000000000082000000000000007a000000000000002400000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000005700000000",
            INIT_2A => X"00000000000000000000002d0000000000000000000000000000003700000000",
            INIT_2B => X"0000004e00000000000000000000000000000000000000000000000100000000",
            INIT_2C => X"00000098000000000000007e0000000000000072000000000000008500000000",
            INIT_2D => X"0000003b000000000000003b0000000000000020000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000082000000000000003000000000",
            INIT_2F => X"0000006a000000000000004c0000000000000000000000000000000000000000",
            INIT_30 => X"000000c100000000000000340000000000000000000000000000004d00000000",
            INIT_31 => X"0000000d00000000000000000000000000000044000000000000005100000000",
            INIT_32 => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_33 => X"000000000000000000000062000000000000006d000000000000001e00000000",
            INIT_34 => X"0000004f00000000000000480000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000002600000000",
            INIT_37 => X"0000000000000000000000000000000000000062000000000000006100000000",
            INIT_38 => X"00000000000000000000005e0000000000000000000000000000000000000000",
            INIT_39 => X"0000002900000000000000070000000000000000000000000000000000000000",
            INIT_3A => X"000000820000000000000079000000000000004d000000000000000400000000",
            INIT_3B => X"0000000000000000000000190000000000000009000000000000008100000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"000000000000000000000000000000000000000d000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000700000000000000150000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"000000000000000000000000000000000000000a000000000000001a00000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"00000000000000000000000e0000000000000018000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000160000000000000013000000000000002000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000001000000000000000030000000000000000000000000000000000000000",
            INIT_59 => X"0000000c00000000000000350000000000000016000000000000002200000000",
            INIT_5A => X"00000005000000000000000e0000000000000016000000000000003300000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000002e00000000000000150000000000000012000000000000000d00000000",
            INIT_5D => X"0000001a00000000000000230000000000000004000000000000002200000000",
            INIT_5E => X"000000000000000000000017000000000000001d000000000000002c00000000",
            INIT_5F => X"0000001400000000000000240000000000000000000000000000000000000000",
            INIT_60 => X"0000001400000000000000020000000000000038000000000000001900000000",
            INIT_61 => X"0000001e000000000000003f0000000000000014000000000000002700000000",
            INIT_62 => X"0000000000000000000000000000000000000011000000000000002200000000",
            INIT_63 => X"0000001900000000000000240000000000000022000000000000002000000000",
            INIT_64 => X"00000013000000000000002e0000000000000019000000000000002b00000000",
            INIT_65 => X"00000020000000000000001b0000000000000036000000000000002f00000000",
            INIT_66 => X"0000003300000000000000030000000000000000000000000000001200000000",
            INIT_67 => X"0000002600000000000000250000000000000026000000000000001a00000000",
            INIT_68 => X"000000100000000000000040000000000000000a000000000000002400000000",
            INIT_69 => X"00000022000000000000001f0000000000000029000000000000002800000000",
            INIT_6A => X"00000023000000000000001a0000000000000028000000000000000000000000",
            INIT_6B => X"00000026000000000000002e0000000000000014000000000000002200000000",
            INIT_6C => X"000000180000000000000020000000000000001e000000000000002200000000",
            INIT_6D => X"000000070000000000000024000000000000001f000000000000002b00000000",
            INIT_6E => X"0000002a0000000000000037000000000000001c000000000000001e00000000",
            INIT_6F => X"0000002e000000000000002d0000000000000016000000000000002b00000000",
            INIT_70 => X"0000000c00000000000000190000000000000022000000000000002400000000",
            INIT_71 => X"0000001100000000000000080000000000000010000000000000003200000000",
            INIT_72 => X"0000001b00000000000000140000000000000028000000000000001100000000",
            INIT_73 => X"0000001700000000000000330000000000000021000000000000001d00000000",
            INIT_74 => X"00000025000000000000000c000000000000001e000000000000002600000000",
            INIT_75 => X"0000002900000000000000150000000000000009000000000000001400000000",
            INIT_76 => X"0000001e00000000000000210000000000000022000000000000001f00000000",
            INIT_77 => X"000000190000000000000012000000000000001a000000000000001d00000000",
            INIT_78 => X"0000001400000000000000140000000000000015000000000000002300000000",
            INIT_79 => X"000000fd000000000000010100000000000000f900000000000000fa00000000",
            INIT_7A => X"000000c800000000000000da00000000000000de00000000000000f000000000",
            INIT_7B => X"00000082000000000000008f00000000000000a400000000000000b800000000",
            INIT_7C => X"000000ed000000000000006e000000000000003f000000000000004200000000",
            INIT_7D => X"000000c700000000000000d400000000000000db00000000000000db00000000",
            INIT_7E => X"000000a000000000000000a900000000000000b500000000000000b700000000",
            INIT_7F => X"0000002100000000000000550000000000000087000000000000009200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE43;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE44 : if BRAM_NAME = "samplegold_layersamples_instance44" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ab00000000000000b3000000000000007d000000000000005000000000",
            INIT_01 => X"0000009c00000000000000a400000000000000a900000000000000ab00000000",
            INIT_02 => X"000000970000000000000099000000000000009b000000000000009f00000000",
            INIT_03 => X"00000073000000000000003a0000000000000023000000000000006700000000",
            INIT_04 => X"000000990000000000000096000000000000008e000000000000008200000000",
            INIT_05 => X"0000009e00000000000000a1000000000000009d000000000000009800000000",
            INIT_06 => X"0000002b000000000000008c0000000000000098000000000000009c00000000",
            INIT_07 => X"0000008500000000000000870000000000000066000000000000002000000000",
            INIT_08 => X"0000009b000000000000009c000000000000009b000000000000009200000000",
            INIT_09 => X"0000008c0000000000000091000000000000009e00000000000000a000000000",
            INIT_0A => X"000000320000000000000007000000000000004b000000000000007500000000",
            INIT_0B => X"0000009b0000000000000082000000000000007e000000000000006d00000000",
            INIT_0C => X"000000930000000000000099000000000000009b000000000000009c00000000",
            INIT_0D => X"0000005e000000000000005c0000000000000062000000000000007800000000",
            INIT_0E => X"0000003d0000000000000000000000000000000b000000000000003a00000000",
            INIT_0F => X"0000009c000000000000009d0000000000000074000000000000005500000000",
            INIT_10 => X"0000004b0000000000000075000000000000008e000000000000009700000000",
            INIT_11 => X"00000020000000000000000f0000000000000002000000000000001500000000",
            INIT_12 => X"0000003400000000000000070000000000000000000000000000003800000000",
            INIT_13 => X"000000860000000000000099000000000000009b000000000000005300000000",
            INIT_14 => X"00000013000000000000002d0000000000000033000000000000006000000000",
            INIT_15 => X"0000001b00000000000000250000000000000016000000000000000000000000",
            INIT_16 => X"00000023000000000000001a0000000000000000000000000000000100000000",
            INIT_17 => X"0000001c000000000000003c0000000000000088000000000000009900000000",
            INIT_18 => X"0000003e00000000000000240000000000000011000000000000000a00000000",
            INIT_19 => X"000000000000000000000001000000000000001a000000000000002900000000",
            INIT_1A => X"000000940000000000000037000000000000001b000000000000003200000000",
            INIT_1B => X"00000000000000000000000d0000000000000000000000000000006500000000",
            INIT_1C => X"0000000c00000000000000210000000000000024000000000000001c00000000",
            INIT_1D => X"0000001d00000000000000000000000000000033000000000000001e00000000",
            INIT_1E => X"0000005000000000000000900000000000000016000000000000001400000000",
            INIT_1F => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000010000000000000002100000000",
            INIT_21 => X"0000000800000000000000000000000000000031000000000000001000000000",
            INIT_22 => X"000000060000000000000002000000000000006c000000000000000100000000",
            INIT_23 => X"0000001d00000000000000170000000000000008000000000000000000000000",
            INIT_24 => X"0000000400000000000000010000000000000000000000000000000f00000000",
            INIT_25 => X"0000000a00000000000000000000000000000007000000000000003500000000",
            INIT_26 => X"00000000000000000000000d0000000000000016000000000000005200000000",
            INIT_27 => X"00000002000000000000001b0000000000000000000000000000000600000000",
            INIT_28 => X"0000000b00000000000000000000000000000015000000000000000000000000",
            INIT_29 => X"0000004800000000000000230000000000000000000000000000002900000000",
            INIT_2A => X"0000001c0000000000000000000000000000001a000000000000002800000000",
            INIT_2B => X"0000000000000000000000140000000000000017000000000000001b00000000",
            INIT_2C => X"0000001d00000000000000000000000000000000000000000000001600000000",
            INIT_2D => X"0000001800000000000000460000000000000019000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000002c00000000000000060000000000000002000000000000000000000000",
            INIT_30 => X"0000000f000000000000000e0000000000000000000000000000000700000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000190000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000029000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"00000000000000000000000c000000000000002a000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_47 => X"0000000000000000000000000000000000000003000000000000002100000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000001a0000000000000018000000000000000d000000000000000600000000",
            INIT_4A => X"0000001800000000000000000000000000000033000000000000002500000000",
            INIT_4B => X"0000000000000000000000000000000000000008000000000000001e00000000",
            INIT_4C => X"0000000f00000000000000070000000000000000000000000000000000000000",
            INIT_4D => X"0000002300000000000000140000000000000000000000000000000000000000",
            INIT_4E => X"0000000d00000000000000000000000000000000000000000000000200000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_50 => X"000000200000000000000024000000000000000d000000000000000b00000000",
            INIT_51 => X"0000000000000000000000000000000000000002000000000000002a00000000",
            INIT_52 => X"0000001600000000000000070000000000000001000000000000000000000000",
            INIT_53 => X"0000002000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000001a0000000000000029000000000000002a000000000000000400000000",
            INIT_55 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_56 => X"00000000000000000000000e0000000000000005000000000000000000000000",
            INIT_57 => X"0000000a000000000000001a0000000000000000000000000000001500000000",
            INIT_58 => X"0000000c000000000000000a0000000000000042000000000000001d00000000",
            INIT_59 => X"0000000000000000000000320000000000000044000000000000000000000000",
            INIT_5A => X"0000000100000000000000000000000000000000000000000000001100000000",
            INIT_5B => X"0000003700000000000000170000000000000006000000000000001a00000000",
            INIT_5C => X"0000001500000000000000000000000000000000000000000000002c00000000",
            INIT_5D => X"000000000000000000000008000000000000004b000000000000001400000000",
            INIT_5E => X"00000023000000000000000c0000000000000000000000000000000e00000000",
            INIT_5F => X"0000002f000000000000000f0000000000000020000000000000000000000000",
            INIT_60 => X"00000005000000000000001c0000000000000000000000000000000000000000",
            INIT_61 => X"000000270000000000000000000000000000003e000000000000002100000000",
            INIT_62 => X"0000000e0000000000000029000000000000000c000000000000000100000000",
            INIT_63 => X"00000025000000000000002b0000000000000033000000000000003c00000000",
            INIT_64 => X"0000000c0000000000000002000000000000002b000000000000000000000000",
            INIT_65 => X"0000000000000000000000220000000000000010000000000000003d00000000",
            INIT_66 => X"0000001b00000000000000160000000000000014000000000000000000000000",
            INIT_67 => X"0000001f000000000000001c000000000000001f000000000000001c00000000",
            INIT_68 => X"000000220000000000000009000000000000000d000000000000004000000000",
            INIT_69 => X"0000000000000000000000000000000000000025000000000000002300000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"00000054000000000000004f000000000000003d000000000000000e00000000",
            INIT_7F => X"0000000000000000000000000000000000000003000000000000000b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE44;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE45 : if BRAM_NAME = "samplegold_layersamples_instance45" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"00000040000000000000004f0000000000000019000000000000000000000000",
            INIT_02 => X"0000002600000000000000ae000000000000003a000000000000002b00000000",
            INIT_03 => X"0000000000000000000000000000000000000010000000000000000200000000",
            INIT_04 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000002500000000000000170000000000000019000000000000000b00000000",
            INIT_06 => X"00000003000000000000006e00000000000000a6000000000000006600000000",
            INIT_07 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_08 => X"00000029000000000000002f000000000000002d000000000000000000000000",
            INIT_09 => X"000000a700000000000000a0000000000000008d000000000000003300000000",
            INIT_0A => X"0000001200000000000000010000000000000018000000000000009b00000000",
            INIT_0B => X"0000001800000000000000000000000000000000000000000000005900000000",
            INIT_0C => X"0000004d000000000000001b000000000000000f000000000000003400000000",
            INIT_0D => X"0000008a000000000000009e00000000000000a100000000000000ae00000000",
            INIT_0E => X"0000006c00000000000000750000000000000054000000000000003700000000",
            INIT_0F => X"0000002e000000000000004d000000000000006b000000000000000000000000",
            INIT_10 => X"000000a10000000000000068000000000000001a000000000000000000000000",
            INIT_11 => X"0000009d000000000000005d000000000000004400000000000000a000000000",
            INIT_12 => X"00000000000000000000003a0000000000000081000000000000008d00000000",
            INIT_13 => X"0000000b000000000000001d0000000000000065000000000000001e00000000",
            INIT_14 => X"0000005d000000000000009b0000000000000084000000000000005400000000",
            INIT_15 => X"0000007b00000000000000500000000000000018000000000000002000000000",
            INIT_16 => X"0000002900000000000000000000000000000000000000000000004900000000",
            INIT_17 => X"0000005e000000000000003b000000000000001b000000000000006b00000000",
            INIT_18 => X"000000300000000000000047000000000000009d000000000000009500000000",
            INIT_19 => X"0000001c0000000000000074000000000000001a000000000000002300000000",
            INIT_1A => X"0000005a00000000000000150000000000000000000000000000000000000000",
            INIT_1B => X"0000008d0000000000000089000000000000006d000000000000003a00000000",
            INIT_1C => X"0000003600000000000000420000000000000043000000000000008d00000000",
            INIT_1D => X"0000000000000000000000040000000000000033000000000000000c00000000",
            INIT_1E => X"0000001800000000000000220000000000000000000000000000000000000000",
            INIT_1F => X"0000001200000000000000180000000000000018000000000000001500000000",
            INIT_20 => X"0000000000000000000000230000000000000031000000000000000900000000",
            INIT_21 => X"000000b300000000000000030000000000000000000000000000000000000000",
            INIT_22 => X"000000ac00000000000000b400000000000000ae00000000000000b200000000",
            INIT_23 => X"0000007b00000000000000910000000000000093000000000000009c00000000",
            INIT_24 => X"0000001e00000000000000560000000000000071000000000000006a00000000",
            INIT_25 => X"00000097000000000000009e0000000000000055000000000000002d00000000",
            INIT_26 => X"00000074000000000000007c0000000000000089000000000000008f00000000",
            INIT_27 => X"0000006a00000000000000680000000000000071000000000000007200000000",
            INIT_28 => X"00000032000000000000003a0000000000000042000000000000005700000000",
            INIT_29 => X"00000069000000000000006c000000000000006c000000000000005500000000",
            INIT_2A => X"0000006700000000000000670000000000000069000000000000006900000000",
            INIT_2B => X"000000250000000000000068000000000000006a000000000000006b00000000",
            INIT_2C => X"00000058000000000000004b000000000000003a000000000000001e00000000",
            INIT_2D => X"0000006300000000000000620000000000000062000000000000005f00000000",
            INIT_2E => X"0000006600000000000000620000000000000067000000000000006700000000",
            INIT_2F => X"0000002a0000000000000029000000000000005c000000000000006a00000000",
            INIT_30 => X"0000005c0000000000000061000000000000005c000000000000005700000000",
            INIT_31 => X"0000006200000000000000620000000000000062000000000000006200000000",
            INIT_32 => X"0000004a0000000000000052000000000000004d000000000000005900000000",
            INIT_33 => X"0000003400000000000000190000000000000021000000000000003300000000",
            INIT_34 => X"0000006100000000000000620000000000000057000000000000005500000000",
            INIT_35 => X"0000003b00000000000000570000000000000060000000000000006000000000",
            INIT_36 => X"0000000400000000000000000000000000000006000000000000001200000000",
            INIT_37 => X"0000002e0000000000000018000000000000002c000000000000000000000000",
            INIT_38 => X"0000005f00000000000000610000000000000062000000000000004c00000000",
            INIT_39 => X"000000100000000000000018000000000000002c000000000000005600000000",
            INIT_3A => X"0000000000000000000000110000000000000016000000000000001800000000",
            INIT_3B => X"0000002a0000000000000008000000000000001d000000000000001600000000",
            INIT_3C => X"000000260000000000000044000000000000005f000000000000006100000000",
            INIT_3D => X"000000160000000000000016000000000000001a000000000000001300000000",
            INIT_3E => X"0000000900000000000000000000000000000000000000000000001600000000",
            INIT_3F => X"0000005e0000000000000009000000000000001e000000000000002100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000d000000000000000c000000000000001f000000000000005000000000",
            INIT_41 => X"0000000000000000000000000000000000000019000000000000001000000000",
            INIT_42 => X"00000018000000000000003c0000000000000000000000000000000000000000",
            INIT_43 => X"0000000d000000000000005c0000000000000000000000000000000800000000",
            INIT_44 => X"00000010000000000000001c0000000000000004000000000000001300000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000100000000000000000000000000000040000000000000000000000000",
            INIT_48 => X"000000000000000000000008000000000000001e000000000000000500000000",
            INIT_49 => X"00000004000000000000001d0000000000000000000000000000000000000000",
            INIT_4A => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000001300000000000000000000000000000014000000000000003b00000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_4D => X"000000030000000000000013000000000000000c000000000000000c00000000",
            INIT_4E => X"000000310000000000000024000000000000000b000000000000000000000000",
            INIT_4F => X"0000000000000000000000130000000000000000000000000000000900000000",
            INIT_50 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"00000000000000000000000f000000000000000b000000000000000400000000",
            INIT_52 => X"0000001200000000000000310000000000000019000000000000001e00000000",
            INIT_53 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_54 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_55 => X"0000001e000000000000000d0000000000000018000000000000000e00000000",
            INIT_56 => X"0000000a00000000000000160000000000000028000000000000001500000000",
            INIT_57 => X"0000000d00000000000000060000000000000007000000000000000800000000",
            INIT_58 => X"0000000600000000000000090000000000000014000000000000001000000000",
            INIT_59 => X"0000001800000000000000180000000000000019000000000000001c00000000",
            INIT_5A => X"00000005000000000000000c0000000000000000000000000000000000000000",
            INIT_5B => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_5D => X"000000030000000000000000000000000000002d000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_60 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_61 => X"00000003000000000000000d0000000000000000000000000000003600000000",
            INIT_62 => X"0000000100000000000000050000000000000000000000000000000600000000",
            INIT_63 => X"0000000800000000000000000000000000000000000000000000000100000000",
            INIT_64 => X"0000001900000000000000000000000000000000000000000000000100000000",
            INIT_65 => X"000000040000000000000007000000000000000a000000000000000000000000",
            INIT_66 => X"0000000000000000000000020000000000000006000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000018000000000000003f00000000",
            INIT_69 => X"0000000000000000000000040000000000000005000000000000000900000000",
            INIT_6A => X"00000007000000000000000d0000000000000001000000000000000d00000000",
            INIT_6B => X"0000000f00000000000000000000000000000000000000000000000100000000",
            INIT_6C => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000001800000000000000000000000000000000000000000000000100000000",
            INIT_6E => X"0000002600000000000000000000000000000001000000000000001700000000",
            INIT_6F => X"0000004500000000000000000000000000000000000000000000000b00000000",
            INIT_70 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_71 => X"0000002f00000000000000150000000000000012000000000000000000000000",
            INIT_72 => X"000000a7000000000000001a0000000000000000000000000000000600000000",
            INIT_73 => X"0000002600000000000000000000000000000000000000000000005d00000000",
            INIT_74 => X"0000000d00000000000000000000000000000006000000000000000800000000",
            INIT_75 => X"00000000000000000000001b0000000000000000000000000000000000000000",
            INIT_76 => X"0000000200000000000000390000000000000000000000000000000000000000",
            INIT_77 => X"0000001d000000000000001b0000000000000000000000000000000000000000",
            INIT_78 => X"0000002200000000000000000000000000000014000000000000000100000000",
            INIT_79 => X"0000006600000000000000780000000000000036000000000000000000000000",
            INIT_7A => X"000000000000000000000000000000000000000e000000000000001600000000",
            INIT_7B => X"0000001f00000000000000170000000000000014000000000000001000000000",
            INIT_7C => X"0000000000000000000000260000000000000000000000000000003f00000000",
            INIT_7D => X"0000000f000000000000003100000000000000c8000000000000003e00000000",
            INIT_7E => X"000000000000000000000000000000000000004f000000000000000000000000",
            INIT_7F => X"0000004700000000000000600000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE45;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE46 : if BRAM_NAME = "samplegold_layersamples_instance46" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003b00000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"000000000000000000000000000000000000001700000000000000a900000000",
            INIT_02 => X"00000000000000000000000000000000000000dd000000000000005900000000",
            INIT_03 => X"00000000000000000000000e000000000000002a000000000000000000000000",
            INIT_04 => X"0000009f00000000000000540000000000000019000000000000000000000000",
            INIT_05 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_06 => X"000000000000000000000000000000000000002c00000000000000a400000000",
            INIT_07 => X"000000000000000000000022000000000000001b000000000000001e00000000",
            INIT_08 => X"0000000500000000000000540000000000000000000000000000004200000000",
            INIT_09 => X"000000110000000000000000000000000000003a000000000000000000000000",
            INIT_0A => X"0000000f00000000000000220000000000000000000000000000007400000000",
            INIT_0B => X"00000068000000000000000c000000000000001f000000000000001f00000000",
            INIT_0C => X"0000000000000000000000570000000000000064000000000000006400000000",
            INIT_0D => X"0000003100000000000000000000000000000000000000000000005c00000000",
            INIT_0E => X"0000000000000000000000050000000000000013000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000004900000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000500000000000000010000000000000000000000000000000000000000",
            INIT_12 => X"0000000100000000000000000000000000000000000000000000001300000000",
            INIT_13 => X"0000001600000000000000170000000000000017000000000000001200000000",
            INIT_14 => X"0000000e0000000000000031000000000000001a000000000000001300000000",
            INIT_15 => X"000000000000000000000025000000000000002a000000000000000400000000",
            INIT_16 => X"00000018000000000000000e0000000000000000000000000000001100000000",
            INIT_17 => X"0000000c000000000000000e0000000000000014000000000000001900000000",
            INIT_18 => X"0000000300000000000000000000000000000000000000000000000600000000",
            INIT_19 => X"0000003100000000000000000000000000000000000000000000000400000000",
            INIT_1A => X"000000090000000000000010000000000000001a000000000000003200000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"000000000000000000000015000000000000000b000000000000000000000000",
            INIT_1D => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000014000000000000003000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"000000000000000000000000000000000000007f000000000000005900000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000004b00000000000000700000000000000066000000000000005d00000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_2C => X"000000000000000000000000000000000000000f000000000000003800000000",
            INIT_2D => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_30 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000001400000000000000370000000000000024000000000000003c00000000",
            INIT_32 => X"0000000000000000000000100000000000000008000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"00000004000000000000001f0000000000000023000000000000001300000000",
            INIT_36 => X"00000000000000000000008a0000000000000055000000000000000000000000",
            INIT_37 => X"0000001f00000000000000120000000000000000000000000000000000000000",
            INIT_38 => X"000000140000000000000000000000000000000e00000000000000a200000000",
            INIT_39 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000002200000000000000a20000000000000061000000000000007400000000",
            INIT_3B => X"0000000a00000000000000290000000000000071000000000000003400000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"00000012000000000000001f000000000000004e000000000000000000000000",
            INIT_3F => X"00000000000000000000000d0000000000000020000000000000000300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"00000012000000000000002f0000000000000059000000000000000600000000",
            INIT_43 => X"0000005a00000000000000470000000000000019000000000000000000000000",
            INIT_44 => X"000000ec00000000000000e800000000000000d4000000000000009000000000",
            INIT_45 => X"00000005000000000000001d000000000000001c000000000000008c00000000",
            INIT_46 => X"0000000000000000000000080000000000000023000000000000004700000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"000000000000000000000018000000000000002f000000000000002f00000000",
            INIT_4A => X"000000ea00000000000000f90000000000000000000000000000000000000000",
            INIT_4B => X"000000c700000000000000dd00000000000000f000000000000000f800000000",
            INIT_4C => X"00000069000000000000009f00000000000000ac00000000000000c700000000",
            INIT_4D => X"0000002900000000000000210000000000000067000000000000006d00000000",
            INIT_4E => X"000000c700000000000000d200000000000000dd000000000000005a00000000",
            INIT_4F => X"00000099000000000000009500000000000000a400000000000000b300000000",
            INIT_50 => X"0000007800000000000000760000000000000082000000000000008900000000",
            INIT_51 => X"0000006500000000000000530000000000000000000000000000004800000000",
            INIT_52 => X"0000008100000000000000860000000000000081000000000000009500000000",
            INIT_53 => X"000000810000000000000083000000000000007e000000000000008100000000",
            INIT_54 => X"0000001900000000000000600000000000000085000000000000008100000000",
            INIT_55 => X"0000006c000000000000006a0000000000000078000000000000003d00000000",
            INIT_56 => X"00000084000000000000007a000000000000007a000000000000007700000000",
            INIT_57 => X"000000930000000000000094000000000000008b000000000000008500000000",
            INIT_58 => X"0000006100000000000000150000000000000000000000000000008a00000000",
            INIT_59 => X"0000007b00000000000000750000000000000062000000000000006900000000",
            INIT_5A => X"000000900000000000000085000000000000007a000000000000007b00000000",
            INIT_5B => X"00000086000000000000009c000000000000008b000000000000008a00000000",
            INIT_5C => X"0000006600000000000000690000000000000050000000000000001a00000000",
            INIT_5D => X"0000007b000000000000007b000000000000007a000000000000006500000000",
            INIT_5E => X"000000b2000000000000008c000000000000007c000000000000007700000000",
            INIT_5F => X"000000710000000000000036000000000000008600000000000000a800000000",
            INIT_60 => X"0000005a000000000000005a0000000000000026000000000000002900000000",
            INIT_61 => X"000000720000000000000074000000000000007b000000000000007d00000000",
            INIT_62 => X"000000000000000000000000000000000000003d000000000000007d00000000",
            INIT_63 => X"0000000e000000000000009c000000000000003d000000000000000000000000",
            INIT_64 => X"0000007c000000000000003f0000000000000015000000000000001800000000",
            INIT_65 => X"0000002800000000000000760000000000000075000000000000007900000000",
            INIT_66 => X"000000a500000000000000400000000000000013000000000000003b00000000",
            INIT_67 => X"00000000000000000000000c000000000000008600000000000000e600000000",
            INIT_68 => X"0000007300000000000000780000000000000063000000000000001100000000",
            INIT_69 => X"0000000700000000000000000000000000000014000000000000003800000000",
            INIT_6A => X"00000073000000000000009000000000000000c3000000000000004400000000",
            INIT_6B => X"0000007c000000000000003d0000000000000000000000000000005300000000",
            INIT_6C => X"0000000e00000000000000c20000000000000079000000000000008300000000",
            INIT_6D => X"00000060000000000000000c0000000000000000000000000000001100000000",
            INIT_6E => X"0000003e000000000000004b0000000000000063000000000000007100000000",
            INIT_6F => X"0000003f000000000000005f000000000000008f000000000000006700000000",
            INIT_70 => X"000000010000000000000000000000000000002e000000000000008c00000000",
            INIT_71 => X"000000620000000000000081000000000000001e000000000000000000000000",
            INIT_72 => X"0000002c00000000000000010000000000000000000000000000002700000000",
            INIT_73 => X"000000480000000000000000000000000000001f000000000000002f00000000",
            INIT_74 => X"0000000a00000000000000000000000000000016000000000000000600000000",
            INIT_75 => X"00000000000000000000006f0000000000000072000000000000003b00000000",
            INIT_76 => X"00000021000000000000003a0000000000000000000000000000000700000000",
            INIT_77 => X"0000001200000000000000320000000000000000000000000000000000000000",
            INIT_78 => X"0000005f000000000000004b0000000000000000000000000000002000000000",
            INIT_79 => X"0000002800000000000000000000000000000057000000000000008c00000000",
            INIT_7A => X"00000000000000000000001b0000000000000011000000000000001500000000",
            INIT_7B => X"0000000400000000000000150000000000000033000000000000000e00000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"00000000000000000000001b0000000000000000000000000000000000000000",
            INIT_7E => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000c0000000000000000000000000000000a000000000000003a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE46;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE47 : if BRAM_NAME = "samplegold_layersamples_instance47" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000030000000000000004000000000000000200000000",
            INIT_01 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_02 => X"0000001d00000000000000080000000000000000000000000000000000000000",
            INIT_03 => X"00000027000000000000001f0000000000000016000000000000002700000000",
            INIT_04 => X"0000000f00000000000000240000000000000012000000000000001e00000000",
            INIT_05 => X"00000018000000000000000d000000000000001f000000000000001f00000000",
            INIT_06 => X"0000001b00000000000000130000000000000014000000000000000000000000",
            INIT_07 => X"000000170000000000000017000000000000001b000000000000002200000000",
            INIT_08 => X"00000016000000000000000f0000000000000016000000000000000e00000000",
            INIT_09 => X"00000000000000000000002c0000000000000019000000000000000000000000",
            INIT_0A => X"0000001300000000000000240000000000000019000000000000000f00000000",
            INIT_0B => X"000000100000000000000011000000000000000f000000000000001700000000",
            INIT_0C => X"00000000000000000000000a0000000000000010000000000000000f00000000",
            INIT_0D => X"0000001e0000000000000000000000000000000b000000000000003600000000",
            INIT_0E => X"00000013000000000000000f000000000000000c000000000000000b00000000",
            INIT_0F => X"0000000900000000000000080000000000000011000000000000000c00000000",
            INIT_10 => X"00000000000000000000004c0000000000000009000000000000000b00000000",
            INIT_11 => X"0000000a00000000000000190000000000000015000000000000001200000000",
            INIT_12 => X"0000000900000000000000150000000000000011000000000000000f00000000",
            INIT_13 => X"0000000000000000000000080000000000000004000000000000000500000000",
            INIT_14 => X"0000000000000000000000000000000000000027000000000000000100000000",
            INIT_15 => X"00000012000000000000000f000000000000000b000000000000000e00000000",
            INIT_16 => X"0000000000000000000000000000000000000013000000000000001300000000",
            INIT_17 => X"00000063000000000000002c0000000000000015000000000000000000000000",
            INIT_18 => X"000000150000000000000000000000000000008d000000000000001900000000",
            INIT_19 => X"0000001b0000000000000015000000000000000f000000000000000900000000",
            INIT_1A => X"0000003a000000000000001b0000000000000000000000000000000400000000",
            INIT_1B => X"000000000000000000000000000000000000000f000000000000003b00000000",
            INIT_1C => X"000000010000000000000000000000000000000e00000000000000e600000000",
            INIT_1D => X"0000000000000000000000000000000000000019000000000000001200000000",
            INIT_1E => X"00000000000000000000002a0000000000000000000000000000001700000000",
            INIT_1F => X"000000da00000000000000300000000000000000000000000000000000000000",
            INIT_20 => X"0000001600000000000000000000000000000000000000000000006b00000000",
            INIT_21 => X"0000004500000000000000000000000000000005000000000000000000000000",
            INIT_22 => X"0000003c00000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000c0000000000000007d000000000000004900000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000460000000000000000000000000000009f00000000",
            INIT_26 => X"0000006d00000000000000310000000000000008000000000000000000000000",
            INIT_27 => X"0000002800000000000000000000000000000066000000000000003f00000000",
            INIT_28 => X"0000008a00000000000000270000000000000000000000000000004800000000",
            INIT_29 => X"000000000000000000000000000000000000001c000000000000001b00000000",
            INIT_2A => X"0000000000000000000000870000000000000080000000000000002200000000",
            INIT_2B => X"0000009900000000000000530000000000000069000000000000000000000000",
            INIT_2C => X"0000004e00000000000000030000000000000008000000000000000000000000",
            INIT_2D => X"0000003400000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"00000000000000000000000e000000000000000000000000000000ed00000000",
            INIT_2F => X"00000000000000000000000c000000000000009a000000000000001100000000",
            INIT_30 => X"0000000000000000000000430000000000000000000000000000000000000000",
            INIT_31 => X"000000d700000000000000310000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000028000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000008f00000000",
            INIT_34 => X"0000002600000000000000000000000000000038000000000000001600000000",
            INIT_35 => X"0000000000000000000000900000000000000043000000000000003400000000",
            INIT_36 => X"000000170000000000000000000000000000002c000000000000003700000000",
            INIT_37 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000002a00000000",
            INIT_3B => X"00000051000000000000004e000000000000004f000000000000004100000000",
            INIT_3C => X"0000004a00000000000000400000000000000049000000000000005700000000",
            INIT_3D => X"000000270000000000000039000000000000003c000000000000002d00000000",
            INIT_3E => X"0000004a00000000000000240000000000000011000000000000002800000000",
            INIT_3F => X"0000003b000000000000003f000000000000004d000000000000004f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002a0000000000000033000000000000002e000000000000003500000000",
            INIT_41 => X"0000002e00000000000000300000000000000012000000000000002b00000000",
            INIT_42 => X"0000004400000000000000390000000000000024000000000000000000000000",
            INIT_43 => X"0000002600000000000000250000000000000030000000000000003700000000",
            INIT_44 => X"0000001f00000000000000250000000000000027000000000000002600000000",
            INIT_45 => X"0000000a0000000000000020000000000000004f000000000000000800000000",
            INIT_46 => X"00000020000000000000001e0000000000000022000000000000003100000000",
            INIT_47 => X"0000002900000000000000260000000000000020000000000000002400000000",
            INIT_48 => X"0000004e0000000000000020000000000000002b000000000000002d00000000",
            INIT_49 => X"0000002e0000000000000029000000000000002a000000000000000000000000",
            INIT_4A => X"000000260000000000000021000000000000001f000000000000001b00000000",
            INIT_4B => X"0000003500000000000000290000000000000024000000000000001f00000000",
            INIT_4C => X"0000000700000000000000510000000000000054000000000000002e00000000",
            INIT_4D => X"0000001e000000000000001f000000000000002c000000000000002f00000000",
            INIT_4E => X"0000001300000000000000260000000000000025000000000000002200000000",
            INIT_4F => X"0000004e0000000000000045000000000000001b000000000000000700000000",
            INIT_50 => X"0000000000000000000000a8000000000000006b000000000000008600000000",
            INIT_51 => X"0000002600000000000000200000000000000021000000000000004100000000",
            INIT_52 => X"0000002700000000000000030000000000000017000000000000002d00000000",
            INIT_53 => X"000000000000000000000033000000000000005b000000000000006200000000",
            INIT_54 => X"0000000f00000000000000140000000000000144000000000000002200000000",
            INIT_55 => X"0000000a000000000000002a0000000000000023000000000000002100000000",
            INIT_56 => X"000000440000000000000016000000000000003c000000000000002100000000",
            INIT_57 => X"0000008a00000000000000000000000000000000000000000000001200000000",
            INIT_58 => X"000000000000000000000000000000000000007d000000000000012100000000",
            INIT_59 => X"00000022000000000000001a000000000000000f000000000000002600000000",
            INIT_5A => X"0000001100000000000000000000000000000000000000000000005b00000000",
            INIT_5B => X"000000fd00000000000000e400000000000000ae000000000000009100000000",
            INIT_5C => X"00000009000000000000002f0000000000000000000000000000000200000000",
            INIT_5D => X"00000053000000000000000200000000000000be000000000000000000000000",
            INIT_5E => X"0000008c00000000000000600000000000000000000000000000000000000000",
            INIT_5F => X"0000003b00000000000000b7000000000000007f00000000000000ae00000000",
            INIT_60 => X"0000003400000000000000000000000000000089000000000000006c00000000",
            INIT_61 => X"000000000000000000000025000000000000003200000000000000cb00000000",
            INIT_62 => X"000000a300000000000000d50000000000000076000000000000000000000000",
            INIT_63 => X"0000009400000000000000ac0000000000000000000000000000000000000000",
            INIT_64 => X"000000400000000000000019000000000000000000000000000000ae00000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000006000000000",
            INIT_66 => X"0000002500000000000000100000000000000132000000000000008600000000",
            INIT_67 => X"0000002000000000000000c20000000000000053000000000000000000000000",
            INIT_68 => X"0000006000000000000000220000000000000007000000000000000000000000",
            INIT_69 => X"0000008b00000000000000090000000000000024000000000000000000000000",
            INIT_6A => X"00000000000000000000004b0000000000000000000000000000011f00000000",
            INIT_6B => X"00000000000000000000000000000000000000a5000000000000000000000000",
            INIT_6C => X"00000000000000000000003e0000000000000027000000000000000300000000",
            INIT_6D => X"000000b50000000000000060000000000000004f000000000000003c00000000",
            INIT_6E => X"00000000000000000000003b0000000000000058000000000000000000000000",
            INIT_6F => X"0000001700000000000000110000000000000000000000000000002600000000",
            INIT_70 => X"0000000000000000000000000000000000000019000000000000001100000000",
            INIT_71 => X"0000000000000000000000070000000000000007000000000000000500000000",
            INIT_72 => X"0000000000000000000000000000000000000033000000000000003800000000",
            INIT_73 => X"0000008c00000000000000770000000000000064000000000000000000000000",
            INIT_74 => X"0000007b000000000000007e000000000000008a000000000000009100000000",
            INIT_75 => X"0000003b00000000000000400000000000000059000000000000006e00000000",
            INIT_76 => X"0000002700000000000000240000000000000002000000000000002a00000000",
            INIT_77 => X"00000076000000000000007a0000000000000079000000000000008d00000000",
            INIT_78 => X"00000054000000000000005d000000000000005f000000000000006c00000000",
            INIT_79 => X"000000100000000000000038000000000000003f000000000000004800000000",
            INIT_7A => X"0000005c000000000000002d000000000000000f000000000000000000000000",
            INIT_7B => X"0000004b0000000000000054000000000000005f000000000000005e00000000",
            INIT_7C => X"0000003b00000000000000400000000000000045000000000000004300000000",
            INIT_7D => X"0000000600000000000000120000000000000000000000000000003800000000",
            INIT_7E => X"0000003e00000000000000400000000000000025000000000000001700000000",
            INIT_7F => X"0000003e0000000000000040000000000000003e000000000000003d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE47;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE48 : if BRAM_NAME = "samplegold_layersamples_instance48" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000270000000000000038000000000000003c000000000000004100000000",
            INIT_01 => X"0000002e000000000000001c0000000000000004000000000000000000000000",
            INIT_02 => X"0000003e000000000000003d0000000000000037000000000000003600000000",
            INIT_03 => X"0000003300000000000000390000000000000040000000000000003d00000000",
            INIT_04 => X"0000000000000000000000080000000000000030000000000000003a00000000",
            INIT_05 => X"0000003100000000000000370000000000000035000000000000000300000000",
            INIT_06 => X"0000003d000000000000003d000000000000003d000000000000003900000000",
            INIT_07 => X"000000000000000000000000000000000000001d000000000000003500000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000003d000000000000002c0000000000000028000000000000000d00000000",
            INIT_0A => X"0000000c00000000000000360000000000000038000000000000003c00000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000003b000000000000003d000000000000002c000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000009000000000000002a00000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"00000000000000000000002b000000000000003a000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000003000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"00000099000000000000007f0000000000000000000000000000000000000000",
            INIT_2C => X"0000009e00000000000000a600000000000000aa00000000000000a100000000",
            INIT_2D => X"00000088000000000000008a0000000000000090000000000000009700000000",
            INIT_2E => X"00000039000000000000004b0000000000000052000000000000006a00000000",
            INIT_2F => X"0000009f0000000000000089000000000000009d000000000000004e00000000",
            INIT_30 => X"00000085000000000000008c000000000000009800000000000000a200000000",
            INIT_31 => X"0000004b00000000000000660000000000000073000000000000007d00000000",
            INIT_32 => X"0000005900000000000000250000000000000022000000000000004000000000",
            INIT_33 => X"00000088000000000000008e000000000000009c000000000000009300000000",
            INIT_34 => X"0000006800000000000000720000000000000073000000000000007b00000000",
            INIT_35 => X"00000026000000000000002b0000000000000056000000000000006200000000",
            INIT_36 => X"0000006e0000000000000059000000000000002d000000000000001400000000",
            INIT_37 => X"0000006c000000000000006f0000000000000070000000000000007000000000",
            INIT_38 => X"0000004c00000000000000540000000000000061000000000000006d00000000",
            INIT_39 => X"000000470000000000000027000000000000004a000000000000004700000000",
            INIT_3A => X"0000007300000000000000690000000000000064000000000000006a00000000",
            INIT_3B => X"0000005b000000000000006d0000000000000075000000000000007700000000",
            INIT_3C => X"00000000000000000000000a0000000000000048000000000000005300000000",
            INIT_3D => X"0000005900000000000000490000000000000005000000000000000000000000",
            INIT_3E => X"0000007300000000000000740000000000000071000000000000005f00000000",
            INIT_3F => X"000000000000000000000008000000000000005d000000000000007200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000340000000000000035000000000000000000000000",
            INIT_41 => X"0000005900000000000000390000000000000026000000000000001700000000",
            INIT_42 => X"0000005b00000000000000740000000000000075000000000000007300000000",
            INIT_43 => X"0000006600000000000000540000000000000058000000000000002c00000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000004100000000",
            INIT_45 => X"0000007500000000000000470000000000000031000000000000000c00000000",
            INIT_46 => X"00000022000000000000001b0000000000000038000000000000007200000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_48 => X"0000001d00000000000000380000000000000000000000000000000000000000",
            INIT_49 => X"0000004900000000000000770000000000000000000000000000000100000000",
            INIT_4A => X"0000001a00000000000000280000000000000014000000000000003800000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000040000000000000000800000000",
            INIT_4D => X"000000090000000000000000000000000000004e000000000000000000000000",
            INIT_4E => X"00000000000000000000000b000000000000002a000000000000000400000000",
            INIT_4F => X"0000001c000000000000003b0000000000000000000000000000000000000000",
            INIT_50 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000130000000000000011000000000000005c000000000000003d00000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_53 => X"0000000f000000000000004b0000000000000060000000000000003100000000",
            INIT_54 => X"0000005000000000000000730000000000000028000000000000000e00000000",
            INIT_55 => X"0000000000000000000000160000000000000000000000000000000800000000",
            INIT_56 => X"0000002d00000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000190000000000000001000000000000000000000000",
            INIT_58 => X"0000000300000000000000390000000000000012000000000000003a00000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_5B => X"0000004300000000000000170000000000000017000000000000000000000000",
            INIT_5C => X"0000002c0000000000000019000000000000002f000000000000002200000000",
            INIT_5D => X"0000008a000000000000007f0000000000000054000000000000003a00000000",
            INIT_5E => X"0000001b00000000000000060000000000000062000000000000009100000000",
            INIT_5F => X"0000001100000000000000200000000000000035000000000000001d00000000",
            INIT_60 => X"0000000000000000000000000000000000000013000000000000002500000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"00000022000000000000002c0000000000000016000000000000000400000000",
            INIT_63 => X"0000000000000000000000000000000000000006000000000000000600000000",
            INIT_64 => X"0000001b00000000000000190000000000000016000000000000000800000000",
            INIT_65 => X"000000180000000000000018000000000000001d000000000000001d00000000",
            INIT_66 => X"0000002100000000000000030000000000000001000000000000000500000000",
            INIT_67 => X"00000019000000000000001c0000000000000000000000000000001a00000000",
            INIT_68 => X"0000001e00000000000000230000000000000024000000000000002000000000",
            INIT_69 => X"0000000700000000000000120000000000000016000000000000001b00000000",
            INIT_6A => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_6B => X"0000002200000000000000270000000000000033000000000000000000000000",
            INIT_6C => X"0000000a000000000000000c0000000000000012000000000000001e00000000",
            INIT_6D => X"0000001e00000000000000000000000000000002000000000000000400000000",
            INIT_6E => X"0000000400000000000000000000000000000000000000000000001d00000000",
            INIT_6F => X"0000000700000000000000090000000000000009000000000000000c00000000",
            INIT_70 => X"0000000000000000000000030000000000000006000000000000000700000000",
            INIT_71 => X"0000000000000000000000010000000000000005000000000000000000000000",
            INIT_72 => X"0000000800000000000000050000000000000000000000000000000000000000",
            INIT_73 => X"0000000c000000000000000b000000000000000c000000000000000a00000000",
            INIT_74 => X"0000000000000000000000000000000000000015000000000000001500000000",
            INIT_75 => X"0000001b00000000000000050000000000000000000000000000000000000000",
            INIT_76 => X"0000000b0000000000000007000000000000000a000000000000000f00000000",
            INIT_77 => X"000000000000000000000005000000000000000c000000000000000c00000000",
            INIT_78 => X"000000520000000000000077000000000000005a000000000000001500000000",
            INIT_79 => X"0000001a000000000000001c0000000000000000000000000000000000000000",
            INIT_7A => X"0000000e000000000000000a000000000000000a000000000000000b00000000",
            INIT_7B => X"0000000600000000000000270000000000000022000000000000000600000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_7D => X"00000023000000000000001c0000000000000000000000000000000000000000",
            INIT_7E => X"000000160000000000000006000000000000000b000000000000000c00000000",
            INIT_7F => X"000000000000000000000000000000000000000b000000000000000500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE48;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE49 : if BRAM_NAME = "samplegold_layersamples_instance49" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000f00000000000000000000000000000000000000000000000600000000",
            INIT_02 => X"00000009000000000000000c0000000000000004000000000000000000000000",
            INIT_03 => X"0000001500000000000000040000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000004000000000000000000000000000000000000000000000000e00000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_09 => X"00000007000000000000003f0000000000000020000000000000001700000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"000000050000000000000000000000000000001c000000000000000000000000",
            INIT_0C => X"00000013000000000000001d0000000000000011000000000000001f00000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000001500000000000000040000000000000000000000000000000000000000",
            INIT_14 => X"0000000400000000000000000000000000000005000000000000000700000000",
            INIT_15 => X"0000004200000000000000360000000000000029000000000000001d00000000",
            INIT_16 => X"000000030000000000000025000000000000004d000000000000004c00000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000002300000000000000040000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000001200000000000000100000000000000004000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000003000000000000001200000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"00000010000000000000000d0000000000000006000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_27 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_28 => X"0000001300000000000000110000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000034000000000000003200000000",
            INIT_2C => X"000000000000000000000010000000000000002a000000000000000600000000",
            INIT_2D => X"0000000000000000000000010000000000000000000000000000000200000000",
            INIT_2E => X"0000000a00000000000000010000000000000000000000000000000300000000",
            INIT_2F => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000d00000000000000000000000000000000000000000000003c00000000",
            INIT_31 => X"0000000900000000000000090000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000400000000000000120000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_35 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_36 => X"0000000000000000000000090000000000000001000000000000000000000000",
            INIT_37 => X"0000000000000000000000350000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000011000000000000000d00000000",
            INIT_39 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_3A => X"00000000000000000000002b0000000000000022000000000000000f00000000",
            INIT_3B => X"0000000000000000000000180000000000000000000000000000000900000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_3D => X"0000004000000000000000000000000000000000000000000000000d00000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_3F => X"0000000900000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_44 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000002a00000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000e000000000000000e0000000000000012000000000000000000000000",
            INIT_48 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000050000000000000021000000000000000800000000",
            INIT_4C => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_50 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_51 => X"0000000c00000000000000080000000000000000000000000000000000000000",
            INIT_52 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_54 => X"0000009500000000000000860000000000000094000000000000000000000000",
            INIT_55 => X"0000007f000000000000009d0000000000000097000000000000009200000000",
            INIT_56 => X"0000003e00000000000000530000000000000060000000000000007200000000",
            INIT_57 => X"0000000c00000000000000140000000000000015000000000000002700000000",
            INIT_58 => X"0000006800000000000000870000000000000083000000000000009000000000",
            INIT_59 => X"0000007000000000000000870000000000000086000000000000008000000000",
            INIT_5A => X"0000004e000000000000004f0000000000000057000000000000005400000000",
            INIT_5B => X"00000080000000000000004f0000000000000058000000000000005100000000",
            INIT_5C => X"0000005c000000000000004d0000000000000057000000000000007e00000000",
            INIT_5D => X"0000007d000000000000006f0000000000000065000000000000005a00000000",
            INIT_5E => X"0000007f00000000000000940000000000000098000000000000009d00000000",
            INIT_5F => X"0000008200000000000000760000000000000051000000000000006f00000000",
            INIT_60 => X"0000005e000000000000004d000000000000002b000000000000005c00000000",
            INIT_61 => X"00000095000000000000007a0000000000000073000000000000006300000000",
            INIT_62 => X"000000670000000000000079000000000000009000000000000000a800000000",
            INIT_63 => X"000000de000000000000010600000000000000d7000000000000005400000000",
            INIT_64 => X"000000ac00000000000000940000000000000048000000000000003400000000",
            INIT_65 => X"0000008c00000000000000770000000000000079000000000000007d00000000",
            INIT_66 => X"0000007f00000000000000880000000000000095000000000000009600000000",
            INIT_67 => X"0000003b00000000000001050000000000000148000000000000013f00000000",
            INIT_68 => X"0000008a00000000000000ac00000000000000ac000000000000006400000000",
            INIT_69 => X"0000008b0000000000000075000000000000007c000000000000008c00000000",
            INIT_6A => X"0000012a000000000000009100000000000000a4000000000000009c00000000",
            INIT_6B => X"0000005c0000000000000076000000000000011d000000000000012600000000",
            INIT_6C => X"000000a800000000000000920000000000000097000000000000009500000000",
            INIT_6D => X"0000008e00000000000000800000000000000076000000000000008d00000000",
            INIT_6E => X"00000131000000000000011e000000000000006e000000000000009200000000",
            INIT_6F => X"0000008900000000000000a500000000000000fc000000000000012a00000000",
            INIT_70 => X"000000aa00000000000000c30000000000000098000000000000009800000000",
            INIT_71 => X"000000760000000000000083000000000000006f000000000000007f00000000",
            INIT_72 => X"000001a900000000000001800000000000000149000000000000006a00000000",
            INIT_73 => X"000000d300000000000000e3000000000000014f000000000000013d00000000",
            INIT_74 => X"0000009400000000000000b500000000000000bb000000000000009d00000000",
            INIT_75 => X"0000004600000000000000700000000000000085000000000000007900000000",
            INIT_76 => X"0000018200000000000001e6000000000000021400000000000001ea00000000",
            INIT_77 => X"000000a300000000000000d5000000000000010b000000000000014900000000",
            INIT_78 => X"0000008500000000000000b000000000000000bc00000000000000b300000000",
            INIT_79 => X"0000023a00000000000000170000000000000040000000000000007500000000",
            INIT_7A => X"000000bc00000000000000ef0000000000000113000000000000020c00000000",
            INIT_7B => X"000000ac0000000000000087000000000000009500000000000000ab00000000",
            INIT_7C => X"00000065000000000000008200000000000000a100000000000000af00000000",
            INIT_7D => X"0000014800000000000001900000000000000026000000000000006100000000",
            INIT_7E => X"00000055000000000000006d00000000000000c900000000000000dd00000000",
            INIT_7F => X"0000009200000000000000700000000000000052000000000000009100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE49;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE50 : if BRAM_NAME = "samplegold_layersamples_instance50" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000720000000000000056000000000000009d00000000000000a900000000",
            INIT_01 => X"000000bc00000000000000c200000000000000c8000000000000004600000000",
            INIT_02 => X"000000850000000000000067000000000000009200000000000000b400000000",
            INIT_03 => X"000000d600000000000000b20000000000000074000000000000006e00000000",
            INIT_04 => X"0000006c0000000000000050000000000000006b00000000000000ac00000000",
            INIT_05 => X"000000680000000000000091000000000000009b000000000000009700000000",
            INIT_06 => X"000000660000000000000059000000000000006a000000000000005300000000",
            INIT_07 => X"0000009400000000000000a10000000000000073000000000000005700000000",
            INIT_08 => X"0000006a000000000000004b000000000000003c000000000000006d00000000",
            INIT_09 => X"000000320000000000000025000000000000003b000000000000004a00000000",
            INIT_0A => X"00000027000000000000003b000000000000005a000000000000006900000000",
            INIT_0B => X"00000038000000000000004d000000000000003f000000000000003000000000",
            INIT_0C => X"0000000000000000000000000000000000000021000000000000002100000000",
            INIT_0D => X"0000000000000000000000000000000000000004000000000000000300000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"000000000000000000000035000000000000002a000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"00000000000000000000001b0000000000000033000000000000003700000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"000000230000000000000000000000000000000a000000000000000000000000",
            INIT_27 => X"00000000000000000000000d0000000000000025000000000000002700000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000003000000000000000280000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000080000000000000000000000000000001b00000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000007e00000000000000600000000000000040000000000000000000000000",
            INIT_2F => X"0000000c00000000000000020000000000000038000000000000002400000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000002b0000000000000010000000000000007c000000000000008800000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000008200000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000011000000000000006500000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000001900000000000000210000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000007000000000000001300000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"00000000000000000000000a000000000000000d000000000000000c00000000",
            INIT_46 => X"0000000a00000000000000060000000000000000000000000000000000000000",
            INIT_47 => X"0000000f000000000000000e000000000000000c000000000000000800000000",
            INIT_48 => X"0000000b000000000000000c0000000000000013000000000000001100000000",
            INIT_49 => X"000000000000000000000000000000000000000b000000000000000600000000",
            INIT_4A => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000a00000000000000090000000000000009000000000000000700000000",
            INIT_4C => X"00000005000000000000000b000000000000000a000000000000000a00000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000700000000000000060000000000000003000000000000000000000000",
            INIT_50 => X"00000000000000000000000e000000000000000a000000000000000900000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000d00000000000000020000000000000008000000000000000400000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000400000000000000040000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000004000000000000000400000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000e000000000000000b0000000000000009000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000b00000000000000000000000000000008000000000000000800000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000400000000000000020000000000000000000000000000000000000000",
            INIT_63 => X"000000000000000000000000000000000000000d000000000000000a00000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"00000003000000000000000b0000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000d0000000000000005000000000000000d000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000170000000000000013000000000000000300000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"000000000000000000000003000000000000000b000000000000000700000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000001c000000000000001d0000000000000014000000000000001500000000",
            INIT_7E => X"0000001c00000000000000230000000000000028000000000000002700000000",
            INIT_7F => X"0000001200000000000000160000000000000017000000000000001500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE50;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE51 : if BRAM_NAME = "samplegold_layersamples_instance51" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001400000000000000100000000000000014000000000000001100000000",
            INIT_01 => X"0000002c000000000000001e000000000000001c000000000000001200000000",
            INIT_02 => X"0000002300000000000000320000000000000035000000000000004000000000",
            INIT_03 => X"0000001f000000000000001b000000000000001b000000000000001a00000000",
            INIT_04 => X"0000001500000000000000150000000000000020000000000000002200000000",
            INIT_05 => X"0000003a000000000000002e000000000000001e000000000000001c00000000",
            INIT_06 => X"0000002d000000000000003c0000000000000047000000000000004300000000",
            INIT_07 => X"00000028000000000000002c000000000000002e000000000000002a00000000",
            INIT_08 => X"0000000b00000000000000160000000000000016000000000000002600000000",
            INIT_09 => X"0000003c0000000000000034000000000000002d000000000000002600000000",
            INIT_0A => X"0000003900000000000000460000000000000051000000000000005000000000",
            INIT_0B => X"0000002e0000000000000027000000000000002a000000000000003600000000",
            INIT_0C => X"00000019000000000000001e0000000000000024000000000000001c00000000",
            INIT_0D => X"00000040000000000000003b000000000000003c000000000000003200000000",
            INIT_0E => X"000000430000000000000051000000000000004f000000000000005000000000",
            INIT_0F => X"0000002d0000000000000040000000000000003c000000000000003e00000000",
            INIT_10 => X"0000002400000000000000150000000000000011000000000000002b00000000",
            INIT_11 => X"0000004300000000000000330000000000000039000000000000004100000000",
            INIT_12 => X"00000050000000000000004a000000000000004d000000000000004900000000",
            INIT_13 => X"0000002300000000000000260000000000000043000000000000004c00000000",
            INIT_14 => X"0000003e00000000000000330000000000000000000000000000002100000000",
            INIT_15 => X"0000003b00000000000000420000000000000040000000000000003200000000",
            INIT_16 => X"00000048000000000000004a000000000000004f000000000000004500000000",
            INIT_17 => X"0000002d00000000000000290000000000000024000000000000003100000000",
            INIT_18 => X"0000003500000000000000310000000000000014000000000000003300000000",
            INIT_19 => X"0000003f00000000000000330000000000000043000000000000004900000000",
            INIT_1A => X"0000002f000000000000003a0000000000000041000000000000004400000000",
            INIT_1B => X"000000290000000000000023000000000000002c000000000000002c00000000",
            INIT_1C => X"00000043000000000000003b0000000000000029000000000000003000000000",
            INIT_1D => X"0000003e00000000000000380000000000000031000000000000004000000000",
            INIT_1E => X"000000320000000000000041000000000000003e000000000000004400000000",
            INIT_1F => X"0000004a00000000000000180000000000000042000000000000003c00000000",
            INIT_20 => X"0000003b0000000000000038000000000000004f000000000000003300000000",
            INIT_21 => X"0000003d000000000000003a000000000000003a000000000000003400000000",
            INIT_22 => X"0000002d00000000000000320000000000000040000000000000003500000000",
            INIT_23 => X"000000410000000000000031000000000000002a000000000000000a00000000",
            INIT_24 => X"0000003e0000000000000040000000000000003a000000000000003b00000000",
            INIT_25 => X"00000040000000000000003d0000000000000035000000000000003d00000000",
            INIT_26 => X"00000009000000000000001c000000000000002a000000000000004600000000",
            INIT_27 => X"00000038000000000000002c000000000000001c000000000000002000000000",
            INIT_28 => X"0000003700000000000000380000000000000031000000000000002300000000",
            INIT_29 => X"0000003d00000000000000570000000000000043000000000000003700000000",
            INIT_2A => X"000000290000000000000021000000000000001e000000000000001800000000",
            INIT_2B => X"0000002a0000000000000044000000000000002d000000000000002700000000",
            INIT_2C => X"0000003b0000000000000030000000000000003d000000000000003600000000",
            INIT_2D => X"00000022000000000000004f0000000000000054000000000000003f00000000",
            INIT_2E => X"0000003b00000000000000380000000000000035000000000000002c00000000",
            INIT_2F => X"00000037000000000000003a0000000000000036000000000000003a00000000",
            INIT_30 => X"00000040000000000000002d0000000000000035000000000000003b00000000",
            INIT_31 => X"0000003700000000000000320000000000000056000000000000005000000000",
            INIT_32 => X"0000004c000000000000004e0000000000000042000000000000003c00000000",
            INIT_33 => X"0000004200000000000000490000000000000047000000000000003f00000000",
            INIT_34 => X"0000005200000000000000420000000000000040000000000000004100000000",
            INIT_35 => X"00000020000000000000001f000000000000001f000000000000005100000000",
            INIT_36 => X"0000002200000000000000270000000000000030000000000000001b00000000",
            INIT_37 => X"0000001f0000000000000022000000000000001d000000000000001d00000000",
            INIT_38 => X"0000001b000000000000001f000000000000001f000000000000001e00000000",
            INIT_39 => X"000000250000000000000024000000000000001e000000000000001f00000000",
            INIT_3A => X"0000003000000000000000320000000000000047000000000000003800000000",
            INIT_3B => X"0000001b000000000000001e0000000000000020000000000000001e00000000",
            INIT_3C => X"0000002200000000000000140000000000000017000000000000001900000000",
            INIT_3D => X"00000043000000000000002a0000000000000026000000000000002000000000",
            INIT_3E => X"00000026000000000000004e0000000000000056000000000000004d00000000",
            INIT_3F => X"00000016000000000000001b000000000000001b000000000000001f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002100000000000000220000000000000014000000000000001400000000",
            INIT_41 => X"00000055000000000000004f000000000000003d000000000000001000000000",
            INIT_42 => X"0000003700000000000000470000000000000053000000000000005200000000",
            INIT_43 => X"0000001300000000000000100000000000000021000000000000002d00000000",
            INIT_44 => X"0000001400000000000000170000000000000019000000000000001500000000",
            INIT_45 => X"00000043000000000000004e0000000000000050000000000000001e00000000",
            INIT_46 => X"0000005100000000000000510000000000000052000000000000004900000000",
            INIT_47 => X"000000120000000000000010000000000000001c000000000000003100000000",
            INIT_48 => X"0000001b00000000000000000000000000000013000000000000001400000000",
            INIT_49 => X"00000048000000000000004d0000000000000058000000000000003600000000",
            INIT_4A => X"0000004c00000000000000530000000000000052000000000000004f00000000",
            INIT_4B => X"00000013000000000000000b000000000000000e000000000000002e00000000",
            INIT_4C => X"0000004600000000000000000000000000000009000000000000000f00000000",
            INIT_4D => X"00000049000000000000004f000000000000003f000000000000004800000000",
            INIT_4E => X"000000330000000000000057000000000000004e000000000000004700000000",
            INIT_4F => X"000000140000000000000017000000000000000b000000000000001a00000000",
            INIT_50 => X"0000003d00000000000000000000000000000000000000000000001600000000",
            INIT_51 => X"000000440000000000000049000000000000004c000000000000003b00000000",
            INIT_52 => X"0000002800000000000000410000000000000054000000000000004e00000000",
            INIT_53 => X"00000000000000000000000c0000000000000016000000000000001500000000",
            INIT_54 => X"000000260000000000000011000000000000000b000000000000001500000000",
            INIT_55 => X"0000004d0000000000000049000000000000004f000000000000003c00000000",
            INIT_56 => X"000000140000000000000031000000000000004f000000000000005000000000",
            INIT_57 => X"0000000000000000000000040000000000000001000000000000000400000000",
            INIT_58 => X"000000310000000000000040000000000000000a000000000000003300000000",
            INIT_59 => X"0000004e000000000000004d000000000000004e000000000000005000000000",
            INIT_5A => X"00000000000000000000000c0000000000000023000000000000004e00000000",
            INIT_5B => X"00000043000000000000003d0000000000000000000000000000000000000000",
            INIT_5C => X"0000004e000000000000003c0000000000000049000000000000004000000000",
            INIT_5D => X"00000042000000000000004a0000000000000047000000000000004d00000000",
            INIT_5E => X"0000000b0000000000000007000000000000000c000000000000001700000000",
            INIT_5F => X"0000005300000000000000380000000000000016000000000000000000000000",
            INIT_60 => X"0000004e0000000000000053000000000000002c000000000000003f00000000",
            INIT_61 => X"00000024000000000000002e0000000000000042000000000000004400000000",
            INIT_62 => X"0000001a000000000000001a0000000000000017000000000000000200000000",
            INIT_63 => X"0000003f0000000000000029000000000000000f000000000000001b00000000",
            INIT_64 => X"00000040000000000000004f000000000000004c000000000000002b00000000",
            INIT_65 => X"0000001200000000000000230000000000000023000000000000004700000000",
            INIT_66 => X"0000001e00000000000000240000000000000021000000000000001e00000000",
            INIT_67 => X"000000380000000000000027000000000000001a000000000000001900000000",
            INIT_68 => X"000000460000000000000046000000000000004c000000000000003c00000000",
            INIT_69 => X"0000001f000000000000001f000000000000001b000000000000003b00000000",
            INIT_6A => X"000000190000000000000015000000000000001b000000000000001c00000000",
            INIT_6B => X"00000019000000000000001a0000000000000021000000000000001d00000000",
            INIT_6C => X"0000002100000000000000330000000000000037000000000000002400000000",
            INIT_6D => X"00000036000000000000003b0000000000000011000000000000001900000000",
            INIT_6E => X"0000002600000000000000320000000000000037000000000000003700000000",
            INIT_6F => X"000000250000000000000028000000000000002c000000000000002a00000000",
            INIT_70 => X"000000110000000000000015000000000000001c000000000000002100000000",
            INIT_71 => X"000000350000000000000035000000000000003a000000000000000b00000000",
            INIT_72 => X"0000001700000000000000210000000000000021000000000000002600000000",
            INIT_73 => X"00000013000000000000001d000000000000001d000000000000001800000000",
            INIT_74 => X"0000000c000000000000000c000000000000000a000000000000000d00000000",
            INIT_75 => X"00000018000000000000002d0000000000000035000000000000003800000000",
            INIT_76 => X"0000000300000000000000090000000000000009000000000000001500000000",
            INIT_77 => X"0000001b000000000000001b000000000000001f000000000000000600000000",
            INIT_78 => X"0000002e0000000000000013000000000000001a000000000000001800000000",
            INIT_79 => X"0000000b000000000000000a0000000000000019000000000000002f00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_7B => X"00000018000000000000001e0000000000000025000000000000001e00000000",
            INIT_7C => X"00000036000000000000002e0000000000000005000000000000001400000000",
            INIT_7D => X"0000001600000000000000080000000000000000000000000000003600000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_7F => X"000000010000000000000011000000000000000d000000000000000c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE51;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE52 : if BRAM_NAME = "samplegold_layersamples_instance52" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000049000000000000005b0000000000000052000000000000000000000000",
            INIT_01 => X"0000002600000000000000220000000000000007000000000000000200000000",
            INIT_02 => X"0000000000000000000000000000000000000004000000000000000e00000000",
            INIT_03 => X"000000000000000000000000000000000000000b000000000000000800000000",
            INIT_04 => X"0000000a000000000000004e0000000000000058000000000000005c00000000",
            INIT_05 => X"0000000f00000000000000150000000000000021000000000000001e00000000",
            INIT_06 => X"0000000300000000000000000000000000000008000000000000001400000000",
            INIT_07 => X"0000005300000000000000100000000000000010000000000000000900000000",
            INIT_08 => X"000000030000000000000029000000000000004f000000000000005000000000",
            INIT_09 => X"0000001c0000000000000005000000000000000b000000000000001000000000",
            INIT_0A => X"0000001000000000000000000000000000000003000000000000001900000000",
            INIT_0B => X"000000550000000000000051000000000000000a000000000000001100000000",
            INIT_0C => X"00000025000000000000003b000000000000003a000000000000005100000000",
            INIT_0D => X"0000002300000000000000240000000000000003000000000000001a00000000",
            INIT_0E => X"0000000b00000000000000100000000000000004000000000000000d00000000",
            INIT_0F => X"0000008600000000000000780000000000000065000000000000000000000000",
            INIT_10 => X"0000002b0000000000000038000000000000005b000000000000005f00000000",
            INIT_11 => X"0000001900000000000000270000000000000020000000000000000700000000",
            INIT_12 => X"000000000000000000000000000000000000000c000000000000000900000000",
            INIT_13 => X"0000006000000000000000550000000000000097000000000000009b00000000",
            INIT_14 => X"0000000d000000000000001f0000000000000031000000000000003b00000000",
            INIT_15 => X"000000080000000000000015000000000000001e000000000000001800000000",
            INIT_16 => X"0000009600000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000001d0000000000000030000000000000003f000000000000008600000000",
            INIT_18 => X"0000001b000000000000000c0000000000000017000000000000000c00000000",
            INIT_19 => X"00000000000000000000000f0000000000000018000000000000001900000000",
            INIT_1A => X"00000047000000000000004d0000000000000000000000000000000000000000",
            INIT_1B => X"000000070000000000000015000000000000002f000000000000003f00000000",
            INIT_1C => X"000000200000000000000013000000000000000c000000000000001500000000",
            INIT_1D => X"000000000000000000000000000000000000001f000000000000002e00000000",
            INIT_1E => X"000000240000000000000028000000000000002e000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000004000000000000001500000000",
            INIT_20 => X"0000002f000000000000001b0000000000000000000000000000000900000000",
            INIT_21 => X"0000000000000000000000000000000000000002000000000000001d00000000",
            INIT_22 => X"000000000000000000000000000000000000000a000000000000001a00000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"00000028000000000000001a0000000000000019000000000000001a00000000",
            INIT_27 => X"0000001e00000000000000250000000000000031000000000000003800000000",
            INIT_28 => X"00000020000000000000001f0000000000000021000000000000001e00000000",
            INIT_29 => X"0000001a00000000000000190000000000000021000000000000001e00000000",
            INIT_2A => X"000000460000000000000035000000000000002a000000000000001a00000000",
            INIT_2B => X"0000002300000000000000330000000000000048000000000000004b00000000",
            INIT_2C => X"000000240000000000000029000000000000002a000000000000002c00000000",
            INIT_2D => X"0000001f000000000000001b000000000000001b000000000000002400000000",
            INIT_2E => X"0000005f00000000000000560000000000000044000000000000002900000000",
            INIT_2F => X"00000029000000000000002d0000000000000053000000000000006700000000",
            INIT_30 => X"0000002600000000000000210000000000000028000000000000002c00000000",
            INIT_31 => X"000000360000000000000026000000000000001e000000000000001f00000000",
            INIT_32 => X"00000065000000000000005f0000000000000059000000000000004e00000000",
            INIT_33 => X"0000003e000000000000003d000000000000004f000000000000006500000000",
            INIT_34 => X"0000002100000000000000310000000000000029000000000000002e00000000",
            INIT_35 => X"0000004b0000000000000041000000000000001b000000000000001e00000000",
            INIT_36 => X"0000006b0000000000000060000000000000004e000000000000004700000000",
            INIT_37 => X"0000004000000000000000560000000000000066000000000000006e00000000",
            INIT_38 => X"0000001a0000000000000019000000000000003c000000000000003b00000000",
            INIT_39 => X"000000460000000000000041000000000000003d000000000000001e00000000",
            INIT_3A => X"00000069000000000000005f000000000000005c000000000000005200000000",
            INIT_3B => X"0000003d00000000000000510000000000000062000000000000006f00000000",
            INIT_3C => X"0000001f000000000000001a0000000000000016000000000000003600000000",
            INIT_3D => X"00000056000000000000003c0000000000000031000000000000003300000000",
            INIT_3E => X"0000006600000000000000580000000000000057000000000000006100000000",
            INIT_3F => X"0000002a00000000000000350000000000000050000000000000006600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000031000000000000001f0000000000000020000000000000001f00000000",
            INIT_41 => X"0000005b000000000000004b000000000000003c000000000000003800000000",
            INIT_42 => X"0000006700000000000000630000000000000055000000000000005500000000",
            INIT_43 => X"0000002000000000000000390000000000000044000000000000005400000000",
            INIT_44 => X"0000002b00000000000000320000000000000023000000000000002100000000",
            INIT_45 => X"0000005600000000000000590000000000000038000000000000003400000000",
            INIT_46 => X"0000005b0000000000000065000000000000005f000000000000005300000000",
            INIT_47 => X"0000000d0000000000000015000000000000003e000000000000004b00000000",
            INIT_48 => X"0000003700000000000000310000000000000021000000000000001300000000",
            INIT_49 => X"000000560000000000000059000000000000005e000000000000003f00000000",
            INIT_4A => X"0000004f000000000000005f0000000000000066000000000000005c00000000",
            INIT_4B => X"00000035000000000000000c000000000000000c000000000000003f00000000",
            INIT_4C => X"0000005200000000000000510000000000000040000000000000003400000000",
            INIT_4D => X"0000005a00000000000000590000000000000056000000000000005200000000",
            INIT_4E => X"000000410000000000000048000000000000005f000000000000006300000000",
            INIT_4F => X"0000002600000000000000250000000000000018000000000000000d00000000",
            INIT_50 => X"0000004100000000000000490000000000000052000000000000003f00000000",
            INIT_51 => X"00000055000000000000004d0000000000000056000000000000004600000000",
            INIT_52 => X"0000002200000000000000450000000000000046000000000000005e00000000",
            INIT_53 => X"0000003400000000000000290000000000000024000000000000001e00000000",
            INIT_54 => X"00000048000000000000004a000000000000003f000000000000003900000000",
            INIT_55 => X"0000005a00000000000000500000000000000043000000000000004e00000000",
            INIT_56 => X"0000002b00000000000000280000000000000042000000000000004e00000000",
            INIT_57 => X"0000003a0000000000000041000000000000003b000000000000003100000000",
            INIT_58 => X"0000004b0000000000000053000000000000004c000000000000004200000000",
            INIT_59 => X"0000005300000000000000540000000000000053000000000000004600000000",
            INIT_5A => X"000000420000000000000039000000000000002e000000000000004600000000",
            INIT_5B => X"00000043000000000000003c0000000000000041000000000000004300000000",
            INIT_5C => X"0000004b000000000000004b000000000000004d000000000000004e00000000",
            INIT_5D => X"00000044000000000000004b0000000000000050000000000000004f00000000",
            INIT_5E => X"0000000200000000000000150000000000000000000000000000000100000000",
            INIT_5F => X"0000000000000000000000000000000000000001000000000000000900000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000100000000000000000000000000000005000000000000000000000000",
            INIT_62 => X"000000000000000000000006000000000000000d000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000100000000000000040000000000000000000000000000000000000000",
            INIT_66 => X"000000050000000000000000000000000000001c000000000000000000000000",
            INIT_67 => X"000000000000000000000008000000000000000a000000000000000c00000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000070000000000000004000000000000000000000000",
            INIT_6A => X"000000060000000000000005000000000000000b000000000000000100000000",
            INIT_6B => X"0000000700000000000000160000000000000009000000000000000b00000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_6E => X"0000000000000000000000000000000000000028000000000000000c00000000",
            INIT_6F => X"0000000000000000000000120000000000000002000000000000000000000000",
            INIT_70 => X"0000000b00000000000000000000000000000000000000000000000300000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_72 => X"0000000100000000000000000000000000000000000000000000002e00000000",
            INIT_73 => X"0000001900000000000000190000000000000000000000000000000000000000",
            INIT_74 => X"00000007000000000000000e0000000000000000000000000000000000000000",
            INIT_75 => X"0000003c00000000000000160000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000060000000000000003000000000000000000000000",
            INIT_77 => X"000000110000000000000003000000000000001d000000000000000000000000",
            INIT_78 => X"000000000000000000000008000000000000000c000000000000000000000000",
            INIT_79 => X"0000000000000000000000130000000000000000000000000000000000000000",
            INIT_7A => X"000000000000000000000000000000000000000b000000000000000d00000000",
            INIT_7B => X"0000000000000000000000090000000000000006000000000000000100000000",
            INIT_7C => X"0000000000000000000000000000000000000015000000000000001200000000",
            INIT_7D => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_7F => X"0000000000000000000000000000000000000004000000000000001100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE52;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE53 : if BRAM_NAME = "samplegold_layersamples_instance53" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001100000000000000000000000000000000000000000000000200000000",
            INIT_01 => X"0000000a00000000000000000000000000000018000000000000000000000000",
            INIT_02 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000180000000000000000000000000000000000000000",
            INIT_05 => X"00000006000000000000000b0000000000000012000000000000001300000000",
            INIT_06 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000040000000000000007000000000000000000000000",
            INIT_08 => X"0000001d00000000000000170000000000000000000000000000000000000000",
            INIT_09 => X"0000000200000000000000190000000000000023000000000000000000000000",
            INIT_0A => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_0B => X"000000030000000000000006000000000000000f000000000000000500000000",
            INIT_0C => X"00000000000000000000001f0000000000000000000000000000000000000000",
            INIT_0D => X"000000000000000000000000000000000000002b000000000000000c00000000",
            INIT_0E => X"000000070000000000000007000000000000000b000000000000000000000000",
            INIT_0F => X"0000001100000000000000040000000000000003000000000000000800000000",
            INIT_10 => X"0000000d00000000000000010000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000020000000000000002c00000000",
            INIT_12 => X"0000000900000000000000020000000000000018000000000000000100000000",
            INIT_13 => X"00000011000000000000001b0000000000000000000000000000000900000000",
            INIT_14 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000900000000000000000000000000000017000000000000001c00000000",
            INIT_16 => X"0000000500000000000000010000000000000000000000000000000400000000",
            INIT_17 => X"000000000000000000000001000000000000000b000000000000000b00000000",
            INIT_18 => X"0000000700000000000000010000000000000000000000000000000400000000",
            INIT_19 => X"0000000000000000000000000000000000000002000000000000000600000000",
            INIT_1A => X"0000001200000000000000040000000000000000000000000000000100000000",
            INIT_1B => X"00000000000000000000000c0000000000000021000000000000000200000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_1D => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"00000010000000000000001a0000000000000014000000000000000600000000",
            INIT_1F => X"0000000000000000000000090000000000000014000000000000000a00000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"000000000000000000000000000000000000000c000000000000000500000000",
            INIT_22 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_23 => X"0000002200000000000000100000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000004000000000000000500000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000010000000000000008000000000000000000000000",
            INIT_27 => X"0000001400000000000000080000000000000003000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000300000000000000070000000000000000000000000000000000000000",
            INIT_2B => X"0000001500000000000000040000000000000000000000000000000000000000",
            INIT_2C => X"0000001200000000000000000000000000000000000000000000000500000000",
            INIT_2D => X"0000000b00000000000000000000000000000000000000000000000e00000000",
            INIT_2E => X"0000000000000000000000020000000000000012000000000000003900000000",
            INIT_2F => X"0000000e00000000000000100000000000000001000000000000000000000000",
            INIT_30 => X"000000000000000000000000000000000000001e000000000000001d00000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000a000000000000000f0000000000000007000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_37 => X"000000200000000000000009000000000000000b000000000000000000000000",
            INIT_38 => X"0000000100000000000000160000000000000000000000000000000000000000",
            INIT_39 => X"00000000000000000000000b0000000000000000000000000000002900000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_3B => X"0000000000000000000000010000000000000008000000000000001000000000",
            INIT_3C => X"00000040000000000000004e000000000000003a000000000000000000000000",
            INIT_3D => X"0000000d0000000000000030000000000000002c000000000000004f00000000",
            INIT_3E => X"0000000000000000000000010000000000000010000000000000000f00000000",
            INIT_3F => X"0000007f00000000000000850000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002000000000000000000000000000000000000000000000001600000000",
            INIT_41 => X"0000001100000000000000220000000000000000000000000000000000000000",
            INIT_42 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000001200000000000000280000000000000030000000000000000000000000",
            INIT_44 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000400000000000000010000000000000000000000000000000000000000",
            INIT_47 => X"0000003000000000000000130000000000000000000000000000000500000000",
            INIT_48 => X"0000000400000000000000000000000000000000000000000000002600000000",
            INIT_49 => X"000000110000000000000041000000000000002c000000000000001100000000",
            INIT_4A => X"0000001b0000000000000012000000000000000e000000000000000c00000000",
            INIT_4B => X"0000000600000000000000000000000000000018000000000000003000000000",
            INIT_4C => X"0000000100000000000000050000000000000000000000000000000400000000",
            INIT_4D => X"0000000f000000000000001d0000000000000011000000000000000000000000",
            INIT_4E => X"0000002e0000000000000032000000000000000d000000000000000700000000",
            INIT_4F => X"0000004900000000000000450000000000000031000000000000003800000000",
            INIT_50 => X"0000002500000000000000260000000000000027000000000000003700000000",
            INIT_51 => X"00000013000000000000000d0000000000000010000000000000001800000000",
            INIT_52 => X"00000035000000000000002c0000000000000030000000000000001000000000",
            INIT_53 => X"0000004d0000000000000059000000000000004d000000000000002e00000000",
            INIT_54 => X"0000002f00000000000000290000000000000024000000000000004500000000",
            INIT_55 => X"000000380000000000000040000000000000003d000000000000003600000000",
            INIT_56 => X"0000002f00000000000000240000000000000029000000000000002b00000000",
            INIT_57 => X"0000006700000000000000610000000000000059000000000000004500000000",
            INIT_58 => X"0000005000000000000000550000000000000057000000000000005800000000",
            INIT_59 => X"0000002d00000000000000290000000000000036000000000000004400000000",
            INIT_5A => X"0000004d00000000000000400000000000000024000000000000003200000000",
            INIT_5B => X"000000700000000000000080000000000000006f000000000000005f00000000",
            INIT_5C => X"0000003700000000000000480000000000000056000000000000005100000000",
            INIT_5D => X"0000007e0000000000000066000000000000003c000000000000003800000000",
            INIT_5E => X"0000006f00000000000000590000000000000036000000000000006300000000",
            INIT_5F => X"00000075000000000000007c000000000000007b000000000000008000000000",
            INIT_60 => X"000000590000000000000055000000000000005f000000000000006e00000000",
            INIT_61 => X"000000380000000000000071000000000000007a000000000000005f00000000",
            INIT_62 => X"0000006c00000000000000800000000000000053000000000000003a00000000",
            INIT_63 => X"0000007d00000000000000830000000000000079000000000000006900000000",
            INIT_64 => X"0000005b0000000000000066000000000000006b000000000000006f00000000",
            INIT_65 => X"0000003500000000000000540000000000000058000000000000005c00000000",
            INIT_66 => X"0000007100000000000000610000000000000062000000000000005000000000",
            INIT_67 => X"0000007c00000000000000750000000000000075000000000000007600000000",
            INIT_68 => X"0000006000000000000000340000000000000052000000000000006800000000",
            INIT_69 => X"00000052000000000000005f000000000000006f000000000000006e00000000",
            INIT_6A => X"0000007d00000000000000840000000000000075000000000000007500000000",
            INIT_6B => X"0000005d00000000000000740000000000000073000000000000006f00000000",
            INIT_6C => X"0000008d000000000000007d0000000000000040000000000000004900000000",
            INIT_6D => X"00000071000000000000008900000000000000a5000000000000009e00000000",
            INIT_6E => X"0000006b00000000000000740000000000000081000000000000007300000000",
            INIT_6F => X"0000005a000000000000006b0000000000000071000000000000007500000000",
            INIT_70 => X"000000a100000000000000d000000000000000ca000000000000003800000000",
            INIT_71 => X"000000780000000000000055000000000000007c000000000000006000000000",
            INIT_72 => X"0000007a00000000000000720000000000000074000000000000006f00000000",
            INIT_73 => X"00000037000000000000003d0000000000000066000000000000007100000000",
            INIT_74 => X"00000035000000000000002c000000000000009100000000000000a900000000",
            INIT_75 => X"0000005c000000000000005b0000000000000045000000000000005400000000",
            INIT_76 => X"00000068000000000000006b0000000000000072000000000000007600000000",
            INIT_77 => X"0000004700000000000000480000000000000055000000000000006300000000",
            INIT_78 => X"00000044000000000000004f0000000000000034000000000000002100000000",
            INIT_79 => X"0000005300000000000000460000000000000064000000000000005200000000",
            INIT_7A => X"0000005e00000000000000720000000000000072000000000000006600000000",
            INIT_7B => X"00000034000000000000002d0000000000000048000000000000006400000000",
            INIT_7C => X"0000005f000000000000004a000000000000004d000000000000003700000000",
            INIT_7D => X"0000007b00000000000000620000000000000044000000000000006200000000",
            INIT_7E => X"0000005f00000000000000610000000000000070000000000000007400000000",
            INIT_7F => X"00000049000000000000004c000000000000003a000000000000005500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE53;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE54 : if BRAM_NAME = "samplegold_layersamples_instance54" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005300000000000000480000000000000032000000000000003400000000",
            INIT_01 => X"0000004b000000000000005b0000000000000056000000000000005600000000",
            INIT_02 => X"0000005900000000000000520000000000000060000000000000005d00000000",
            INIT_03 => X"000000400000000000000035000000000000002c000000000000003a00000000",
            INIT_04 => X"0000004b00000000000000540000000000000056000000000000005100000000",
            INIT_05 => X"0000004c000000000000004e0000000000000049000000000000004c00000000",
            INIT_06 => X"0000000e00000000000000460000000000000051000000000000004600000000",
            INIT_07 => X"0000000b00000000000000180000000000000001000000000000001100000000",
            INIT_08 => X"0000001000000000000000140000000000000018000000000000000e00000000",
            INIT_09 => X"000000090000000000000010000000000000000f000000000000000b00000000",
            INIT_0A => X"00000013000000000000000e0000000000000002000000000000000000000000",
            INIT_0B => X"00000000000000000000000c000000000000000e000000000000000400000000",
            INIT_0C => X"0000000600000000000000130000000000000011000000000000001900000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_0E => X"00000019000000000000000f000000000000000d000000000000000900000000",
            INIT_0F => X"0000000000000000000000000000000000000004000000000000000500000000",
            INIT_10 => X"0000000c00000000000000040000000000000000000000000000000000000000",
            INIT_11 => X"0000001b00000000000000180000000000000012000000000000000e00000000",
            INIT_12 => X"00000000000000000000001e0000000000000003000000000000000800000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"00000020000000000000000d0000000000000001000000000000000000000000",
            INIT_15 => X"0000000000000000000000110000000000000017000000000000001200000000",
            INIT_16 => X"000000000000000000000031000000000000003a000000000000000000000000",
            INIT_17 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_18 => X"0000000b000000000000000b0000000000000000000000000000000000000000",
            INIT_19 => X"000000210000000000000012000000000000000f000000000000001500000000",
            INIT_1A => X"0000000000000000000000000000000000000029000000000000006900000000",
            INIT_1B => X"000000000000000000000000000000000000000d000000000000000700000000",
            INIT_1C => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000003100000000000000290000000000000023000000000000001a00000000",
            INIT_1E => X"0000001e00000000000000000000000000000000000000000000005f00000000",
            INIT_1F => X"0000000300000000000000020000000000000000000000000000000000000000",
            INIT_20 => X"0000002600000000000000080000000000000003000000000000000000000000",
            INIT_21 => X"0000003900000000000000270000000000000013000000000000001500000000",
            INIT_22 => X"0000000000000000000000090000000000000000000000000000005900000000",
            INIT_23 => X"0000000000000000000000070000000000000014000000000000000000000000",
            INIT_24 => X"0000000e00000000000000100000000000000002000000000000000000000000",
            INIT_25 => X"0000002f00000000000000270000000000000014000000000000000700000000",
            INIT_26 => X"0000000000000000000000130000000000000005000000000000003d00000000",
            INIT_27 => X"0000000000000000000000010000000000000003000000000000000c00000000",
            INIT_28 => X"0000001e0000000000000002000000000000002e000000000000000800000000",
            INIT_29 => X"00000062000000000000001e000000000000009d000000000000005900000000",
            INIT_2A => X"000000000000000000000000000000000000002c000000000000000000000000",
            INIT_2B => X"0000001e0000000000000000000000000000000f000000000000000400000000",
            INIT_2C => X"000000b000000000000000640000000000000044000000000000000c00000000",
            INIT_2D => X"00000005000000000000002c0000000000000013000000000000002800000000",
            INIT_2E => X"0000001000000000000000020000000000000000000000000000000a00000000",
            INIT_2F => X"00000017000000000000000a0000000000000000000000000000000800000000",
            INIT_30 => X"00000032000000000000004d0000000000000066000000000000007c00000000",
            INIT_31 => X"0000001e00000000000000000000000000000000000000000000002600000000",
            INIT_32 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000002c000000000000002e0000000000000000000000000000001200000000",
            INIT_34 => X"0000002f0000000000000013000000000000001b000000000000002500000000",
            INIT_35 => X"0000000000000000000000190000000000000000000000000000001100000000",
            INIT_36 => X"0000001f000000000000000d0000000000000005000000000000000000000000",
            INIT_37 => X"0000000b000000000000000d0000000000000008000000000000000000000000",
            INIT_38 => X"000000090000000000000019000000000000002d000000000000001e00000000",
            INIT_39 => X"0000000000000000000000040000000000000007000000000000000200000000",
            INIT_3A => X"00000010000000000000000c000000000000000c000000000000000500000000",
            INIT_3B => X"0000001300000000000000240000000000000021000000000000000000000000",
            INIT_3C => X"0000001000000000000000000000000000000000000000000000000d00000000",
            INIT_3D => X"000000000000000000000003000000000000000b000000000000001900000000",
            INIT_3E => X"0000000900000000000000020000000000000016000000000000000700000000",
            INIT_3F => X"00000040000000000000002a000000000000003a000000000000003900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003800000000000000420000000000000043000000000000003c00000000",
            INIT_41 => X"000000260000000000000028000000000000002c000000000000003200000000",
            INIT_42 => X"000000390000000000000015000000000000000e000000000000001c00000000",
            INIT_43 => X"00000040000000000000002f000000000000002e000000000000003e00000000",
            INIT_44 => X"0000002f000000000000003a000000000000004e000000000000002a00000000",
            INIT_45 => X"0000001b00000000000000200000000000000024000000000000002a00000000",
            INIT_46 => X"0000003800000000000000340000000000000025000000000000001a00000000",
            INIT_47 => X"0000002a00000000000000390000000000000025000000000000003b00000000",
            INIT_48 => X"0000002e0000000000000023000000000000002d000000000000002a00000000",
            INIT_49 => X"0000003c0000000000000036000000000000003b000000000000003a00000000",
            INIT_4A => X"0000004d000000000000002c000000000000002f000000000000003c00000000",
            INIT_4B => X"0000002200000000000000220000000000000023000000000000001000000000",
            INIT_4C => X"000000420000000000000033000000000000002d000000000000002800000000",
            INIT_4D => X"00000033000000000000003b0000000000000039000000000000004f00000000",
            INIT_4E => X"0000004f00000000000000800000000000000033000000000000002800000000",
            INIT_4F => X"0000004800000000000000380000000000000015000000000000001600000000",
            INIT_50 => X"00000044000000000000002e0000000000000033000000000000003400000000",
            INIT_51 => X"0000005600000000000000380000000000000041000000000000003500000000",
            INIT_52 => X"0000002b000000000000004a00000000000000ba000000000000006900000000",
            INIT_53 => X"0000003300000000000000540000000000000047000000000000000100000000",
            INIT_54 => X"0000002e00000000000000270000000000000036000000000000003900000000",
            INIT_55 => X"0000006e00000000000000680000000000000049000000000000004600000000",
            INIT_56 => X"0000001d00000000000000120000000000000095000000000000007a00000000",
            INIT_57 => X"000000470000000000000030000000000000003c000000000000005d00000000",
            INIT_58 => X"00000038000000000000003c0000000000000019000000000000004400000000",
            INIT_59 => X"00000070000000000000005b000000000000005a000000000000004e00000000",
            INIT_5A => X"000000490000000000000000000000000000008c000000000000007800000000",
            INIT_5B => X"00000049000000000000005b0000000000000033000000000000002c00000000",
            INIT_5C => X"00000039000000000000002c0000000000000035000000000000002e00000000",
            INIT_5D => X"00000079000000000000007d000000000000005c000000000000005700000000",
            INIT_5E => X"0000004e00000000000000520000000000000088000000000000008e00000000",
            INIT_5F => X"00000042000000000000004a0000000000000056000000000000003100000000",
            INIT_60 => X"0000006b000000000000004a0000000000000032000000000000002100000000",
            INIT_61 => X"0000006b000000000000010800000000000000b1000000000000008500000000",
            INIT_62 => X"00000033000000000000006f000000000000003600000000000000ba00000000",
            INIT_63 => X"000000290000000000000050000000000000004a000000000000004500000000",
            INIT_64 => X"000000d600000000000000b60000000000000028000000000000004700000000",
            INIT_65 => X"0000006c000000000000005b000000000000007e00000000000000f100000000",
            INIT_66 => X"00000043000000000000003a0000000000000044000000000000003e00000000",
            INIT_67 => X"00000037000000000000002f000000000000004c000000000000004f00000000",
            INIT_68 => X"0000009c00000000000000b400000000000000c7000000000000002f00000000",
            INIT_69 => X"0000001c0000000000000021000000000000005a000000000000006a00000000",
            INIT_6A => X"00000036000000000000002a000000000000001d000000000000004400000000",
            INIT_6B => X"0000005500000000000000180000000000000041000000000000004f00000000",
            INIT_6C => X"0000004900000000000000510000000000000054000000000000006800000000",
            INIT_6D => X"00000051000000000000001d0000000000000036000000000000005f00000000",
            INIT_6E => X"00000055000000000000004c0000000000000015000000000000001d00000000",
            INIT_6F => X"0000003f00000000000000330000000000000023000000000000005a00000000",
            INIT_70 => X"00000037000000000000004e0000000000000047000000000000003900000000",
            INIT_71 => X"0000002600000000000000340000000000000026000000000000003700000000",
            INIT_72 => X"00000046000000000000004b000000000000003b000000000000001800000000",
            INIT_73 => X"0000004000000000000000410000000000000018000000000000003200000000",
            INIT_74 => X"00000024000000000000000e000000000000002c000000000000003400000000",
            INIT_75 => X"000000220000000000000025000000000000003c000000000000003900000000",
            INIT_76 => X"0000001f000000000000003b000000000000002b000000000000001400000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000010000000000000001000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000c00000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE54;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE55 : if BRAM_NAME = "samplegold_layersamples_instance55" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000130000000000000016000000000000001100000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000001400000000000000120000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000110000000000000020000000000000001c00000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000900000000000000090000000000000009000000000000000e00000000",
            INIT_08 => X"0000000e00000000000000190000000000000022000000000000002000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_0A => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000001c00000000000000070000000000000000000000000000000600000000",
            INIT_0C => X"0000001100000000000000200000000000000028000000000000001a00000000",
            INIT_0D => X"0000000000000000000000000000000000000003000000000000000200000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000800000000000000120000000000000013000000000000000f00000000",
            INIT_10 => X"0000000900000000000000150000000000000020000000000000001a00000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000e00000000000000040000000000000017000000000000000d00000000",
            INIT_14 => X"0000000000000000000000070000000000000018000000000000001e00000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"00000018000000000000000d0000000000000006000000000000001400000000",
            INIT_18 => X"0000000500000000000000000000000000000007000000000000001700000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000001900000000000000040000000000000000000000000000000000000000",
            INIT_1B => X"0000001700000000000000110000000000000009000000000000000500000000",
            INIT_1C => X"00000000000000000000000b0000000000000009000000000000000a00000000",
            INIT_1D => X"0000000900000000000000040000000000000000000000000000000000000000",
            INIT_1E => X"000000100000000000000020000000000000000d000000000000001200000000",
            INIT_1F => X"0000000c000000000000001a0000000000000015000000000000000a00000000",
            INIT_20 => X"0000000000000000000000000000000000000004000000000000000500000000",
            INIT_21 => X"00000019000000000000000b0000000000000000000000000000000000000000",
            INIT_22 => X"0000001100000000000000170000000000000002000000000000000000000000",
            INIT_23 => X"0000000800000000000000100000000000000011000000000000000b00000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_25 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000040000000000000005000000000000000400000000",
            INIT_27 => X"0000000b000000000000000c0000000000000014000000000000000f00000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000700000000000000040000000000000002000000000000000700000000",
            INIT_2A => X"0000001200000000000000070000000000000005000000000000000b00000000",
            INIT_2B => X"00000000000000000000000c0000000000000016000000000000001400000000",
            INIT_2C => X"0000000c000000000000000d000000000000000c000000000000000400000000",
            INIT_2D => X"0000001100000000000000140000000000000009000000000000000300000000",
            INIT_2E => X"00000014000000000000000e0000000000000009000000000000000b00000000",
            INIT_2F => X"0000000000000000000000000000000000000010000000000000001700000000",
            INIT_30 => X"0000000000000000000000010000000000000002000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000050000000000000007000000000000000400000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000b00000000000000120000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000190000000000000010000000000000000300000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000400000000000000070000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000006000000000000000600000000",
            INIT_3F => X"0000000000000000000000000000000000000006000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000001500000000000000120000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000006000000000000000400000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000250000000000000017000000000000000200000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000500000000000000000000000000000000000000000000003c00000000",
            INIT_52 => X"0000000000000000000000000000000000000002000000000000000300000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000002400000000000000170000000000000000000000000000000000000000",
            INIT_55 => X"00000024000000000000004a0000000000000000000000000000000000000000",
            INIT_56 => X"000000090000000000000007000000000000001d000000000000001500000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000004d000000000000001e0000000000000000000000000000000000000000",
            INIT_59 => X"0000000300000000000000000000000000000005000000000000004700000000",
            INIT_5A => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_5B => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"000000120000000000000014000000000000001a000000000000001200000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_5F => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000001900000000000000000000000000000000000000000000001300000000",
            INIT_61 => X"000000030000000000000009000000000000002f000000000000003800000000",
            INIT_62 => X"00000008000000000000000e0000000000000008000000000000000500000000",
            INIT_63 => X"0000002a00000000000000240000000000000007000000000000000000000000",
            INIT_64 => X"00000024000000000000002c000000000000003c000000000000002600000000",
            INIT_65 => X"0000002700000000000000160000000000000018000000000000002200000000",
            INIT_66 => X"00000023000000000000001a0000000000000017000000000000002500000000",
            INIT_67 => X"000000000000000000000032000000000000002c000000000000002500000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000110000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE55;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE56 : if BRAM_NAME = "samplegold_layersamples_instance56" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000800000000000000060000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000012000000000000001b00000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000020000000000000008000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"000000000000000000000004000000000000000e000000000000003600000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000005000000000000000200000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000030000000000000008000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"000000000000000000000034000000000000005c000000000000000000000000",
            INIT_21 => X"0000000500000000000000000000000000000002000000000000000000000000",
            INIT_22 => X"00000019000000000000005d0000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000c0000000000000000000000000000005c000000000000002f00000000",
            INIT_25 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_26 => X"000000000000000000000000000000000000009b000000000000000000000000",
            INIT_27 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"000000000000000000000030000000000000000e000000000000008900000000",
            INIT_29 => X"0000000200000000000000000000000000000002000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000004000000000000004a00000000",
            INIT_2B => X"0000008600000000000000660000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000031000000000000000000000000",
            INIT_2D => X"00000001000000000000003d000000000000000c000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_2F => X"000000000000000000000000000000000000002e000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000004d00000000",
            INIT_31 => X"000000320000000000000016000000000000001a000000000000000b00000000",
            INIT_32 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_33 => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"00000000000000000000003e000000000000000b000000000000002400000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000600000000000000000000000000000021000000000000000000000000",
            INIT_38 => X"0000000c00000000000000000000000000000001000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000039000000000000000e00000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000006300000000",
            INIT_3C => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_3E => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000008000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000000000000000000000b0000000000000000000000000000000f00000000",
            INIT_41 => X"00000000000000000000001d0000000000000000000000000000001e00000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000c00000000000000010000000000000000000000000000002500000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_48 => X"0000000000000000000000010000000000000010000000000000000000000000",
            INIT_49 => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_4D => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_4E => X"00000000000000000000001b0000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000000000000000000009000000000000000d000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_53 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000006000000000000001100000000",
            INIT_55 => X"000000000000000000000000000000000000001d000000000000000000000000",
            INIT_56 => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000b00000000000000000000000000000002000000000000000000000000",
            INIT_58 => X"0000012d000000000000006b0000000000000000000000000000000000000000",
            INIT_59 => X"00000120000000000000011a000000000000010f000000000000011500000000",
            INIT_5A => X"000000eb0000000000000077000000000000011a000000000000012d00000000",
            INIT_5B => X"0000014e0000000000000159000000000000015c000000000000016c00000000",
            INIT_5C => X"0000011300000000000001130000000000000025000000000000000000000000",
            INIT_5D => X"0000015a0000000000000133000000000000011f000000000000015700000000",
            INIT_5E => X"000001a3000000000000014e00000000000000b7000000000000015600000000",
            INIT_5F => X"00000000000000000000016d000000000000017b000000000000018a00000000",
            INIT_60 => X"00000192000000000000011300000000000000f8000000000000000000000000",
            INIT_61 => X"000000ff00000000000000fe00000000000000d9000000000000012900000000",
            INIT_62 => X"000001b800000000000001b2000000000000018f000000000000010a00000000",
            INIT_63 => X"0000008d000000000000006b00000000000001ac00000000000001ba00000000",
            INIT_64 => X"000001770000000000000188000000000000011b000000000000015c00000000",
            INIT_65 => X"0000012e00000000000000d200000000000000db000000000000011800000000",
            INIT_66 => X"000001c000000000000001eb00000000000001d6000000000000019a00000000",
            INIT_67 => X"00000193000000000000016d000000000000015b00000000000001c300000000",
            INIT_68 => X"00000162000000000000018e0000000000000165000000000000010600000000",
            INIT_69 => X"00000195000000000000011c00000000000000dd00000000000000e800000000",
            INIT_6A => X"00000196000000000000019900000000000001fe00000000000001fe00000000",
            INIT_6B => X"0000012e00000000000001940000000000000190000000000000019400000000",
            INIT_6C => X"000000e400000000000001400000000000000178000000000000017400000000",
            INIT_6D => X"0000020400000000000001790000000000000129000000000000010a00000000",
            INIT_6E => X"0000019a000000000000017e00000000000001b4000000000000021300000000",
            INIT_6F => X"0000015200000000000001640000000000000142000000000000018800000000",
            INIT_70 => X"00000146000000000000011e0000000000000136000000000000015500000000",
            INIT_71 => X"0000021600000000000001fe0000000000000172000000000000014b00000000",
            INIT_72 => X"0000017c000000000000018d00000000000001a9000000000000020200000000",
            INIT_73 => X"0000017100000000000001800000000000000190000000000000010f00000000",
            INIT_74 => X"00000141000000000000014c000000000000011c000000000000015000000000",
            INIT_75 => X"000001f600000000000001f60000000000000171000000000000015a00000000",
            INIT_76 => X"0000015e0000000000000157000000000000018200000000000001d500000000",
            INIT_77 => X"0000017e00000000000001bd00000000000001af000000000000018700000000",
            INIT_78 => X"0000014d000000000000011c000000000000011a000000000000013100000000",
            INIT_79 => X"000001bb000000000000016c000000000000013800000000000000e700000000",
            INIT_7A => X"00000190000000000000019d000000000000017800000000000001ae00000000",
            INIT_7B => X"0000018900000000000001ab00000000000001a700000000000001a100000000",
            INIT_7C => X"000001130000000000000123000000000000013c000000000000012800000000",
            INIT_7D => X"000001c80000000000000137000000000000012a000000000000011400000000",
            INIT_7E => X"000001b000000000000001af00000000000001aa000000000000017b00000000",
            INIT_7F => X"0000017f000000000000018f0000000000000180000000000000016b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE56;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE57 : if BRAM_NAME = "samplegold_layersamples_instance57" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000140000000000000012c00000000000000fe000000000000012700000000",
            INIT_01 => X"0000018100000000000001c000000000000000f9000000000000011300000000",
            INIT_02 => X"0000016100000000000001b200000000000001c800000000000001aa00000000",
            INIT_03 => X"000000f800000000000001700000000000000184000000000000018800000000",
            INIT_04 => X"00000118000000000000014a0000000000000126000000000000011500000000",
            INIT_05 => X"0000019a000000000000017e00000000000001ae00000000000000ef00000000",
            INIT_06 => X"0000017b00000000000000f8000000000000016e00000000000001be00000000",
            INIT_07 => X"0000010e00000000000000e4000000000000013a000000000000016500000000",
            INIT_08 => X"000000fc0000000000000105000000000000010c000000000000010600000000",
            INIT_09 => X"000001c60000000000000175000000000000015e000000000000019800000000",
            INIT_0A => X"000001210000000000000149000000000000013a000000000000018200000000",
            INIT_0B => X"000000ef00000000000000f600000000000000c300000000000000f100000000",
            INIT_0C => X"0000015c000000000000011200000000000000eb00000000000000cd00000000",
            INIT_0D => X"0000019800000000000001b70000000000000138000000000000015300000000",
            INIT_0E => X"000000b700000000000000f000000000000000f8000000000000016200000000",
            INIT_0F => X"000000da00000000000000f000000000000000de00000000000000b900000000",
            INIT_10 => X"00000033000000000000000000000000000000ff00000000000000e800000000",
            INIT_11 => X"00000027000000000000001d000000000000001c000000000000003800000000",
            INIT_12 => X"0000000000000000000000000000000000000021000000000000001a00000000",
            INIT_13 => X"00000029000000000000002c0000000000000033000000000000003e00000000",
            INIT_14 => X"0000005300000000000000070000000000000000000000000000002600000000",
            INIT_15 => X"0000003a000000000000001f000000000000002a000000000000003300000000",
            INIT_16 => X"0000004f00000000000000000000000000000037000000000000003600000000",
            INIT_17 => X"0000003400000000000000360000000000000038000000000000003d00000000",
            INIT_18 => X"0000002b000000000000004b0000000000000000000000000000000000000000",
            INIT_19 => X"000000510000000000000028000000000000000a000000000000006800000000",
            INIT_1A => X"00000058000000000000004d000000000000001e000000000000003f00000000",
            INIT_1B => X"00000000000000000000003b0000000000000048000000000000004a00000000",
            INIT_1C => X"0000007c000000000000001c000000000000002e000000000000000000000000",
            INIT_1D => X"0000001800000000000000000000000000000000000000000000002e00000000",
            INIT_1E => X"0000005f000000000000006b0000000000000055000000000000005300000000",
            INIT_1F => X"0000002100000000000000050000000000000062000000000000005400000000",
            INIT_20 => X"0000005c00000000000000670000000000000000000000000000003900000000",
            INIT_21 => X"0000004700000000000000240000000000000008000000000000003b00000000",
            INIT_22 => X"000000290000000000000063000000000000006f000000000000005e00000000",
            INIT_23 => X"0000003e0000000000000046000000000000003a000000000000005200000000",
            INIT_24 => X"0000003200000000000000550000000000000055000000000000000e00000000",
            INIT_25 => X"00000054000000000000003a000000000000001d000000000000001100000000",
            INIT_26 => X"00000029000000000000001d0000000000000061000000000000008300000000",
            INIT_27 => X"0000003b000000000000002d000000000000003d000000000000003700000000",
            INIT_28 => X"0000003700000000000000280000000000000047000000000000003400000000",
            INIT_29 => X"0000007c0000000000000050000000000000003e000000000000002a00000000",
            INIT_2A => X"0000003200000000000000180000000000000045000000000000006a00000000",
            INIT_2B => X"0000003c00000000000000720000000000000009000000000000004600000000",
            INIT_2C => X"00000047000000000000002c0000000000000039000000000000004300000000",
            INIT_2D => X"00000084000000000000008a0000000000000042000000000000003f00000000",
            INIT_2E => X"00000039000000000000001a000000000000004f000000000000006500000000",
            INIT_2F => X"0000003f000000000000004d0000000000000060000000000000003300000000",
            INIT_30 => X"00000021000000000000004b0000000000000014000000000000003000000000",
            INIT_31 => X"0000006100000000000000760000000000000000000000000000003600000000",
            INIT_32 => X"00000054000000000000002c0000000000000028000000000000007400000000",
            INIT_33 => X"0000006400000000000000760000000000000060000000000000004700000000",
            INIT_34 => X"0000002b000000000000003a0000000000000000000000000000002c00000000",
            INIT_35 => X"0000004900000000000000240000000000000018000000000000002900000000",
            INIT_36 => X"0000004b0000000000000060000000000000002a000000000000004500000000",
            INIT_37 => X"000000630000000000000065000000000000002d000000000000004c00000000",
            INIT_38 => X"0000002e0000000000000024000000000000002a000000000000003f00000000",
            INIT_39 => X"0000004d00000000000000260000000000000021000000000000003700000000",
            INIT_3A => X"0000005900000000000000630000000000000069000000000000002200000000",
            INIT_3B => X"00000042000000000000004b0000000000000047000000000000003e00000000",
            INIT_3C => X"0000004100000000000000310000000000000030000000000000000700000000",
            INIT_3D => X"0000002b0000000000000040000000000000000c000000000000001e00000000",
            INIT_3E => X"00000047000000000000003c0000000000000061000000000000005900000000",
            INIT_3F => X"000000120000000000000037000000000000004b000000000000005d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002d000000000000003e0000000000000028000000000000003400000000",
            INIT_41 => X"00000047000000000000001c0000000000000037000000000000001900000000",
            INIT_42 => X"0000003b0000000000000025000000000000002e000000000000006500000000",
            INIT_43 => X"0000002700000000000000100000000000000023000000000000003500000000",
            INIT_44 => X"000000280000000000000029000000000000000e000000000000001f00000000",
            INIT_45 => X"000000730000000000000032000000000000001b000000000000003400000000",
            INIT_46 => X"0000002a0000000000000023000000000000003b000000000000004500000000",
            INIT_47 => X"0000001f000000000000001c0000000000000014000000000000000700000000",
            INIT_48 => X"00000019000000000000002c000000000000001f000000000000000800000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000010000000000000000200000000",
            INIT_4C => X"0000000f00000000000000190000000000000000000000000000000000000000",
            INIT_4D => X"00000000000000000000000d0000000000000002000000000000000000000000",
            INIT_4E => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000120000000000000018000000000000000000000000",
            INIT_51 => X"000000060000000000000012000000000000000f000000000000000000000000",
            INIT_52 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000018000000000000000400000000",
            INIT_55 => X"000000060000000000000012000000000000001b000000000000000a00000000",
            INIT_56 => X"000000020000000000000000000000000000000a000000000000000b00000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_58 => X"0000000300000000000000010000000000000000000000000000000000000000",
            INIT_59 => X"0000000e000000000000000d000000000000000c000000000000001200000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000e00000000000000000000000000000004000000000000000000000000",
            INIT_5D => X"00000012000000000000000c000000000000001a000000000000000d00000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000c00000000000000180000000000000004000000000000000000000000",
            INIT_61 => X"0000000a000000000000000b0000000000000008000000000000001c00000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_64 => X"00000009000000000000001b0000000000000009000000000000000800000000",
            INIT_65 => X"0000000000000000000000000000000000000006000000000000000a00000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"000000120000000000000000000000000000000c000000000000000000000000",
            INIT_68 => X"00000000000000000000000e0000000000000014000000000000000c00000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000600000000000000010000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000040000000000000019000000000000001500000000",
            INIT_6D => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_6E => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000200000000000000030000000000000002000000000000000300000000",
            INIT_70 => X"000000080000000000000000000000000000000c000000000000000900000000",
            INIT_71 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_72 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"000000040000000000000000000000000000000f000000000000000200000000",
            INIT_74 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_75 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_76 => X"0000000100000000000000050000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_78 => X"0000000000000000000000020000000000000000000000000000000100000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_7A => X"00000006000000000000000c0000000000000002000000000000000000000000",
            INIT_7B => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000020000000000000001000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000008000000000000000400000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE57;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE58 : if BRAM_NAME = "samplegold_layersamples_instance58" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_01 => X"000000540000000000000063000000000000004f000000000000001000000000",
            INIT_02 => X"0000005a000000000000005b000000000000005b000000000000004700000000",
            INIT_03 => X"0000005e0000000000000048000000000000001e000000000000003c00000000",
            INIT_04 => X"0000001100000000000000660000000000000066000000000000006500000000",
            INIT_05 => X"0000002d00000000000000500000000000000068000000000000002f00000000",
            INIT_06 => X"0000004c000000000000004f000000000000004b000000000000003a00000000",
            INIT_07 => X"00000054000000000000004d0000000000000057000000000000001d00000000",
            INIT_08 => X"0000001b0000000000000014000000000000005e000000000000005b00000000",
            INIT_09 => X"00000012000000000000003a000000000000004c000000000000006400000000",
            INIT_0A => X"0000002d000000000000003f0000000000000048000000000000003200000000",
            INIT_0B => X"00000044000000000000003e0000000000000040000000000000004500000000",
            INIT_0C => X"000000560000000000000029000000000000000f000000000000004800000000",
            INIT_0D => X"00000020000000000000001f0000000000000045000000000000004100000000",
            INIT_0E => X"0000003800000000000000460000000000000031000000000000002800000000",
            INIT_0F => X"00000044000000000000003a000000000000003f000000000000004800000000",
            INIT_10 => X"0000002900000000000000400000000000000042000000000000003300000000",
            INIT_11 => X"0000001f000000000000002c0000000000000030000000000000004600000000",
            INIT_12 => X"0000004e00000000000000430000000000000039000000000000002c00000000",
            INIT_13 => X"0000003f000000000000004c0000000000000033000000000000003b00000000",
            INIT_14 => X"000000440000000000000030000000000000003f000000000000004400000000",
            INIT_15 => X"00000028000000000000001f0000000000000026000000000000003300000000",
            INIT_16 => X"0000003a000000000000004e0000000000000037000000000000003000000000",
            INIT_17 => X"0000004100000000000000420000000000000040000000000000002900000000",
            INIT_18 => X"00000027000000000000002d000000000000003e000000000000004200000000",
            INIT_19 => X"0000002d000000000000002f000000000000002e000000000000002300000000",
            INIT_1A => X"0000003400000000000000400000000000000051000000000000003500000000",
            INIT_1B => X"000000330000000000000045000000000000003e000000000000003200000000",
            INIT_1C => X"00000023000000000000002c0000000000000033000000000000006100000000",
            INIT_1D => X"0000003600000000000000400000000000000035000000000000002a00000000",
            INIT_1E => X"00000036000000000000003f0000000000000050000000000000006100000000",
            INIT_1F => X"000000590000000000000040000000000000003e000000000000002d00000000",
            INIT_20 => X"0000001d0000000000000022000000000000002d000000000000002d00000000",
            INIT_21 => X"00000029000000000000003e0000000000000032000000000000005200000000",
            INIT_22 => X"0000003400000000000000520000000000000041000000000000005b00000000",
            INIT_23 => X"0000003c00000000000000350000000000000044000000000000003b00000000",
            INIT_24 => X"000000200000000000000026000000000000002c000000000000003900000000",
            INIT_25 => X"0000003e00000000000000480000000000000044000000000000003e00000000",
            INIT_26 => X"0000002d0000000000000039000000000000004b000000000000004400000000",
            INIT_27 => X"0000002c00000000000000370000000000000039000000000000003f00000000",
            INIT_28 => X"0000004100000000000000300000000000000038000000000000004000000000",
            INIT_29 => X"000000390000000000000042000000000000004a000000000000003c00000000",
            INIT_2A => X"00000048000000000000002b000000000000003d000000000000004100000000",
            INIT_2B => X"0000004500000000000000380000000000000038000000000000003800000000",
            INIT_2C => X"0000004a0000000000000030000000000000003a000000000000003e00000000",
            INIT_2D => X"0000003600000000000000390000000000000042000000000000004000000000",
            INIT_2E => X"000000340000000000000049000000000000003b000000000000003900000000",
            INIT_2F => X"00000044000000000000004b0000000000000041000000000000002a00000000",
            INIT_30 => X"0000003b00000000000000470000000000000033000000000000003d00000000",
            INIT_31 => X"000000380000000000000039000000000000003d000000000000004500000000",
            INIT_32 => X"0000003200000000000000360000000000000047000000000000003700000000",
            INIT_33 => X"0000003d0000000000000042000000000000004d000000000000004000000000",
            INIT_34 => X"0000003500000000000000390000000000000043000000000000003900000000",
            INIT_35 => X"000000360000000000000038000000000000003f000000000000004400000000",
            INIT_36 => X"0000003a000000000000002e000000000000003b000000000000004300000000",
            INIT_37 => X"0000003a00000000000000350000000000000046000000000000003b00000000",
            INIT_38 => X"000000420000000000000036000000000000003e000000000000003f00000000",
            INIT_39 => X"0000001e000000000000004b000000000000001a000000000000004200000000",
            INIT_3A => X"00000008000000000000000d0000000000000010000000000000000000000000",
            INIT_3B => X"0000002700000000000000000000000000000000000000000000000800000000",
            INIT_3C => X"0000000300000000000000060000000000000003000000000000001500000000",
            INIT_3D => X"00000000000000000000003c0000000000000039000000000000001a00000000",
            INIT_3E => X"0000000b000000000000000b000000000000000f000000000000000000000000",
            INIT_3F => X"00000009000000000000003b0000000000000000000000000000000500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001800000000000000010000000000000006000000000000000400000000",
            INIT_41 => X"000000060000000000000005000000000000004c000000000000002600000000",
            INIT_42 => X"0000000800000000000000230000000000000010000000000000000000000000",
            INIT_43 => X"0000000400000000000000140000000000000030000000000000000000000000",
            INIT_44 => X"0000001c00000000000000050000000000000000000000000000000300000000",
            INIT_45 => X"0000000000000000000000120000000000000001000000000000004200000000",
            INIT_46 => X"00000021000000000000000f0000000000000000000000000000000000000000",
            INIT_47 => X"0000000200000000000000000000000000000011000000000000001100000000",
            INIT_48 => X"0000001900000000000000180000000000000000000000000000000d00000000",
            INIT_49 => X"0000000000000000000000000000000000000023000000000000000000000000",
            INIT_4A => X"0000001b0000000000000014000000000000000d000000000000000000000000",
            INIT_4B => X"0000002a00000000000000060000000000000005000000000000001b00000000",
            INIT_4C => X"0000000000000000000000130000000000000014000000000000000a00000000",
            INIT_4D => X"0000000000000000000000000000000000000001000000000000001000000000",
            INIT_4E => X"00000025000000000000001a0000000000000011000000000000000d00000000",
            INIT_4F => X"0000001400000000000000260000000000000005000000000000000d00000000",
            INIT_50 => X"000000080000000000000002000000000000000e000000000000001100000000",
            INIT_51 => X"0000000400000000000000000000000000000000000000000000000600000000",
            INIT_52 => X"0000000e00000000000000270000000000000018000000000000000b00000000",
            INIT_53 => X"0000000f0000000000000015000000000000000a000000000000000300000000",
            INIT_54 => X"0000000100000000000000000000000000000018000000000000000000000000",
            INIT_55 => X"000000120000000000000004000000000000000c000000000000000000000000",
            INIT_56 => X"0000001000000000000000120000000000000030000000000000001100000000",
            INIT_57 => X"000000000000000000000015000000000000000b000000000000000b00000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_59 => X"0000000e00000000000000000000000000000028000000000000000000000000",
            INIT_5A => X"0000002a000000000000001b0000000000000044000000000000000000000000",
            INIT_5B => X"000000000000000000000009000000000000000d000000000000000c00000000",
            INIT_5C => X"000000000000000000000000000000000000000c000000000000001300000000",
            INIT_5D => X"00000008000000000000000a000000000000000c000000000000000000000000",
            INIT_5E => X"000000100000000000000028000000000000000f000000000000000400000000",
            INIT_5F => X"0000000000000000000000050000000000000011000000000000000800000000",
            INIT_60 => X"0000000000000000000000040000000000000017000000000000000000000000",
            INIT_61 => X"00000007000000000000000f0000000000000001000000000000000a00000000",
            INIT_62 => X"000000040000000000000018000000000000000e000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_64 => X"0000000000000000000000040000000000000000000000000000000b00000000",
            INIT_65 => X"0000000000000000000000090000000000000007000000000000001b00000000",
            INIT_66 => X"0000001e00000000000000180000000000000018000000000000000000000000",
            INIT_67 => X"0000000f00000000000000000000000000000000000000000000000300000000",
            INIT_68 => X"0000001900000000000000000000000000000000000000000000000500000000",
            INIT_69 => X"0000000600000000000000030000000000000015000000000000000500000000",
            INIT_6A => X"0000000d0000000000000024000000000000001e000000000000001500000000",
            INIT_6B => X"00000007000000000000000b0000000000000000000000000000000000000000",
            INIT_6C => X"0000000a00000000000000180000000000000004000000000000000500000000",
            INIT_6D => X"00000017000000000000000a0000000000000018000000000000000500000000",
            INIT_6E => X"0000000000000000000000180000000000000022000000000000001f00000000",
            INIT_6F => X"0000000200000000000000090000000000000000000000000000000700000000",
            INIT_70 => X"0000000300000000000000100000000000000011000000000000001600000000",
            INIT_71 => X"0000001a00000000000000080000000000000010000000000000001600000000",
            INIT_72 => X"00000010000000000000001f0000000000000013000000000000001f00000000",
            INIT_73 => X"0000000a00000000000000110000000000000013000000000000000d00000000",
            INIT_74 => X"000000130000000000000014000000000000002d000000000000002800000000",
            INIT_75 => X"0000003400000000000000110000000000000008000000000000001000000000",
            INIT_76 => X"0000003100000000000000360000000000000046000000000000001d00000000",
            INIT_77 => X"0000003f000000000000000a000000000000003b000000000000003300000000",
            INIT_78 => X"00000020000000000000002a0000000000000034000000000000004600000000",
            INIT_79 => X"000000200000000000000032000000000000000b000000000000000500000000",
            INIT_7A => X"0000004400000000000000370000000000000045000000000000006700000000",
            INIT_7B => X"0000006500000000000000640000000000000025000000000000003b00000000",
            INIT_7C => X"0000000000000000000000450000000000000050000000000000005600000000",
            INIT_7D => X"0000006d00000000000000320000000000000043000000000000000500000000",
            INIT_7E => X"0000002e0000000000000028000000000000002a000000000000005300000000",
            INIT_7F => X"0000006d000000000000006b000000000000006b000000000000004800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE58;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE59 : if BRAM_NAME = "samplegold_layersamples_instance59" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003c00000000000000330000000000000069000000000000006f00000000",
            INIT_01 => X"0000006a00000000000000630000000000000025000000000000005900000000",
            INIT_02 => X"0000004600000000000000370000000000000031000000000000005400000000",
            INIT_03 => X"0000005a00000000000000770000000000000078000000000000006500000000",
            INIT_04 => X"0000005b000000000000005a0000000000000054000000000000006100000000",
            INIT_05 => X"0000005300000000000000640000000000000059000000000000002d00000000",
            INIT_06 => X"0000006100000000000000490000000000000042000000000000003000000000",
            INIT_07 => X"00000051000000000000005a000000000000007f000000000000008300000000",
            INIT_08 => X"0000004000000000000000420000000000000050000000000000005400000000",
            INIT_09 => X"0000003a0000000000000052000000000000005b000000000000005600000000",
            INIT_0A => X"0000008100000000000000600000000000000057000000000000005300000000",
            INIT_0B => X"0000005600000000000000500000000000000070000000000000008100000000",
            INIT_0C => X"00000059000000000000004e000000000000001e000000000000004e00000000",
            INIT_0D => X"0000004d000000000000004c0000000000000054000000000000006000000000",
            INIT_0E => X"000000780000000000000069000000000000005b000000000000004d00000000",
            INIT_0F => X"0000004b00000000000000530000000000000068000000000000008100000000",
            INIT_10 => X"0000006300000000000000630000000000000053000000000000003200000000",
            INIT_11 => X"0000002f000000000000003f0000000000000049000000000000005b00000000",
            INIT_12 => X"00000066000000000000005f0000000000000019000000000000004700000000",
            INIT_13 => X"0000005d000000000000004a000000000000005c000000000000006900000000",
            INIT_14 => X"0000006e000000000000007e0000000000000072000000000000005500000000",
            INIT_15 => X"0000003d000000000000003b0000000000000031000000000000005400000000",
            INIT_16 => X"000000490000000000000034000000000000001e000000000000002700000000",
            INIT_17 => X"0000006100000000000000690000000000000059000000000000006900000000",
            INIT_18 => X"0000006700000000000000660000000000000058000000000000005e00000000",
            INIT_19 => X"0000003200000000000000260000000000000041000000000000005500000000",
            INIT_1A => X"0000006c000000000000002d000000000000002f000000000000003c00000000",
            INIT_1B => X"00000069000000000000006e000000000000006d000000000000005800000000",
            INIT_1C => X"0000005400000000000000530000000000000050000000000000004100000000",
            INIT_1D => X"000000430000000000000039000000000000002e000000000000002500000000",
            INIT_1E => X"0000005800000000000000660000000000000023000000000000002f00000000",
            INIT_1F => X"00000028000000000000005f0000000000000074000000000000006400000000",
            INIT_20 => X"000000220000000000000041000000000000004c000000000000005200000000",
            INIT_21 => X"0000003000000000000000410000000000000030000000000000003500000000",
            INIT_22 => X"00000056000000000000004c000000000000005e000000000000002900000000",
            INIT_23 => X"00000042000000000000001f000000000000004f000000000000007700000000",
            INIT_24 => X"0000002f000000000000001a000000000000002b000000000000003700000000",
            INIT_25 => X"0000002f000000000000002a0000000000000023000000000000002a00000000",
            INIT_26 => X"0000007e00000000000000490000000000000048000000000000005300000000",
            INIT_27 => X"00000026000000000000002c0000000000000052000000000000006000000000",
            INIT_28 => X"0000002b0000000000000027000000000000001a000000000000001b00000000",
            INIT_29 => X"0000001400000000000000320000000000000028000000000000001d00000000",
            INIT_2A => X"00000028000000000000003f0000000000000033000000000000001700000000",
            INIT_2B => X"00000037000000000000003c0000000000000041000000000000003c00000000",
            INIT_2C => X"0000004600000000000000310000000000000024000000000000003000000000",
            INIT_2D => X"000000140000000000000015000000000000004c000000000000004800000000",
            INIT_2E => X"000000240000000000000012000000000000003e000000000000002200000000",
            INIT_2F => X"0000003b00000000000000330000000000000030000000000000002800000000",
            INIT_30 => X"0000003e000000000000003a000000000000002e000000000000001400000000",
            INIT_31 => X"0000001600000000000000140000000000000018000000000000004100000000",
            INIT_32 => X"00000021000000000000001b000000000000000a000000000000003a00000000",
            INIT_33 => X"0000001200000000000000280000000000000025000000000000001f00000000",
            INIT_34 => X"0000002c0000000000000026000000000000002a000000000000002900000000",
            INIT_35 => X"0000003600000000000000130000000000000030000000000000003400000000",
            INIT_36 => X"0000002200000000000000220000000000000018000000000000000b00000000",
            INIT_37 => X"0000002000000000000000140000000000000018000000000000001e00000000",
            INIT_38 => X"0000003a000000000000002a0000000000000020000000000000001c00000000",
            INIT_39 => X"000000110000000000000040000000000000002b000000000000002800000000",
            INIT_3A => X"000000170000000000000022000000000000001a000000000000001200000000",
            INIT_3B => X"0000002600000000000000200000000000000019000000000000001600000000",
            INIT_3C => X"0000002f00000000000000340000000000000036000000000000003c00000000",
            INIT_3D => X"000000130000000000000017000000000000003e000000000000002f00000000",
            INIT_3E => X"0000001400000000000000110000000000000027000000000000001b00000000",
            INIT_3F => X"0000003c0000000000000026000000000000001d000000000000001600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000040000000000000003a000000000000003a000000000000004100000000",
            INIT_41 => X"00000017000000000000001c0000000000000022000000000000002a00000000",
            INIT_42 => X"0000001b00000000000000130000000000000012000000000000001a00000000",
            INIT_43 => X"0000003c000000000000002f000000000000002b000000000000001d00000000",
            INIT_44 => X"00000016000000000000003a0000000000000035000000000000003a00000000",
            INIT_45 => X"0000001300000000000000190000000000000012000000000000001e00000000",
            INIT_46 => X"00000029000000000000001d000000000000002b000000000000001d00000000",
            INIT_47 => X"0000003a0000000000000035000000000000002a000000000000002700000000",
            INIT_48 => X"0000001c00000000000000170000000000000029000000000000003500000000",
            INIT_49 => X"00000027000000000000001a0000000000000018000000000000001300000000",
            INIT_4A => X"0000002c000000000000003b0000000000000023000000000000003400000000",
            INIT_4B => X"0000003500000000000000380000000000000031000000000000003200000000",
            INIT_4C => X"00000016000000000000001f0000000000000020000000000000001d00000000",
            INIT_4D => X"000000260000000000000026000000000000001c000000000000001400000000",
            INIT_4E => X"0000002c00000000000000320000000000000031000000000000002b00000000",
            INIT_4F => X"0000002000000000000000320000000000000031000000000000002d00000000",
            INIT_50 => X"0000001a00000000000000280000000000000023000000000000002300000000",
            INIT_51 => X"0000003200000000000000280000000000000021000000000000001e00000000",
            INIT_52 => X"0000002b000000000000002f0000000000000023000000000000002700000000",
            INIT_53 => X"0000001900000000000000210000000000000035000000000000003100000000",
            INIT_54 => X"00000027000000000000001e000000000000002f000000000000001b00000000",
            INIT_55 => X"0000002a00000000000000290000000000000037000000000000002400000000",
            INIT_56 => X"000000330000000000000030000000000000002d000000000000002100000000",
            INIT_57 => X"0000001e000000000000001b000000000000002f000000000000003d00000000",
            INIT_58 => X"0000002e000000000000002e000000000000001c000000000000003800000000",
            INIT_59 => X"00000024000000000000002d0000000000000027000000000000003300000000",
            INIT_5A => X"000000410000000000000037000000000000002c000000000000002c00000000",
            INIT_5B => X"0000002600000000000000230000000000000019000000000000003900000000",
            INIT_5C => X"0000003600000000000000320000000000000032000000000000002700000000",
            INIT_5D => X"00000029000000000000002f000000000000002d000000000000002800000000",
            INIT_5E => X"0000003d000000000000003c0000000000000039000000000000002a00000000",
            INIT_5F => X"0000003200000000000000240000000000000022000000000000001100000000",
            INIT_60 => X"0000002c000000000000002d0000000000000031000000000000002e00000000",
            INIT_61 => X"0000002a00000000000000280000000000000030000000000000002a00000000",
            INIT_62 => X"00000000000000000000003000000000000000b0000000000000000000000000",
            INIT_63 => X"0000000400000000000000000000000000000013000000000000000000000000",
            INIT_64 => X"0000000800000000000000860000000000000000000000000000000000000000",
            INIT_65 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"00000000000000000000001d000000000000006b000000000000006c00000000",
            INIT_67 => X"0000000000000000000000130000000000000019000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000090000000000000000000000000",
            INIT_69 => X"0000002800000000000000020000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000320000000000000017000000000000009b00000000",
            INIT_6B => X"00000014000000000000000c0000000000000038000000000000000900000000",
            INIT_6C => X"000000000000000000000000000000000000001f000000000000003700000000",
            INIT_6D => X"00000047000000000000001f0000000000000000000000000000000000000000",
            INIT_6E => X"000000000000000000000000000000000000005a000000000000000000000000",
            INIT_6F => X"000000090000000000000062000000000000000b000000000000000000000000",
            INIT_70 => X"0000002400000000000000000000000000000000000000000000003f00000000",
            INIT_71 => X"000000000000000000000000000000000000001b000000000000000000000000",
            INIT_72 => X"000000000000000000000000000000000000000c000000000000005900000000",
            INIT_73 => X"0000003a000000000000002c0000000000000048000000000000001600000000",
            INIT_74 => X"00000000000000000000002b0000000000000000000000000000000000000000",
            INIT_75 => X"0000002b00000000000000000000000000000000000000000000000900000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_77 => X"000000000000000000000052000000000000002c000000000000003200000000",
            INIT_78 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000001600000000000000000000000000000015000000000000000000000000",
            INIT_7A => X"0000001e00000000000000000000000000000025000000000000000000000000",
            INIT_7B => X"000000000000000000000006000000000000004b000000000000002300000000",
            INIT_7C => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000010000000000000000000000000000006400000000",
            INIT_7E => X"0000000100000000000000100000000000000025000000000000000000000000",
            INIT_7F => X"0000000c0000000000000000000000000000004d000000000000005e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE59;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE60 : if BRAM_NAME = "samplegold_layersamples_instance60" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002d00000000000000000000000000000015000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000004a00000000",
            INIT_03 => X"000000000000000000000060000000000000001b000000000000007100000000",
            INIT_04 => X"0000001700000000000000000000000000000008000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000009000000000000001400000000",
            INIT_06 => X"00000009000000000000000a0000000000000000000000000000001900000000",
            INIT_07 => X"0000000000000000000000000000000000000039000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000002d00000000",
            INIT_09 => X"0000000000000000000000000000000000000016000000000000003700000000",
            INIT_0A => X"000000000000000000000009000000000000000f000000000000000e00000000",
            INIT_0B => X"0000004600000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000001100000000000000000000000000000000000000000000000300000000",
            INIT_0D => X"0000003200000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000011000000000000000100000000",
            INIT_0F => X"00000003000000000000003a0000000000000000000000000000000000000000",
            INIT_10 => X"0000000400000000000000240000000000000025000000000000000000000000",
            INIT_11 => X"0000000200000000000000290000000000000000000000000000000000000000",
            INIT_12 => X"000000000000000000000000000000000000000c000000000000000b00000000",
            INIT_13 => X"0000000000000000000000150000000000000041000000000000000000000000",
            INIT_14 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_15 => X"000000000000000000000005000000000000001a000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000008000000000000002c00000000",
            INIT_17 => X"0000000000000000000000000000000000000039000000000000002c00000000",
            INIT_18 => X"000000250000000000000000000000000000000d000000000000000000000000",
            INIT_19 => X"0000001100000000000000000000000000000008000000000000000e00000000",
            INIT_1A => X"0000000000000000000000260000000000000000000000000000001300000000",
            INIT_1B => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_1C => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"00000015000000000000001e000000000000001c000000000000000100000000",
            INIT_1F => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000010000000000000000c00000000",
            INIT_23 => X"000000450000000000000040000000000000001c000000000000000000000000",
            INIT_24 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"00000000000000000000001d0000000000000001000000000000000000000000",
            INIT_27 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_2C => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000020000000000000003000000000000000000000000",
            INIT_2F => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_36 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_37 => X"000000040000000000000038000000000000006f000000000000000700000000",
            INIT_38 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000010000000000000013000000000000000000000000",
            INIT_3B => X"0000002f00000000000000530000000000000051000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000080000000000000021000000000000000400000000",
            INIT_3E => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000270000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"00000000000000000000000c000000000000000d000000000000000000000000",
            INIT_42 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_44 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_47 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"00000003000000000000002d0000000000000000000000000000000000000000",
            INIT_49 => X"0000000600000000000000070000000000000011000000000000000e00000000",
            INIT_4A => X"000000000000000000000019000000000000001d000000000000000900000000",
            INIT_4B => X"00000000000000000000001d0000000000000000000000000000000000000000",
            INIT_4C => X"0000001400000000000000040000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000017000000000000001400000000",
            INIT_4E => X"0000002100000000000000000000000000000006000000000000000000000000",
            INIT_4F => X"00000000000000000000000e0000000000000020000000000000000000000000",
            INIT_50 => X"0000000e0000000000000019000000000000001e000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000007000000000000000200000000",
            INIT_52 => X"0000006c0000000000000000000000000000000f000000000000000000000000",
            INIT_53 => X"000000980000000000000089000000000000008300000000000000a100000000",
            INIT_54 => X"000000460000000000000081000000000000009e000000000000009c00000000",
            INIT_55 => X"000000b500000000000000b500000000000000b7000000000000007c00000000",
            INIT_56 => X"00000092000000000000003e000000000000000000000000000000af00000000",
            INIT_57 => X"000000890000000000000088000000000000007c000000000000007500000000",
            INIT_58 => X"000000bd0000000000000035000000000000008c000000000000009c00000000",
            INIT_59 => X"000000ae00000000000000b200000000000000af00000000000000b100000000",
            INIT_5A => X"00000089000000000000008d0000000000000016000000000000000400000000",
            INIT_5B => X"0000006400000000000000510000000000000056000000000000008100000000",
            INIT_5C => X"0000009c00000000000000b0000000000000005f000000000000005100000000",
            INIT_5D => X"0000005100000000000000b100000000000000b000000000000000a500000000",
            INIT_5E => X"00000079000000000000007b00000000000000d3000000000000006800000000",
            INIT_5F => X"00000057000000000000005a0000000000000077000000000000006b00000000",
            INIT_60 => X"000000b100000000000000b20000000000000086000000000000008a00000000",
            INIT_61 => X"000000b9000000000000008b000000000000009b000000000000009600000000",
            INIT_62 => X"000000780000000000000086000000000000005d000000000000009d00000000",
            INIT_63 => X"0000007300000000000000530000000000000044000000000000007000000000",
            INIT_64 => X"0000008900000000000000ad00000000000000c2000000000000009100000000",
            INIT_65 => X"00000093000000000000009c000000000000009800000000000000a300000000",
            INIT_66 => X"000000570000000000000078000000000000008d000000000000007800000000",
            INIT_67 => X"0000008a00000000000000780000000000000066000000000000004300000000",
            INIT_68 => X"000000a1000000000000009800000000000000b300000000000000bc00000000",
            INIT_69 => X"00000083000000000000007c0000000000000097000000000000009f00000000",
            INIT_6A => X"0000006a000000000000005f0000000000000069000000000000006e00000000",
            INIT_6B => X"000000c000000000000000880000000000000072000000000000007000000000",
            INIT_6C => X"0000009800000000000000ac00000000000000b000000000000000b500000000",
            INIT_6D => X"0000008700000000000000a3000000000000006a000000000000009300000000",
            INIT_6E => X"000000650000000000000074000000000000005a000000000000007700000000",
            INIT_6F => X"000000a2000000000000008e0000000000000076000000000000008100000000",
            INIT_70 => X"00000084000000000000008900000000000000a400000000000000a300000000",
            INIT_71 => X"00000099000000000000008500000000000000ac000000000000008200000000",
            INIT_72 => X"0000006b00000000000000880000000000000053000000000000008300000000",
            INIT_73 => X"000000680000000000000081000000000000006b000000000000007d00000000",
            INIT_74 => X"00000098000000000000009d000000000000009900000000000000aa00000000",
            INIT_75 => X"00000075000000000000007b000000000000008b000000000000008900000000",
            INIT_76 => X"0000006d00000000000000870000000000000087000000000000007a00000000",
            INIT_77 => X"0000008500000000000000850000000000000086000000000000007500000000",
            INIT_78 => X"0000009c000000000000008f000000000000008800000000000000a100000000",
            INIT_79 => X"0000007f00000000000000810000000000000072000000000000009b00000000",
            INIT_7A => X"0000008b00000000000000610000000000000073000000000000007500000000",
            INIT_7B => X"000000a100000000000000700000000000000067000000000000008400000000",
            INIT_7C => X"000000910000000000000095000000000000009f000000000000007e00000000",
            INIT_7D => X"00000082000000000000008c000000000000009b000000000000007500000000",
            INIT_7E => X"0000007e00000000000000750000000000000089000000000000005400000000",
            INIT_7F => X"0000008a000000000000009c0000000000000060000000000000007300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE60;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE61 : if BRAM_NAME = "samplegold_layersamples_instance61" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005f0000000000000066000000000000008a000000000000009b00000000",
            INIT_01 => X"0000005800000000000000690000000000000082000000000000008c00000000",
            INIT_02 => X"0000005d00000000000000660000000000000068000000000000007800000000",
            INIT_03 => X"0000009600000000000000870000000000000094000000000000006a00000000",
            INIT_04 => X"0000007f00000000000000a0000000000000007a000000000000009000000000",
            INIT_05 => X"0000006f0000000000000051000000000000005d000000000000006e00000000",
            INIT_06 => X"00000075000000000000006e0000000000000053000000000000006500000000",
            INIT_07 => X"0000008800000000000000880000000000000082000000000000007900000000",
            INIT_08 => X"00000064000000000000005c0000000000000080000000000000008200000000",
            INIT_09 => X"0000006900000000000000630000000000000061000000000000004900000000",
            INIT_0A => X"0000000000000000000000670000000000000075000000000000005f00000000",
            INIT_0B => X"00000014000000000000002d0000000000000000000000000000000000000000",
            INIT_0C => X"0000003900000000000000100000000000000020000000000000000f00000000",
            INIT_0D => X"00000025000000000000000d0000000000000000000000000000004900000000",
            INIT_0E => X"000000000000000000000000000000000000002d000000000000002500000000",
            INIT_0F => X"00000023000000000000001c000000000000001a000000000000000000000000",
            INIT_10 => X"000000860000000000000037000000000000001b000000000000001900000000",
            INIT_11 => X"00000029000000000000002e0000000000000029000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000003000000000",
            INIT_13 => X"0000002500000000000000780000000000000003000000000000000700000000",
            INIT_14 => X"0000000000000000000000180000000000000036000000000000000400000000",
            INIT_15 => X"0000002f0000000000000026000000000000002f000000000000001b00000000",
            INIT_16 => X"0000004a00000000000000000000000000000000000000000000002600000000",
            INIT_17 => X"00000035000000000000003e0000000000000057000000000000000000000000",
            INIT_18 => X"00000000000000000000002a0000000000000000000000000000000700000000",
            INIT_19 => X"000000490000000000000027000000000000005b000000000000004100000000",
            INIT_1A => X"00000000000000000000006f0000000000000027000000000000000000000000",
            INIT_1B => X"0000000a0000000000000066000000000000004f000000000000002f00000000",
            INIT_1C => X"000000430000000000000001000000000000000a000000000000000000000000",
            INIT_1D => X"000000260000000000000038000000000000000d000000000000006e00000000",
            INIT_1E => X"000000380000000000000004000000000000004b000000000000003c00000000",
            INIT_1F => X"000000000000000000000009000000000000003c000000000000005c00000000",
            INIT_20 => X"0000006800000000000000420000000000000000000000000000000c00000000",
            INIT_21 => X"00000059000000000000002e0000000000000037000000000000002500000000",
            INIT_22 => X"000000480000000000000012000000000000002c000000000000001a00000000",
            INIT_23 => X"0000000900000000000000120000000000000036000000000000001300000000",
            INIT_24 => X"00000046000000000000004f000000000000003b000000000000000000000000",
            INIT_25 => X"000000000000000000000073000000000000002b000000000000004200000000",
            INIT_26 => X"0000002d00000000000000420000000000000036000000000000004500000000",
            INIT_27 => X"000000120000000000000039000000000000001f000000000000002200000000",
            INIT_28 => X"0000005b00000000000000350000000000000054000000000000002200000000",
            INIT_29 => X"0000003c00000000000000000000000000000035000000000000001b00000000",
            INIT_2A => X"000000000000000000000065000000000000003c000000000000003100000000",
            INIT_2B => X"0000000000000000000000410000000000000026000000000000004200000000",
            INIT_2C => X"00000026000000000000004a0000000000000000000000000000003d00000000",
            INIT_2D => X"000000360000000000000025000000000000003b000000000000002300000000",
            INIT_2E => X"00000004000000000000003c000000000000004e000000000000004300000000",
            INIT_2F => X"000000280000000000000010000000000000001d000000000000004a00000000",
            INIT_30 => X"00000010000000000000004e000000000000003a000000000000000b00000000",
            INIT_31 => X"0000000a00000000000000630000000000000031000000000000003000000000",
            INIT_32 => X"0000002300000000000000510000000000000056000000000000002f00000000",
            INIT_33 => X"000000220000000000000040000000000000001e000000000000000a00000000",
            INIT_34 => X"000000380000000000000000000000000000005e000000000000003400000000",
            INIT_35 => X"0000003400000000000000180000000000000060000000000000004800000000",
            INIT_36 => X"0000002b00000000000000000000000000000069000000000000004300000000",
            INIT_37 => X"0000003b0000000000000038000000000000003b000000000000001c00000000",
            INIT_38 => X"0000006d00000000000000370000000000000007000000000000004800000000",
            INIT_39 => X"00000051000000000000003c0000000000000012000000000000002b00000000",
            INIT_3A => X"00000026000000000000002b0000000000000002000000000000004700000000",
            INIT_3B => X"0000004500000000000000450000000000000028000000000000002c00000000",
            INIT_3C => X"0000001e000000000000005e0000000000000023000000000000000000000000",
            INIT_3D => X"0000002e000000000000003d0000000000000035000000000000003e00000000",
            INIT_3E => X"000000000000000000000035000000000000001f000000000000000800000000",
            INIT_3F => X"0000000a00000000000000330000000000000042000000000000001800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005500000000000000460000000000000049000000000000000e00000000",
            INIT_41 => X"0000001600000000000000000000000000000042000000000000002700000000",
            INIT_42 => X"0000001c00000000000000080000000000000028000000000000001600000000",
            INIT_43 => X"0000006d00000000000000520000000000000000000000000000000400000000",
            INIT_44 => X"0000005f000000000000006f000000000000005f000000000000006600000000",
            INIT_45 => X"0000006700000000000000000000000000000073000000000000008800000000",
            INIT_46 => X"000000010000000000000081000000000000007a000000000000007d00000000",
            INIT_47 => X"0000006c000000000000004d0000000000000020000000000000000000000000",
            INIT_48 => X"0000008500000000000000680000000000000064000000000000006b00000000",
            INIT_49 => X"00000091000000000000008f000000000000000000000000000000be00000000",
            INIT_4A => X"000000000000000000000004000000000000008d000000000000008a00000000",
            INIT_4B => X"000000c600000000000000530000000000000044000000000000000000000000",
            INIT_4C => X"00000059000000000000007a0000000000000049000000000000005d00000000",
            INIT_4D => X"000000900000000000000097000000000000007f000000000000003100000000",
            INIT_4E => X"0000000000000000000000000000000000000050000000000000009600000000",
            INIT_4F => X"0000008400000000000000b3000000000000003c000000000000008a00000000",
            INIT_50 => X"00000087000000000000000a0000000000000040000000000000006e00000000",
            INIT_51 => X"0000008800000000000000bc00000000000000a6000000000000005f00000000",
            INIT_52 => X"000000b40000000000000086000000000000004000000000000000a300000000",
            INIT_53 => X"000000a000000000000000a40000000000000086000000000000001b00000000",
            INIT_54 => X"0000006900000000000000620000000000000026000000000000004400000000",
            INIT_55 => X"00000098000000000000006800000000000000d500000000000000b800000000",
            INIT_56 => X"0000004a0000000000000099000000000000009d000000000000007c00000000",
            INIT_57 => X"0000004d000000000000007700000000000000a9000000000000008400000000",
            INIT_58 => X"000000b90000000000000061000000000000005c000000000000003100000000",
            INIT_59 => X"000000860000000000000099000000000000008500000000000000de00000000",
            INIT_5A => X"000000650000000000000077000000000000007300000000000000a500000000",
            INIT_5B => X"00000056000000000000007c000000000000004b000000000000009a00000000",
            INIT_5C => X"000000c900000000000000ad0000000000000061000000000000005a00000000",
            INIT_5D => X"000000c3000000000000008000000000000000a400000000000000a900000000",
            INIT_5E => X"0000009100000000000000800000000000000098000000000000002100000000",
            INIT_5F => X"00000084000000000000005a000000000000006d000000000000006e00000000",
            INIT_60 => X"000000a100000000000000c50000000000000085000000000000005700000000",
            INIT_61 => X"000000390000000000000093000000000000006d00000000000000c200000000",
            INIT_62 => X"000000ba000000000000008e000000000000008e000000000000009b00000000",
            INIT_63 => X"00000080000000000000007e0000000000000082000000000000002100000000",
            INIT_64 => X"000000b700000000000000580000000000000099000000000000001a00000000",
            INIT_65 => X"0000007b0000000000000092000000000000007d000000000000007900000000",
            INIT_66 => X"0000008c00000000000000a3000000000000009e000000000000009100000000",
            INIT_67 => X"000000510000000000000066000000000000008d000000000000005700000000",
            INIT_68 => X"000000a900000000000000a5000000000000004c000000000000007100000000",
            INIT_69 => X"000000b40000000000000091000000000000008d000000000000006d00000000",
            INIT_6A => X"0000009600000000000000b40000000000000082000000000000005c00000000",
            INIT_6B => X"0000008700000000000000670000000000000050000000000000006500000000",
            INIT_6C => X"0000004b00000000000000c3000000000000009b000000000000006300000000",
            INIT_6D => X"0000006a00000000000000ab00000000000000a7000000000000009a00000000",
            INIT_6E => X"0000002f00000000000000ad0000000000000097000000000000008500000000",
            INIT_6F => X"000000750000000000000082000000000000006a000000000000006d00000000",
            INIT_70 => X"00000098000000000000005700000000000000ab00000000000000a200000000",
            INIT_71 => X"0000008a000000000000006b000000000000005d00000000000000cd00000000",
            INIT_72 => X"0000006a00000000000000430000000000000086000000000000009d00000000",
            INIT_73 => X"000000a60000000000000069000000000000006d000000000000006400000000",
            INIT_74 => X"000000c10000000000000087000000000000004a00000000000000a400000000",
            INIT_75 => X"00000080000000000000007d0000000000000084000000000000006a00000000",
            INIT_76 => X"0000006e000000000000005d0000000000000045000000000000005f00000000",
            INIT_77 => X"000000930000000000000098000000000000005f000000000000003400000000",
            INIT_78 => X"0000009d00000000000000a7000000000000006a000000000000004a00000000",
            INIT_79 => X"00000030000000000000007a0000000000000062000000000000009600000000",
            INIT_7A => X"0000004200000000000000620000000000000055000000000000004d00000000",
            INIT_7B => X"0000000f00000000000000000000000000000000000000000000005700000000",
            INIT_7C => X"0000000f0000000000000014000000000000000e000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_7E => X"0000000c000000000000000a0000000000000009000000000000000000000000",
            INIT_7F => X"00000000000000000000000b0000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE61;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE62 : if BRAM_NAME = "samplegold_layersamples_instance62" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"00000000000000000000000a0000000000000007000000000000000200000000",
            INIT_03 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000d000000000000000d0000000000000000000000000000000000000000",
            INIT_34 => X"00000006000000000000000c000000000000000a000000000000000500000000",
            INIT_35 => X"0000001100000000000000000000000000000000000000000000000500000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"000000110000000000000018000000000000000c000000000000000500000000",
            INIT_38 => X"0000000300000000000000000000000000000000000000000000000400000000",
            INIT_39 => X"00000000000000000000000c0000000000000002000000000000000000000000",
            INIT_3A => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000016000000000000000d00000000",
            INIT_3C => X"0000002e00000000000000260000000000000003000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000003400000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"00000000000000000000000d0000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"000000000000000000000000000000000000001d000000000000000000000000",
            INIT_4F => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_50 => X"000000000000000000000032000000000000000d000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000b00000000000000070000000000000000000000000000000000000000",
            INIT_54 => X"0000002900000000000000280000000000000009000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_57 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000002000000000000000000000000000000000000000000000000600000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_5B => X"000000000000000000000009000000000000001d000000000000000000000000",
            INIT_5C => X"00000000000000000000000e000000000000000f000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000200000000000000000000000000000000000000000000000800000000",
            INIT_5F => X"0000000000000000000000080000000000000000000000000000001800000000",
            INIT_60 => X"0000000000000000000000000000000000000007000000000000000600000000",
            INIT_61 => X"00000032000000000000001c0000000000000000000000000000000000000000",
            INIT_62 => X"00000019000000000000001c000000000000000f000000000000000300000000",
            INIT_63 => X"000000140000000000000021000000000000000d000000000000000400000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_65 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"00000005000000000000001a0000000000000022000000000000001b00000000",
            INIT_67 => X"0000000000000000000000070000000000000014000000000000000a00000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_69 => X"0000001d000000000000002a0000000000000006000000000000000000000000",
            INIT_6A => X"00000004000000000000000d0000000000000004000000000000002500000000",
            INIT_6B => X"0000000000000000000000110000000000000001000000000000000100000000",
            INIT_6C => X"0000000300000000000000000000000000000002000000000000001000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000017000000000000001100000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000200000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE62;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE63 : if BRAM_NAME = "samplegold_layersamples_instance63" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000002900000000000000040000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000002000000000000000700000000",
            INIT_0E => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000002900000000000000090000000000000003000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_2C => X"0000002000000000000000300000000000000000000000000000000000000000",
            INIT_2D => X"0000001200000000000000030000000000000000000000000000000f00000000",
            INIT_2E => X"000000000000000000000000000000000000000b000000000000004000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_30 => X"000000000000000000000000000000000000006a000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000002e00000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000003d00000000",
            INIT_35 => X"0000003e00000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"00000006000000000000001d0000000000000000000000000000000a00000000",
            INIT_37 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000005000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_3D => X"00000000000000000000000c0000000000000012000000000000000000000000",
            INIT_3E => X"0000003800000000000000000000000000000000000000000000000700000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000006d000000000000000f0000000000000009000000000000000000000000",
            INIT_42 => X"0000000000000000000000450000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000002f00000000",
            INIT_44 => X"000000410000000000000003000000000000004f000000000000005a00000000",
            INIT_45 => X"0000000000000000000000400000000000000000000000000000006700000000",
            INIT_46 => X"000000010000000000000000000000000000000e000000000000000000000000",
            INIT_47 => X"00000000000000000000001d0000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000071000000000000000000000000",
            INIT_4A => X"0000000300000000000000000000000000000000000000000000000c00000000",
            INIT_4B => X"00000000000000000000002f0000000000000000000000000000003100000000",
            INIT_4C => X"0000003b00000000000000000000000000000047000000000000000200000000",
            INIT_4D => X"0000002200000000000000000000000000000000000000000000003100000000",
            INIT_4E => X"0000000100000000000000000000000000000000000000000000002800000000",
            INIT_4F => X"0000000300000000000000000000000000000052000000000000000000000000",
            INIT_50 => X"0000006600000000000000000000000000000000000000000000000800000000",
            INIT_51 => X"0000000500000000000000200000000000000000000000000000000000000000",
            INIT_52 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"00000000000000000000000000000000000000bc000000000000001200000000",
            INIT_54 => X"00000005000000000000007b000000000000001e000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000002100000000000000150000000000000005000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_58 => X"0000000000000000000000000000000000000057000000000000003d00000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000d000000000000000b000000000000000b000000000000000000000000",
            INIT_5B => X"0000003000000000000000000000000000000000000000000000000800000000",
            INIT_5C => X"000001e000000000000001e900000000000001ef000000000000009600000000",
            INIT_5D => X"0000019e000000000000017e0000000000000172000000000000017000000000",
            INIT_5E => X"000001e90000000000000201000000000000020200000000000001cc00000000",
            INIT_5F => X"0000019c00000000000001c700000000000001d400000000000001f700000000",
            INIT_60 => X"0000012100000000000002020000000000000223000000000000022300000000",
            INIT_61 => X"00000147000000000000012b000000000000012e000000000000011c00000000",
            INIT_62 => X"000001f100000000000001be00000000000001ac000000000000017e00000000",
            INIT_63 => X"0000022900000000000001d300000000000001b900000000000001f600000000",
            INIT_64 => X"000000f500000000000000e300000000000001f3000000000000022800000000",
            INIT_65 => X"0000010900000000000001100000000000000118000000000000012000000000",
            INIT_66 => X"000001d10000000000000201000000000000019e000000000000011c00000000",
            INIT_67 => X"00000219000000000000022700000000000001aa000000000000018100000000",
            INIT_68 => X"00000194000000000000014200000000000000f800000000000001d400000000",
            INIT_69 => X"00000155000000000000014b0000000000000149000000000000015a00000000",
            INIT_6A => X"0000019b00000000000001db00000000000001cf000000000000016b00000000",
            INIT_6B => X"0000017200000000000002110000000000000224000000000000016200000000",
            INIT_6C => X"0000011c000000000000012c000000000000012300000000000000ca00000000",
            INIT_6D => X"00000168000000000000014b0000000000000144000000000000012a00000000",
            INIT_6E => X"000001c700000000000001f3000000000000020e00000000000001bd00000000",
            INIT_6F => X"000000a9000000000000015700000000000001e8000000000000020200000000",
            INIT_70 => X"000000dc00000000000000e300000000000000f000000000000000ba00000000",
            INIT_71 => X"00000160000000000000011a000000000000010100000000000000e300000000",
            INIT_72 => X"000001c0000000000000022a000000000000022a000000000000020600000000",
            INIT_73 => X"000000d600000000000000da000000000000012c000000000000017300000000",
            INIT_74 => X"000000d100000000000000b800000000000000dd00000000000000eb00000000",
            INIT_75 => X"00000183000000000000010200000000000000c400000000000000f300000000",
            INIT_76 => X"000000d00000000000000185000000000000022700000000000001c100000000",
            INIT_77 => X"000000a500000000000000b20000000000000106000000000000012500000000",
            INIT_78 => X"00000052000000000000004a0000000000000064000000000000008f00000000",
            INIT_79 => X"0000010d00000000000000b4000000000000004c000000000000004400000000",
            INIT_7A => X"0000012100000000000000b80000000000000183000000000000020600000000",
            INIT_7B => X"000000e500000000000000cb00000000000000ba000000000000007500000000",
            INIT_7C => X"000000fc00000000000000f900000000000000d800000000000000c800000000",
            INIT_7D => X"000001c80000000000000111000000000000010d00000000000000d500000000",
            INIT_7E => X"0000003100000000000000cb000000000000009700000000000001a200000000",
            INIT_7F => X"000000c50000000000000080000000000000006c000000000000008100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE63;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE64 : if BRAM_NAME = "samplegold_layersamples_instance64" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000f200000000000000f400000000000000fb000000000000010f00000000",
            INIT_01 => X"000001ac000000000000016300000000000000a7000000000000011400000000",
            INIT_02 => X"000000220000000000000056000000000000008d00000000000000a800000000",
            INIT_03 => X"000000c1000000000000005f00000000000000b3000000000000005500000000",
            INIT_04 => X"0000008f00000000000000fb00000000000000aa00000000000000b300000000",
            INIT_05 => X"0000006e0000000000000196000000000000014500000000000000d600000000",
            INIT_06 => X"00000014000000000000003500000000000000c3000000000000009500000000",
            INIT_07 => X"000000d1000000000000008d0000000000000023000000000000005800000000",
            INIT_08 => X"000000840000000000000044000000000000010900000000000000f400000000",
            INIT_09 => X"000000c400000000000000f70000000000000177000000000000010b00000000",
            INIT_0A => X"00000000000000000000000d000000000000006d00000000000000f300000000",
            INIT_0B => X"0000017500000000000001480000000000000036000000000000000a00000000",
            INIT_0C => X"00000114000000000000004e000000000000001b00000000000000f600000000",
            INIT_0D => X"000000d400000000000000e80000000000000157000000000000017500000000",
            INIT_0E => X"000000200000000000000008000000000000002a000000000000009100000000",
            INIT_0F => X"000000cc000000000000011b00000000000000e9000000000000005800000000",
            INIT_10 => X"000001570000000000000116000000000000005b000000000000000000000000",
            INIT_11 => X"0000007c00000000000000880000000000000103000000000000013f00000000",
            INIT_12 => X"0000004f000000000000003c000000000000002f000000000000004400000000",
            INIT_13 => X"0000000e00000000000000a500000000000000b1000000000000007800000000",
            INIT_14 => X"0000005300000000000000570000000000000137000000000000005600000000",
            INIT_15 => X"000000440000000000000046000000000000003a000000000000005b00000000",
            INIT_16 => X"00000067000000000000005e000000000000003c000000000000003a00000000",
            INIT_17 => X"000000440000000000000038000000000000006d000000000000005f00000000",
            INIT_18 => X"0000006c00000000000000750000000000000076000000000000002500000000",
            INIT_19 => X"0000007a0000000000000075000000000000005f000000000000002900000000",
            INIT_1A => X"000000620000000000000084000000000000009d000000000000008d00000000",
            INIT_1B => X"0000006000000000000000450000000000000070000000000000007700000000",
            INIT_1C => X"0000000000000000000000680000000000000085000000000000008300000000",
            INIT_1D => X"0000002800000000000000380000000000000042000000000000004a00000000",
            INIT_1E => X"00000073000000000000007c0000000000000058000000000000004000000000",
            INIT_1F => X"0000008200000000000000690000000000000037000000000000006000000000",
            INIT_20 => X"000000820000000000000009000000000000006c000000000000007d00000000",
            INIT_21 => X"00000060000000000000006f0000000000000050000000000000007a00000000",
            INIT_22 => X"0000005900000000000000980000000000000056000000000000005e00000000",
            INIT_23 => X"0000007600000000000000850000000000000035000000000000002d00000000",
            INIT_24 => X"0000007800000000000000740000000000000026000000000000005e00000000",
            INIT_25 => X"000000720000000000000074000000000000006d000000000000006300000000",
            INIT_26 => X"0000004000000000000000790000000000000089000000000000005d00000000",
            INIT_27 => X"0000003000000000000000730000000000000095000000000000002d00000000",
            INIT_28 => X"000000510000000000000052000000000000005f000000000000000500000000",
            INIT_29 => X"0000007e000000000000006b000000000000005f000000000000005e00000000",
            INIT_2A => X"00000084000000000000008300000000000000a7000000000000007d00000000",
            INIT_2B => X"000000110000000000000059000000000000005a000000000000008200000000",
            INIT_2C => X"0000003600000000000000480000000000000054000000000000002800000000",
            INIT_2D => X"00000061000000000000002c0000000000000055000000000000004e00000000",
            INIT_2E => X"00000064000000000000009200000000000000aa000000000000009f00000000",
            INIT_2F => X"00000048000000000000001a000000000000005d000000000000002900000000",
            INIT_30 => X"000000380000000000000027000000000000002e000000000000002400000000",
            INIT_31 => X"000000660000000000000042000000000000002a000000000000003200000000",
            INIT_32 => X"00000000000000000000004700000000000000c0000000000000007500000000",
            INIT_33 => X"0000004200000000000000400000000000000017000000000000005900000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_35 => X"0000004500000000000000180000000000000000000000000000000000000000",
            INIT_36 => X"000000500000000000000000000000000000005200000000000000b400000000",
            INIT_37 => X"000000380000000000000011000000000000003e000000000000000000000000",
            INIT_38 => X"00000060000000000000006c0000000000000051000000000000006c00000000",
            INIT_39 => X"000000a2000000000000002b0000000000000070000000000000006000000000",
            INIT_3A => X"0000000000000000000000090000000000000000000000000000006800000000",
            INIT_3B => X"000000000000000000000016000000000000001c000000000000000000000000",
            INIT_3C => X"000000360000000000000028000000000000001f000000000000005300000000",
            INIT_3D => X"0000006d000000000000007c0000000000000030000000000000001d00000000",
            INIT_3E => X"0000000000000000000000070000000000000033000000000000000000000000",
            INIT_3F => X"0000005d00000000000000000000000000000051000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000660000000000000030000000000000003300000000",
            INIT_41 => X"0000000000000000000000700000000000000084000000000000004800000000",
            INIT_42 => X"000000000000000000000000000000000000003c000000000000000800000000",
            INIT_43 => X"0000005d00000000000000010000000000000000000000000000000000000000",
            INIT_44 => X"0000000400000000000000000000000000000000000000000000002b00000000",
            INIT_45 => X"000000250000000000000060000000000000006b000000000000007300000000",
            INIT_46 => X"000000000000000000000000000000000000001a000000000000003000000000",
            INIT_47 => X"00000077000000000000006e0000000000000007000000000000000000000000",
            INIT_48 => X"00000075000000000000001b0000000000000000000000000000001500000000",
            INIT_49 => X"00000012000000000000002a0000000000000053000000000000006800000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_4B => X"0000001f000000000000004c0000000000000020000000000000000000000000",
            INIT_4C => X"0000000d000000000000007a0000000000000011000000000000000000000000",
            INIT_4D => X"00000015000000000000000e000000000000000b000000000000000900000000",
            INIT_4E => X"0000000100000000000000090000000000000013000000000000001900000000",
            INIT_4F => X"0000000d00000000000000080000000000000000000000000000000600000000",
            INIT_50 => X"0000001100000000000000120000000000000005000000000000000000000000",
            INIT_51 => X"00000034000000000000002a0000000000000027000000000000000d00000000",
            INIT_52 => X"0000000d0000000000000021000000000000002f000000000000003a00000000",
            INIT_53 => X"0000000000000000000000040000000000000003000000000000000500000000",
            INIT_54 => X"0000001900000000000000140000000000000014000000000000000000000000",
            INIT_55 => X"0000006000000000000000580000000000000058000000000000003b00000000",
            INIT_56 => X"0000001d000000000000003c0000000000000055000000000000005c00000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_58 => X"0000003f00000000000000230000000000000010000000000000001400000000",
            INIT_59 => X"00000066000000000000004e000000000000004b000000000000004800000000",
            INIT_5A => X"0000001200000000000000260000000000000061000000000000006400000000",
            INIT_5B => X"0000001400000000000000000000000000000000000000000000001300000000",
            INIT_5C => X"00000049000000000000005b0000000000000024000000000000001300000000",
            INIT_5D => X"0000005c00000000000000620000000000000065000000000000005400000000",
            INIT_5E => X"0000001200000000000000270000000000000054000000000000005f00000000",
            INIT_5F => X"0000001200000000000000150000000000000014000000000000001500000000",
            INIT_60 => X"0000005e000000000000004c0000000000000043000000000000003d00000000",
            INIT_61 => X"00000055000000000000005a000000000000005a000000000000005d00000000",
            INIT_62 => X"0000001400000000000000190000000000000038000000000000004c00000000",
            INIT_63 => X"00000023000000000000001d0000000000000015000000000000001400000000",
            INIT_64 => X"00000061000000000000005c000000000000004e000000000000005000000000",
            INIT_65 => X"0000004400000000000000490000000000000059000000000000005d00000000",
            INIT_66 => X"0000001800000000000000270000000000000020000000000000003300000000",
            INIT_67 => X"00000018000000000000002b0000000000000023000000000000000f00000000",
            INIT_68 => X"00000042000000000000004f0000000000000054000000000000005300000000",
            INIT_69 => X"00000031000000000000003a0000000000000042000000000000003a00000000",
            INIT_6A => X"0000001c00000000000000200000000000000047000000000000004300000000",
            INIT_6B => X"0000003d000000000000003d000000000000000b000000000000003200000000",
            INIT_6C => X"0000003500000000000000480000000000000048000000000000003500000000",
            INIT_6D => X"0000002d000000000000002e0000000000000031000000000000003800000000",
            INIT_6E => X"0000002d00000000000000210000000000000025000000000000003900000000",
            INIT_6F => X"0000003f0000000000000031000000000000003b000000000000001900000000",
            INIT_70 => X"00000045000000000000003b0000000000000046000000000000003800000000",
            INIT_71 => X"0000004d00000000000000380000000000000043000000000000004500000000",
            INIT_72 => X"00000022000000000000003e0000000000000022000000000000003600000000",
            INIT_73 => X"00000046000000000000003b000000000000002f000000000000003200000000",
            INIT_74 => X"00000040000000000000003b0000000000000040000000000000002b00000000",
            INIT_75 => X"000000350000000000000042000000000000003b000000000000003e00000000",
            INIT_76 => X"00000032000000000000002e000000000000003a000000000000003300000000",
            INIT_77 => X"0000004000000000000000240000000000000022000000000000003100000000",
            INIT_78 => X"00000017000000000000002d0000000000000037000000000000001c00000000",
            INIT_79 => X"0000004300000000000000450000000000000023000000000000004800000000",
            INIT_7A => X"0000003f000000000000002a000000000000002b000000000000005300000000",
            INIT_7B => X"0000003100000000000000260000000000000022000000000000002800000000",
            INIT_7C => X"0000002e000000000000001f0000000000000022000000000000002000000000",
            INIT_7D => X"0000003f000000000000003c0000000000000039000000000000003500000000",
            INIT_7E => X"000000320000000000000039000000000000002a000000000000004100000000",
            INIT_7F => X"0000001c00000000000000260000000000000026000000000000002300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE64;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE65 : if BRAM_NAME = "samplegold_layersamples_instance65" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002b0000000000000033000000000000002d000000000000004000000000",
            INIT_01 => X"00000040000000000000004b0000000000000049000000000000004500000000",
            INIT_02 => X"0000002900000000000000320000000000000032000000000000003b00000000",
            INIT_03 => X"000000330000000000000031000000000000002e000000000000002b00000000",
            INIT_04 => X"00000042000000000000002a000000000000002d000000000000003800000000",
            INIT_05 => X"000000260000000000000028000000000000002a000000000000002900000000",
            INIT_06 => X"0000002f000000000000002d000000000000002e000000000000002b00000000",
            INIT_07 => X"0000003500000000000000330000000000000032000000000000003700000000",
            INIT_08 => X"0000002d00000000000000240000000000000037000000000000002200000000",
            INIT_09 => X"00000010000000000000000b000000000000002c000000000000002d00000000",
            INIT_0A => X"0000002300000000000000190000000000000011000000000000000b00000000",
            INIT_0B => X"0000003600000000000000380000000000000032000000000000002b00000000",
            INIT_0C => X"0000002d000000000000002c000000000000003e000000000000002e00000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"000000280000000000000032000000000000003c000000000000002700000000",
            INIT_10 => X"000000210000000000000027000000000000002b000000000000004800000000",
            INIT_11 => X"0000000000000000000000110000000000000017000000000000000000000000",
            INIT_12 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"00000038000000000000002e000000000000002d000000000000003600000000",
            INIT_14 => X"0000000000000000000000100000000000000029000000000000002f00000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_16 => X"0000002f00000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"000000380000000000000027000000000000001c000000000000003200000000",
            INIT_18 => X"0000000a00000000000000000000000000000004000000000000002800000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000003300000000000000100000000000000000000000000000000000000000",
            INIT_1B => X"00000022000000000000003a000000000000002d000000000000002c00000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000002600000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000002e000000000000002c0000000000000012000000000000000000000000",
            INIT_1F => X"0000003300000000000000170000000000000038000000000000002e00000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_21 => X"0000000000000000000000010000000000000005000000000000000000000000",
            INIT_22 => X"0000003900000000000000020000000000000011000000000000001000000000",
            INIT_23 => X"0000000b000000000000003c0000000000000007000000000000002e00000000",
            INIT_24 => X"000000000000000000000009000000000000001d000000000000000800000000",
            INIT_25 => X"0000000300000000000000000000000000000013000000000000000500000000",
            INIT_26 => X"0000002100000000000000450000000000000012000000000000001900000000",
            INIT_27 => X"000000180000000000000000000000000000002d000000000000000000000000",
            INIT_28 => X"0000000400000000000000110000000000000003000000000000000000000000",
            INIT_29 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"000000000000000000000026000000000000002d000000000000000000000000",
            INIT_2B => X"0000000f00000000000000040000000000000000000000000000001a00000000",
            INIT_2C => X"00000000000000000000000f0000000000000000000000000000000100000000",
            INIT_2D => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_2E => X"0000001c00000000000000000000000000000015000000000000002f00000000",
            INIT_2F => X"00000020000000000000000a0000000000000000000000000000000900000000",
            INIT_30 => X"000000120000000000000012000000000000003c000000000000000000000000",
            INIT_31 => X"00000020000000000000001d0000000000000000000000000000002c00000000",
            INIT_32 => X"00000010000000000000000d0000000000000000000000000000000c00000000",
            INIT_33 => X"0000000d000000000000000d0000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000210000000000000036000000000000001300000000",
            INIT_35 => X"0000000e00000000000000260000000000000010000000000000000300000000",
            INIT_36 => X"00000002000000000000000d0000000000000000000000000000000800000000",
            INIT_37 => X"000000140000000000000011000000000000000c000000000000000000000000",
            INIT_38 => X"000000000000000000000000000000000000000c000000000000002d00000000",
            INIT_39 => X"000000000000000000000002000000000000001e000000000000001a00000000",
            INIT_3A => X"0000000000000000000000050000000000000004000000000000000000000000",
            INIT_3B => X"0000000e000000000000000b0000000000000008000000000000000800000000",
            INIT_3C => X"0000001400000000000000000000000000000002000000000000001400000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"000000060000000000000003000000000000000f000000000000000500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000160000000000000000000000000000000300000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000a00000000000000050000000000000000000000000000000000000000",
            INIT_43 => X"00000011000000000000000d0000000000000014000000000000000e00000000",
            INIT_44 => X"000000000000000000000012000000000000000a000000000000000200000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"000000040000000000000008000000000000001a000000000000001800000000",
            INIT_48 => X"000000000000000000000000000000000000002d000000000000000700000000",
            INIT_49 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"000000000000000000000000000000000000001c000000000000001900000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_52 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000300000000000000000000000000000000000000000000001600000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000002700000000000000180000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000070000000000000004000000000000000000000000",
            INIT_5A => X"0000000200000000000000060000000000000010000000000000000a00000000",
            INIT_5B => X"0000002200000000000000000000000000000000000000000000002000000000",
            INIT_5C => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000002600000000000000000000000000000002000000000000000000000000",
            INIT_5F => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_60 => X"0000000900000000000000100000000000000000000000000000001400000000",
            INIT_61 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_62 => X"0000000000000000000000260000000000000000000000000000000000000000",
            INIT_63 => X"0000000800000000000000000000000000000013000000000000000000000000",
            INIT_64 => X"0000000800000000000000000000000000000000000000000000000700000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_67 => X"0000001400000000000000000000000000000000000000000000000400000000",
            INIT_68 => X"00000000000000000000003e0000000000000000000000000000002e00000000",
            INIT_69 => X"000000230000000000000000000000000000001e000000000000000000000000",
            INIT_6A => X"0000000400000000000000000000000000000000000000000000001800000000",
            INIT_6B => X"0000001200000000000000050000000000000000000000000000000000000000",
            INIT_6C => X"00000000000000000000001e0000000000000013000000000000001300000000",
            INIT_6D => X"0000001f00000000000000070000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000001400000000000000100000000000000000000000000000000000000000",
            INIT_70 => X"000000000000000000000000000000000000002f000000000000000c00000000",
            INIT_71 => X"00000000000000000000000f0000000000000017000000000000000000000000",
            INIT_72 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000b000000000000000b0000000000000009000000000000000000000000",
            INIT_74 => X"000000000000000000000000000000000000000c000000000000000b00000000",
            INIT_75 => X"0000007700000000000000790000000000000019000000000000001300000000",
            INIT_76 => X"0000005c000000000000005c000000000000005e000000000000007c00000000",
            INIT_77 => X"0000008300000000000000820000000000000066000000000000005d00000000",
            INIT_78 => X"0000006d00000000000000690000000000000081000000000000007f00000000",
            INIT_79 => X"0000008d000000000000008f000000000000008f000000000000005e00000000",
            INIT_7A => X"000000820000000000000084000000000000007a000000000000005900000000",
            INIT_7B => X"0000007a00000000000000890000000000000099000000000000009100000000",
            INIT_7C => X"00000071000000000000006e0000000000000082000000000000008600000000",
            INIT_7D => X"0000004600000000000000880000000000000099000000000000009800000000",
            INIT_7E => X"0000007800000000000000780000000000000083000000000000007600000000",
            INIT_7F => X"000000860000000000000078000000000000008b000000000000008400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE65;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE66 : if BRAM_NAME = "samplegold_layersamples_instance66" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000097000000000000006f0000000000000061000000000000007a00000000",
            INIT_01 => X"00000090000000000000005a0000000000000083000000000000009700000000",
            INIT_02 => X"0000009800000000000000a6000000000000008e000000000000008b00000000",
            INIT_03 => X"00000072000000000000008c0000000000000094000000000000009000000000",
            INIT_04 => X"0000009400000000000000950000000000000054000000000000005b00000000",
            INIT_05 => X"0000009c00000000000000930000000000000060000000000000007b00000000",
            INIT_06 => X"0000009c00000000000000a2000000000000009e000000000000008f00000000",
            INIT_07 => X"000000700000000000000085000000000000008d000000000000009800000000",
            INIT_08 => X"00000055000000000000008e000000000000008d000000000000005500000000",
            INIT_09 => X"000000860000000000000081000000000000007b000000000000005a00000000",
            INIT_0A => X"0000009b0000000000000095000000000000008d000000000000008b00000000",
            INIT_0B => X"00000098000000000000009800000000000000a2000000000000009700000000",
            INIT_0C => X"00000042000000000000005f000000000000006c000000000000007f00000000",
            INIT_0D => X"0000006d000000000000007f0000000000000080000000000000005c00000000",
            INIT_0E => X"000000730000000000000061000000000000007e000000000000007200000000",
            INIT_0F => X"00000062000000000000009c0000000000000094000000000000009a00000000",
            INIT_10 => X"0000006d000000000000004b0000000000000048000000000000003d00000000",
            INIT_11 => X"00000059000000000000005c0000000000000064000000000000006600000000",
            INIT_12 => X"00000072000000000000005a0000000000000055000000000000005500000000",
            INIT_13 => X"00000020000000000000005600000000000000aa000000000000008200000000",
            INIT_14 => X"00000053000000000000005e0000000000000039000000000000005c00000000",
            INIT_15 => X"0000002b00000000000000260000000000000034000000000000005100000000",
            INIT_16 => X"00000069000000000000004e000000000000001f000000000000002900000000",
            INIT_17 => X"000000560000000000000030000000000000006a000000000000009900000000",
            INIT_18 => X"0000005c00000000000000480000000000000055000000000000001300000000",
            INIT_19 => X"000000820000000000000083000000000000007e000000000000006100000000",
            INIT_1A => X"00000082000000000000005b0000000000000084000000000000007e00000000",
            INIT_1B => X"0000002b000000000000003f0000000000000023000000000000007400000000",
            INIT_1C => X"000000440000000000000041000000000000003a000000000000002900000000",
            INIT_1D => X"00000062000000000000005f000000000000005d000000000000006200000000",
            INIT_1E => X"00000082000000000000006f0000000000000058000000000000004f00000000",
            INIT_1F => X"0000001c0000000000000043000000000000003d000000000000003100000000",
            INIT_20 => X"000000520000000000000029000000000000005a000000000000002600000000",
            INIT_21 => X"0000002400000000000000780000000000000058000000000000004c00000000",
            INIT_22 => X"0000003800000000000000870000000000000064000000000000006500000000",
            INIT_23 => X"00000016000000000000002e000000000000006b000000000000003e00000000",
            INIT_24 => X"0000005d0000000000000026000000000000001c000000000000001500000000",
            INIT_25 => X"0000002a000000000000001f000000000000004f000000000000005c00000000",
            INIT_26 => X"0000006000000000000000820000000000000085000000000000006800000000",
            INIT_27 => X"00000011000000000000001e000000000000004a000000000000005f00000000",
            INIT_28 => X"00000080000000000000007c0000000000000028000000000000001b00000000",
            INIT_29 => X"000000700000000000000035000000000000000d000000000000006600000000",
            INIT_2A => X"000000480000000000000069000000000000007d000000000000008a00000000",
            INIT_2B => X"00000025000000000000001d0000000000000028000000000000004800000000",
            INIT_2C => X"0000005300000000000000600000000000000045000000000000003000000000",
            INIT_2D => X"0000001800000000000000780000000000000034000000000000001100000000",
            INIT_2E => X"0000001500000000000000210000000000000012000000000000001700000000",
            INIT_2F => X"0000000e000000000000000e0000000000000011000000000000000b00000000",
            INIT_30 => X"00000020000000000000001b000000000000001d000000000000001700000000",
            INIT_31 => X"0000000d000000000000000c000000000000002e000000000000002200000000",
            INIT_32 => X"0000000000000000000000000000000000000015000000000000000d00000000",
            INIT_33 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000002b000000000000001c0000000000000014000000000000002500000000",
            INIT_35 => X"0000000f000000000000000b000000000000000b000000000000002c00000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000002b000000000000002b000000000000001a000000000000001200000000",
            INIT_39 => X"0000000400000000000000120000000000000009000000000000000b00000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000c00000000000000290000000000000025000000000000001d00000000",
            INIT_3D => X"0000000000000000000000000000000000000007000000000000000b00000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000500000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000a00000000000000090000000000000019000000000000001500000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000001000000000000000130000000000000006000000000000000a00000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"00000000000000000000000d000000000000001d000000000000001000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"00000000000000000000001a0000000000000000000000000000001c00000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000001a000000000000000e0000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"00000000000000000000001f0000000000000006000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000003000000000000000300000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_58 => X"0000000b00000000000000000000000000000002000000000000000400000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000600000000000000060000000000000009000000000000000900000000",
            INIT_5D => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000007000000000000000d00000000",
            INIT_61 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000600000000000000020000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_65 => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000300000000000000000000000000000000000000000000000300000000",
            INIT_68 => X"0000000e00000000000000000000000000000000000000000000001200000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000004d000000000000003d0000000000000041000000000000003c00000000",
            INIT_6C => X"0000000600000000000000220000000000000015000000000000004400000000",
            INIT_6D => X"0000000400000000000000020000000000000022000000000000000000000000",
            INIT_6E => X"00000000000000000000002a0000000000000000000000000000000000000000",
            INIT_6F => X"0000003000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000011000000000000007700000000",
            INIT_71 => X"0000000000000000000000000000000000000002000000000000004d00000000",
            INIT_72 => X"000000000000000000000025000000000000006a000000000000000000000000",
            INIT_73 => X"0000001800000000000000050000000000000001000000000000000d00000000",
            INIT_74 => X"0000000d00000000000000000000000000000000000000000000006400000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_76 => X"0000001900000000000000000000000000000035000000000000004d00000000",
            INIT_77 => X"0000006100000000000000000000000000000021000000000000001d00000000",
            INIT_78 => X"0000003400000000000000000000000000000000000000000000002200000000",
            INIT_79 => X"0000005400000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000001c00000000000000180000000000000000000000000000002000000000",
            INIT_7B => X"0000006b0000000000000055000000000000002a000000000000002c00000000",
            INIT_7C => X"0000000000000000000000290000000000000004000000000000000000000000",
            INIT_7D => X"0000000e00000000000000030000000000000000000000000000000800000000",
            INIT_7E => X"0000000e000000000000001f0000000000000000000000000000000000000000",
            INIT_7F => X"0000005c0000000000000074000000000000005b000000000000000300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE66;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE67 : if BRAM_NAME = "samplegold_layersamples_instance67" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005700000000000000000000000000000000000000000000002900000000",
            INIT_01 => X"0000000400000000000000000000000000000002000000000000000000000000",
            INIT_02 => X"000000090000000000000029000000000000001f000000000000000000000000",
            INIT_03 => X"0000009b000000000000005c0000000000000072000000000000003500000000",
            INIT_04 => X"00000000000000000000004e0000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000010000000000000014000000000000003200000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000ab0000000000000000000000000000000b00000000",
            INIT_08 => X"0000003d00000000000000000000000000000040000000000000000000000000",
            INIT_09 => X"00000003000000000000006f000000000000003c000000000000000000000000",
            INIT_0A => X"0000002a00000000000000260000000000000014000000000000003700000000",
            INIT_0B => X"00000000000000000000000000000000000000cc000000000000000000000000",
            INIT_0C => X"0000003400000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000680000000000000000000000000000002600000000",
            INIT_0E => X"0000001d0000000000000000000000000000002f000000000000000300000000",
            INIT_0F => X"0000004700000000000000000000000000000000000000000000009400000000",
            INIT_10 => X"00000064000000000000001b0000000000000000000000000000000000000000",
            INIT_11 => X"00000004000000000000000c0000000000000091000000000000000000000000",
            INIT_12 => X"000000ce00000000000000390000000000000000000000000000002900000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_14 => X"0000001700000000000000070000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000085000000000000002f00000000",
            INIT_16 => X"0000001100000000000000b50000000000000032000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000002e00000000000000120000000000000000000000000000000000000000",
            INIT_19 => X"000000000000000000000000000000000000004a000000000000007000000000",
            INIT_1A => X"000000000000000000000000000000000000009f000000000000005000000000",
            INIT_1B => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_1C => X"0000002300000000000000150000000000000006000000000000000000000000",
            INIT_1D => X"0000003f00000000000000000000000000000000000000000000003d00000000",
            INIT_1E => X"000000000000000000000000000000000000000000000000000000ae00000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"00000087000000000000006c0000000000000051000000000000004800000000",
            INIT_24 => X"0000000000000000000000230000000000000054000000000000007a00000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"000000000000000000000000000000000000001d000000000000000b00000000",
            INIT_29 => X"0000000000000000000000000000000000000029000000000000000e00000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000032000000000000000000000000",
            INIT_2D => X"0000003700000000000000000000000000000000000000000000000600000000",
            INIT_2E => X"0000002c00000000000000200000000000000007000000000000002700000000",
            INIT_2F => X"00000000000000000000000e0000000000000007000000000000000600000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000002000000000000001400000000",
            INIT_32 => X"000000210000000000000000000000000000000b000000000000003e00000000",
            INIT_33 => X"0000002900000000000000340000000000000015000000000000002900000000",
            INIT_34 => X"0000000700000000000000000000000000000000000000000000000400000000",
            INIT_35 => X"0000000000000000000000000000000000000027000000000000002400000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"00000069000000000000003a000000000000001c000000000000001100000000",
            INIT_38 => X"0000003d00000000000000070000000000000008000000000000006900000000",
            INIT_39 => X"0000000000000000000000220000000000000000000000000000000e00000000",
            INIT_3A => X"0000004d000000000000004c000000000000000c000000000000000000000000",
            INIT_3B => X"000000340000000000000067000000000000005b000000000000002d00000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_3D => X"00000000000000000000000a0000000000000000000000000000006400000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000003000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000400000000000000000000000000000000000000000",
            INIT_41 => X"0000004500000000000000380000000000000017000000000000003400000000",
            INIT_42 => X"00000046000000000000004a000000000000003f000000000000003800000000",
            INIT_43 => X"0000000000000000000000260000000000000032000000000000003c00000000",
            INIT_44 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000002c00000000000000000000000000000000000000000000002300000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"000000110000000000000005000000000000000c000000000000000000000000",
            INIT_48 => X"0000001300000000000000000000000000000000000000000000002800000000",
            INIT_49 => X"00000030000000000000003a0000000000000041000000000000006b00000000",
            INIT_4A => X"00000050000000000000003b0000000000000022000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000003000000000000003a00000000",
            INIT_4C => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000007000000000000000800000000",
            INIT_4E => X"0000000000000000000000080000000000000008000000000000000000000000",
            INIT_4F => X"0000000400000000000000000000000000000008000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000200000000000000530000000000000051000000000000000000000000",
            INIT_52 => X"0000000c00000000000000150000000000000008000000000000000700000000",
            INIT_53 => X"0000000700000000000000130000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000110000000000000027000000000000000900000000",
            INIT_56 => X"000000a6000000000000009f0000000000000000000000000000000500000000",
            INIT_57 => X"0000008400000000000000720000000000000071000000000000009200000000",
            INIT_58 => X"000000a400000000000000bd00000000000000b9000000000000009600000000",
            INIT_59 => X"000000b20000000000000097000000000000009d00000000000000a000000000",
            INIT_5A => X"0000009500000000000000a800000000000000a6000000000000008800000000",
            INIT_5B => X"00000031000000000000002a000000000000002c000000000000003500000000",
            INIT_5C => X"00000081000000000000006e0000000000000045000000000000002c00000000",
            INIT_5D => X"000000a2000000000000008f000000000000009a00000000000000a200000000",
            INIT_5E => X"0000000b000000000000007f000000000000009f000000000000009e00000000",
            INIT_5F => X"0000001f00000000000000220000000000000026000000000000000b00000000",
            INIT_60 => X"000000a5000000000000008b0000000000000039000000000000001a00000000",
            INIT_61 => X"0000009e000000000000009f0000000000000076000000000000009600000000",
            INIT_62 => X"0000004700000000000000000000000000000079000000000000009400000000",
            INIT_63 => X"0000001800000000000000090000000000000022000000000000005000000000",
            INIT_64 => X"0000008900000000000000890000000000000067000000000000002d00000000",
            INIT_65 => X"00000090000000000000009d000000000000008b000000000000009600000000",
            INIT_66 => X"0000001e00000000000000220000000000000000000000000000004500000000",
            INIT_67 => X"0000001a00000000000000190000000000000008000000000000000000000000",
            INIT_68 => X"0000009100000000000000aa000000000000009b000000000000002400000000",
            INIT_69 => X"00000044000000000000007d000000000000009200000000000000b300000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000a00000000000000010000000000000000000000000000000000000000",
            INIT_6C => X"0000009f000000000000009e000000000000009d000000000000004100000000",
            INIT_6D => X"0000000500000000000000450000000000000049000000000000008800000000",
            INIT_6E => X"0000000000000000000000000000000000000013000000000000002900000000",
            INIT_6F => X"0000003700000000000000110000000000000014000000000000001100000000",
            INIT_70 => X"0000007200000000000000980000000000000067000000000000005900000000",
            INIT_71 => X"000000000000000000000040000000000000005f000000000000001900000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"00000029000000000000007f0000000000000097000000000000002800000000",
            INIT_75 => X"0000003300000000000000100000000000000000000000000000007600000000",
            INIT_76 => X"00000082000000000000006a0000000000000020000000000000002500000000",
            INIT_77 => X"000000430000000000000079000000000000006b000000000000005c00000000",
            INIT_78 => X"0000002b0000000000000009000000000000006e000000000000009000000000",
            INIT_79 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_7A => X"000000000000000000000011000000000000000a000000000000002400000000",
            INIT_7B => X"0000007200000000000000000000000000000018000000000000000300000000",
            INIT_7C => X"0000000000000000000000310000000000000003000000000000007200000000",
            INIT_7D => X"0000000d00000000000000240000000000000000000000000000000000000000",
            INIT_7E => X"0000002800000000000000000000000000000005000000000000000100000000",
            INIT_7F => X"0000005b00000000000000790000000000000021000000000000000700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE67;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE68 : if BRAM_NAME = "samplegold_layersamples_instance68" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000700000000000000360000000000000014000000000000000000000000",
            INIT_01 => X"0000004800000000000000000000000000000000000000000000000300000000",
            INIT_02 => X"00000000000000000000004d0000000000000035000000000000001900000000",
            INIT_03 => X"0000001f000000000000003d000000000000004f000000000000000000000000",
            INIT_04 => X"0000000300000000000000000000000000000022000000000000005d00000000",
            INIT_05 => X"0000008900000000000000100000000000000000000000000000000000000000",
            INIT_06 => X"0000000b0000000000000000000000000000002c000000000000007e00000000",
            INIT_07 => X"00000011000000000000002e0000000000000053000000000000006b00000000",
            INIT_08 => X"000000080000000000000000000000000000000a000000000000001800000000",
            INIT_09 => X"0000001b00000000000000310000000000000027000000000000001300000000",
            INIT_0A => X"0000004e00000000000000210000000000000000000000000000000000000000",
            INIT_0B => X"00000003000000000000001d000000000000002a000000000000002b00000000",
            INIT_0C => X"0000000f000000000000000f0000000000000000000000000000000500000000",
            INIT_0D => X"0000000000000000000000150000000000000011000000000000001000000000",
            INIT_0E => X"0000003b00000000000000620000000000000014000000000000000100000000",
            INIT_0F => X"0000002e000000000000005d0000000000000042000000000000003000000000",
            INIT_10 => X"0000002000000000000000150000000000000027000000000000002500000000",
            INIT_11 => X"0000005000000000000000360000000000000043000000000000004200000000",
            INIT_12 => X"000000410000000000000045000000000000004a000000000000002700000000",
            INIT_13 => X"0000001c0000000000000030000000000000009a000000000000005b00000000",
            INIT_14 => X"0000002d000000000000002a0000000000000035000000000000002400000000",
            INIT_15 => X"0000005c0000000000000042000000000000001f000000000000003a00000000",
            INIT_16 => X"0000006e00000000000000450000000000000048000000000000001b00000000",
            INIT_17 => X"00000018000000000000000e000000000000000000000000000000bd00000000",
            INIT_18 => X"0000000000000000000000000000000000000014000000000000002700000000",
            INIT_19 => X"00000000000000000000005e000000000000004e000000000000002700000000",
            INIT_1A => X"000000cc00000000000000550000000000000053000000000000004800000000",
            INIT_1B => X"0000003a000000000000006f0000000000000030000000000000000000000000",
            INIT_1C => X"0000000000000000000000170000000000000026000000000000003a00000000",
            INIT_1D => X"00000044000000000000002f0000000000000050000000000000004e00000000",
            INIT_1E => X"00000000000000000000009c0000000000000083000000000000005900000000",
            INIT_1F => X"00000028000000000000002c000000000000005b000000000000001c00000000",
            INIT_20 => X"0000002800000000000000000000000000000042000000000000002f00000000",
            INIT_21 => X"0000006d0000000000000028000000000000001d000000000000006100000000",
            INIT_22 => X"0000002100000000000000000000000000000097000000000000007900000000",
            INIT_23 => X"0000001b00000000000000350000000000000032000000000000002e00000000",
            INIT_24 => X"0000004a00000000000000000000000000000010000000000000002e00000000",
            INIT_25 => X"00000045000000000000007d0000000000000022000000000000004600000000",
            INIT_26 => X"0000004b0000000000000024000000000000000b000000000000006f00000000",
            INIT_27 => X"0000003c00000000000000320000000000000010000000000000002e00000000",
            INIT_28 => X"0000003200000000000000250000000000000000000000000000000000000000",
            INIT_29 => X"0000006e00000000000000000000000000000084000000000000005300000000",
            INIT_2A => X"0000002e00000000000000170000000000000039000000000000004000000000",
            INIT_2B => X"0000001c0000000000000021000000000000002a000000000000002d00000000",
            INIT_2C => X"0000004b00000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000900000000000000000000000000000008b00000000",
            INIT_2E => X"00000000000000000000004b0000000000000039000000000000001a00000000",
            INIT_2F => X"000000000000000000000000000000000000003f000000000000000000000000",
            INIT_30 => X"000000a7000000000000005f0000000000000000000000000000002a00000000",
            INIT_31 => X"0000002c00000000000000000000000000000050000000000000000200000000",
            INIT_32 => X"00000011000000000000004d0000000000000000000000000000000000000000",
            INIT_33 => X"0000005700000000000000220000000000000027000000000000003b00000000",
            INIT_34 => X"0000000500000000000000c30000000000000044000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000016000000000000002e00000000",
            INIT_36 => X"0000001900000000000000330000000000000000000000000000004300000000",
            INIT_37 => X"0000000000000000000000000000000000000047000000000000000000000000",
            INIT_38 => X"00000009000000000000000000000000000000ca000000000000004900000000",
            INIT_39 => X"0000006600000000000000000000000000000000000000000000004d00000000",
            INIT_3A => X"0000000b0000000000000020000000000000003f000000000000000000000000",
            INIT_3B => X"0000003f00000000000000000000000000000003000000000000009000000000",
            INIT_3C => X"0000004800000000000000280000000000000000000000000000007e00000000",
            INIT_3D => X"0000000000000000000000000000000000000001000000000000002700000000",
            INIT_3E => X"0000004600000000000000870000000000000041000000000000000000000000",
            INIT_3F => X"0000005800000000000000250000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004d00000000000000220000000000000037000000000000006100000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"000000000000000000000033000000000000008a000000000000001100000000",
            INIT_43 => X"00000051000000000000003e0000000000000043000000000000000000000000",
            INIT_44 => X"00000004000000000000002f0000000000000019000000000000004900000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000030000000000000005700000000",
            INIT_47 => X"000000ae00000000000000af000000000000009900000000000000a500000000",
            INIT_48 => X"0000006b00000000000000750000000000000072000000000000008100000000",
            INIT_49 => X"0000009f00000000000000aa00000000000000ac000000000000007e00000000",
            INIT_4A => X"000000b200000000000000a4000000000000008800000000000000b900000000",
            INIT_4B => X"0000006a00000000000000cf00000000000000c800000000000000af00000000",
            INIT_4C => X"0000007a0000000000000074000000000000005b000000000000005c00000000",
            INIT_4D => X"000000a90000000000000089000000000000009b000000000000008800000000",
            INIT_4E => X"000000b400000000000000b7000000000000008100000000000000c500000000",
            INIT_4F => X"00000042000000000000002600000000000000f300000000000000d400000000",
            INIT_50 => X"000000390000000000000049000000000000005f000000000000004b00000000",
            INIT_51 => X"000000be00000000000000b50000000000000090000000000000004200000000",
            INIT_52 => X"000000b200000000000000c200000000000000b7000000000000005800000000",
            INIT_53 => X"0000009500000000000000650000000000000000000000000000010500000000",
            INIT_54 => X"0000005a00000000000000570000000000000070000000000000006e00000000",
            INIT_55 => X"0000007300000000000000b400000000000000b3000000000000006600000000",
            INIT_56 => X"000000c900000000000000c100000000000000c800000000000000b000000000",
            INIT_57 => X"00000054000000000000008b0000000000000045000000000000001900000000",
            INIT_58 => X"0000003a0000000000000089000000000000005b000000000000005900000000",
            INIT_59 => X"0000008c000000000000008a00000000000000d5000000000000008d00000000",
            INIT_5A => X"0000000800000000000000b000000000000000bb00000000000000d300000000",
            INIT_5B => X"00000053000000000000004e0000000000000057000000000000004600000000",
            INIT_5C => X"00000056000000000000004d000000000000005a000000000000004600000000",
            INIT_5D => X"000000cd000000000000007800000000000000b400000000000000b800000000",
            INIT_5E => X"0000003d00000000000000200000000000000099000000000000008100000000",
            INIT_5F => X"0000004f000000000000002e0000000000000044000000000000006e00000000",
            INIT_60 => X"0000007c00000000000000430000000000000020000000000000005600000000",
            INIT_61 => X"0000002f00000000000000af000000000000009e00000000000000a200000000",
            INIT_62 => X"000000330000000000000056000000000000005400000000000000a000000000",
            INIT_63 => X"00000035000000000000002e0000000000000032000000000000004c00000000",
            INIT_64 => X"00000037000000000000002d0000000000000007000000000000002200000000",
            INIT_65 => X"000000a2000000000000001a00000000000000af00000000000000a000000000",
            INIT_66 => X"0000006a00000000000000500000000000000036000000000000001800000000",
            INIT_67 => X"0000002b0000000000000073000000000000000d000000000000002100000000",
            INIT_68 => X"000000b70000000000000006000000000000004f000000000000000000000000",
            INIT_69 => X"000000030000000000000067000000000000003200000000000000d000000000",
            INIT_6A => X"00000078000000000000000a0000000000000015000000000000004a00000000",
            INIT_6B => X"00000062000000000000005c0000000000000072000000000000004900000000",
            INIT_6C => X"000000f1000000000000009c0000000000000000000000000000007800000000",
            INIT_6D => X"0000000700000000000000210000000000000047000000000000002400000000",
            INIT_6E => X"0000005c0000000000000006000000000000005b000000000000000f00000000",
            INIT_6F => X"00000032000000000000005f0000000000000027000000000000004400000000",
            INIT_70 => X"0000001400000000000000f30000000000000098000000000000000000000000",
            INIT_71 => X"0000000000000000000000050000000000000060000000000000003700000000",
            INIT_72 => X"0000004c00000000000000640000000000000000000000000000008100000000",
            INIT_73 => X"00000000000000000000001800000000000000a4000000000000003a00000000",
            INIT_74 => X"0000005e000000000000001900000000000000c7000000000000008200000000",
            INIT_75 => X"0000000000000000000000080000000000000039000000000000006e00000000",
            INIT_76 => X"000000c600000000000000770000000000000000000000000000000000000000",
            INIT_77 => X"0000006b00000000000000000000000000000000000000000000004c00000000",
            INIT_78 => X"0000004200000000000000690000000000000096000000000000009700000000",
            INIT_79 => X"0000000000000000000000000000000000000006000000000000006700000000",
            INIT_7A => X"0000004400000000000000d1000000000000004f000000000000000000000000",
            INIT_7B => X"0000007b000000000000007e0000000000000000000000000000000000000000",
            INIT_7C => X"0000004800000000000000360000000000000065000000000000008e00000000",
            INIT_7D => X"00000013000000000000000d0000000000000010000000000000001500000000",
            INIT_7E => X"00000000000000000000003a0000000000000086000000000000001c00000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE68;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE69 : if BRAM_NAME = "samplegold_layersamples_instance69" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000003800000000000000260000000000000028000000000000002b00000000",
            INIT_3D => X"0000000000000000000000180000000000000036000000000000004900000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000001100000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_43 => X"0000000000000000000000190000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_47 => X"0000001000000000000000000000000000000024000000000000002c00000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_4B => X"000000060000000000000000000000000000001b000000000000001f00000000",
            INIT_4C => X"000000150000000000000009000000000000001b000000000000001600000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_4E => X"000000000000000000000028000000000000002b000000000000000300000000",
            INIT_4F => X"0000000200000000000000070000000000000000000000000000000000000000",
            INIT_50 => X"00000018000000000000001c0000000000000009000000000000000000000000",
            INIT_51 => X"0000001a0000000000000000000000000000001d000000000000002f00000000",
            INIT_52 => X"0000001e000000000000000d0000000000000000000000000000005500000000",
            INIT_53 => X"0000004500000000000000280000000000000010000000000000001700000000",
            INIT_54 => X"0000003100000000000000480000000000000033000000000000003c00000000",
            INIT_55 => X"0000001100000000000000000000000000000000000000000000001b00000000",
            INIT_56 => X"000000010000000000000000000000000000005b000000000000000300000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000002500000000000000310000000000000000000000000000000000000000",
            INIT_5A => X"0000002c000000000000001f000000000000001a000000000000001a00000000",
            INIT_5B => X"0000003700000000000000250000000000000034000000000000001300000000",
            INIT_5C => X"000000000000000000000033000000000000001d000000000000002c00000000",
            INIT_5D => X"0000000a00000000000000030000000000000013000000000000000000000000",
            INIT_5E => X"000000220000000000000000000000000000000e000000000000001d00000000",
            INIT_5F => X"0000000000000000000000050000000000000008000000000000000700000000",
            INIT_60 => X"0000000300000000000000000000000000000000000000000000001e00000000",
            INIT_61 => X"0000000b00000000000000000000000000000000000000000000004e00000000",
            INIT_62 => X"00000012000000000000003c000000000000004b000000000000001f00000000",
            INIT_63 => X"00000047000000000000001e0000000000000000000000000000001800000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000003c00000000",
            INIT_65 => X"0000000900000000000000000000000000000002000000000000000000000000",
            INIT_66 => X"000000000000000000000001000000000000000d000000000000001100000000",
            INIT_67 => X"0000000000000000000000280000000000000000000000000000000000000000",
            INIT_68 => X"0000000b000000000000000d0000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000110000000000000008000000000000000c00000000",
            INIT_6A => X"0000002100000000000000300000000000000000000000000000000000000000",
            INIT_6B => X"000000000000000000000000000000000000001a000000000000002c00000000",
            INIT_6C => X"0000002100000000000000000000000000000000000000000000000500000000",
            INIT_6D => X"000000000000000000000000000000000000000c000000000000000d00000000",
            INIT_6E => X"00000019000000000000001d000000000000000b000000000000000200000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000002800000000000000280000000000000014000000000000000000000000",
            INIT_75 => X"00000025000000000000003a0000000000000038000000000000003000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000500000000000000010000000000000019000000000000001600000000",
            INIT_7D => X"0000000600000000000000080000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000600000000000000100000000000000013000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE69;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE70 : if BRAM_NAME = "samplegold_layersamples_instance70" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000b00000000000000060000000000000012000000000000001300000000",
            INIT_01 => X"00000000000000000000000a0000000000000000000000000000000e00000000",
            INIT_02 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"000000000000000000000007000000000000000e000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000001300000000000000120000000000000000000000000000000000000000",
            INIT_08 => X"0000001b000000000000002f000000000000001b000000000000000b00000000",
            INIT_09 => X"0000000100000000000000250000000000000026000000000000001f00000000",
            INIT_0A => X"0000000500000000000000010000000000000007000000000000000700000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_0C => X"00000028000000000000000e0000000000000006000000000000001500000000",
            INIT_0D => X"000000000000000000000003000000000000000d000000000000000d00000000",
            INIT_0E => X"000000050000000000000006000000000000000b000000000000000400000000",
            INIT_0F => X"0000000000000000000000000000000000000011000000000000001b00000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000100000000000000000000000000000011000000000000000a00000000",
            INIT_12 => X"0000000200000000000000070000000000000003000000000000001500000000",
            INIT_13 => X"0000000200000000000000090000000000000023000000000000000000000000",
            INIT_14 => X"0000000300000000000000140000000000000003000000000000000c00000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"000000000000000000000000000000000000000c000000000000000a00000000",
            INIT_1A => X"0000000a00000000000000200000000000000008000000000000000000000000",
            INIT_1B => X"0000002900000000000000000000000000000023000000000000002a00000000",
            INIT_1C => X"0000000000000000000000080000000000000005000000000000002000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000300000000000000000000000000000001000000000000000100000000",
            INIT_20 => X"0000000200000000000000020000000000000004000000000000000000000000",
            INIT_21 => X"0000000000000000000000010000000000000001000000000000000000000000",
            INIT_22 => X"0000000d000000000000000e0000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_24 => X"0000000000000000000000000000000000000001000000000000000300000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE70;

MEM_EMPTY_36Kb : if BRAM_NAME(1 to 7) = "default" generate
    BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
    generic map (
        BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
        DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
        DO_REG => 0,                     -- Optional output register (0 or 1)
        INIT => X"000000000000000000",   -- Initial values on output port
        INIT_FILE => "NONE",
        WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        SRVAL => X"000000000000000000",  -- Set/Reset value for port output
        WRITE_MODE => "WRITE_FIRST"      -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
    )
    port map (
        DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
        ADDR => bram_addr,  -- Input address, width defined by read/write port depth
        CLK => CLK,    -- 1-bit input clock
        DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
        EN => EN,      -- 1-bit input RAM enable
        REGCE => '1', -- 1-bit input output register enable
        RST => RST,    -- 1-bit input reset
        WE => bram_wr_en       -- Input write enable, width defined by write port depth
    );
-- End of BRAM_SINGLE_MACRO_inst instantiation
end generate;


end a1;