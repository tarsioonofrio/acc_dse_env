LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE gold_package is
		type padroes is array(0 to 4000000) of integer;
		constant gold: padroes := ( 0, 0, 0, 
		17, 0, 133, 
		32, 0, 0, 
		
		28, 0, 148, 
		0, 0, 0, 
		0, 0, 26, 
		
		0, 0, 0, 
		0, 0, 0, 
		84, 0, 79, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 113, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		6, 29, 184, 
		30, 52, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		41, 108, 4, 
		41, 0, 0, 
		15, 95, 80, 
		
		20, 77, 67, 
		54, 156, 100, 
		49, 0, 15, 
		
		0, 0, 0, 
		0, 0, 0, 
		65, 0, 0, 
		
		0, 0, 37, 
		4, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 24, 
		43, 23, 0, 
		
		0, 0, 0, 
		0, 63, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		74, 0, 14, 
		119, 45, 0, 
		0, 49, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		240, 0, 0, 
		74, 0, 0, 
		
		0, 0, 67, 
		0, 30, 149, 
		3, 0, 38, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		95, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		154, 2, 58, 
		0, 210, 162, 
		0, 69, 17, 
		
		42, 30, 184, 
		85, 98, 0, 
		7, 70, 47, 
		
		212, 147, 142, 
		48, 0, 17, 
		0, 0, 0, 
		
		88, 11, 0, 
		171, 0, 0, 
		0, 0, 0, 
		
		153, 0, 142, 
		0, 0, 0, 
		104, 0, 0, 
		
		0, 66, 7, 
		0, 111, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 19, 0, 
		147, 0, 0, 
		0, 50, 127, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		112, 0, 180, 
		192, 87, 209, 
		29, 214, 203, 
		
		40, 0, 62, 
		31, 13, 115, 
		76, 215, 252, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		8, 76, 106, 
		0, 0, 0, 
		
		3, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 11, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 9, 
		0, 0, 0, 
		
		5, 0, 134, 
		46, 8, 0, 
		0, 0, 129, 
		
		0, 0, 177, 
		0, 38, 141, 
		79, 0, 120, 
		
		75, 0, 0, 
		0, 4, 42, 
		0, 74, 2, 
		
		0, 0, 0, 
		12, 0, 0, 
		0, 40, 94, 
		
		7, 0, 0, 
		46, 9, 188, 
		42, 0, 0, 
		
		0, 58, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		143, 89, 218, 
		14, 172, 172, 
		0, 0, 0, 
		
		103, 0, 36, 
		0, 0, 0, 
		0, 0, 44, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		others=>0 );
END gold_package;
