LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE gold_package is
		type padroes is array(0 to 4000000) of integer;
		constant gold: padroes := ( 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		123, 232, 28, 4, 179, 221, 130, 
		94, 160, 121, 232, 137, 56, 45, 
		112, 12, 58, 165, 133, 0, 69, 
		131, 16, 6, 73, 32, 182, 147, 
		125, 253, 251, 195, 120, 218, 45, 
		159, 60, 187, 171, 77, 71, 76, 
		106, 83, 23, 138, 41, 70, 126, 
		
		0, 0, 0, 0, 202, 30, 168, 
		218, 0, 0, 0, 89, 113, 156, 
		247, 247, 0, 0, 230, 0, 0, 
		18, 0, 0, 23, 108, 0, 0, 
		0, 14, 159, 0, 0, 38, 0, 
		0, 29, 230, 0, 66, 0, 0, 
		254, 0, 193, 0, 0, 31, 0, 
		
		0, 0, 192, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 169, 0, 0, 142, 
		0, 130, 0, 0, 0, 62, 0, 
		0, 0, 0, 0, 0, 0, 108, 
		
		0, 117, 0, 0, 0, 0, 0, 
		0, 0, 0, 44, 0, 53, 225, 
		0, 0, 0, 0, 0, 49, 0, 
		0, 163, 0, 0, 0, 203, 0, 
		0, 0, 90, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 119, 0, 
		0, 156, 0, 0, 0, 78, 30, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		231, 66, 147, 17, 4, 39, 52, 
		119, 22, 0, 126, 93, 38, 31, 
		198, 118, 227, 235, 165, 177, 47, 
		207, 222, 148, 36, 230, 27, 248, 
		121, 47, 142, 219, 241, 8, 174, 
		218, 137, 21, 7, 0, 7, 91, 
		45, 3, 34, 201, 149, 191, 121, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 214, 60, 
		123, 38, 70, 72, 87, 31, 152, 
		133, 79, 36, 0, 144, 0, 93, 
		0, 0, 0, 72, 63, 154, 103, 
		0, 26, 0, 0, 0, 65, 0, 
		95, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 168, 129, 113, 41, 
		22, 7, 116, 78, 0, 205, 0, 
		0, 0, 0, 39, 0, 166, 16, 
		55, 163, 0, 0, 39, 11, 0, 
		0, 0, 91, 0, 182, 235, 0, 
		82, 0, 175, 76, 3, 0, 182, 
		28, 246, 47, 0, 2, 22, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 35, 0, 0, 0, 
		0, 0, 0, 152, 34, 0, 0, 
		11, 0, 0, 0, 0, 0, 0, 
		30, 0, 58, 129, 41, 50, 0, 
		0, 62, 184, 142, 26, 42, 115, 
		0, 21, 68, 8, 27, 13, 126, 
		
		134, 77, 201, 176, 28, 229, 129, 
		191, 88, 103, 153, 98, 78, 159, 
		238, 38, 174, 154, 119, 1, 124, 
		78, 82, 24, 97, 66, 236, 41, 
		98, 157, 147, 215, 84, 217, 8, 
		220, 125, 240, 116, 100, 20, 248, 
		176, 134, 189, 186, 120, 67, 205, 
		
		0, 149, 141, 0, 0, 0, 73, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 18, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 119, 
		62, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 94, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 76, 0, 2, 19, 89, 
		89, 14, 0, 59, 73, 32, 136, 
		154, 0, 79, 104, 0, 0, 88, 
		165, 65, 42, 39, 116, 200, 0, 
		13, 100, 0, 70, 147, 159, 115, 
		0, 0, 49, 1, 66, 195, 227, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 15, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 51, 90, 
		0, 0, 0, 82, 81, 118, 74, 
		
		0, 99, 108, 31, 145, 77, 5, 
		192, 123, 22, 237, 43, 95, 0, 
		224, 0, 17, 0, 0, 9, 0, 
		87, 92, 0, 18, 0, 0, 0, 
		0, 9, 92, 125, 215, 78, 199, 
		212, 0, 204, 95, 211, 22, 0, 
		79, 201, 137, 0, 0, 15, 69, 
		
		24, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 28, 55, 0, 
		0, 228, 176, 0, 0, 0, 0, 
		50, 0, 97, 22, 0, 116, 35, 
		71, 39, 103, 10, 0, 128, 51, 
		158, 0, 87, 34, 118, 31, 17, 
		161, 68, 98, 148, 29, 115, 35, 
		
		145, 38, 194, 38, 246, 0, 96, 
		0, 0, 112, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 60, 9, 
		0, 0, 0, 0, 0, 102, 0, 
		0, 0, 0, 0, 0, 0, 59, 
		0, 215, 199, 0, 35, 0, 0, 
		
		97, 0, 61, 100, 103, 144, 81, 
		146, 186, 114, 176, 215, 234, 138, 
		208, 152, 108, 200, 140, 152, 6, 
		237, 34, 52, 63, 193, 50, 239, 
		75, 147, 24, 15, 92, 33, 6, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		54, 58, 167, 223, 174, 73, 106, 
		0, 56, 87, 32, 0, 144, 138, 
		16, 79, 0, 35, 0, 40, 30, 
		0, 5, 0, 0, 0, 49, 0, 
		32, 0, 0, 0, 104, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		4, 37, 0, 6, 0, 0, 6, 
		11, 0, 0, 0, 0, 42, 192, 
		0, 0, 0, 62, 0, 0, 0, 
		0, 0, 0, 0, 57, 40, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 178, 0, 
		0, 0, 59, 117, 0, 13, 0, 
		143, 0, 50, 0, 0, 0, 0, 
		111, 0, 0, 124, 0, 0, 0, 
		29, 0, 97, 231, 92, 148, 154, 
		3, 113, 0, 0, 105, 122, 127, 
		
		139, 189, 127, 231, 137, 41, 75, 
		9, 69, 105, 234, 198, 0, 145, 
		110, 22, 172, 3, 242, 153, 31, 
		1, 179, 155, 123, 243, 72, 201, 
		231, 37, 175, 192, 140, 69, 159, 
		253, 14, 0, 0, 0, 0, 127, 
		0, 107, 0, 11, 149, 44, 111, 
		
		0, 0, 0, 51, 23, 62, 0, 
		0, 0, 0, 107, 0, 188, 108, 
		18, 0, 0, 110, 0, 17, 160, 
		71, 238, 0, 0, 0, 23, 0, 
		144, 0, 0, 234, 162, 0, 0, 
		0, 0, 0, 0, 55, 0, 138, 
		131, 0, 0, 0, 92, 72, 0, 
		
		239, 241, 84, 112, 91, 6, 47, 
		243, 135, 241, 134, 1, 125, 91, 
		136, 31, 26, 96, 189, 21, 59, 
		151, 189, 139, 44, 24, 0, 248, 
		136, 213, 156, 24, 136, 179, 59, 
		149, 232, 12, 66, 115, 169, 187, 
		29, 13, 97, 157, 0, 190, 67, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 32, 251, 173, 209, 59, 
		112, 142, 228, 224, 190, 143, 107, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 123, 0, 26, 126, 
		225, 71, 0, 17, 0, 129, 153, 
		21, 215, 24, 59, 159, 0, 112, 
		25, 0, 110, 0, 0, 187, 0, 
		0, 0, 15, 0, 164, 139, 0, 
		0, 0, 0, 0, 134, 153, 12, 
		
		0, 0, 0, 0, 0, 0, 0, 
		105, 0, 0, 0, 0, 0, 30, 
		0, 34, 0, 0, 64, 0, 0, 
		0, 100, 0, 0, 0, 18, 0, 
		0, 0, 0, 0, 0, 6, 0, 
		0, 0, 0, 0, 242, 0, 0, 
		139, 0, 64, 102, 175, 46, 0, 
		
		0, 0, 0, 0, 62, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 129, 0, 0, 76, 
		160, 198, 0, 0, 0, 0, 0, 
		118, 34, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 57, 184, 0, 
		0, 0, 0, 0, 18, 163, 0, 
		
		174, 21, 115, 120, 124, 46, 98, 
		19, 167, 95, 0, 0, 0, 182, 
		0, 13, 0, 0, 0, 0, 0, 
		0, 9, 0, 0, 24, 0, 129, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 62, 0, 
		0, 0, 0, 165, 96, 157, 184, 
		153, 0, 53, 83, 85, 31, 215, 
		
		others=>0 );
END gold_package;
