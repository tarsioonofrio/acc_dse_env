-gN_BRAM_IWGHT=30 -gN_BRAM_IFMAP=6