library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -- layer=2
    -4793, -4705, -405, 3023, 7547, -6642, 11021, -7940, 6175, -4770,

    -- weights
    -- layer=2 filter=0 channel=0
    19, -3, 16, -65, -29, -17, 8, 2, 0, -42, 5, 5, -51, 1, 7, -1, -13, 3, -6, 34, 49, 1, 1, -9, -24, -3, -42, 0, -38, 12, -34, 4, -5, -32, -33, 18, -18, 6, -11, -60, -27, 23, -41, -34, 24, -1, 3, 18, 9, 13, 50, -50, -40, 2, 17, 0, -48, 29, 1, -12, -3, -13, -3, 19, -15, 24, -60, 20, -23, 25, 3, -7, -8, 39, 25, 11, 62, 10, 9, -6, -74, 7, -45, 0, -43, 11, 7, -16, 3, 2, 16, 8, 32, 15, -6, 3, 6, 14, 12, 33, -5, -39, -1, -65, 5, 7, -10, -59, -1, 1, 22, 22, -16, -1, 1, 17, -2, -15, -33, 0, 4, 4, -55, 20, -10, 57, -30, -7, 8, -5, 1, -60, -18, -10, 0, 2, 4, -18, 20, -4, -19, -4, 9, 6, -10, -17, 26, 13, 28, -1, -4, -13, 5, 6, -34, -8, -63, 42, 24, 0, -16, -3, 13, 14, -41, 6, 19, -3, -46, 8, -28, -35, 16, -2, -3, -6, 23, -9, 31, 7, -15, -13, -20, -5, 12, 6, -25, 21, -4, -42, -8, 9, -16, 2, -52, 5, -26, 21, -14, -6, 24, 30, -9, -17, 36, -3, -10, 22, 1, 10, 32, 15, -19, 17, -35, -16, -28, 1, -5, 34, 15, 11, 0, -42, 2, 9, 7, 16, 7, -15, -5, 32, 0, 21, 9, -39, -1, 7, 9, 1, -5, 5, 23, 3, 2, -41, -19, 7, 0, -1, -48, 24, -19, 20, -27, 7, -1, -6, -3, -47, -4, -25, -42, 2, 10, -19, 18, 0, 27, -19, 8, -8, -13, -3, -1, -14, -11, 2, -3, -37, -30, -2, -16, -3, -27, 4, 11, 4, 0, 23, -6, -2, 9, 20, 15, -6, -62, -1, -19, -23, 10, -2, 3, -3, 9, -18, 12, -55, -20, 28, -9, -3, 3, -68, -15, 36, 2, -11, 2, 15, -8, -22, -29, -30, -21, 4, 2, 0, 6, -5, -6, -17, 14, 2, 21, 16, -5, -24, 8, 19, 4, -13, 50, -5, 4, 2, -12, 10, 8, 0, 6, -6, -3, 2, 3, 8, 35, -32, 7, 17, -7, -2, 18, -48, -3, 4, -4, 13, -5, 17, 2, 3, 1, -45, 7, -26, 0, -6, -55, -11, -10, -43, -25, -2, 3, 0, -9, -23, -19, -9, -24, 9, -6, -6, 21, 0, 36, -9, 8, -8, -9, 2, 8, 14, 62, 0, 0, -27, -31, 2, -10, -7, -2, 22, 9, 0, -12, 21, 34, 3, -33, 14, -6, -16, -5, 11, -28, 16, 23, -3, 2, 18, 11, 30, -4, -49, -16, 51, 18, -5, 20, 26, -28, 12, -12, -38, 1, 24, -7, 0, -19, 17, 9, -11, -23, -1, -25, -12, 13, 4, -6, 8, 49, -6, 41, 37, -23, 18, -15, -10, 31, -10, -21, -2, -7, 1, 18, 9, 3, -37, -5, 3, 12, 37, 0, -39, 2, -2, -7, -7, -8, -31, -5, -7, 3, 11, 4, 9, 14, 14, -25, -36, -6, 6, 11, -2, 18, -23, 5, -39, -2, 7, 0, -5, 10, 32, -26, -32, -4, 22, -17, 27, -14, -4, -41, -4, 13, 1, -7, 19, 23, -1, -23, 4, -4, -28, -25, 6, -2, 9, -5, -10, 34, 6, 11, 12, 9, -6, -3, -19, 4, 34, -62, -2, -36, -42, 0, -10, 4, -28, 24, -1, 15, -51, -42, 46, 4, -3, -7, 17, -4, -12, -11, -40, 19, 19, -14, -9, 0, 23, 10, 7, -12, -1, 7, 13, 7, -39, 11, -4, 3, 20, 0, 0, 24, 27, -16, 0, 88, -8, -1, -3, 11, 9, 8, 0, -7, -60, 2, 0, 5, 36, -1, -45, -3, 30, 4, 19, -22, -46, -2, 0, 2, 12, -11, 8, 19, -7, -22, -52, 3, -15, 8, -5, 38, -30, 11, -24, -9, -34, 4, -7, -7, 9, 0, -24, -21, 16, 3, -42, 23, -7, 5, -3, 11, -3, -4, -10, 22, -34, 13, 1, -5, -29, -11, 3, -23, 0, 31, 5, -1, -3, -31, 1, 0, -4, -21, -24, 2, 32, -35, 3, -55, -3, 4, 3, -4, -26, 2, -23, 5, -44, -21, -13, 0, -5, -32, 6, -10, 12, -14, -31, 1, 26, -17, 5, -40, 9, -25, -5, -18, -1, 62, -93, 8, -4, 30, 6, -33, 16, 4, -15, -8, -6, -9, -16, -35, -13, 8, 2, -4, 30, 9, 3, -3, -13, 0, 3, 3, -17, 15, -79, 3, -1, 3, 16, -10, -35, -5, 7, 6, -1, 5, 34, -1, 0, -21, -33, -41, -30, 11, 3, 11, -14, -4, 57, 0, 22, 0, 1, 4, 8, 9, -23, -27, 20, 2, -18, -35, 6, 8, 12, 9, -4, 1, -24, 4, -1, -9, 0, -4, -13, -12, 3, -6, -2, 58, 21, -20, 4, -15, 2, -52, -10, 27, -11, -10, -9, -47, 14, -68, -11, 2, -6, 0, -24, 13, 9, -31, -101, 2, 32, 24, -8, 5, 20, -42, -14, -3, -25, 14, 19, 21, 10, -99, 23, -13, -22, 34, -1, 30, -86, 2, -23, 18, -2, -3, -3, 0, 10, 14, -2, -38, -17, -40, -7, -20, -6, 17, 2, -5, 14, -4, -33, 2, -7, 10, 43, 41, -84, -1, -18, 0, -1, -2, -77, 7, -4, -14, 6, 4, 32, -1, -4, -23, -8, -98, -18, -8, 8, 17, 31, 13, -16, -14, 21, 8, -6, 19, -68, -2, 0, -25, -4, 5, -37, -71, 3, 7, -11, 13, 0, 0, -6, 1, 11, 27, 0, 4, 0, -26, -2, 12, 3, -48, 21, 22, 7, 3, 16, -15, -17, -8, -22, -6, 26, -26, -4, 8, -3, 11, -5, 10, 7, 6, -15, 16, -21, -26, 9, 1, -7, -5, 29, 0, 19, 3, -5, -27, 10, -3, 20, -42, -22, 13, 19, -1, -6, -10, 55, -26, -31, 2, 7, -24, 0, -15, -12, -3, 3, -14, -6, 8, 0, 3, -6, -2, -2, 32, 3, -6, -4, 3, 7, 11, 0, 20, -29, -6, -43, -6, 0, 2, -24, 7, -3, 18, 7, 1, 11, -50, -1, 10, 7, -2, 24, -9, 0, -49, 52, -8, 22, -27, -36, -2, 6, 13, -59, 16, 13, -5, 0, -1, 5, 19, 0, 6, -9, 13, 1, -9, -5, 56, 7, -49, -4, 5, -5, -18, 7, -14, -2, -33, 41, 31, -2, 0, 1, 14, 11, -16, -17, 3, -27, -19, -11, 12, -28, 8, 1, 7, 44, 1, 56, 29, -30, -1, -14, -14, -7, 26, 49, -37, 0, -8, -33, -21, 7, 6, -5, -27, -2, 13, 0, -12, 6, -27, 65, -24, 45, 31, 0, 34, 39, -1, 6, -24, 0, 9, -3, 34, -14, 10, -7, 4, -16, 7, -8, -1, -27, -9, 16, 2, -4, 17, 3, 3, 24, 2, 6, 21, 9, 2, -2, 12, -11, 0, -8, 3, 0, -19, -8, 15, 6, 12, 2, -32, 0, 0, 11, -30, -25, -1, -7, 33, -37, -22, 1, -42, 21, 7, 24, 32, -8, 29, -5, 12, 0, -7, -10, 10, -1, 23, -3, 4, -8, -1, -5, 11, -2, 2, 13, 33, -3, 12, -5, -11, -14, -12, 51, -1, 2, -14, -9, -10, -31, 4, 0, -4, 5, -3, -11, -14, 8, 1, -40, 9, 2, -23, 28, -5, 16, -7, 45, 7, 9, -6, 0, 11, -38, -13, 3, -23, 3, -15, 74, 15, 26, 29, 7, 49, 23, 4, -7, 7, 6, -14, -5, 44, -15, 19, -4, -13, 16, 23, 8, 4, -41, 0, 1, 2, -11, 14, -9, 6, 20, 6, 16, 32, 5, 2, -2, 6, 12, 7, 23, 1, -3, -6, 14, 17, 12, 21, -4, -19, -26, -8, -29, -6, -19, 9, -2, 1, 18, -1, -13, 6, -21, -3, -3, -21, -3, -29, -12, 7, -7, 0, 3, 18, -13, 27, 0, -3, -5, 6, -3, -26, -2, -2, 1, 31, 5, -20, -11, -15, -24, 0, 18, -6, -11, 14, 2, 15, -25, 3, -10, 6, -13, -19, 10, 36, 2, 3, -6, 13, -9, 33, 18, -11, -3, 1, -17, 1, 13, 4, 29, 16, -4, 13, 6, -27, -2, -33, 26, -10, 30, -11, -3, 27, 11, -55, 9, -5, 46, -13, 0, 46, -24, -28, 0, -6, -3, 16, -2, 7, -31, 0, 3, 13, 0, 0, -17, -2, 47, -4, 9, -11, -6, 6, -7, 5, 9, 12, -6, 2, 4, -17, -23, 9, 5, -8, 3, 4, -40, 5, -8, -22, -47, 4, -7, 17, 33, 1, 11, -6, -2, 0, 33, -2, 5, 20, -32, 15, -6, -12, -16, 51, -12, 8, 4, 0, -3, -5, 3, 4, -1, 13, -11, -1, -6, -1, -13, 17, -23, 28, -10, 8, 1, -13, -8, 11, -44, 8, -3, 2, 21, 22, -74, 10, -17, -6, 36, 0, 4, 5, -9, -18, -15, -2, 19, -3, -11, 28, 9, 16, 6, -4, 10, 8, 4, -8, -16, -2, 4, -10, -3, 30, 48, -43, -9, -3, 26, 0, -5, -4, 11, -11, -5, 8, -2, 23, 12, 1, -42, -5, 0, 10, 5, 11, -4, 3, 44, -1, -2, -6, -9, 0, -4, -14, 14, 15, 6, 27, 0, -9, 18, -4, 15, 3, 8, 29, 11, 15, 16, -3, -1, 10, 6, 18, 60, -25, -10, 7, -9, 10, 33, 35, -8, 39, -32, 14, 1, -6, -11, 12, -35, -34, 5, 3, -20, -18, 2, 14, -6, 49, 16, 27, 0, -9, -16, -34, -29, 4, -20, -1, 17, -3, -23, 18, -10, -3, 2, -3, -1, -1, -44, 11, -16, -4, 44, -1, -8, -6, 22, 43, -19, 0, -8, -7, 0, 8, 20, -14, 0, 24, 14, 30, 0, -15, -37, 17, -27, 3, 0, 86, 34, 26, 13, -11, 26, 7, 0, -10, -21, -14, 5, 9, -7, 26, 2, 0, -22, 0, -15, 14, -2, 17, -31, -1, 46, -7, -7, -8, -21, 0, -1, -2, 3, 3, 37, 1, -4, 1, 26, 1, -26, -30, 0, 26, 9, 4, -14, 35, 6, -1, 7, 17, 14, -36, -37, -8, -15, 13, 22, 18, -9, -7, -27, 8, -1, -6, -14, -5, -28, -32, -5, 3, -9, -18, -3, 2, 4, 78, -11, -26, 1, 21, 12, -41, -15, 43, -7, 9, 37, -18, 12, -46, -42, 9, 0, -3, -5, -14, 33, -1, 7, 12, 29, 13, -4, 19, 29, 43, -17, -18, -1, -12, -23, -25, 3, -36, -4, -29, 15, -2, -6, 22, -81, -15, -57, 0, 0, -30, 45, -8, -9, -14, -10, -9, -7, -19, 0, -11, 0, -15, 19, 0, -2, 0, -20, 2, -6, 7, 11, 20, -25, 4, 43, 1, 5, -15, -45, 3, 0, -2, -26, -29, 13, -22, -8, 12, 3, 23, -40, -15, 6, 42, 26, 8, 60, -3, -40, -14, 4, -6, -81, 8, 39, 18, -4, -8, -5, -70, 0, -25, -16, 5, 0, -3, 10, 0, 34, 49, -6, 5, 9, -25, -1, 12, 3, -55, 21, 38, 6, 9, 22, -37, -11, 10, 3, 3, -62, -35, 0, 5, 12, 11, 0, -4, 49, 7, -48, 50, -3, -31, 14, 3, -2, -22, 37, 4, 41, -2, 28, -8, 28, 17, 2, -11, -24, -22, 8, 4, -4, 5, 79, 5, 6, 31, 1, -44, 18, 24, -40, 23, 4, -1, 5, 10, 12, -2, 0, 18, -5, 15, -3, 7, 23, -7, -9, 3, 14, 3, 24, -5, 24, 3, 37, 9, -17, -5, -5, -2, 16, -17, 8, -69, -7, 5, 29, 14, -44, -46, 0, -45, -29, -33, 11, 0, 0, 1, -6, 6, -62, 6, 67, 9, -24, 0, -31, -48, 0, -8, 24, 15, -6, 0, 22, 35, -1, 41, -4, -9, 1, 2, -7, 1, 5, -46, 40, 25, 1, -11, 25, 22, 12, -28, 11, -5, -51, -27, -23, 29, 5, 18, 4, 4, 36, 39, -9, 41, 15, -29, 8, -9, -3, 17, 8, -24, 5, 0, 6, -2, 10, 4, -7, 0, 7, 26, 12, -11, -1, 9, 33, -12, 38, 12, 8, 40, -5, 5, -9, -14, 8, -7, 1, 39, -13, -2, -2, 11, -7, -5, 18, -2, -2, -4, -26, 16, 6, -1, 45, -6, -7, 5, -13, 11, 16, 2, 2, -9, 9, 31, -12, 9, 0, 5, 11, 2, 24, 0, 1, -47, -38, -25, 23, 5, -15, 5, 7, 23, -40, 20, 19, -31, -23, -5, -10, 10, -4, -24, -31, 11, 7, -6, 16, 8, 11, 0, 2, 5, -8, 6, 2, -35, 2, 7, -13, -16, 0, -4, -11, 3, 19, 23, -47, 17, -12, -20, -5, 11, -14, -4, -11, -2, 13, 17, 31, 42, 30, -2, -48, -4, -3, 56, 20, -27, -44, -1, 17, -13, -14, -2, 15, 0, -46, 20, 39, 6, -7, -33, 36, -10, 0, 19, 8, 37, -12, -49, 0, 6, 30, -5, 1, 39, 2, 17, -2, 25, 15, 23, 15, 4, 8, -4, 22, -3, 12, 8, 8, -1, 26, -3, 0, 11, -1, 2, 3, 2, -3, 3, 5, -9, 14, 5, -23, 1, 35, 11, -5, -18, -1, 19, 13, -45, -57, 30, -3, 39, -4, 15, -5, -28, 3, 5, -61, 19, -4, -16, -40, 7, -7, -11, 7, -30, -26, 60, 3, 5, -12, -4, 4, -28, 6, 11, -56, -3, 0, -21, -12, 8, 4, -14, -25, 24, -6, 6, 24, 3, -4, 31, 2, -4, -10, -3, 5, 14, -18, -35, -35, 29, -6, 28, -57, -35, -4, 0, 14, 5, -16, -6, 24, 5, -13, -3, 26, -28, 1, 13, 23, -14, 26, -7, 5, 25, 11, -29, -9, 0, 2, 26, 19, 15, -5, 21, -4, -6, 13, 3, 11, 0, -15, 3, 4, 14, -50, 22, -16, 4, 32, 5, -6, -25, 19, -6, 7, -10, 20, 23, -12, -9, 17, 10, -25, -20, -5, 66, 0, 15, 1, 15, 55, 2, -24, 3, 7, 3, 17, 28, 10, 11, 10, 0, -30, -30, 2, -23, -25, 13, 7, -7, -4, 10, -27, 6, -5, -3, -24, 13, 2, 0, 5, 18, -35, 0, -2, -22, -20, -8, 26, -16, 14, 29, 41, -13, -15, 1, -37, -2, -7, 7, -8, 16, 32, -4, -16, -15, -19, 36, 4, -13, -6, -6, -48, -8, 0, 28, -11, -3, 12, 17, -25, -11, -3, 4, 3, 5, 9, -22, -16, -1, 7, 21, 25, -45, 2, -49, 26, -7, 14, 10, -10, -9, 3, -13, -8, 0, 10, 0, -42, 1, 16, 11, -31, 28, 2, 4, -27, 3, -15, -20, 22, -6, 1, -12, 14, -3, -18, 40, -23, -17, -32, -45, 12, 48, 3, 26, 12, 1, -23, 16, -39, 4, 1, 27, 68, 21, -8, 0, 35, -19, -37, 31, -8, -10, -5, 21, 0, 0, 0, -34, -31, 0, 0, 3, -22, 13, -2, -17, 5, 65, -13, -28, -1, 1, -37, -32, 0, 42, 2, 31, 36, 26, 4, -19, -5, -10, 8, -5, 43, 0, 77, 23, 3, 17, -40, 16, 4, 7, 17, 45, -29, -15, 56, 34, 5, 23, -15, -11, -3, -11, 33, 17, 1, 16, -34, 17, -74, 41, 6, 2, 19, -2, -20, -18, 22, -14, 10, -5, -1, 5, 0, -14, 26, -9, -13, -3, -23, 4, 3, 7, 56, -15, 8, 2, 67, 0, 28, -11, 4, 2, -5, -18, 2, 15, 35, -47, 2, 13, 0, -65, -33, 8, 8, 48, 16, -30, -26, -26, 2, -20, 0, 8, 4, 7, 2, 10, -9, -7, 14, 10, -3, 12, -17, 11, 1, -8, 12, -55, -35, 16, -2, -7, 14, -18, 0, -27, -5, 23, 14, 23, -2, 0, 0, -76, -10, 33, 11, 15, 42, 8, 9, -28, -8, 14, 1, 2, 27, 16, 20, -36, -7, -38, 58, -7, -6, 6, 0, 3, 1, -8, 39, 13, 21, 32, -11, -69, -3, -7, 11, 41, -5, 30, -20, -28, -16, 23, 2, 57, -3, 25, -37, 16, 0, -31, -7, 0, -3, 8, 0, 20, 23, 0, -1, -2, 1, 3, -22, 15, 10, 1, 24, 4, 58, 4, 19, 28, -61, -1, 4, -4, 14, -4, 9, -58, -11, -18, -16, -39, -14, -65, 0, 67, -15, 6, -11, -34, 37, -4, -5, 6, -68, -23, 28, 16, 6, -3, -25, -21, 0, 10, -17, 5, -2, 0, 2, 32, -11, -15, -1, 1, 15, -10, 1, 16, 2, -12, 25, 16, 0, -1, -25, -27, 0, -2, 8, -19, -91, -21, -28, 0, -34, -30, -6, 7, 26, -3, 1, -6, 15, -6, 61, -4, 1, 10, 44, -14, 22, -6, 3, -27, -1, -7, 3, -27, -16, 3, 17, -44, -5, 23, 24, -10, -29, 19, 6, -36, -7, -1, 3, -29, 1, -29, 8, -7, 3, -62, 4, 1, 0, 25, 5, -3, 0, -1, 18, 9, 29, -33, 24, 7, -37, -1, 17, -7, -18, 1, 0, 5, 17, -23, 9, -13, -1, -6, -9, 17, -30, -5, -6, -38, -40, -22, 24, -24, -24, -25, -6, 0, 28, 19, 45, 38, 6, 0, 9, 1, -1, 9, 12, 15, 6, -9, 7, -8, 9, 0, 0, 1, -21, -9, -2, -6, -3, 8, 43, -9, 2, -31, -16, -16, 7, 9, -27, 18, -3, -38, -45, 14, -33, 1, -9, 7, 22, 0, 1, 25, 0, 9, -18, 37, -5, 26, 22, -10, -2, -7, 14, -4, -26, 16, -34, -32, 10, 12, 4, -2, 7, -12, 17, 7, -16, 27, 6, 6, 29, 11, -14, -1, 18, -24, 3, 10, 0, 12, 5, -2, 18, -29, 23, 1, -20, -4, 3, 6, 25, 5, 45, 6, 5, 5, 42, -14, 2, 6, 1, 10, -25, -17, -41, -14, -7, -15, 9, -2, 40, 29, 7, -7, -5, -19, 30, -8, -3, 3, -1, 3, 17, 34, 9, 24, -3, -13, -18, 7, 0, -16, -2, 5, 2, -2, 4, -27, 1, 50, -5, -5, 3, -4, 3, 12, -6, -25, -50, -39, -1, -42, -20, -1, 19, 28, -34, 24, -6, 28, -24, -22, 2, -32, -1, 0, -12, 18, -2, 46, -11, 20, 13, -37, -3, -1, 13, -6, -61, -14, 32, 16, -4, -20, 14, -2, -17, -8, -25, 7, 7, -2, 1, 9, 25, 23, 3, 59, 3, -79, -11, -38, -23, -20, 22, 11, -16, 48, -5, -23, 26, -42, 1, 5, -30, 4, 26, 16, -25, -18, 2, 6, 36, -4, 5, -43, 21, 0, 6, 34, -6, -11, -26, -31, -2, -13, -22, -25, 67, 51, 5, 5, -8, -10, -22, -49, -29, 61, 0, 37, 19, 26, -13, -10, 12, -12, -38, -7, -4, 19, 0, 5, 8, -2, 36, 48, 18, 59, -6, 2, 9, -5, 0, -27, -3, -36, -31, -71, 6, -77, -57, -29, 26, 6, 0, 4, 5, 39, -43, 20, 25, -18, -9, 6, 16, 7, 2, -25, -27, -14, -24, 10, 0, -9, -43, -3, -58, -2, 11, 19, 18, 12, 53, -22, 5, -5, -53, 11, 5, -27, 5, 44, 4, -15, -3, 45, -30, -41, -9, -12, -18, -59, 56, 33, -8, 17, 3, 29, 24, 7, 39, -6, -10, -6, -9, 19, -12, -32, 4, 3, -9, 0, 22, -16, 31, -5, -6, 27, 48, 27, 9, 7, 6, -6, -13, -40, -2, 51, -3, 11, -34, 16, -40, 3, 7, 11, -6, -10, -4, -8, 38, 2, 1, -2, -84, 27, 0, -38, -1, 2, 0, -8, 11, -19, 6, 43, 3, 4, -29, -25, 0, 19, 3, -5, -25, -9, 2, -71, -41, -1, 21, 7, -5, 4, -8, 46, -20, -21, -31, -18, -8, 7, 2, -8, 37, 50, -16, -20, -36, -16, -8, -3, 10, -14, -32, 0, 1, 28, -5, 20, 10, -5, 22, -11, 14, 0, -5, -40, 3, 4, 0, 3, 2, 43, 30, -54, 21, 22, -2, -41, 36, 25, -6, 9, 0, -6, 7, -15, -19, -6, -18, -4, -7, 11, -17, -38, 26, 2, 6, -5, 23, -25, 44, -4, -4, -16, 25, -18, -2, 14, -15, -3, -38, -47, 11, 38, 8, 20, -8, -29, -16, -21, -8, 0, -5, -12, 11, 31, 20, 20, 4, 7, -9, -11, 8, -34, 27, 18, 3, 3, -32, -17, -3, -32, -2, -8, -7, -16, 4, -26, 2, 19, -31, -70, 4, -13, -7, -53, 0, 33, -41, 4, 47, -2, -20, -36, -9, -48, 3, 8, -17, -1, 28, -13, -15, 0, 0, 0, -6, 34, -22, 20, -36, 4, 21, 13, -3, 21, -15, -33, -17, 22, 39, 11, -1, 14, -1, 0, -3, 9, -1, 17, 7, -60, -4, -19, 19, -38, 17, 20, 9, -6, -7, -8, -6, -54, -29, -5, -20, -5, -24, 10, -5, -40, 21, 1, 36, -2, 28, -48, 7, 5, 3, 1, -2, 4, -15, -10, -23, -21, -23, 3, 4, -11, -3, 44, 20, -3, -40, -61, -5, -8, 1, -6, 8, 26, 23, 29, -28, 6, 22, 35, 0, 28, 1, 14, 1, 4, -1, -12, -19, 56, -3, -5, -35, -11, -5, 35, -5, 30, -13, -30, 3, 9, 26, -61, 4, 2, -21, -11, 15, -36, 24, -26, -6, -15, 3, 7, 47, -4, 7, 18, -35, -4, 2, -4, -6, 12, 26, 5, 23, 9, 0, -5, -3, 43, -18, -36, 40, 5, -12, 12, -3, -18, 0, 8, -14, 47, 7, 8, 11, -12, -42, -7, -13, -16, -24, 3, 1, -1, 2, 39, -19, -33, -17, -1, -32, -5, -9, 18, -38, -45, 11, -4, -28, 5, 12, 8, -20, -7, 0, -1, -17, 2, 28, -59, 5, -17, -1, 30, -10, -20, 5, 33, 4, -20, -69, -36, -15, -10, 0, 7, -10, 28, 26, 24, 2, 0, -22, 43, -8, -7, -20, 5, -5, -6, -11, 24, 0, -53, 3, 0, -5, -12, 5, -6, 0, 6, 9, -30, 7, 0, 9, -12, -3, 9, -10, -6, -60, 39, -6, -10, -44, -18, -3, 0, 3, 25, 15, 3, -5, -12, 39, 18, 1, 5, 53, -12, 13, 4, -1, 5, 19, 6, 10, -10, -14, 10, -14, -11, 0, -7, 21, 23, 25, 26, -4, -33, -19, -5, -11, -24, 20, -49, 3, -40, -7, -5, -5, 7, 10, -11, -9, -4, -1, -7, 46, 15, 40, -3, -3, 1, 22, -7, 30, 34, -1, -2, 5, 0, 34, -4, 16, -34, 34, -15, -12, 33, 13, -11, 2, -5, -6, 8, 63, -29, -31, -7, -7, -1, -14, 5, 7, 16, -3, 6, 6, 20, -1, -9, 3, 14, 3, -8, 11, -20, 1, 18, -1, 5, -10, -12, 1, 15, -5, 12, 31, -32, 1, 14, -1, -16, -9, -20, -71, 0, -1, -50, -20, -22, -45, -35, -2, -11, 21, 7, 0, 11, -22, -17, 9, 47, 3, -12, 15, -25, -15, -7, -6, 19, 42, 16, -12, -4, -5, -6, 3, 0, 4, 3, -4, 6, -47, -11, 1, -14, -2, 19, -17, 0, -20, 6, 13, -22, -11, 12, -2, -1, 11, -9, 1, 6, -17, 5, -1, 6, 33, 5, 34, 7, -9, -7, 41, -7, 0, -1, -5, -28, 17, -15, 15, -37, 4, -8, 13, 9, -5, -50, 7, -3, 12, -24, 6, 18, -11, 5, -4, 47, 13, 16, 5, 32, 16, 9, -2, -47, 1, 10, -11, 9, -5, -9, -6, -45, 26, 64, -1, -5, -48, -7, -3, 7, 0, 8, -38, -55, 1, -5, -26, -25, 15, 18, -78, -16, -13, -49, 24, -45, 16, -57, 2, 2, -27, 32, -7, 1, -27, 6, 44, 2, 4, 48, 10, -1, -66, 0, 18, -7, -1, 22, -8, -10, 15, -20, 22, -5, 0, -17, -10, 13, -14, 16, 0, -15, -9, -13, -34, -2, -41, -11, 28, -28, -19, 20, -1, 11, -3, -20, -26, 3, -25, -4, -15, 14, -36, -67, 5, -2, 26, -4, 9, -36, 17, 0, 2, 11, 45, -21, -21, -12, 4, 21, 1, -57, 13, -28, 0, 26, 15, 17, -32, 23, 15, 2, -1, -6, 62, 19, 9, -8, -31, 21, -33, 8, -8, -11, -10, 4, 1, -7, -26, 32, 24, 20, -3, -2, 15, -16, -6, -34, -14, 28, -36, -67, -7, -19, -39, 14, 33, 15, -13, -4, 15, -24, 0, -47, 10, -11, -3, 4, 33, 5, -8, -11, -15, -51, -16, -32, -1, -4, -40, -16, -58, -3, 4, 0, -14, 7, -4, 21, 9, 29, -10, -6, 3, -32, -6, 27, -9, -20, -3, -29, -28, -19, 16, 9, 15, -22, 12, 9, 8, 33, 3, -9, 9, 12, -9, -4, 18, -2, 2, 8, 0, -23, 11, 6, -51, 3, 8, -41, 40, 7, -5, -49, 27, 14, 1, 37, 7, 27, 6, -34, 13, 5, -5, 14, -9, 15, -21, -5, -6, -4, 3, 4, 12, -37, 36, 19, -18, 22, -29, -5, -3, -56, 17, 0, -3, -16, -10, -1, 2, 23, -4, -3, 16, -18, 2, -16, -7, -6, -37, -27, -3, -13, 8, -22, 27, -31, 1, -14, -9, 39, -8, -41, -8, -15, 6, 1, 6, 13, -27, -12, -16, -30, 45, -51, 3, -6, -8, -16, -35, -1, 3, -1, -22, 0, 3, -3, 0, 22, -18, -47, 5, -30, 27, -26, -4, -19, -3, -1, -7, 0, -8, -23, 4, -32, 2, 0, -3, -8, 2, 13, 5, -30, -1, -1, -8, 0, -35, 15, -18, -27, -11, -6, -9, -7, 14, -23, 32, 5, -6, -60, -27, -8, 5, 50, -28, -29, -37, 8, 9, 38, 7, -17, 20, -18, -1, 9, -37, -11, 4, -30, -16, 12, 38, -8, 12, 13, -27, 11, -1, -46, 20, 6, -2, -3, -10, -37, -3, -5, -3, -5, -47, -7, 2, 23, -3, 4, -17, -26, -7, -6, 10, -40, 14, -46, 13, 27, -17, -48, 1, -30, -7, -27, -2, 1, -14, 15, 34, 9, -2, -33, 15, 23, 5, 0, -29, -1, -4, 2, -1, 8, 4, 16, -26, -13, -5, 39, 22, 14, -1, -6, -21, -13, 2, -4, -2, 24, 22, 4, -22, -64, 2, -26, 12, -43, 5, 0, 7, -37, 14, -25, -8, 6, -43, -3, -22, 2, -14, -33, 4, -2, 26, -1, 29, -20, -2, -4, 5, 17, -11, 7, -39, 25, 2, -20, -12, 28, 16, 27, 0, 14, 29, 0, 2, -43, 7, -20, 0, 5, -16, 8, 14, 44, 11, 6, -7, -72, -4, -16, 11, 2, 4, -13, -2, 6, -6, 24, 8, -4, -13, 8, -6, 3, -1, -7, -21, 0, -3, 12, 23, -64, -4, -16, 31, 24, 7, -88, 2, -41, -72, 11, -9, 12, 0, 14, 35, 8, -31, -30, -26, 41, 3, -15, 20, -23, 23, 4, 10, 4, 21, 15, 15, -12, 21, -28, 15, 16, -7, -7, -31, -16, 32, 62, -3, -4, 46, 24, -2, -3, 13, -11, 0, -2, 1, 12, -5, 16, -9, -15, 13, -1, -31, 6, 16, 20, 0, -13, 5, 2, 40, 5, 31, 16, -19, 1, -3, 9, -1, -19, 9, -41, 10, -1, -5, -15, -6, 1, -5, 3, 9, 30, 13, -26, 7, -17, -8, -9, -27, -17, 34, -4, -15, 0, 23, -4, -4, 41, 4, 9, 7, -3, 9, -12, 5, 3, 3, 1, -51, -25, -1, -20, -4, 30, 12, 18, 7, 7, 27, -33, -34, -7, 14, -2, -20, 33, 13, -20, 62, 0, 0, -5, -7, -3, 32, 16, -36, -7, -34, 22, -3, -19, 55, 1, -12, 3, 25, 5, 14, 11, 51, -4, -21, 20, 3, 0, -3, -13, -26, 7, -67, 8, -5, 23, 48, 11, 40, 10, -3, -12, -34, -6, -14, -25, -4, 4, -6, -26, 13, -2, -17, -2, -6, 13, 38, 4, -12, -5, 32, 1, 37, -4, -23, 1, -6, -11, 4, -19, 25, -11, 28, -28, 5, 1, 18, -4, -4, 19, 46, 26, -1, -40, 28, 14, 0, -4, 6, -10, 0, 24, 14, -2, 73, 25, 0, 8, -3, 13, 0, -4, 1, -30, -14, -5, -4, -9, -29, -21, -7, 4, 5, 54, -16, -18, -7, 12, 10, -37, -43, 7, -24, -17, -36, -44, -7, -45, -9, -10, -2, -6, -19, -1, 57, 17, -15, 11, 15, 17, -6, 15, 32, 23, -36, -2, -2, -18, 10, -6, 17, -12, 10, 8, 31, -26, 0, -31, -36, -17, -18, 12, 4, 25, 8, -13, 36, -1, -20, -3, -7, 42, -14, -8, -1, -14, 4, 10, 12, -6, -35, -7, -4, 10, -6, 11, -16, 6, 43, 2, 7, -29, 0, 7, -2, -14, -10, 13, 19, -20, 16, 0, 26, 41, -6, -5, 8, 54, 17, 16, -66, -9, 17, -22, 2, -3, 16, 8, -12, -7, 22, -5, 16, 14, -8, -10, -33, 10, -3, -1, -10, -24, 15, 13, 9, -3, -16, 0, 5, -14, -5, 24, 6, 22, -2, -17, 18, 17, -14, 9, -48, -11, -34, -24, 10, -3, 12, -40, -2, -4, 0, -28, 19, 15, -22, -4, -7, 21, -8, -5, -20, 0, -15, -7, -11, -29, 12, 10, -1, 16, -14, 2, -4, 9, 2, 12, 6, -7, 2, -23, -1, -9, -43, -35, 39, -2, -14, 20, -3, -24, -23, 0, -6, 0, -12, -29, -9, -3, -5, -2, 1, 13, 8, -27, -3, 1, -6, 3, 8, -12, 14, 7, -7, -10, 24, -8, 27, -3, 26, 16, 14, 10, 1, -22, 6, 58, 13, 9, 34, -25, 21, 8, -11, -20, 44, -7, 21, 18, -17, 5, 22, 37, -3, -19, -41, 1, -4, 1, 25, -14, 8, 24, 0, -5, -6, 0, 3, 8, -5, 21, 2, 14, 0, 12, -39, 30, 10, -13, -9, -18, 13, -24, 19, -22, 10, -16, -5, 0, -18, 0, -29, -2, -43, -9, -32, 16, 2, 5, 53, -19, -5, 3, -20, 0, 15, 19, -28, 11, 4, 9, 13, -1, 0, -22, 0, -4, 20, 6, -4, -8, -41, -29, 57, 22, 2, -3, 2, -4, -14, 3, 0, -4, -9, 11, -26, -6, -12, 4, 2, -1, 34, 4, 2, -5, 41, 6, 10, -36, 26, -4, -10, -26, 5, 19, 9, 68, 35, 30, -21, -3, 27, 15, 2, 16, 19, 23, 5, 0, -8, 7, 0, 35, -24, -26, 12, -1, 6, -16, 17, -9, 2, 35, -33, 3, -7, -2, -12, 43, -25, -10, -2, 4, -9, -9, -1, -3, -3, -3, 30, 4, 7, 3, -10, -10, 18, -11, -12, 31, -39, 8, 0, -3, -36, -10, 0, -7, -10, -9, -66, 2, 35, 0, 17, 6, 4, -25, 46, 8, 17, -10, 16, 0, 23, 0, -10, -3, -30, 2, -4, -14, -2, -19, 8, 3, -14, 20, 11, -9, -33, 37, -10, -2, 15, -1, 19, -23, -4, 11, -4, 13, 19, 28, 27, -7, 14, 0, 0, 5, -1, 53, 28, 3, -21, -5, 0, 1, 6, -6, 2, 5, 8, 5, 48, 45, 25, -11, -11, 1, -40, 5, 0, -1, -4, 29, 59, 26, -11, 9, 5, -10, -56, -27, 19, -1, 8, -4, -3, 29, 7, 28, -11, 9, 6, -7, 2, -9, 20, 34, -6, 2, -5, -21, 7, -5, -5, -1, -9, -16, 2, 16, 10, -21, 9, -40, 28, 4, -2, -53, 28, -28, -33, 18, 3, -1, 30, 10, -57, 19, -32, -37, 25, 8, 5, -45, -17, -20, -11, -17, 32, -4, -2, 11, 0, 8, -2, 3, -18, -15, -5, -66, 27, 24, -20, -16, 6, 54, 3, -28, -42, 4, -16, -47, 18, -18, -4, -14, 7, -21, 0, -12, 8, 1, -14, 6, -6, 5, -13, 12, 26, 0, 6, 4, 12, -14, 41, 5, 2, 6, -11, -7, -22, 50, 43, -4, 26, 21, -29, -3, -5, 4, 6, -6, -12, -1, -37, -11, 4, -1, -74, -1, 33, 24, 0, -10, -15, -32, -5, -2, -27, 12, -2, -2, 35, 23, 9, 71, 5, 6, -21, -18, -6, -10, -4, -47, 20, -27, -6, -17, 35, -60, 16, -86, 41, 42, 30, -43, -17, 1, -49, 15, -5, 9, -17, 14, 27, 41, -20, -43, 58, 14, 0, 3, -63, -1, 13, -1, -21, -5, 1, -25, 26, -12, -19, -21, 20, -57, -5, -13, -20, 0, 29, -15, 0, 26, 31, 31, -29, 20, 24, 6, -16, 25, -14, -31, -2, 4, 14, 11, 28, 2, 4, 6, -5, 5, -22, 8, 14, -4, 5, -7, 26, 24, 4, 5, -2, 13, 9, 12, 3, 29, 18, 1, -41, 27, 15, 18, 6, -39, -24, 0, 5, 7, -30, -10, -6, -23, 20, -25, -14, -8, -4, -3, -5, -41, 1, 40, -4, 9, -9, 0, -2, -14, -14, -26, 6, -7, -17, -8, 3, 0, -6, -5, 0, -12, -4, -9, 2, -1, -34, -1, -21, 1, -4, -5, -6, -61, 17, 11, 0, -3, -23, -17, -46, 19, -91, -24, 52, 9, -1, 23, -21, -49, 7, -4, 1, -16, -6, 17, 25, 3, -29, 44, 23, 14, -6, -16, -57, -8, -63, 10, -3, 33, 4, -4, 21, -2, 15, -12, -62, -47, -13, 5, 1, 10, -9, 2, -6, -5, -40, 5, -27, 9, 21, 22, -49, -4, 8, -1, -2, -1, -20, 4, 0, -3, 24, 0, 11, -13, 19, 13, -6, -7, 6, 8, 4, 27, 23, 13, -34, -11, -32, -10, -1, 6, 27, 3, 6, -4, 20, -5, 48, 4, 0, -8, 0, 12, -4, -7, -15, -5, -22, -21, 3, -6, -34, -14, 5, -39, -6, 19, 9, 23, 0, 11, -13, -26, 0, 1, 1, -3, 11, -38, -1, -67, -5, -17, 0, 3, -20, -12, 22, -3, -33, 2, 36, 20, -8, 16, 5, 6, -15, -3, -1, 0, -4, -8, 16, 0, -38, -4, 28, -14, -1, 25, -89, 12, -24, -2, 3, -32, -26, 12, 35, -20, 4, 1, -6, -10, -4, 12, -5, 16, -9, -20, -6, 0, -42, 3, 4, -3, 38, -26, -17, 6, -9, 5, 8, -14, -14, 7, 0, 0, 0, 5, 30, -8, 25, 12, -10, -1, -6, 16, 5, 39, -1, 28, -18, -9, 1, 9, 4, -7, 18, -42, -20, 5, 2, 0, 15, -26, 4, 0, 1, 8, 7, -12, 1, 2, -21, -29, -2, 1, 26, -15, -3, -8, -8, 30, 0, 2, 5, 29, -23, -10, -20, -26, 9, -7, 7, 10, 13, -22, 20, -6, -5, -5, -6, -13, 17, -10, -46, 24, 2, 46, -8, -24, 40, -8, -10, -1, 11, -14, -1, -11, 3, 18, -5, -6, 44, 27, -4, 18, -9, 26, 0, 10, -3, 9, -22, -15, 20, 38, -1, 22, -14, 21, -24, 13, 6, -14, -9, 8, 2, 1, -42, 1, 3, 8, 8, -25, -9, 2, -28, 1, 15, 3, 39, 2, -3, 7, 40, 12, 21, 14, 30, 41, -5, 15, -47, -26, 2, 61, 33, 25, -63, -10, -26, 17, -3, -27, 45, -11, -39, -25, -13, 1, -13, 26, 2, -40, 3, 16, -4, -5, -8, -16, -1, -56, 0, 4, 21, -5, -10, -3, -1, -18, -4, 5, 6, 47, -20, 2, -17, -3, -8, 8, 4, -1, 30, -8, -44, -7, -9, 5, -35, -10, -2, 4, -28, -5, 22, 14, -2, 27, 36, -37, 11, 10, -1, 14, -17, -24, 7, 8, -20, -16, 24, -2, -4, 48, 25, 6, -16, -13, 5, 51, -36, -31, 23, 13, -4, 6, -9, 46, 1, 2, 4, 35, -11, 2, 7, -3, -2, -8, 38, 2, 11, -15, -20, -6, 40, 2, -11, -3, 13, -2, -4, -6, 8, 64, 35, 14, 31, 47, -25, -3, -7, -23, -1, 13, 0, 18, 16, 0, -2, 9, -1, -1, -38, -32, 9, 0, 16, 1, 0, 31, -6, 27, -8, 11, -4, -8, 3, -43, 17, -27, -7, 4, 7, 3, 0, 1, -6, 35, 32, 32, 0, 35, -30, -4, -1, -30, 3, 17, 15, -18, 1, -17, -34, -18, -8, -3, 1, 27, -35, 0, -8, -22, 43, 3, 2, 0, 6, 8, 10, 1, 1, 8, 0, -15, -31, -6, 20, -26, 19, -32, 3, -12, 49, 1, -53, 0, -3, 47, -5, -8, 12, 7, -11, -32, 19, 17, -9, 17, -7, 9, -23, -10, -8, -4, -36, 4, 39, 4, 29, -19, 4, 3, 41, -4, -2, -2, 12, 1, 3, 15, 6, 24, 6, -11, -1, 43, -14, 7, 0, 14, -5, 0, -2, 20, 1, 17, -20, 7, 3, -7, -44, -27, 8, 3, 22, 1, -1, 28, -3, 35, -16, 5, -3, -4, 25, -5, 10, -29, 2, -2, -6, -15, -5, -7, 0, -36, 7, 36, -2, -3, -7, -15, 1, -37, 48, -10, -14, -25, -15, 4, -8, 6, 1, 7, -20, 19, -16, 14, -29, -21, 19, 9, -5, -10, 3, 9, 16, 0, -16, 0, -37, -34, 1, 28, -24, -15, 8, -41, -2, -9, 26, 28, 6, -35, 5, 23, -4, 2, 19, -13, -1, -3, -22, -16, -11, 1, 1, 1, -10, -6, 39, 0, -36, 1, -5, 10, 24, -24, -15, 5, 49, 7, 13, 21, 11, 0, 5, 8, -6, 10, -12, 60, 6, -4, 1, 45, -28, 13, -2, -17, -34, 15, 5, 34, 1, -9, -6, -17, -48, 9, 44, -6, -9, -4, 37, -42, 0, 9, -19, 14, 4, 1, 18, -8, 42, 72, -7, 5, -15, -1, -4, -14, 6, -101, 40, 26, 6, -10, 7, -32, -31, -68, 70, 5, 21, -17, 6, 13, -12, 4, 0, 8, 6, -14, 31, 28, -42, -66, 26, 22, 4, -21, -60, 6, 2, -4, -33, -8, -10, 1, 10, -25, -40, -10, -4, -35, -3, -49, 45, -16, 32, -21, 0, -88, -3, 43, -14, -19, 24, 10, -12, -22, -19, 9, -5, -2, -29, -6, 16, -6, 1, 6, 13, 21, 27, -3, 15, 2, -21, 2, 42, 2, -15, 4, -2, 23, 19, -32, -5, -2, 3, 10, 0, 32, 19, -11, -1, -41, 6, -3, -14, 12, -63,
    -- layer=2 filter=0 channel=1
    -26, 6, -11, 21, 4, 40, 38, -16, 5, 32, 11, -2, 39, 19, -12, 0, 3, 0, -9, -17, 4, -4, 0, -5, -8, -3, 33, 6, -4, 44, 23, 3, 1, -11, 19, -28, -24, 26, 0, -15, -8, 0, 19, 7, 26, -3, -2, -17, -13, -51, 8, -2, -19, -18, 3, -9, 17, 11, -18, 25, -1, 25, -19, -10, 30, -1, 1, -3, -27, -20, 39, -2, 5, 1, -13, 0, 0, 2, 2, 14, 33, 32, 66, -16, -9, -22, 14, 12, 4, 6, -9, -6, 14, -25, 1, -2, -9, -8, -1, 31, 15, 42, 3, -3, -1, -11, 12, 2, -6, 4, -11, 0, -25, 32, 1, 0, -10, 34, 23, 0, -28, 0, 0, 49, -9, -36, 13, 36, -15, -8, 0, 15, 7, 16, 2, -14, 8, 12, -48, -2, 18, -14, -10, -2, 3, 19, 14, -17, 17, -2, 0, -5, 1, 2, -2, -1, 1, 5, 36, -1, 5, -2, -10, -21, 1, -18, -35, -12, 0, -2, 23, 6, 17, 2, 5, 7, -6, -35, 5, -21, 4, 21, -25, 7, 22, 0, 2, 10, 0, -2, 7, 0, -3, -16, -2, -30, 5, -42, 20, -6, 16, -31, -1, -45, -17, 2, 0, -14, -19, -3, 12, -30, -1, -39, 11, -3, 16, 0, -5, -22, 10, -6, 0, 23, 0, -10, -11, 26, 39, 10, -3, -10, 0, -12, 7, 0, -6, 4, 14, 32, 10, 40, 1, -5, 0, 16, 2, 3, 1, 5, -13, -19, 7, -36, -4, 16, 1, -6, 18, -20, -18, 4, 9, 5, 13, 24, -1, 0, 25, 0, -6, 3, 3, -16, -27, -1, 34, -2, 0, -9, 10, -3, -25, -2, 24, 37, 48, -6, -26, -5, -11, -17, 17, 8, 2, -8, -40, 7, 0, 66, 28, 2, 8, -22, -23, 18, 0, -12, 4, -90, 9, -2, 46, 36, -8, 8, 7, 17, 11, 5, -4, 1, 12, 18, 1, -2, 11, -8, -33, -13, 3, -37, 22, -3, -36, 9, 29, -2, 31, 13, 2, 9, -46, -6, 32, -3, -10, 18, -2, -11, 0, 0, 4, -23, 1, 12, 20, 8, 4, -8, 2, 15, -19, -3, -3, 5, 14, 26, 5, 57, 3, 6, -28, 17, -24, 21, 22, -5, 5, 2, -28, 10, 0, 43, 2, -2, 33, -6, -19, 16, 58, -10, 2, 17, 3, 2, 19, -9, -6, -3, -9, -14, -4, 7, 22, 7, 1, 11, 8, -4, -3, -5, 41, 31, -9, 4, -11, -2, 16, 6, -1, -22, -22, -24, 0, -6, -22, 13, 26, 3, 4, -32, -4, 0, -33, -11, -1, -51, -8, 6, 9, -25, 37, 4, 8, 35, -4, 16, 27, -26, 14, 0, -29, -11, 11, -2, -25, -12, 9, 6, 9, -8, 17, 3, 3, 4, 7, -29, -13, 31, -42, -8, -6, -5, 2, 7, -21, -4, 1, -38, -4, -46, 0, -9, 9, 17, 0, -11, -2, 5, -10, -4, -5, 2, 18, -8, -14, -13, -1, -12, -41, 5, -9, -44, 23, 0, 12, 13, -37, 6, -24, -14, -9, 0, 9, -53, 22, 31, 10, -14, 12, 32, -10, -5, 16, -4, -2, -3, 0, 8, -29, -8, -42, -2, -3, 0, 8, -2, 19, 2, -33, 15, -8, -3, -18, 2, 39, 29, -19, -25, -11, -35, 5, -2, 31, -14, 12, -8, 0, 1, 11, -9, 8, 28, 2, 19, 8, 3, 50, 4, -11, -41, 6, 22, 0, 22, -6, -2, -15, 4, -12, -31, -20, -6, -31, 19, 22, 10, -4, -8, -87, 0, 22, 17, 5, 16, -9, 29, 40, -5, -2, -6, -25, -3, -18, -12, -2, -4, 2, -10, -10, 29, 28, 46, 3, -21, 0, -9, -6, -14, -6, -2, -25, 2, -6, 35, 16, -1, -18, -19, 1, 12, 13, -5, -17, 4, -18, -6, -18, 4, -15, -1, -10, -40, 18, 7, -6, -18, -3, 27, 30, -9, 24, -11, -11, 0, -3, 11, 4, -36, -55, 5, 2, -7, 16, -8, -7, 4, -37, -8, 12, 4, -10, 11, -36, 16, 7, -35, 0, -23, -3, 8, 22, 64, 13, 3, 8, 0, -3, 29, 8, 11, 17, -3, 0, -4, 13, -3, 39, -10, -1, 0, -1, 5, -23, 4, -34, -17, -2, -38, -12, 0, -6, -6, -18, -6, -14, -3, -17, -19, 32, -4, 33, -4, -5, 2, -2, -2, 1, -11, -14, -5, 1, -28, 3, 1, -5, 0, -8, 0, 17, 25, 5, 20, 7, -15, 5, -1, -2, 0, 3, 25, -10, 20, 16, 18, -37, 25, 11, 32, -7, 7, -32, 3, -21, 23, -5, 3, -22, 2, 1, 17, 19, 29, 19, -28, 1, 12, -39, -5, 37, -5, -7, -8, 4, -4, -31, 4, 36, -1, 8, -16, 7, 2, 12, 5, -30, -9, -26, -6, -2, 4, 4, -29, 13, -47, -11, 28, -9, -17, 11, 38, 0, 5, 3, 25, 14, 34, 0, 18, -2, -9, -11, 7, 29, 17, 32, -11, 5, 28, -25, -24, 2, 16, 2, 12, 3, 5, 6, 3, 22, -29, -20, -28, 19, -9, -9, 21, 26, -20, 13, -9, -13, -28, 13, -8, -25, -8, -35, -3, -9, -40, 5, -2, 5, 16, 7, -37, -19, 27, 4, -2, 1, 19, 0, -9, -1, -1, -9, -6, -23, 44, -15, -23, -37, 68, 56, 42, 29, -4, -34, 23, 12, -12, -14, 24, -13, -3, -18, -25, 29, 5, -11, -17, 4, 11, -33, 2, -19, 4, -10, 3, -3, -17, -21, 5, -50, -6, -5, -34, 0, 1, -16, -3, -32, 10, 0, -1, 1, 0, -7, -29, 5, -17, -2, 11, -34, 5, -4, 0, -5, -2, -8, 21, 2, -28, -3, -21, -42, 29, 13, -6, 29, 48, -9, 15, -1, 20, -9, -9, -18, 17, 7, -21, 13, -5, -3, 2, 13, -18, 16, -37, 11, -4, 17, 11, 8, 2, -14, 13, 10, -27, -17, 7, -4, -6, -7, 6, -28, -14, -7, -49, -5, 13, -6, -2, 11, -9, 1, -5, 1, 0, -23, 0, -6, -6, 15, 23, -21, 9, -21, 23, -22, 18, 5, 47, 4, 1, 13, 8, 13, 15, 3, 8, -1, 0, -5, 6, -5, 11, -4, -5, -2, -14, -5, 4, -15, -9, -19, 4, -5, -10, -3, -5, -18, 8, -5, 0, -1, 0, 9, -3, -9, -37, -33, 6, 13, -10, -10, 0, 8, -33, -21, 7, -6, -9, -20, 36, -9, -9, -4, 7, 12, -35, 19, -10, -45, -43, -33, 1, -12, 14, -1, 3, 7, -26, 1, -14, -13, 8, 1, 28, 8, 3, 10, 0, 2, -22, 22, -41, -25, -4, 5, -11, 9, 14, 14, -21, 2, -37, -22, -8, 3, -6, -12, 2, -8, 9, -2, 4, -9, -31, -6, -29, 14, 8, -4, -11, 6, -20, -19, 0, -2, -8, -6, 31, 27, 13, -3, 0, 11, 7, 7, -20, -4, 4, -2, 16, -6, 25, 5, 14, -1, -8, -15, 20, 2, -15, 8, -8, -7, -22, 2, 0, -20, -28, -3, 2, 4, -28, -13, -4, 11, 2, 7, -28, 7, 3, -54, -6, -4, 17, 0, 0, 6, -29, -4, -3, -8, -60, -22, -3, -32, -11, 25, 0, 5, -5, 7, 12, -11, 5, -2, 5, -2, 60, -13, 9, 1, -3, 16, -22, 1, -4, 17, -28, 3, 13, -24, 54, -27, -5, -13, 2, -15, -29, 12, -47, 8, -5, 13, -13, 13, 14, 3, -33, -18, 11, -64, 0, -36, 1, 22, -5, 24, 5, 3, -29, 4, -15, 3, 14, 0, 3, 5, -12, -4, -1, -32, 14, 5, 4, -15, 25, 15, -24, -13, -12, -1, 11, -32, -29, -41, 1, 4, 19, 0, -10, 37, 39, 6, -2, 21, 9, 0, 1, 6, -27, -5, -32, 27, -3, -1, -26, -12, -6, -7, -14, -9, 6, 10, 3, 6, -18, -12, 2, -18, 0, -27, 10, -28, 4, -10, -33, -41, 27, 9, -44, -4, 3, -9, -9, 6, 3, -29, 2, -4, 23, -8, -20, 31, 11, -4, 5, 5, -4, -17, 16, 24, -32, 3, -7, 19, 8, 1, -17, -2, 40, -26, -28, -7, 3, -39, -5, 31, -47, -16, -2, -88, -10, -13, 22, 30, -23, -26, 18, -32, 9, 20, 7, 23, 20, -43, 6, -6, 12, -1, -10, -12, 0, -2, -11, 5, 21, -6, 28, -59, 19, 0, 1, -5, 29, -6, -23, 3, -18, -23, -25, -7, -31, -9, 6, 0, -15, -17, -11, 6, 0, 20, -6, 23, -19, 1, 32, 25, 4, -8, -18, -6, 6, -13, -18, -4, -9, 0, 13, 28, 9, -26, 3, -7, -1, -9, -2, -23, -6, -5, 0, -22, 0, 22, -14, -14, 32, -10, -15, 0, -33, -49, -10, 4, 1, -5, -7, 1, 13, 33, -35, 41, 5, 3, 15, 19, -10, -41, 0, -16, 4, 2, -8, 19, 20, 7, 21, -8, 24, -9, -4, -6, 3, 18, 9, 13, 0, -29, -6, -65, -14, -8, 0, 4, -16, -10, 18, 23, 7, 34, 0, 7, 10, -35, 13, -7, 5, -2, 1, -14, -18, -2, 4, 1, -16, -7, 1, -36, 0, 2, 2, 5, 44, 4, -34, -6, 8, -10, 15, -7, 1, 0, 2, -1, 1, 41, -34, 40, -26, 11, 6, 3, 20, 24, 31, 21, -12, 1, -21, 14, 1, 5, -33, -1, 0, 3, -3, -10, 4, 16, -9, 3, -6, -2, 5, -10, 1, -39, -4, 6, 7, 13, -7, 9, 37, 11, -5, -2, -17, -49, 15, 1, -9, 12, -14, 1, -24, 20, 15, -6, 13, -4, -7, -2, 9, 32, -16, 29, 19, 8, 0, 5, 32, 0, -19, -4, -6, -20, 4, -19, 0, 35, 5, -6, -15, 16, 3, -40, 0, -22, 21, 3, 8, -9, 23, -23, -7, 4, -5, -26, -10, 7, 3, 1, 0, 2, -15, 0, 16, -11, -6, -5, 53, 0, 0, -35, 0, -1, 1, 15, 31, 15, 0, 19, 19, 13, -16, 9, 4, -5, -7, -18, 16, -26, 19, 12, 15, -5, 0, 9, 14, 10, 9, 20, -12, 0, 0, 12, 0, -4, -28, -5, -4, 2, 4, -35, 15, 11, 2, 1, -3, 3, -8, 2, 2, -35, 16, 11, -2, 21, 17, 12, -17, 9, 12, -13, 34, -32, 0, -12, -11, 2, -13, -8, 25, 2, 8, 0, -15, -15, 21, -31, 0, 11, -4, 1, 16, -3, 27, 0, 15, 5, 6, 0, 6, 8, -5, 36, 0, 47, 0, -32, -23, -16, -7, 16, 0, -10, -32, 24, -2, 1, -14, -48, 5, -31, 1, -27, -39, -2, -9, 7, 1, -3, -27, -6, -32, 11, 33, -6, -20, -3, -6, 23, -5, -7, -3, 6, 29, 0, 28, -28, 24, -1, 33, 1, 29, -18, 5, -4, -7, 10, 39, 2, 33, -21, 2, 17, -8, 33, 0, -18, -13, 3, 28, -16, -2, 3, 17, -21, 0, -1, 2, -15, 38, -1, -2, 4, -50, -23, 2, -16, -4, -9, 15, 33, -3, 16, -23, 5, -24, 10, 3, -34, -3, -28, 12, -14, -17, -11, -2, 4, 7, -14, -7, -14, -14, -57, 11, 10, -7, -7, 24, -6, 11, 1, 39, 12, -10, 3, -4, -36, -10, -23, 11, 9, 5, 37, -18, -14, -28, -15, 2, 16, 10, 15, -4, -29, -18, -5, -30, -51, 13, -7, -1, 20, -39, -12, -3, -4, -22, 6, 7, -2, 21, -1, -6, -1, 9, -4, -27, -6, -8, 0, -5, -16, 21, -19, -31, 19, -6, 7, 13, 5, 10, -4, 7, 3, 39, -8, 12, 28, 48, 0, -1, 29, -5, 29, -13, 35, -17, 3, 9, -40, -5, 3, -3, -13, 2, -3, 1, 21, 28, -17, -4, -2, -40, -17, 2, 11, 4, -20, 40, 64, -2, -19, -20, 22, 1, 14, -3, -17, 25, -7, 11, -30, 16, -22, 0, 0, 3, -5, 14, 18, -62, 1, -29, -1, 0, 18, -1, 4, 31, -1, 10, 17, -7, 0, -6, 18, -26, -8, 11, 2, 3, 30, -6, 28, -56, -7, -4, -18, 20, 9, 0, -24, -13, -12, 12, -54, 6, 19, 0, 29, -13, -4, -12, 0, -25, -4, 2, -1, 14, 12, 4, -3, 9, 4, 7, 15, 31, -2, 5, -43, 11, -17, 14, 23, -34, 33, -14, -16, 17, -7, -2, -34, 31, 0, -37, 29, 28, 25, 2, -4, -10, 6, -37, 35, 13, 6, -16, -68, -4, -22, -6, -5, -3, 2, -3, 40, -5, 0, -2, 6, -46, -2, 3, -28, 5, -15, -15, 23, 2, -20, -37, 3, 13, -3, -12, -2, 19, -18, -17, -16, 43, -11, 2, -3, -13, 18, 75, 24, -47, -14, -11, 14, -6, -36, -17, 10, 25, 14, -23, 18, -36, 13, 16, 0, 10, -11, -11, -9, 5, -12, -62, 22, -35, 2, 1, 4, 22, -15, -31, 28, 11, -22, 26, -26, 16, 37, -5, 10, 0, -20, 43, -4, 0, 0, 28, -5, -53, -41, -9, 0, 37, 4, 13, -28, 20, -2, -1, 16, -3, 26, -12, 0, -19, 25, -1, -17, 6, -14, -4, -28, -8, 30, 5, 8, 15, 18, -5, 16, 10, -3, -10, 61, -21, 3, -10, -28, 9, -53, -12, -12, -7, -7, 21, -45, 0, 9, -6, -3, -47, -9, -1, 1, 0, -15, -1, -29, 3, -69, -73, 3, 26, -8, -17, 44, 24, -9, -2, 9, -6, -54, 0, -2, 12, 41, 30, 42, 31, -10, -28, -2, -8, -30, 32, -9, -22, 4, 3, -4, -30, -8, 26, -30, 24, -3, -6, -8, -5, -25, -19, 29, 18, 15, -6, -2, 0, -34, -39, -14, 36, -37, 44, -48, -18, 29, 2, 26, 31, -41, 42, 4, -29, 3, 23, -17, -82, -63, -13, -8, -19, 0, 7, -17, 17, -7, -4, 4, 4, 21, -68, -16, -35, 5, -6, -7, -11, -2, 0, -24, 25, -13, -22, 2, -25, 8, -2, -24, -7, 45, -27, 35, -21, -3, 14, 11, -7, -10, 9, -11, -8, 4, -7, 18, 33, 34, -1, 6, -47, -3, 6, -1, 1, -49, -3, 16, 6, -12, -41, 5, 15, -5, -18, 42, 32, -25, 17, 23, -14, -69, 1, -5, 2, 29, 26, -4, -1, -56, -20, -15, -8, 5, -15, -20, 12, -5, -1, 6, -19, 5, -28, -24, 21, -14, 25, -7, -5, -40, 0, 17, -43, -27, -4, 37, -4, -49, -8, 39, 27, -23, 38, -85, -3, 42, 4, -12, 27, -32, 17, -1, -5, -5, 20, -2, -44, -13, 2, -1, 14, 2, 19, -1, 3, -7, -1, -16, -4, 27, -61, 32, 4, -13, -13, -22, 20, -16, 0, -41, 22, 44, -20, -31, -21, -7, -1, -8, -28, 17, -9, 55, -60, -19, -15, -7, 2, 10, 12, -6, -7, -6, 9, -9, 26, 8, 2, -8, -25, -5, 5, 0, 2, -21, -38, 44, -2, -7, 11, 13, -2, 8, -19, -7, 52, 0, 22, -10, -20, 6, 1, 8, 4, 17, -44, -34, -2, -26, -4, -22, 4, 27, -18, -5, 2, -1, 16, -17, -6, 11, -7, 3, 28, -2, -19, 10, -2, 33, 42, 5, -33, 3, 5, 13, -6, 7, -37, -9, -36, 3, 32, -57, 2, 34, -6, 1, -27, -3, 12, 6, 3, -6, 36, 3, -53, 4, -3, -3, -32, 1, 10, 11, -1, -1, 3, -4, -19, 0, -51, -7, -24, -8, -23, 27, 24, -51, -9, 0, 59, 15, -8, -9, -36, -23, 1, -36, -26, 13, 9, -20, -56, -5, 31, -24, -4, -9, -3, 1, 4, 2, 17, -36, 23, 29, 2, 8, -19, 3, 0, 43, -2, -34, -12, -26, -2, 3, 12, 23, -36, -7, -18, -20, 10, -12, 30, 0, -14, 22, 3, 5, 16, -7, 16, 0, 8, -28, -8, 0, 3, 18, -1, 11, -10, 3, 22, 18, -17, 1, 16, -13, 25, 10, 8, 12, 0, 48, 35, -20, -13, -1, 7, -1, 4, -2, -6, -12, -65, 3, -6, -57, -2, -13, -5, -58, -30, -8, 8, 5, -20, -2, 30, -13, -11, -4, 29, -7, -50, -3, -26, 28, 5, 0, 5, -11, 23, -2, -17, -15, 43, -11, 34, 29, 18, 3, 3, 0, 27, -8, -52, -24, -7, -34, 4, 16, 8, -4, 31, -28, -23, -8, 0, -56, 7, 25, 20, -9, 3, 4, 15, 16, 10, -18, 7, 1, -22, 0, 5, 8, -3, 30, 4, 26, 7, 6, 21, 6, -48, 34, -4, -57, 31, -45, -7, -33, 0, -3, -2, -3, 8, -42, -2, 9, 4, -29, 13, -44, 7, 8, -17, 31, 11, 1, -1, -32, -8, -12, -28, 8, 2, 4, -10, 3, 2, 13, 21, 3, -4, -6, -5, -52, 3, 15, -12, -9, -5, 21, -35, -1, 7, 3, 4, 17, -39, 4, -73, -1, -8, -6, -5, -7, -49, 25, -14, 2, -33, 1, -24, 22, 9, -8, 4, -26, 0, -22, -7, 66, -16, 20, 18, -39, 2, -31, 7, 32, 21, -26, 13, 33, 25, -9, -7, 33, -28, -11, 24, -7, -4, -16, -8, -58, 0, -15, 49, -10, 5, -5, 18, 72, -7, 19, 7, 0, -24, 15, 0, 0, 4, -26, 14, 24, 5, -8, 11, -26, 4, -34, 53, 15, 5, -37, 1, -29, -41, -35, -2, 5, -29, 16, -9, -3, -59, -47, 35, -9, -6, -15, -6, -7, -25, -5, -4, 30, -15, -1, 11, -6, 15, 6, 12, 1, 1, 9, -5, 52, 41, 32, -7, -14, -3, 15, 24, -37, -6, -34, 2, -65, 0, 6, 7, 6, 22, -9, -25, -7, -21, -8, 15, -9, 9, -21, -23, 3, 8, 7, 9, 5, -4, 2, 2, -20, 2, 17, -35, 35, 8, -1, -21, -9, 30, 5, 1, -12, 33, -24, 8, -13, -3, -11, 4, 9, 35, 14, 2, 31, -56, -20, -41, -41, -3, -34, 9, -9, -5, 5, 13, 16, 12, -10, 0, 6, -42, 4, -3, 8, -2, -8, -18, 17, 0, -25, 6, 10, 4, 8, 14, 42, 3, 33, 18, -33, -72, -54, 2, 4, -25, 25, 21, 43, -88, -31, 44, 21, 2, 5, -2, -23, 5, 6, -12, 25, -2, 23, 12, -7, 17, 4, -14, 22, 1, -18, 0, 64, -15, 10, 2, 22, -7, 1, 16, 12, 28, -18, 25, -49, -6, -4, 4, 19, 1, -80, -18, 3, -23, -4, 33, 7, 15, -29, -16, 7, -33, -2, -18, 14, -20, 4, -2, -21, 7, 10, -65, 12, -7, 0, -20, -6, 16, -1, 0, 18, 45, 5, -11, -4, 13, -11, 0, 22, 17, 18, -4, 12, 1, 2, -13, -53, -3, -40, 24, -4, -4, -3, 20, 22, 5, 17, 5, -5, -41, 0, -6, 12, 7, 22, -36, 23, -2, -44, -14, 7, 40, 19, 43, 23, 6, -3, -11, -3, -26, -41, 0, 1, 7, 43, -2, 22, 10, -43, -46, -20, 1, -10, -4, 33, 7, 0, 31, 8, -17, 17, 32, -16, 34, 11, 2, 13, -7, -62, -3, 34, -10, 38, -1, 40, 11, -7, -15, -16, 24, -43, 41, -50, 3, 42, 1, 27, -12, -46, -13, 3, -49, -6, 67, -10, -26, -32, 5, -3, 13, 5, -12, 10, 1, -7, 1, -34, 26, 23, -78, 27, -47, 24, -15, -16, 19, 28, 0, 20, 31, 12, -7, -33, -23, -22, -8, 3, 21, 58, 0, 41, 22, 3, -10, -66, 3, -37, 15, -2, 2, 3, 9, -38, 15, 5, 0, -9, -41, 15, -2, 0, -2, -10, -19, -9, 4, 12, 5, 9, 40, 10, 17, 16, 36, -30, 15, -12, -38, -36, -2, 6, -7, 25, -50, 6, -65, -65, 21, 46, 3, 8, -33, 7, 21, 0, -14, 1, -10, -9, 5, 7, 35, 0, 6, 13, -8, -47, -7, 38, -34, 2, 8, 61, 1, -42, -56, -21, 11, -1, 31, -103, 11, 17, -4, 19, 3, -54, 39, 5, -61, 0, 35, -17, -52, -53, 0, 0, -57, 7, -22, 2, -6, -2, -6, 6, 13, 13, -98, -40, -43, 38, -10, -5, 53, -30, 0, 7, 11, 17, -64, -30, -27, -29, 7, 25, 17, 40, -17, 25, -4, 4, -4, -22, 4, -10, 24, -5, 0, 3, 12, -41, 24, -7, -4, 4, -56, 13, 0, -2, -4, -19, -2, 8, 6, 13, -8, -8, 16, -12, 13, 16, 4, 46, -11, -34, -47, -5, 0, 1, -4, 7, 10, 33, -57, -60, -63, 48, -3, 22, -32, -19, -22, -6, 15, 26, -48, 15, -20, 10, 4, -1, -7, 15, 0, 17, 8, 19, -36, 3, -6, 24, -1, -3, -6, -27, 18, 18, 14, -54, -18, 24, 1, -4, 20, -62, 11, -1, -47, -2, 0, -3, 6, -2, -16, 7, -91, 0, -9, 11, -3, 2, -7, 16, -23, -7, -13, -40, 0, 52, -26, -19, 24, -7, 5, 32, -7, -9, 0, -22, -19, -13, 5, 11, -13, 16, 0, -32, -13, 11, -8, -54, 1, 15, -10, 0, 0, 0, 29, -44, 22, 31, 4, 0, -20, 6, -5, 17, 4, 17, -22, 34, -5, 36, -7, 35, -21, 28, -3, -17, -14, 2, 7, 9, -23, 13, 5, 6, -9, -2, -5, 29, -16, 1, -1, -4, -4, -17, 15, 7, 0, -11, 29, -9, -77, 6, 2, 9, -8, 9, 47, 7, -5, 12, 17, -59, -22, -44, 8, 37, -14, -14, -4, 3, -70, -7, 4, -72, 3, 22, -3, -13, -22, -6, -32, 1, -24, 9, -7, -15, 8, -21, 6, 2, 13, -6, -36, 11, -1, 0, 5, -27, 2, -2, -1, 7, 29, 14, 25, 14, -4, 5, -9, -23, 5, -12, -10, 26, 3, -9, -1, -56, -33, -4, 25, -24, -62, 1, 31, -13, 7, -2, -2, -4, 0, 2, -2, -41, 28, -27, 2, 3, -2, 38, 3, 18, 3, 20, -29, 20, 2, 44, 12, 56, -47, -7, -29, -125, -26, -36, -7, -53, -16, -17, 3, 3, -4, -58, 2, -10, -13, -52, 38, -44, 5, -48, 3, -5, -18, -1, -32, -13, -51, 14, -33, 32, -3, 1, -38, -8, 5, 0, 27, -44, -35, -14, -1, -30, -64, 54, -4, 8, -73, 8, -42, -3, 0, -8, 5, 3, -53, 2, -22, 5, 18, 7, -26, 2, -48, -9, 0, -1, -32, -3, -24, -19, 5, -2, 2, 9, -8, -15, -11, -23, -17, 0, 37, 2, -17, -11, 6, 6, 23, -13, -30, 33, -16, 34, -4, 14, -60, -6, 20, 12, -47, 12, -6, -70, 3, -42, 39, -3, -2, 0, 27, 51, 19, -21, -5, 1, -11, -10, 3, -7, 4, -25, 56, 40, -6, 7, 0, 64, 36, -7, 27, -17, -20, -32, -46, 1, -7, -49, 3, -1, 8, 22, -49, 45, -24, -62, 17, -30, -1, 8, 31, -29, -29, -4, 52, 40, -48, 24, -59, -19, 0, 33, 3, -5, -2, -20, 10, 35, 31, 36, 4, 41, 22, 3, 0, 20, -11, -27, 26, -31, 7, 10, 7, 19, 13, -41, 32, 3, -10, 0, -4, -7, 4, -13, 21, 0, 12, 6, 14, -29, -7, 5, -6, 57, -42, -23, -11, 27, -50, -13, -19, -45, 2, 17, -6, 3, 8, 15, -36, 22, -25, 35, 1, -38, -17, 2, -16, -36, -25, -4, -20, -32, 1, 11, 8, -4, -1, 4, -14, 7, 12, -10, -1, -9, 16, 8, -1, 0, 0, 10, -26, 17, 6, 0, -3, 45, 13, 9, 32, 0, 6, 0, -25, 1, 16, -55, -6, 6, -35, -3, 19, 30, -42, -19, 11, 23, -7, 6, 28, -3, -27, 2, -5, 7, -42, -15, -75, -40, -8, 13, -4, 1, -2, -2, 8, 29, -22, -14, 7, 76, -29, 18, -4, 5, -40, -7, 14, 51, 1, 31, 3, 5, 28, -27, 24, -4, -11, -6, 33, -1, 20, 6, -7, -6, 32, -5, -8, -1, 12, 4, 1, 3, -21, 49, -59, -23, -17, 11, -40, -26, 21, 12, -4, 9, -6, 11, -53, 0, -6, -14, -4, -9, -32, 17, 4, -11, 34, 12, -60, -88, 4, 11, 19, -7, -2, 0, 18, -78, 30, 73, -6, 4, -16, -7, 4, -7, 5, 23, 29, 31, -5, 5, -5, 23, 39, 36, 38, 35, 50, -30, -8, 12, 33, -40, -2, 0, -3, 2, 6, 40, -5, -22, -14, 36, 0, -24, -18, 10, -15, 4, 14, 20, -8, -4, 4, -6, 50, 1, 4, -3, -8, -43, -4, 30, 6, 1, 6, 63, 20, -25, -3, 13, -2, -20, 27, -4, 5, 20, -6, 10, 33, -43, -5, -6, 13, -3, 31, -4, 12, 17, -3, 3, -7, 3, 23, -4, -9, 0, 4, -1, -26, 2, -13, -34, -21, 56, -26, -46, 23, 38, 5, 13, 12, 6, -78, 6, -36, -8, 4, -8, 4, 8, 5, -31, 6, -4, -43, -34, 10, 28, 16, -3, -7, -7, 40, 15, 21, 43, 6, 6, -5, -13, 4, 18, 0, -8, 11, 3, -5, -12, -15, 15, 38, 28, 37, 26, 31, -29, 0, 46, -27, -13, 0, -4, 1, 25, -3, 32, -2, -33, -8, 45, -3, 12, -3, 14, -24, 0, -5, 39, -43, 3, -23, -4, -11, 4, 38, -18, -9, -70, 18, 37, -41, -12, -6, 71, -7, -26, 24, -17, -1, -6, 31, 22, 5, -6, -4, -9, 9, -29, 19, 4, 22, 4, -2, -6, -10, 7, 16, 0, -29, -6, -7, 4, 0, -3, 3, 36, -35, 19, -6, 2, -22, 58, -35, -39, 16, 30, -4, -28, -10, 5, -25, 14, 10, 23, 4, 42, 10, 6, 7, -11, 21, -6, -39, -91, 1, -2, 10, -7, 1, -6, -12, 0, -1, 23, 8, 1, -5, -2, -1, -10, 2, 35, -6, -17, 6, -7, -15, 22, 11, 5, -17, 30, 53, 7, 0, -54, -36, -52, -1, -3, -17, 26, 12, 10, -53, -56, -25, -17, -2, 15, -16, -15, -30, 8, 6, 23, -54, 16, -27, -21, 32, 7, 40, 2, 0, 6, 17, 31, -62, 9, 8, 18, -28, 2, 27, -9, -4, 4, 9, -15, 0, 29, 2, 7, 21, -99, 36, -4, 43, 3, 34, 3, 17, 2, -21, -3, 31, -6, 8, -16, 1, -3, 0, 10, -55, 23, 24, -36, -31, 49, -21, -55, 3, -9, -4, -13, 9, -18, 50, -11, 12, -27, 1, -36, 2, -7, 0, -12, -46, -1, 35, -56, 3, -23, -40, -11, -8, 2, 0, -69, 31, -25, -5, 0, -2, 0, -5, -14, -3, -13, -72, 17, 0, 19, -18, -11, -12, 6, -59, -71, 10, 15, -10, -9, 13, -62, -6, -2, 37, 4, 5, 35, -48, -35, 36, -49, -2, -10, 12, -6, -14, 3, 32, -6, -91, 35, -50, -15, 17, -12, -59, 24, 4, 39, 35, -33, -15, -4, -6, 34, -69, -25, -61, -22, -104, -15, -24, -85, -10, 22, -4, 28, -39, -57, 0, 6, -18, 0, -11, -14, 10, -50, 8, -8, -34, 4, -16, -25, 2, -6, 0, -47, -10, 37, -4, -18, -9, 3, 18, 8, -18, -110, -2, 7, 32, 11, -33, -26, 9, 0, 0, 0, -56, -6, 31, -46, -46, 4, -6, -12, -3, -10, 1, 0, 2, 3, -11, 8, 29, -36, -3, 2, 0, 0, -2, 6, -7, -74, -4, -25, -1, 1, 10, 8, -13, 26, -26, -67, -29, -63, -7, -13, -44, 33, 3, -2, 27, -28, -85, 3, 2, -61, 54, -67, 10, -12, -6, 6, 0, 5, -1, -33, 27, 10, -31, 31, -16, -40, -31, 0, -1, 15, 34, -22, 11, -14, -2, 0, -70, -13, -35, -53, -2, -28, 0, 7, -22, -17, -5, -2, -67, 44, -30, 1, 10, 7, -5, -8, -59, 15, -3, -2, -72, 5, -22, -28, -7, 3, 2, 4, 51, 35, -29, 20, 31, -37, -8, 17, 6, -55, 5, -15, -6, -33, 7, 19, -35, 3, 4, 2, -27, -3, 36, 0, -57, -1, -28, -32, 0, -1, 31, -9, 0, -8, 4, 23, 24, -3, -6, 4, 33, -8, -6, 10, 1, -6, 30, 28, -7, -29, -31, 45, 64, 3, 5, 5, 4, 4, -7, -27, 7, 5, 8, 5, 33, 27, 44, 47, -9, -78, -22, -74, 5, -14, -35, -32, 9, 9, -10, -2, -46, 35, -60, -10, 22, 9, -48, 13, -3, -48, 15, -6, -23, 8, 6, 61, 6, -14, -45, 54, 7, -23, 20, -10, 9, 50, 1, -9, -1, 26, -3, 6, 16, 2, 0, -8, -20, 28, 16, -7, -71, -7, 19, -21, 19, -1, 0, -30, 21, -16, -29, 39, -19, 18, 11, -33, -26, -36, 1, -34, 7, -19, -15, 14, -35, -23, -8, 16, -20, -28, 19, -6, 11, 9, -24, -48, -2, 30, 21, -5, 3, -1, 9, -9, 5, -4, -6, 2, 24, 9, -4, -6, 1, -8, -1, -55, -5, 12, -24, 20, 33, -12, 9, 22, 24, 26, -20, 2, 17, 0, 5, -8, 10, 1, 24, 8, 7, -43, -11, 17, 4, -13, 3, -35, -42, 2, -6, 20, -66, 19, -16, -4, 21, 33, 16, -4, 2, -42, 13, -23, 33, 26, -1, 50, 40, -17, 9, 24, -6, -11, -2, -21, -2, 25, 5, -9, 16, -21, -18, -4, 26, 7, 39, 9, 15, 56, 2, 0, -41, -5, 23, -14, 36, -4, -5, -37, -26, 25, 17, -12, -48, 59, -11, -32, -3, 5, -8, -19, -17, -34, -29, 18, -29, -59, 5, -29, 14, -12, -20, -12, 23, 8, -33, -40, -11, 25, 33, -20, -3, 0, -19, -8, -4, 57, 6, -1, 37, -15, 1, -2, -1, -2, -8, -34, -6, -16, -3, 18, -5, 4, 13, 56, 23, 0, 14, -9, 38, -17, -6, 0, 6, -6, 43, -5, -13, -37, -31, 33, -5, -65, -19, -35, -35, -5, -13, 5, -43, -9, -19, -43, 4, 16, -3, -6, 0, -70, 6, 0, -30, -15, -4, 46, 26, -8, 27, 48, 39, -15, -19, 50, 10, -2, 0, 17, 42, -33, -33, 7, 76, 5, -3, -18, -4, 0, -12, 5, -25, 0, 1, -31, 5, -6, -4, -16, 14, -57, 23, -22, -19, 33, -18, -56, 15, -16, 0, -18, -11, -6, -53, 34, 0, -11, -4, -43, 22, -18, 3, -5, 11, 3, -64, -14, 1, 3, 27, -13, -5, -5, -13, -3, 9, 27, 7, -1, 19, 0, -5, -23, -1, 15, -47, -29, -2, 27, -1, 17, 6, 26, 21, 34, 30, 0, -2, -2, 20, -49, 3, 3, 5, 11, 13, -4, -36, -47, 0, 39, 0, -41, -16, -5, -6, -3, -29, 15, -38, 14, -31, -9, 14, 43, 30, 18, -9, 5, -15, 4, -16, 22, -7, -9, 25, -13, 39, 36, 39, 10, -11, -14, 2, 12, -2, -6, 41, -83, -49, 2, 34, 4, 16, -8, 31, 11, -17, -3, -8, -3, 9, -17, -7, 5, -2, -28, -8, 45, 56, -15, -42, 46, -23, -48, -7, 4, 3, 21, 21, -16, -56, 7, -7, -27, -6, -17, 27, -33, -10, 15, 10, 12, -27, -43, -5, -1, 29, -9, -1, 4, -9, -1, 19, -25, 4, 3, -24, -4, 3, -27, 0, 25, -42, 11, -8, -12, 0, 28, 0, -17, 16, -1, 39, -2, -28, -11, -2, -7, 0, 1, 0, 17, 20, -8, -38, -21, 4, 14, -1, 24, 20, -46, -17, 0, 12, 4, -14, 20, -9, -37, 23, 18, -34, 1, -4, 26, -54, 13, -34, 27, -5, 50, 20, -11, -11, -4, -16, -6, -31, -10, 9, 51, -2, -7, 37, -11, -1, 7, -4, -5, 23, -4, 6, -35, -14, 0, 0, -5, 11, -14, 1, 6, -6, -55, 32, 11, 33, -5, -16, 39, -25, -67, -5, 30, -7, 48, -11, -15, 24, -6, 0, -33, 2, -3, 19, -45, 6, -37, -36, -4, 0, -42, 9, 12, -26, -11, -3, -4, -8, -14, 27, -30, 2, -3, -11, -3, -2, -17, -3, 13, -36, 37, -5, -17, 0, -27, -10, 1, -19, -26, 21, 44, -22, -2, 28, 24, -3, -1, 6, 4, -24, -69, -42, 2, -53, -13, -2, -60, 27, -41, 15, -11, 19, -7, 6, 25, -74, -32, -1, 16, -55, 30, 1, -12, 10, -36, -82, 4, -1, 12, -33, -18, -13, -14, 9, -31, -32, -45, -12, 32, 1, 29, -4, 7, -5, 6, 0, 6, 16, -13, 25, -14, -3, -6, -26, -1, -21, -3, -12, 3, -6, -33, 44, 12, 37, -29, 12, -13, 9, -37, -22, -27, 4, 28, 11, -38, 6, -13, 8, -9, 1, 2, -54, -35, 3, -13, 0, 13, -31, -67, -12, -22, -6, -6, -7, -8, -9, 62, 27, 36, 0, -1, 23, 6, 3, -4, 5, -69, 0, 4, -7, 3, -12, 26, -87, 42, -34, -56, -21, -49, 14, 16, -38, 22, -1, 5, 3, -44, -40, 10, 12, -33, 38, 19, 7, 29, -22, 8, 16, 0, -3, -58, 50, -17, 0, 23, -30, 2, -16, -52, -2, 32, 85, -11, 40, -31, 0, -46, -36, -28, 11, -66, 26, -43, 1, 40, -6, -3, 1, -18, -29, 47, -26, 2, -43, -4, 16, -8, 28, -41, -30, 6, -19, 1, 6, 4, -8, 0, 4, 5, 78, 15, -20, -5, 39, -5, -25, 16, 49, -48, -1, -7, -2, -13, -13, 13, -51, -35, -4, -18, -47, -28, 15, 13, -4, 3, 1, -66, 1, -50, 28, -12, -8, 0, -12, 54, 35, 47, -4, 6, -14, 17, 6, 6, -2, -3, 17, -8, -2, -5, -10, 5, -15, -38, -19, 12, -6, 24, 25, -6, -84, 25, 4, -6, 36, 3, 59, -1, -10, -42, 38, 21, -5, 1, 45, -8, -19, -10, -11, -28, 17, 58, 18, -29, 13, -3, 5, -9, 0, -23, 31, -12, -7, 40, 3, 50, 13, -45, -14, 1, 12, -33, -2, -13, -15, 1, 5, -4, -2, 26, 0, 1, 5, 6, -5, 6, -12, -24, 13, -6, 78, 3, 34, 0, -1, -4, 0, -50, 47, -29, -13, -16, 45, -23, 17, -3, 21, -44, 0, -10, 15, 5, -32, 10, -51, -47, -3, 11, -2, 2, 25, 19, 11, 6, -23, -30, 5, -25, -4, -8, -1, -3, -27, 46, 61, 58, 6, -3, 41, -5, 2, -9, 2, -86, -8, -26, 1, -14, -14, 27, 21, 24, -22, 34, 14, 26, 19, 28, -25, 8, 4, 4, 52, -4, -22, 1, -16, -30, 21, 44, -4, -7, -14, -49, -11, 0, 4, -20, 41, 50, 12, -21, -1, 25, 1, -3, 4, 5, 3, -20, 14, 29, 5, 14, 8, -35, -6, 15, 54, -20, -25, -3, 2, 18, -6, -16, 35, 32, -5, -3, 50, 7, 31, 3, 13, 29, 20, -2, -61, 7, 37, -13, 9, -4, 0, -27, 69, 19, -1, 7, 28, 6, -22, 6, 26, -14, 1, -42, 33, -2, 14, -12, -57, -35, -1, -13, -38, 6, 24, 21, 44, -5, -17, -14, 0, -12, -16, 0, -7, -1, -14, 21, 8, 53, 7, -5, 2, 5, 4, -9, -2, -13, -15, 1, -3, -19, -4, 17, 11, -24, 0, 39, 16, 38, -3, 25, 0, -2, -8, 0, 24, -13, -13, -15, -18, -29, -29, 45, -6, -32, 28, -53, -12, -6, 6, -40, 28, 33, 27, -61, 16, 56, -6, 6, -4, -30, -16, -12, 0, 39, 6, 37, 4, -10, -12, 31, 61, -45, 5, -3, 5, 57, 1, -2, 39, 27, -10, -6, 7, 5, 20, -6, -13, 5, 1, -3, 20, 6, 11, -27, -8, -2, 1, -57, 94, -8, -28, 14, 22, -11, -16, -17, 21, -42, -4, 0, 10, 15, 7, 7, -16, -46, -6, -30, 42, -15, -15, 25, -1, -3, -23, -60, 3, 2, -13, -11, -2, 2, -31, -7, 5, 59, 7, -4, 31, 8, 3, -7, -8, 11, -37, -22, -6, -21, -10, 7, 16, -8, 1, 32, 26, 26, -15, -13, 4, -33, -2, -4, 23, 5, 26, -6, -41, -43, -3, 28, 5, -33, -13, -53, -5, -3, 6, 30, 32, 25, -13, -21, 15, 36, 4, 16, -5, -43, -13, -12, -30, 22, -2, 20, 38, -19, -27, 40, 60, -37, -10, -15, 4, 4, 0, 5, 34, -28, 0, 2, 10, 0, 33, -3, 3, -48, 11, -3, 30, 0, 19, -18, 23, 5, 0, -46, 32, 19, -6, -13, 0, 3, -35, 1, 32, 9, 5, 24, -12, 25, -2, -5, -17, -48, 1, -7, 24, 10, -28, 9, 3, 2, -4, -33, 0, -11, -7, -18, 4, -8, -10, -25, -9, 9, -2, 5, -13, 8, -2, -2, 5, 29, -45, -45, -5, -4, -11, 9, -24, -11, -16, 15, 13, 1, 9, -95, 5, 5, -5, -4, -22, -6, 4, -4, -48, -36, 28, 8, -3, -39, 7, -26, 12, 6, 8, -9, 51, 35, 1, -40, 18, 0, 4, 8, 0, -36, -66, -6, -65, 36, 2, 55, 12, -11, 10, 29, 53, -35, -10, -84, -7, 31, 1, -26, 14, 3, -39, -4, -21, -5, 14, -4, 25, 7, -17, 0, -7, 7, 5, -20, 2, -7, 0, -69, 47, 10, 30, -34, 7, 27, -15, -25, 21, 0, 5, 28, 2, 13, -4, -25, 18, -39, 4, 32, 29, 8, -42, -11, 13, -3, 11, -32, -6, -10, -43, -15, -1, 3, -46, -5, -32, -22, -3, 8, 40, 15, 4, -9, 6, 43, 6, 26, 0, -44, -32, 4, -39, 14, -41, -15, 30, 53, 14, 19, 41, 49, 1, 2, 50, -47, -32, -32, -42, 4, 54, 24, 6, 14, 53, -58, 27, -6, 46, -31, 64, 16, 0, -43, 19, 12, -23, 32, -2, 29, 0, -11, -30, -1, 0, -29, -26, -3, 6, 7, 26, -31, -14, -16, 11, -8, 6, -10, 9, 65, -30, 1, -30, 7, 23, -16, 44, 9, -22, 3, 41, -1, 21, -4, 7, 0, -7, -58, 69, -18, 50, -30, 21, -1, -3, 12, -22, -18, 3, 60, -13, 3, 30, -24, 18,
    -- layer=2 filter=0 channel=2
    -15, -4, -36, 4, 8, -9, -7, -16, -8, -13, -6, 4, 35, 20, 0, 0, 0, -24, 1, -30, 56, -3, 9, 14, -18, -5, 5, 0, -18, 0, 24, 6, -4, 31, -57, -22, 51, -38, -15, -34, -10, -18, -4, 18, -4, -6, -2, -9, 2, -19, -39, 21, -13, -50, 0, 5, -4, 7, 4, 27, -3, -41, 3, 12, 26, -19, 16, -54, -21, 9, -17, 0, 55, 7, -6, 2, -22, 5, -30, -27, 39, -14, -7, -14, 12, 0, -9, 1, -47, -1, -6, -13, -7, 9, -3, -17, 1, 3, 5, -3, 7, 7, -6, 17, 3, -10, -8, 15, -7, -5, -7, -8, -4, 11, 10, 0, 14, -30, -5, 4, 31, 2, 15, -47, 3, -51, 7, 17, -17, 6, -13, 3, 17, 15, 7, -7, -9, 43, 25, -5, 17, 1, -3, -4, -4, -11, -30, -24, -24, 3, 5, -31, -25, -4, 4, 0, -8, 6, -4, -2, 12, 39, -9, -19, 21, -36, -14, -30, 5, -30, -5, 18, -13, 2, 7, 1, 12, -26, -20, 9, -19, -3, -10, -9, -38, 11, 13, 9, 2, 18, -3, 0, 4, 2, 1, -5, -17, 4, -10, -5, 25, -27, 22, 49, -11, 2, -22, -20, 31, -4, -25, -15, 9, 27, -2, -12, 4, 0, -15, -2, -13, 7, -5, -53, -3, -26, -18, 2, -19, -13, -3, 21, 0, -6, 3, 24, 1, 6, 4, -6, -19, -18, -3, -15, 5, 2, 7, 37, 28, 1, 27, 0, 8, 24, -7, 26, 3, 0, -1, 30, 0, -15, -21, -2, -8, 47, -20, -4, 7, 14, -7, -1, 3, 1, 14, -20, 21, 2, 2, -33, -7, 7, 19, -4, 15, -30, -1, 0, 14, -6, 3, -1, -20, -42, -5, -15, 10, -6, -19, 16, -7, 3, -2, -12, -5, 40, -6, 35, -10, 14, -2, -1, -5, 26, 23, -10, -4, -21, -7, 4, -28, -1, -30, 1, -16, -6, -24, 2, -9, -10, 6, 19, 3, 2, -30, -13, -23, 0, -18, -14, 13, -8, -51, -4, 12, 4, -11, 20, 7, 11, -6, -29, -6, -5, -1, -11, -21, -8, 1, 53, 3, -5, -34, -7, 4, -4, -29, -7, -15, -3, -20, 2, -17, -2, 3, 2, 3, 0, 14, -20, 5, 8, -17, 1, -2, 0, -4, -2, -6, -17, 12, -3, 2, -2, 0, -7, -4, -2, -8, 7, 6, -11, 25, -4, -59, 3, 0, -67, 6, -4, 30, 0, -15, -12, -22, -5, 3, 1, 8, -18, 27, -21, -7, -5, -20, -8, -13, -21, 1, 7, -1, -36, -14, 9, -6, 18, -3, -39, 5, 1, -11, -7, 16, 0, 0, 11, -28, 0, 11, -1, 1, -6, -11, -15, -10, -7, -33, -16, -46, 8, 35, 1, -10, -18, 32, -13, -1, 0, -8, 0, -27, -1, -2, 5, 2, 0, 3, 21, 3, -34, 8, -5, 4, 12, 2, -2, -4, 30, -3, -14, -1, -3, -2, -4, -26, -12, 9, 16, -11, 0, -4, -1, -1, -54, -10, 4, 7, 13, 11, -9, -3, -2, 6, 2, -6, -23, 4, 28, -15, -11, -4, 27, -20, -6, 1, -12, -1, 4, 3, -4, 23, 28, -20, 5, -5, -69, 3, 7, -4, 6, 6, 0, -14, -6, 7, 11, -29, -7, -47, -6, 8, -9, 5, -2, 26, 28, 16, 6, 7, 7, 12, -18, 2, 5, -5, -26, -8, 4, -1, 1, 12, -1, 0, -38, -28, -6, -41, -6, -8, 3, -20, -36, -57, -2, -33, -1, -8, 30, 8, -4, 29, -12, -9, -30, -23, -12, 3, 5, -50, -9, -14, 0, 3, -13, 28, 40, 6, -59, 0, -16, -20, -37, -7, 4, 0, 3, 1, -30, 0, 3, -4, -7, -1, 1, -7, -14, 14, 13, -1, -16, 19, -12, -16, 2, -27, -16, -8, -21, 14, 23, 10, -5, -6, 0, 0, -8, 9, -21, -7, -9, -61, 4, 29, -5, 4, 2, 7, -28, 42, 22, 28, -1, 2, -30, 5, 2, -37, -2, -37, -19, 0, 4, -1, 0, -16, -3, -3, -27, -1, -25, 21, -11, 18, 17, 1, 5, -5, 14, -7, -89, 11, 22, -10, -20, -11, -4, -52, 12, -18, 0, 10, 3, -14, 0, -10, -8, 4, 38, 5, -11, -49, -5, 5, 40, 4, -4, -11, 1, -25, -12, 13, 13, -3, -7, 3, 17, -13, -5, -20, -6, 2, -10, 11, 14, 7, -36, -3, -8, 0, 2, -1, 4, 4, 22, -1, -16, -21, 8, 7, -5, -30, 8, 0, -24, 29, 3, 2, -12, 23, 28, 19, -2, -14, -25, -26, -26, 17, -4, 4, -5, 6, -61, -5, -1, -2, -17, 6, 0, 3, -7, 4, -1, 2, 4, 10, 2, 1, -25, 6, 2, -3, -34, -18, -5, 8, 3, -21, 33, 8, -7, 15, 4, 8, -4, -26, -48, -7, -7, 1, -35, 14, -7, -14, -2, 4, 21, 24, 7, 16, 36, -8, 0, -12, -6, -22, 14, 5, 16, 7, 16, 26, 16, 3, -23, 1, -13, -23, -29, -39, -6, -2, 24, 24, -2, -2, 2, 3, -26, 47, 5, -54, 13, 5, 24, 6, 0, -32, 3, 4, 6, -15, 8, -5, -39, 1, -20, -13, 39, -4, 30, 5, -16, -7, -22, -33, 22, 2, 2, 0, -6, 22, -17, 6, -15, 19, -7, -16, -20, -8, -3, -12, -29, -9, 3, 26, -22, -4, 6, -6, -22, 5, -34, 2, -4, -7, -9, -7, 0, 12, -9, -12, 0, 8, -1, -17, -30, 5, 8, -3, 11, -14, 1, -44, 0, 13, 31, 43, -7, -9, -20, -2, 8, -6, 42, 30, -56, -3, -2, 13, -4, -7, 8, 0, -21, 2, 8, 23, 15, -7, -15, -4, -8, -50, -26, -4, 0, 6, -43, 17, -3, -16, -8, 29, -28, -47, 29, -21, -5, 1, 1, 12, -36, 16, 1, -4, -3, 14, -6, -7, 15, 5, 1, -12, 0, 23, -1, 3, 32, 4, 1, 4, -8, -3, 10, -6, 15, 1, 1, 4, -16, 5, 5, -13, 2, -3, 1, -19, 5, 23, 5, -4, -13, -2, -21, 31, -6, 14, -1, 7, -37, -7, -23, -14, -9, -5, -1, 4, -13, -77, -28, 11, -2, -18, -8, -15, 1, -4, 3, -1, -3, 2, 23, -2, -25, 23, 8, -6, -14, -17, -3, -1, 3, 19, 24, 14, -5, -17, -38, -41, -2, 4, -13, -7, -7, 17, -18, 17, -14, -3, -6, 0, -8, 13, 0, 43, 1, -4, 58, 9, -6, -11, 15, 13, -14, 10, 20, 14, 8, -3, 2, 0, 12, -34, 8, 11, -6, 15, -18, 45, -27, -17, -5, -18, -27, 12, 14, 9, -9, -2, 28, 14, -3, 4, -6, 8, -1, 17, 1, 0, -28, -5, 12, -6, 32, -52, 8, 4, -54, -2, -13, -3, 5, 0, 1, 8, 39, -19, -13, -24, 9, -14, -31, -15, 14, -43, 6, -8, -34, 11, -18, -1, 8, -2, -1, -10, 18, 44, -29, -13, 2, -11, 10, 21, 0, 3, -16, 0, 2, -1, 0, 25, 2, -43, 4, -4, -32, -26, 0, 16, -1, 4, 1, 5, -1, 0, -18, -54, 7, 28, -9, 4, -19, 20, 15, 29, -15, 13, 4, 2, 2, -17, 47, -23, 27, -3, 30, 3, -2, -12, 36, 35, -5, -4, 11, -12, 32, 5, 36, -6, -17, 0, 7, 32, -4, 9, -6, 12, -24, 39, -2, -35, -19, 15, -26, -16, 8, -16, 3, 10, -1, 13, 4, -26, -7, 5, 7, -2, -19, 0, -3, -11, -13, -9, 8, -2, 54, 0, -1, -7, -10, -6, 7, 18, 17, -9, -4, -13, 21, -12, 3, -17, 7, 17, -5, 10, 22, 31, 19, -18, -13, -33, 6, 1, 22, 15, 7, -16, 11, 3, -3, 21, -7, 4, -28, -5, 6, -2, 4, 13, 9, -22, 7, -3, -6, -5, -6, 5, -4, 14, -18, 4, -7, 1, 1, -25, 10, 24, -26, -12, 12, -9, -20, 0, -1, 2, 5, -1, -8, 2, 32, -37, 11, 14, -28, 0, 6, -12, 18, 28, -12, -1, 0, -37, -30, -21, 2, -13, -8, 13, -4, -18, 3, 5, 0, -23, 15, 37, -4, 9, -20, -10, -11, -19, -3, 0, -18, 6, -8, 10, -2, -3, -8, -5, 31, -3, -37, 0, -17, -22, -5, -14, -13, -5, 21, -7, 4, 35, -7, -1, 2, 11, -21, 10, 5, 0, -2, 4, 21, 2, -3, 10, -4, 10, -16, 0, 26, -16, 4, -14, 0, -11, 31, 20, 21, -28, -3, -4, -20, 13, 7, -39, -9, -4, 2, -3, 18, 3, 5, -27, -5, 8, -8, -7, 1, 24, -1, -19, 7, -11, -7, -9, 6, -12, -3, 12, -14, 16, 13, 24, 23, 26, -5, -2, 4, -4, 24, -17, 36, -7, 28, 13, -6, 0, 5, -7, -18, 30, 3, -5, -11, -2, -17, 0, -4, -14, -19, 25, -8, 7, 6, -52, -5, -19, 37, 17, 2, 15, -34, -10, -26, -21, -10, -19, 0, 17, 6, 25, 7, -5, 24, 3, -8, 7, -44, 7, 24, -20, -22, -1, 15, -7, 16, 6, -9, 16, 0, -3, -2, 15, 7, -15, 9, -12, 39, -10, -6, -4, 0, -48, 6, -8, -32, 18, 36, -1, -11, -23, 3, -31, -39, -3, 13, 19, -39, -8, -29, -89, 0, -19, 35, -5, -2, 3, 18, -9, -9, 51, 2, -1, 13, 0, 2, 12, 0, 20, -6, -17, 4, 0, 5, -33, 1, 7, -27, 19, -3, -17, 18, 23, -4, 8, 0, -4, 6, 32, -13, -31, 9, 46, -26, 1, 5, 4, 9, -8, 9, 9, 25, -17, 14, -26, 29, 13, 8, -11, 4, -1, -2, 13, 24, -12, 0, 13, 0, 11, 0, -2, -36, 44, -2, 2, 0, 4, -3, 35, 6, 6, 9, 7, -21, -4, -1, -3, 13, -6, -41, 22, 10, -1, 23, -3, -4, 4, 1, 2, 1, -5, 5, -3, 7, 4, 9, -3, -13, 22, 0, -18, -1, -20, -26, -12, 10, -3, 1, 0, -1, -28, -10, -3, 8, -4, -21, -11, 5, -26, 0, 23, 22, -3, -6, -4, -35, -38, -51, 19, 0, -3, -3, -1, 1, 1, -3, 10, -4, 6, 4, 22, -2, -49, -28, -31, -26, 20, -38, 19, 3, -15, 8, -5, -4, -3, 8, 30, -30, 18, 9, 19, -9, 3, 5, -8, -9, -7, 7, 8, -10, 16, 32, 17, -5, -1, -20, 2, 8, -15, -3, 33, -6, 0, -17, -6, 4, 15, -12, 12, -29, -39, 13, 12, 3, 16, 2, -2, 6, -20, -18, -4, 17, 1, -16, -1, -5, -3, 4, 9, 19, 6, -36, -2, -5, -33, 2, -3, 1, 1, -1, 24, 13, -41, -2, 1, -15, -3, -15, -21, -5, -14, -67, 7, -41, 9, -24, 5, -6, 10, -20, -45, -2, -32, 10, 0, 28, 38, -10, 26, -3, 0, 0, 9, 0, 26, -34, -20, 6, 4, 0, 7, 9, -3, 1, 6, 17, -18, 4, 10, 16, -25, 19, -22, 34, 5, 0, -2, -4, 26, 29, 15, 5, -6, -45, -1, 24, 46, 10, 21, 34, 9, -9, 17, -2, 0, -3, 2, -9, 6, -2, -78, 0, 20, 30, -19, 40, -29, -2, 3, -38, 1, 22, -3, 2, 11, -16, -1, 8, 0, -3, 23, -2, -15, 10, 26, -5, 8, 41, 21, 2, -4, -37, 0, 15, -7, 21, 8, -19, -7, 0, 2, -13, 14, 6, 0, 1, 0, 19, 19, 30, 13, 9, 0, -13, 7, -8, -1, -4, -51, -114, 22, 17, -11, 9, 3, -3, 0, -8, -14, -30, -24, 22, -4, -17, -57, 4, 4, -1, -12, -5, -5, -14, -4, -29, -7, -4, -1, -7, -4, -3, 27, 1, 13, -7, 0, 0, 1, -21, -34, -8, -1, 41, -9, 2, -23, 10, 18, -10, 12, -4, -2, -1, -22, 9, 0, 27, 15, 15, -5, -6, -14, -14, 6, -8, -5, 14, 14, 18, -1, 30, -1, -6, -3, 10, 29, -5, -27, 7, -13, 20, 43, 0, -15, -11, -23, 10, 17, 9, 17, 27, -4, -17, 28, -4, 21, 31, 22, 5, -3, 7, 1, 23, -18, 3, -14, -4, -3, 17, 7, 7, -2, -4, 0, -4, 0, 19, -23, 26, -17, 23, 7, -9, -15, -12, -48, -6, -1, -16, 20, -3, 8, -53, 0, -6, 12, 23, 0, -30, -20, 48, -10, -9, -23, -4, 18, -27, -19, -6, 9, -18, 5, 1, -31, 1, 2, -25, -13, 1, 22, 2, 27, 4, 37, 2, -20, -11, -11, 4, 26, -18, -18, 17, -3, -16, 7, -13, 30, -7, 7, -3, 20, 5, 4, 31, 39, 1, 33, 2, -21, -3, 21, 27, -6, 19, -40, 22, -15, -29, -4, 0, 9, 9, 9, 2, 3, -34, -4, 0, 29, -2, -31, -28, -33, 35, 10, 33, 22, 21, 10, -10, 21, -2, -30, 10, 10, -19, 3, -36, -4, 21, -12, 0, 4, -13, 4, -28, 6, 4, 2, 17, 1, 1, -9, 12, 0, 28, -16, 0, 31, 2, -11, -20, -35, 3, 14, 9, -4, 26, -17, -10, -30, -4, -1, -30, 33, 4, -4, 16, -8, -14, -30, 3, -3, -17, -5, -6, 10, -31, 12, 11, -25, 5, -3, -3, 7, 3, 15, 2, 21, -10, 11, -4, 5, 15, -3, -16, 34, 15, -30, 33, -14, -30, 34, -28, 28, -7, 2, 0, 6, -33, -30, 20, 52, 47, -9, -4, -33, 10, 46, 22, -3, 2, -50, -9, -7, -45, -20, 13, 11, -17, 14, 1, 7, -13, 22, -12, 5, 3, 7, -4, 9, -3, -19, -5, -13, -29, -2, 5, -16, -3, 25, 0, 6, -19, 0, -53, 2, 30, -5, -25, 12, -23, 6, -31, 5, 10, 41, -15, -2, 7, 18, -17, 0, 29, 15, -27, -4, -11, 3, -12, -47, 0, 17, 33, 24, -42, 4, -7, -5, -4, -12, -21, 22, 4, -14, 8, 3, -33, -44, 6, -32, -33, -4, -3, 5, 1, 57, 21, -55, 7, 5, -17, -9, -6, 23, -3, 2, -27, -22, 0, 19, -21, -38, 4, -1, 2, -13, 0, -17, -40, 28, -31, 37, 6, 0, 36, -23, -24, 16, 57, 32, -5, 2, 0, -11, -35, 20, 20, 5, 37, -10, -7, 22, -18, -14, 1, 9, 23, 2, -1, -17, 26, -32, 18, 40, 0, 0, -7, -2, -10, -19, 14, -7, -1, 8, 6, -5, -3, 13, -3, 21, -4, -2, -28, 0, 8, -5, -31, -10, -17, -5, -13, 3, -15, 27, 15, 5, 0, 6, 7, 14, 10, 6, 43, -1, -20, 8, 27, -45, 0, 14, 35, 14, 7, 7, -32, 0, 6, 21, -37, -45, -1, -23, 15, 0, 9, -79, 0, -9, -44, -11, -7, -5, -11, 4, -3, -4, 0, -2, -8, -19, -5, -20, 3, 7, -1, 13, -6, 12, -10, -28, 9, 3, -22, -19, 17, -8, 11, 17, -13, 13, 5, -7, -10, -19, -4, 36, 10, 19, 50, 12, -5, -15, -9, -11, 1, -1, 16, -8, 24, -8, 7, -3, -3, -22, 2, 5, 5, -41, -9, -9, 39, 15, -1, 50, -11, -1, 10, 0, -15, 0, 18, -4, 6, 5, -6, -3, 23, 28, 17, -3, -18, -1, -11, -2, -13, -3, -3, -1, -3, -1, 7, -9, 7, -2, 5, 0, 34, -18, 12, 0, 33, 33, -22, -19, 16, -29, -6, 10, -10, 21, -28, 7, -16, -1, 1, -3, 7, -5, -9, -4, -17, 11, 0, -79, -4, 27, 0, 0, -7, -4, -12, -11, -88, -22, 1, 0, 12, -7, -4, -2, -6, 13, 21, 27, 1, 5, 1, -48, -14, 38, 9, 24, 9, 27, -4, 4, 7, -13, -1, 2, -19, -6, -31, -7, 31, 26, -67, 2, -8, 9, 18, 0, 7, -5, 27, 0, 16, -33, -4, -1, 0, -20, 35, -21, -8, 3, -6, -8, -11, 34, -1, -36, 21, 46, -28, 1, 22, 29, 0, 36, 10, -18, -6, -36, -12, 7, -12, 6, 23, 9, 8, 0, -15, 14, 0, -6, 46, 6, -65, -16, 7, -1, -4, -4, 1, 9, 36, -19, 4, 15, -26, -5, -38, -16, 1, -10, -64, 13, -1, 3, -18, 6, 2, 1, 1, -43, -12, 35, 9, -8, 7, -22, 0, 27, 7, -2, 1, 4, 12, 16, -22, -1, 0, 0, -29, -2, 0, 11, -2, -28, 20, 13, 4, 34, 17, -2, -12, -20, -7, 4, -25, -3, -7, 0, 35, 40, 2, -4, -24, 20, -2, -12, -26, -31, -36, 31, 0, -2, 5, -33, 1, 11, -10, -4, 2, -9, 25, 17, 0, 18, 35, -22, -1, 7, 10, -12, 60, 32, 1, 37, 24, 20, 1, -15, 29, 9, -30, 13, 0, 19, -5, 35, 27, 19, 2, 5, 3, 6, -9, 3, 13, 26, -23, 0, 16, -3, 21, 14, -4, 2, 6, -8, 16, -3, 12, 0, 19, 14, -6, -6, -9, 16, -1, -9, -99, 13, -54, 20, -13, 21, -5, -18, -22, -10, -25, -14, 15, 3, -8, -13, 9, 14, -45, 1, 0, 6, 27, 16, -41, -3, 0, -6, -17, 0, 3, 7, -7, -8, -13, 0, -1, -11, -35, 19, 0, 4, -37, -18, -16, -10, 3, -14, 38, 4, 9, -3, 0, -13, -6, 1, 6, 2, -13, 27, -1, -22, -58, -11, -4, -11, -4, 28, 35, -13, 19, 2, -12, -41, -3, 27, 4, -13, 14, 10, 38, 22, 1, 33, -35, -4, 27, 37, -1, 12, 5, 25, 0, -17, -6, 16, 10, 34, -9, -1, -10, 4, 13, -15, 40, 0, 10, 0, 27, -1, -13, 13, 25, 0, 7, -11, 34, 3, 42, -46, 11, 21, 5, -5, -11, -9, -5, 24, -41, 21, -53, 9, -7, -40, 6, -15, 20, -22, -15, -6, 7, 2, 11, -36, -4, -17, -47, -5, 2, -4, 13, 17, 0, 16, -1, 4, -23, -3, 0, -15, 0, 35, -5, -26, 6, -12, 4, 9, 7, 28, -13, -25, -14, -16, -20, 29, 4, 25, 1, 6, 14, -9, -29, -7, 37, 36, -41, 11, 0, 4, -22, 28, -13, 8, 39, -16, -22, -1, 36, 9, 15, -10, -1, 4, 2, -14, 0, -8, 13, 15, 8, 5, 0, -30, 12, 8, -43, -9, 6, -19, 0, 6, -6, 28, -6, 0, 6, 3, -41, -4, -23, -9, 43, 5, 3, 7, 30, -1, 9, 2, 14, -5, 5, -15, -9, -7, 0, 5, -40, 17, 11, 15, 12, -23, -1, 24, 28, -29, -56, -14, -13, -53, 4, -44, 3, -32, 0, -7, -67, 1, 9, -14, -3, -24, -24, -14, -6, 0, -42, -13, -8, 6, 3, 7, -12, -5, 2, 18, -4, 62, 18, 19, 3, -20, 5, 11, -21, 37, 0, 11, 34, -4, -29, 22, -46, 26, -9, -4, 13, 19, -2, 10, 70, 28, 17, 4, 0, -50, -1, 33, 33, -2, 35, -12, 13, -7, -72, -18, -13, -7, 29, -8, -3, 51, 21, -31, 22, 14, -5, 22, -2, 2, 30, 1, -36, 15, 26, -14, -7, 35, -6, -50, -4, 24, -52, -5, -49, 0, 48, 6, 13, 35, -8, 0, -19, 5, -40, 4, -2, -6, -8, -1, -12, 11, 12, 43, -28, -6, -19, 14, -38, 74, 4, 40, 31, -14, 59, -15, -14, -24, -3, -10, -41, -15, 2, -46, -67, -26, 5, -51, 3, -16, -26, -22, 4, 8, -25, -5, 43, -20, -4, -1, -17, 5, -3, -3, 6, 38, -19, 21, 2, 21, 8, 11, 28, 2, 11, 0, 40, -6, -13, 33, -24, 47, 7, 0, 23, 22, -64, -34, 37, 36, 32, -48, 1, -43, 1, 18, 9, -14, -3, -16, -10, 8, -15, 8, -15, -9, 10, -5, -3, -17, 43, -37, 18, 22, 0, 53, -33, -30, -16, -48, -3, 2, -12, -31, -1, 44, -4, 2, -6, 21, 1, 0, -39, -3, 38, -9, -2, -8, -8, -6, -34, 2, -3, 24, 4, -3, -2, 16, -19, 19, 24, 9, 50, -4, -24, 12, -39, -4, 4, -2, 26, 8, 31, 0, -33, 7, -2, 11, -14, -68, -8, 0, -6, -5, -20, 11, -10, 19, -50, -11, -6, 4, 19, 16, 0, -6, 6, 1, -14, -19, 6, 5, -7, 14, 24, 9, -4, -15, 11, -9, 1, 4, 57, 15, 19, -13, 36, 11, -5, 3, 1, -6, 5, 30, -48, -3, 50, 11, 5, 9, 0, -18, -4, 22, 13, 4, -18, 18, 0, -19, -34, 9, 14, -9, -30, -20, 0, -6, 0, 27, 7, -9, 4, 29, -1, 14, 27, -9, 20, -14, 7, -1, 1, -53, 3, 2, -20, 24, 11, 4, -19, 3, 26, -20, 38, 16, -6, -7, 45, 2, -17, 3, -6, 0, 6, 34, 7, 2, 45, 35, 14, 22, -12, 22, -23, -63, 0, -4, -28, 4, 23, 5, 14, 7, 2, 6, -16, 21, -2, 5, -18, 9, -6, 6, 1, 7, 4, 3, 2, -4, 7, 3, -6, -15, 0, -3, 0, 0, -1, -33, 4, 25, 28, 26, 2, 10, 20, -74, 0, -6, 44, 32, 25, 19, 7, -8, -15, 7, 3, 6, -9, 26, 10, -22, -10, 5, 17, 27, -6, 8, -4, -25, 21, 2, -30, 41, 42, -26, -2, 0, 2, -46, 19, -21, -7, 4, 18, -3, -26, -7, -4, 0, 27, 31, -6, 17, 47, 4, -14, 13, 14, -14, -2, -21, 33, 10, 19, 1, -19, -1, -14, 7, 3, 17, 1, -1, 17, -6, 37, -2, 2, 6, -4, 2, 12, 11, 16, -23, 17, 7, -28, 6, -8, -7, -7, -6, -70, -17, 5, -3, 9, 15, 5, 16, 10, -47, -8, 29, 13, 5, 7, -71, 0, 4, -18, -6, 8, -1, 33, 13, -42, -37, 0, -6, -33, -8, -1, -23, 5, -34, 19, -4, 2, 27, 10, -34, -14, -7, -39, -4, -24, -10, 4, -4, 24, 8, 4, 3, -17, 4, 51, -11, -36, -20, -2, 9, 0, 0, -6, -21, 1, -3, -1, 1, 8, -11, 46, 41, -30, -5, 24, -13, -5, 27, -16, 40, 33, 28, 6, -3, 6, 29, -8, 3, 0, 20, 3, 17, 0, -9, -7, 5, 5, 20, 22, 5, 0, 7, -7, 3, 4, 31, -14, 2, 33, -3, 41, 16, 11, -4, 0, -39, 22, 15, 24, -8, 15, 21, -22, 2, 8, -12, 6, 6, -33, 35, -29, 6, -14, 12, 3, 8, -1, -29, 1, 10, 19, 7, 38, -4, 0, -9, -75, -6, -5, -1, 27, 8, -25, -37, 4, -3, -31, -18, -6, -20, -7, 8, 13, -9, 0, 7, 1, 14, -13, -28, -50, -9, -53, 0, 7, 5, 18, 3, -1, 0, 2, -17, 29, -5, -1, -22, -37, 23, -7, -31, -11, -3, -4, 4, -5, 17, -20, 11, 21, 34, -3, -24, 20, 42, 5, -28, 0, 5, 68, 29, 1, 34, -9, -16, 29, 3, 10, 13, 26, 36, 0, -13, -7, -11, -12, 11, 4, 6, -14, -4, -9, -12, 13, -4, -3, 1, -22, -6, 9, 2, 21, -1, -2, -44, 28, 24, -49, 10, 30, 7, 29, -4, 5, -39, -4, 25, -47, 35, -18, 21, -22, -6, 0, 1, 11, 4, 16, 17, 0, -8, 21, -18, 0, -21, -23, -7, -6, -2, 26, 15, 4, -53, 0, 7, -62, -16, -1, -4, 4, 20, -3, 6, 5, 13, 7, 15, -25, 3, -33, 4, 30, -6, -26, -10, -16, 2, -6, 3, 31, 3, -6, 14, 26, -21, -36, 66, -6, -14, -37, 12, 11, 6, 0, -31, -7, -18, 60, 40, -29, -21, 3, -29, 4, 50, -12, -9, 37, 37, -6, -25, -17, -17, 36, -35, 2, 4, 65, 6, 4, -16, 2, -32, 3, 0, 10, -6, -53, 3, -9, -10, 45, 0, 19, -6, -76, -2, 41, 31, 14, 2, -5, -11, -10, 3, -13, 4, 11, -4, 2, 37, 8, -2, 6, 67, 7, -7, 29, -8, -19, -13, 4, -17, 34, 25, -9, -16, -34, 0, 34, -1, -2, -19, -4, -16, 2, -2, -30, 29, 4, -41, 7, 6, -42, -9, -3, 8, 0, 51, -10, -11, 4, 3, 4, -17, -4, -38, -9, 8, 13, 7, 5, -2, -26, 10, -7, 4, -9, -8, 15, 13, 29, 26, 35, 17, 0, -32, 24, 6, -3, 1, 5, -11, -8, -13, 17, -16, -31, -11, 25, -18, -1, 46, 1, -56, 25, 1, -3, 47, -21, -17, 6, -11, -26, 1, 22, -19, -5, -29, -4, -27, 1, 10, -22, -6, -73, -2, 6, -1, 50, -18, -12, -2, 83, 6, -26, -6, 1, -7, 3, 17, 2, 20, 33, 22, -5, -2, 1, 28, 16, -45, 0, -5, 13, -13, 79, -14, -4, -10, -5, -8, 4, 9, 11, -9, -38, -9, 24, 16, 0, 9, -31, -3, -2, 3, -37, -23, -20, 14, -5, -4, -17, 0, 3, -8, -1, 70, -21, 25, -1, -8, 11, -9, -21, -16, -7, 10, 18, 15, -12, 0, -34, 21, -8, 1, 19, 0, -26, -13, 9, 10, -27, -3, -1, -45, 28, 13, 8, -3, 10, 3, 11, -11, -19, 17, 5, -27, -19, -6, -4, 30, 24, -11, 24, -13, -1, 0, 3, -26, -25, -52, 11, -4, -12, -40, 13, 2, 4, 11, -9, 7, -30, -3, -42, 6, 43, -11, 4, -25, 12, 0, 55, 1, 4, 8, 2, 1, 6, 16, 11, -20, 13, -47, 29, -13, 4, 36, -31, -22, 3, 47, 35, 8, 28, -14, -8, 2, -2, 17, 12, 35, 16, 12, -3, 10, 14, -1, -3, -5, -41, 1, 3, 3, 27, 0, -17, 43, 0, 0, -15, -6, 1, -4, -7, 26, -36, -8, -2, -24, -17, -42, -11, 8, -10, 16, 52, 1, 7, 0, -15, -11, 0, -5, 4, 28, 1, 4, 11, -12, 3, 44, 8, 0, -15, 4, 5, -10, 8, -17, -10, -22, 7, 17, -8, -38, 3, 1, 3, -48, 49, 9, -23, 9, -7, 21, 0, -20, -19, 18, 56, -13, -13, -1, 6, 32, -4, -28, 27, -12, -20, -1, -36, -3, 13, -16, -16, -36, 10, 3, 32, -4, -1, -17, 11, 7, 6, -3, 35, 23, 8, -22, 14, -6, -4, 25, -16, -70, -5, 13, -10, 27, 18, -4, 4, 8, 7, 10, 38, -13, 15, -15, 15, -16, -3, -58, 0, 8, -32, 1, -2, 9, 12, 22, -20, 5, -5, 4, -30, -19, 1, -31, 0, 18, 29, -5, -4, 12, -16, -49, 3, 8, 37, 39, 33, -10, 6, -2, -3, 12, 1, -6, 11, 4, -9, -38, 34, -11, -10, 50, -2, 2, -10, 14, 13, -1, 1, 8, 21, -18, 28, -1, -7, -9, 33, -38, -3, -8, 16, 27, 0, 4, -3, 24, 18, -13, 6, -14, 38, 0, 12, -23, 7, -8, -7, -16, -8, -2, 9, 4, -21, -5, -7, 11, 17, 4, -12, 1, 74, 0, -17, -9, 12, -2, 0, -17, 34, 20, 1, -8, 21, 21, -24, -16, -41, -36, 4, 27, -68, -19, 34, 3, 11, 25, -2, 16, 27, -8, 19, 9, -4, -7, 15, -53, -5, 14, -4, -12, 2, 9, 10, 13, -66, -2, 0, 2, -28, 13, -6, -23, 4, -45, 18, 1, -6, 14, 0, 3, 10, -5, -31, 35, -2, 18, 12, 3, 4, -1, 4, 5, 6, 10, 52, -3, -33, -25, 30, 16, 6, -24, -2, -18, 13, -8, 10, 7, 11, -5, 27, 10, 24, 22, 18, -9, 0, -21, -27, -7, 12, -16, -5, 25, 10, -15, 19, 1, 25, 0, -9, -15, 3, -3, 1, 7, -5, -1, 19, 6, -16, 2, 37, -14, 3, -3, -6, -2, 20, -5, -34, -19, 15, -3, -2, 14, -2, 13, 3, -19, 22, 19, 22, -18, 16, 16, -4, 1, -20, 18, 7, -9, -23, 15, -5, 26, 31, -18, -10, -12, 2, -13, 15, -81, 0, -8, -14, -4, -2, 9, 0, 26, -37, -68, -2, 1, -41, 4, -2, -1, -5, -21, 12, -2, -4, -17, -13, 3, -6, -41, 3, 21, 0, -11, 31, -3, 5, -3, 0, 0, 4, 7, 25, 3, -40, -33, -1, 34, 0, 0, -11, -38, -4, -1, 16, 4, 11, 0, 16, 33, -7, -25, 9, -2, 6, -40, -41, -9, 59, -2, -6, 12, -9, -32, 21, -53, 34, 7, 2, -3, 3, -1, -3, 39, -26, 3, 2, 3, 1, 5, 39, -12, -14, -2, -16, -2, 4, -5, -19, -38, 26, -5, -3, -18, 6, 36, -5, 4, 47, 10, -21, 8, 11, -12, 0, 24, -30, 29, 19, -2, -20, 20, 2, 4, -3, -27, 25, 4, -2, -12, 2, -44, -4, 1, 5, -11, -6, 8, -10, 5, -15, -8, 6, 5, -17, -1, -3, 19, -3, 18, 10, -9, -6, -7, -23, -13, 13, -2, 24, -14, -41, 11, 24, 1, -28, 0, 8, 5, 0, 3, -14, -17, -11, -5, -19, 41, 1, 12, 1, -21, -2, -2, 32, -29, -23, -22, 28, 17, -43, -34, 22, -19, 0, -9, 18, 0, 57, 20, 5, 41, -2, -30, -10, -28, -5, -8, 42, 20, -4, -26, -2, -13, 0, 14, -22, 3, -30, -3, -4, -10, 6, -6, 2, 4, 26, -3, 6, -14, 24, 6, -6, 35, -15, -12, 0, -16, 38, 22, -3, 0, 14, -3, 5, 29, -1, -10, -66, -12, 9, -13, -6, 1, -5, -39, 2, 8, -25, -3, -3, -52, -6, -29, -11, -5, -3, 7, -6, -17, -3, -35, 0, 2, -34, 0, 7, 8, -4, 41, 2, 9, -7, 6, 0, -21, -7, -46, 21, 0, -27, -23, -36, -24, -40, 13, -6, -4, -24, 17, 61, 40, -7, 10, -39, -1, 0, -12, 15, 19, 19, -2, 15, -31, 14, -13, 2, 24, -25, -2, 8, -27, 5, 14, -12, -39, -15, 40, 2, -25, 11, 24, -14, 8, -22, 7, 28, 0, -21, 16, 1, -11, -9, 6, -26, 4, -33, -4, 26, -3, 48, -27, 5, 2, 23, 6, 3, -1, 17, 7, 3, 34, -21, 4, 1, -49, 1, 31, 8, 32, -30, 10, 3, 23, 11, 15, 16, 4, 0, -25, -2, -32, -21, 5, 0, -12, -13, -9, 1, -16, 5, -3, -15, -6, 0, 5, -18, 26, 0, -34, 8, -4, -31, -13, 3, -3, 0, -9, -25, 25, -5, -1, -2, -5, -4, -20, 9, -16, 13, 11, 0, -1, 7, 7, 5, 1, -18, -2, -25, 1, -14, 14, 0, 21, 2, 11, 9, 8, 16, -4, -1, 15, -8, -29, -35, 30, -13, -36, 16, -23, -3, 14, -19, -4, 5, -11, -1, 25, -4, -6, -17, -5, -20, 20, -5, -6, 10, 12, -3, -37, -37, 0, -25, 0, -42, -3, 19, -11, 8, -6, 0, 5, 40, 2, 8, -12, 10, -3, 3, 17, -4, -8, 24, -21, 18, 9, -1, 8, -14, -7, 2, 17, 33, 18, 52, 10, -6, 13, 5, -2, -21, 10, 11, -33, 32, 0, -8, -70, 4, 0, -5, -19, -3, 0, -35, 22, -27, -37, -6, 9, -31, -15, 1, -3, 0, 11, -11, -23, 2, 34, 4, -10, 24, 0, -2, 7, 22, -24, -3, -8, 3, -6, -1, 3, 16, 14, 0, 0, -9, -9, -7, 14, 5, -9, -16, -2, -12, 0, 8, 11, -14, -26, 8, 36, 7, -18, 27, -5, 5, 10, 16, 7, -19, -39, 2, -24, -41, 5, -22, -22, 9, 3, 3, -26, 7, -18, 0, 31, -14, 14, 7, -5, -16, 2, 47, -8, -30, -9, 1, 4, -39, 2, 6, 4, 24, -4, 1, -6, 0, 20, 18, -55, 10, 15, 9, 10, -14, 6, -6, 3, -19, 31, 48, 25, 1, -7, 4, -3, 5, 7, 43, -38, 8, 8, -36, -25, -2, 2, -37, -9, 6, 3, 11, 8, -9, 17, -2, -8, -19, -5, 0, -30, -3, 4, -14, -12, 0, -21, -13, -35, 14, -33, -44, 7, -6, 0, 8, 9, 27, -13, -2, 1, -11, 25, -16, 18, -4, -28, 7, 50, -2, -20, 8, -18, 0, 0, -8, 2, 16, 16, 33, -25, -17, -3, 29, -36, 3, -44, 9, -16, 10, 36, 0, 48, -4, 17, 18, -25, 10, 14, 0, 29, 2, -7, 7, 8, 9, 3, 6, -4, -34, 4, -6, -10, 3, 5, -3, 2, -5, -1, 17, -11, 14, -4, -1, -10, 26, 11, 5, 11, 6, 11, -12, -7, 1, 21, 6, 11, -23, 23, -35, 32, 1, 5, 0, -16, 34, 1, 5, 7, -13, -10, 53, 4, 3, 20, -33, -1, 1, -3, 31, -34, -46, 7, -4, 0, -2, -6, 5, -11, -1, 0, 25, -22, 0, 12, 13, -29, 26, 18, -10, -25, 6, 66, -13, 0, 41, -13, -3, 2, -41, -11, 7, 28, -6, -24, -49, -36, -9, 0, -12, -12, -36, 0, 25, -22, -39, -34, -19, -10, 19, 16, 30, 5, -8, -9, -47, -22, -16, 52, -5, 40, 46, 17, 11, 37, -38, 15, -38, -15, 7, -13, -4, -11, -8, -42, -7, 3, 0, -4, -16, 7, -39, 26, 17, 1, -19, 2, 3, -15, 1, -7, -3, -23, -42, 12, 13, 7, -24, 17, 10, -5, 0, 33, -2, 55, -15, -15, 24, 15, 40, 14, 0, -24, 36, -16, -6, -47, -10, -19, 13, -6, 7, 22, -34, -8, 4, 1, -3, -40, -36, -22, 0, -3, -20, -24, 6, -7, 0, 25, -15, -26, 6, 3, 7, -28, 19, 22, 18, 17, 19, 34, 8, -7, 61, 6, -2, 8, -35, -4, 52, 29, -1, -4, -83, 36, -2, 9, 0, 20, 11, -4, 22, -2, 31, -47, -32, 3, -10, -13, -3, 2, -6, -10, 7, -22, 17, 30, 3, -3, 16, -18, -2, -5, -30, 6, -14, 24, 3, 24, 3, -9, 7, -18, -7, 0, -41, 0, 9, -13, -20, 35, -18, 3, 12, -3, 11, -22, 2, 0, 0, 22, -37, -33, 45, 8, -15, 0, -14, -8, -45, 30, -6, 48, -18, -25, 16, -3, 5, 11, -4, -5, 6, -58, -45, -20, -17, -5, -6, 4, 1, 22, 24, -9, 6, 3, 30, -30, -5, -77, -5, 0, 1, -20, 4, 27, 4, 29, 2, -41, -5, 18, 33, -15, -16, 20, 15, -27, -12, -43, -40, 6, 16, 0, -3, 3, -37, -13, -22, 5, -10, 25, -21, -15, -2, 38, -45, 18, 8, 0, 5, 6, -10, -59, -14, -11, 15, -17, 16, 1, 0, 14, 10, -39, 35, -46, -2, 4, 1, -22, 34, 6, -48, -7, -38, 60, 1, -16, -4, -5, -2, -44, -24, -4, 12, -6, 33, 5, 5, 6, -25, -1, 53, -7, -19, 5, -36, 7, 5, 30, -48, -20, 79, -29, -26, -4, -14, -5, -38, 24, 0, -8, -42, -36, 22, 9, 33, -6, -5, -13, 0, -8, 0, -9, -57, -3, 2, 23, 4, 20, 2, -19, 4, 6, 27, -21, 6, -2, 0, 6, 1, -20, 8, 22, -2, 22, 17, -20, -1, 14, 35, 2, -20, 14, 48, -36, -12, 9, -38, -14, 29, 8, 0, -4, -26, 9, 15, -16, -16, -6, -44, -32, 4, 8, -20, -3, 1, 2, -2, -2, 9, -25, -37, -29, 5, 8, -9, 5, 4, -9, -11, -20, 64, -13, -5, 25, 13, 22, -2, -22, -41, 2, -41, 28, -15, 1, 4, -19, 1, -41, -12, 7, 11, -4, -9, -3, 23, 3, -3, -9, -23, 0, 23, 28, -31, 3, 0, 20, -75, -4, 80, -29, -32, -30, 9, 12, -20, 22, 7, -29, -33, 14, 9, -10, 33, -3, -3, 3, -26, -46, 13, -20, -42, 0, -1, 19, -7, 32, -18, -13, -6, -6, -29, 18, -37, -36, -4, -4, 19, -5, 6, 5, -6, -30, 4, -12, 0, 11, 44, -17, 6, 9, 3, -28, -30, 26, -38, 18, 54, 1, -1, 5, -27, -13, -3, -9, 5, 11, 0, -23, -3, 32, 18, 15, 2, 11, -42, -12, -43, -72, -50, -9, -2, -4, -16, -18, 0, 17, 27, -20, 6, 9, 2, 4, 1, 16, 1, 0, -69, 20, -43, 29, -8, -30, -6, -4, 14, 5, 10, -5, 25, 7, 22, -7, 4, 40, -2, -5, 10, -5, 14, 24, -25, 3, 2, -2, -49, -28, 56, -2, -17, -19, 29, 7, -12, 9, 6, -12, -8, -36, -48, 10, 11, 16, -1, -3, -22, -1, 32, -27, -10, 13, -18, -8, -7, 12, 7, -9, 0, 9, 24, 28, -13, -65, 7, 4, 18, -16, 5, 10, 3, -26, 7, 4, 4, 7, 6, -20, 17, 26, 13, 0, 11, 0, -16, 13, 22, 2, 4, 0, -10, -5, -53, 21, 28, -1, -8, -10, 0, 42, 2, -12, -13, -2, -3, -6, -36, -35, -14, -8, -7, -15, 12, -21, -3, 30, 54, 13, 77, 8, 0, -13, 11, 12, -9, -10, -25, 9, -26, 4, -1, -9, -6, -1, 13, -15, -27, 0, 41, 6, 3, -4, -7, 23, 11, -7, -28, 7, 28, -3, -5, 5, 0, -2, -35, 11, 16, -3, -26, -3, 13, -6, 24, 10, -1, -35, -69, -29, -13, 6, -6, 5, 5, -16, -19, -20, 63, 35, -17, 0, -25, -9, -1, 0, 6, -7, -7, 4, 17, -14, -25, 12, 3, -2, -8, -11, -5, 3, 3, -27, 11, 16, -3, 9, 1, -22, 25, 15, -27, 12, -37, -10, -6, -9, 1, -6, 7, 0, -3, 12, -18, 30, 19, -35, -30, -2, -4, 12, 27, -45, -7, 10, -23, 13, -26, 10, -37, -2, -22, -40, -6, -60, 0, -27, 49, -10, 47, 38, -11, 4, 26, 16, -21, 0, -41, 10, -4, -2, -5, 2, -7, 7, -4, -10, 13, 4, 1, 1, 6, -4, 11, 19, 37, 3, 0, 3, 6, -2, 6, -1, 4, 6, -34, -9, -38, 6, -16, 0, -9, -24, 21, 25, 8, -58, -79, 2, -25, 21, -34,
    -- layer=2 filter=0 channel=3
    7, 5, 30, -21, 17, 33, 0, 16, -24, 13, -7, 5, -5, -14, 0, 4, 0, 3, 2, -8, 0, -6, 1, 27, 12, 4, 3, 0, -8, -2, -7, -6, 2, -2, 18, 15, -23, -9, 7, -2, 16, -15, -3, 28, 18, 0, -3, -2, 4, -7, 0, 18, 13, 38, -7, -6, -8, -21, -1, -4, 0, 1, -5, -24, -27, -17, -22, 35, 14, 20, 9, -1, -18, 0, -13, -15, 19, 0, 38, 3, -19, -29, 36, -5, 6, 32, 7, -11, -35, 6, -30, -2, 25, -18, 1, -18, -1, -8, 3, -6, -4, 21, 6, -11, -7, 15, 14, -30, -4, -1, -2, 16, -29, -2, -26, -25, -19, 44, 6, -5, -7, 6, -46, -20, -38, 15, -5, -5, 1, -3, -26, -53, -21, -18, -42, 15, -16, -39, 10, -9, 6, 12, -1, 3, -2, -20, 6, -31, 16, -8, 5, 17, 5, 0, 27, -6, -11, -29, -38, -6, 21, 0, 12, 25, 16, 3, -1, -32, 16, 15, 44, 1, -9, 1, 1, -2, -32, -9, 36, 33, 12, 36, -1, 2, 3, -22, 19, 0, -8, -18, -46, -5, -21, -12, 1, -3, 11, 9, 3, -6, 15, 7, -38, -6, 26, -2, 2, 8, -20, -17, 0, -6, -1, -6, 7, -2, -25, -7, -37, -26, 10, -27, 4, 27, 8, 8, 5, -24, -2, 19, -6, 26, -1, -4, 25, -15, -5, 5, -4, 6, 0, -5, 3, -22, -18, 10, 4, -22, -35, -6, 2, -16, 11, -31, 8, 1, -7, -6, 35, -35, 0, 2, 9, 24, 2, 0, -22, -6, -18, 4, 5, 1, 0, -18, 12, 10, -16, -8, 4, 0, -16, -5, -5, -7, -43, 12, 3, 2, 6, -12, -8, 40, 12, -19, 14, 23, 8, -1, 17, -10, 21, -10, -3, 31, -26, 24, 4, 21, 18, 5, 22, -5, 14, 37, 1, 20, -4, 21, -31, 10, 4, 19, 11, 0, -1, 15, -3, 8, 46, 13, -35, -6, 36, 0, 31, 10, 5, 5, 9, 20, 12, 2, 24, -8, -13, 4, -40, -27, 18, -9, -3, 12, 6, 4, 10, -16, 14, 17, -7, -43, 7, -8, 10, 30, 0, -4, 0, 19, -17, -2, -35, 6, 16, 12, 8, -19, -32, -5, -6, -12, -5, -4, 21, -3, 0, 1, 7, 5, -8, 14, 0, 16, 3, 0, 7, -2, 12, 4, 1, 3, 4, -25, -3, -11, -1, 1, 2, 22, 18, 5, 8, 6, 2, 0, -36, 1, 4, 9, -12, 32, -4, 19, 20, -7, -36, -8, 10, 30, 0, -17, -12, -9, -1, -6, 6, 0, 8, 13, 2, 2, -29, -7, 15, -11, 1, -13, -18, -16, -11, 14, -6, 13, 6, 2, 15, 8, -10, -17, -23, 19, 12, -1, 1, 0, -7, -7, -14, 25, 10, 4, -3, -12, 32, 6, -21, 13, 9, -10, -7, 14, 0, -9, 0, -50, 22, 7, -4, -14, 0, -3, 0, -4, 0, -1, -7, 16, -8, 14, -5, -8, 5, 4, 3, 9, -10, 4, 13, -10, 4, -45, 2, 9, 5, 0, 29, -17, -12, 34, -11, 40, -2, 5, -14, 7, -8, 37, 1, 5, 3, -22, -2, -3, -21, 4, 6, 13, 1, -1, 16, 6, 7, 8, -7, 1, -10, 31, 18, 2, -8, 44, 9, -19, 50, -23, -13, 3, 9, -14, 5, 7, -31, -23, 2, 37, 25, -19, 4, 2, -4, -10, 17, 28, 0, 2, -29, 5, -13, -1, -4, -4, 19, -15, 26, -1, 15, -32, -2, -4, -8, 3, 1, 19, -3, -13, 16, 24, 18, 13, -9, 10, 1, -2, -6, 6, 12, -21, 0, -12, 0, 7, 5, -26, 28, -9, -4, 41, 5, 19, -4, 3, 6, -3, 25, -8, -41, 8, -8, -3, -7, 30, 30, -13, -34, 3, 14, 17, -13, 34, -11, 31, -24, 1, -5, 30, 11, -21, -15, -14, -3, 0, -30, 5, -22, 18, 7, 0, 3, -15, -15, -8, -19, 6, -8, -5, -15, 3, 26, 8, 0, -6, -1, -6, -21, 14, -10, 5, 3, 10, -3, 31, -20, 1, -12, 10, -6, -14, -4, 21, -20, 18, -22, -5, -2, 0, -16, -2, 1, -43, 2, 17, -9, 28, -26, -3, 0, -4, -13, -3, -6, 1, 35, -5, 19, -14, -23, -7, 20, 0, -18, 4, 12, -9, 0, 3, 0, 4, 2, 3, -1, 2, -7, -2, -1, -36, -7, 11, -3, 32, 10, -16, 6, -2, 1, 28, 7, 28, 21, -3, -3, -4, 36, 3, -23, 24, -16, -38, 14, 3, -38, -39, -13, -2, 14, 19, -21, 26, -4, 45, -5, -1, 0, 21, 8, -17, -14, 11, -14, -30, -10, -3, -24, 16, 11, -5, 0, -37, -14, -17, -66, -5, -2, 16, -3, -7, 4, -4, 42, -5, -61, 6, -7, 12, -10, 9, 37, 1, -30, -34, 0, -19, 0, -11, 10, 2, 5, 5, -26, -44, -55, 22, 21, 7, -10, 9, 2, -26, 21, -13, -7, -1, -14, -10, -12, 3, -33, 24, -1, 19, 27, 6, 2, -9, -16, -23, 17, 0, -23, -6, -38, 29, 14, -8, 12, -4, -6, -5, -27, 1, -6, 13, 17, -40, 2, 11, -3, -5, 4, -22, 22, -5, -5, 39, 0, -4, 5, -24, 5, 3, -6, -4, -6, 1, -13, -36, 32, 23, -32, -14, -34, -3, 35, -5, -50, 21, -26, 26, 15, -5, -4, -33, -38, 15, -35, 6, -15, -4, 36, 1, -33, 16, 2, 8, -3, -19, 12, 21, -6, 4, 2, -5, -3, -2, 23, 1, 4, -12, -10, 7, -5, 19, 30, 19, 12, 0, 33, 29, -15, -9, -5, -21, 13, -6, 4, 15, 19, -2, -30, 20, 1, -23, -2, 8, -7, -22, 13, 6, 1, 18, 4, 3, -1, -3, -35, 16, 25, -27, 26, 4, 0, 22, 10, 2, 45, 3, 40, 8, 2, 7, -1, 0, -6, 45, -14, -6, -19, 6, 1, 41, 10, 0, 5, 23, -1, 32, 8, 36, 19, 9, 3, 21, 6, 6, 23, -44, -1, -4, -12, -7, -2, 10, -16, -18, -16, -5, 3, -35, -28, -7, -29, -3, -1, 11, -2, 8, 8, -7, -30, -27, -19, -2, -2, -1, -7, -21, 0, 4, 11, 22, -1, 3, 1, -11, -33, -1, 27, 2, 0, 21, -23, -6, 24, -6, 22, -5, -21, -2, 16, -7, 17, 0, 25, 24, 12, 6, 21, -8, 10, 0, 29, -4, 6, 17, -16, 0, -21, 4, 25, -13, 3, -3, -11, -73, 16, 11, -8, 12, -18, 10, -7, -39, 2, 29, 9, 7, 0, 0, -2, 15, -17, -1, 3, 0, -30, 32, -3, 1, 3, 18, -10, -10, -4, -11, -1, 0, -13, 14, 24, -42, 5, 12, 2, -5, 5, 10, 7, 12, 2, -9, -6, 28, 3, -2, -4, 6, -15, -41, -7, 16, -6, -5, 26, 10, -7, -11, -32, 7, 10, -26, -57, -19, 0, -14, -18, 3, -7, -21, -28, -3, 0, -2, 3, 7, 6, -3, 5, 16, 2, -1, -1, -1, -7, 4, 63, 2, -3, 15, 0, 3, 22, 5, 23, -3, 1, 6, 7, 7, 19, 16, 16, 27, -9, 19, 21, -4, -3, 1, 4, 1, -1, -6, -29, 1, -32, 44, -13, 8, 25, 5, -18, -7, 10, 12, -2, -4, -19, -15, -21, 13, -3, -24, 44, -8, 11, 0, 33, -3, -11, -11, 0, -8, -33, -16, 7, -20, 22, 23, 1, -9, 8, 9, 20, -4, 2, 5, 16, 10, 4, 1, -3, -6, 6, 21, 3, -6, -7, -17, 5, 8, 19, -14, 0, 6, 11, -44, -3, -13, -7, -18, 9, 0, 12, 16, -24, 7, -13, -40, 2, 7, 11, 5, 9, -6, -37, -33, 20, -31, 16, -14, -14, -3, 43, -9, 15, 26, 6, -3, -1, -26, 11, 1, -5, -2, -8, 8, -8, 5, 29, -1, -15, 0, 15, -6, 0, 6, 34, -12, -18, 27, -29, 8, 17, -16, 3, -17, 25, -9, -5, -14, -43, -3, -42, 8, -1, 6, -2, 3, -9, -13, 3, 28, -3, 0, -24, 28, 0, 16, 0, 12, 4, 4, 20, 0, 28, -12, -7, 12, -8, -6, -3, -19, 0, 10, 15, 0, 1, -18, -9, -14, 34, -2, -19, 4, 16, -24, 0, 25, -2, 4, 12, 9, -9, -22, 5, 36, 5, -16, 1, -17, -2, 4, 24, -32, -6, 3, -8, 38, -39, -15, -8, 20, -31, 0, 18, 19, 14, -54, -16, -3, -6, -1, -32, -25, 4, -16, -16, 8, -8, 30, -6, 0, 24, 17, 9, 6, -1, -16, -22, 35, 6, 3, -7, 9, -1, 6, 13, 4, -9, 10, 35, -6, -17, 4, -1, 27, -2, -2, 7, -35, 47, -11, -7, 27, 15, -7, -1, -4, -19, 13, -3, -8, 2, -22, 2, -6, 0, -22, 4, 4, -2, -17, -32, 2, -14, 8, -3, 12, 15, -30, 18, 1, 25, -17, 13, -12, -17, -2, -44, -16, 7, -14, -19, -12, 11, 3, 2, 8, 46, -4, -16, 48, 2, -29, 4, -3, -5, -4, 1, -18, -5, -6, 6, 24, -3, -1, 18, 17, -7, -1, 34, -19, -21, -15, 0, 3, -33, 7, 6, 26, -20, -5, -12, -15, -5, 39, 3, 34, 8, 7, -11, -17, -18, -6, -47, 22, -3, 0, 14, 1, 5, 1, 14, 5, 6, -34, 23, -11, -16, 0, -7, 0, 0, -2, 9, 4, -18, -7, 25, 5, -12, -15, 23, 28, 30, 2, -35, 2, -8, -3, 7, -1, 0, 0, 2, 10, -45, 3, -28, 5, 3, -17, -15, -3, 6, 24, 9, 23, 1, 6, -17, 2, 4, 23, -5, 4, 13, 0, 21, 4, -21, -32, -31, 1, -17, -9, -43, -34, 2, 29, -10, -22, 2, -4, -2, 6, -15, -3, 12, -3, 14, -14, 4, -2, 9, 12, 7, 13, -23, -12, 6, -21, -5, -7, -3, -14, -6, -4, 14, -15, -31, 14, 1, 10, -9, 18, -16, -3, -53, 0, -7, -16, -2, 2, -13, 47, 4, 0, 26, -5, 16, -5, -15, 33, 0, 0, 17, -2, 0, 8, -1, 0, 7, -15, 5, 49, -46, -3, 3, 6, -8, 0, 10, -8, 18, 1, -42, 7, -4, -3, 12, 30, 40, 25, -14, -38, 12, 18, 10, -2, 14, -16, 4, 7, -13, -14, 7, -6, 16, 1, -6, -3, 14, 27, 27, -21, -3, 5, 0, 3, 19, 16, -16, -11, 21, 12, 27, 0, -18, 3, 8, -6, 22, -2, -23, 2, -13, 6, -1, -18, -1, 12, 17, 1, -19, -3, 18, 18, 9, -3, 4, -4, 2, 15, 11, 7, -11, -8, 1, 27, -2, 28, 7, -25, -4, -1, -11, 23, 23, -28, -17, 8, -3, 12, -18, -14, -34, -5, 34, -15, 11, -15, -30, 35, 37, 0, -18, -4, -1, 19, -41, -5, -20, -16, 12, -4, -12, 8, 0, 0, 6, -14, -9, 5, -29, 3, 7, 13, -11, -7, -10, 4, 11, -7, 4, 7, 4, 19, -2, 29, 15, -22, 16, 22, -20, 0, -5, -5, 10, -4, 3, 11, 3, -39, -25, 8, 14, -33, -14, 2, 10, 17, 11, 0, -1, 0, 0, 6, 14, 1, -11, -34, 2, -37, 0, -2, 3, 15, 21, -43, 12, 0, 18, -33, 1, 38, -1, -26, -12, 33, 0, -12, 5, 7, -3, 5, 11, 27, -4, 25, -1, -3, 0, 0, 1, 3, -5, 4, 3, -5, -7, -9, 5, 5, 19, -8, 3, 17, 35, 16, -24, -5, -8, 20, 37, -3, 18, 14, 10, -22, 23, 28, 7, 2, -17, 5, 3, -6, -20, -3, -8, -4, 25, 5, -14, 13, -2, 0, -5, 20, -2, 3, -10, 5, 5, -9, -32, 5, -18, -5, -4, 38, -8, -5, -18, -15, 11, -23, 24, -21, 6, 9, 19, 19, 3, -5, 2, -5, 2, -16, -51, 11, -38, 7, -9, -3, 23, -1, 15, 37, 8, 8, -14, -26, 1, -1, -28, 25, 5, -12, 0, 9, -11, -3, -3, -30, -17, -22, 2, -10, 17, -9, -7, 36, 32, 11, -4, -25, 33, 2, -33, -6, -15, 8, 7, 0, -6, -11, -8, -39, 8, 17, -16, -23, 6, 6, 4, 10, -2, 12, 5, 1, -37, -19, -23, 5, -56, -18, 4, -22, 4, 12, 15, 0, 17, 21, 23, -73, -11, 13, -43, -4, -15, -12, -16, 3, -32, 29, -4, 8, 60, -3, 4, -27, 0, -3, 6, -23, -4, -5, 44, -3, 7, -7, 2, -5, 17, 2, 55, 16, 10, -3, 44, 9, -17, -33, 11, -19, -39, -15, 45, -7, 17, -8, 13, -3, 3, -30, -36, -67, -57, 9, 18, -7, 0, -2, -15, -30, 34, 22, -10, -45, -2, -9, -16, 15, 15, -11, -16, 48, -7, 1, 10, 13, 2, -5, -7, -3, 15, -32, 16, -5, -27, -4, 29, -70, -8, -2, -11, 5, 0, -27, 25, -14, 3, -15, 0, -88, 2, 9, 11, -10, 4, -29, -7, 5, -1, 11, 4, 7, -24, -8, -17, 12, -10, -16, 33, -5, 2, -33, -10, -5, -9, -10, -56, -20, 17, 3, -62, 7, -38, 19, -18, 2, -24, -42, -2, 2, 81, 0, 15, -11, -7, 2, 7, 38, -13, 31, 17, 6, 0, -18, -7, -1, -3, -3, 42, 22, 14, 4, -4, -15, 9, -77, 20, -79, -15, -5, 82, 10, 1, 66, -11, 3, -2, -9, -28, 19, -44, 7, 7, 4, -50, 8, 1, -81, 21, 35, -8, -30, -37, 25, 23, -32, 28, -58, -35, -16, -20, 1, -7, -10, 0, 5, 8, -3, -39, -37, 25, 9, 15, -20, 17, -64, 6, -1, 55, -4, -47, -17, -31, -4, 7, 6, 2, -71, 6, -23, -18, 8, 1, -4, 0, 34, -27, 9, 3, -6, 25, -49, -49, 26, 48, -13, -25, -23, -1, -10, 28, 5, -22, -15, 23, 19, 13, 19, -23, 0, 20, 10, -32, -15, -21, -7, -17, 44, 45, 6, 1, -21, -3, -6, 5, -23, 22, -18, -3, 4, -7, -17, 9, 6, -12, -4, -17, 33, 36, 6, 1, 10, 35, 12, -13, -20, -18, -23, 73, -7, 11, 56, 14, -9, -1, 0, 13, 0, -11, 13, 0, -24, 16, -2, 2, 0, 11, 11, 4, -28, -12, 28, 0, 13, 6, -25, -14, -1, -14, 1, 0, -24, -16, 2, -35, -1, 16, -12, 33, 0, -20, 11, 17, -58, 13, -4, -31, -6, -12, 13, 1, 10, 7, 3, -4, -37, 4, 9, 11, -9, -7, 6, 2, 19, -14, 16, 7, 2, 6, -36, -15, 4, 40, 16, 7, 6, 18, -21, 27, 4, -11, -53, 2, -14, 26, 32, -28, -6, -36, -39, 14, 19, -46, -10, -7, 9, -17, 5, -22, -8, 8, 4, -4, 14, -9, -17, -15, 4, -3, -3, 14, 4, 4, -1, 3, -9, 20, 0, 16, -6, -16, 31, -2, -32, -12, -25, 30, 8, 6, 26, -6, -4, -6, 3, -21, -9, -36, 11, -15, 2, 13, 0, -16, -30, -18, 11, -6, -26, 19, 29, -24, 25, 17, 15, 13, 19, -30, -6, -4, 5, -30, -51, -12, -4, 6, 9, -5, 0, 27, -4, 26, -8, 4, -11, -7, -3, -39, -22, 11, -64, 7, 5, 0, -4, 0, -11, 8, 3, 4, 28, 7, 4, -10, 0, 5, 7, 16, -17, -10, -8, 28, -13, 2, 16, 8, 0, -49, 0, 3, -40, -29, 25, -37, 18, 20, -6, 1, -14, -32, 27, -63, 3, -10, -15, 19, 5, -8, -3, 0, -6, 7, 36, 39, 22, 24, 5, 5, -4, -3, -1, 11, -9, -55, 4, -11, -5, -4, -14, 6, 61, 18, -24, -17, -52, 15, 14, 5, -18, 11, -9, 4, 32, -8, 4, 7, 5, -3, -16, -32, -2, 18, 0, 26, -10, 1, -21, -20, -11, 14, -27, 12, -23, 8, 7, 10, -4, 11, -12, 14, -1, 11, -4, 13, -27, -5, 7, 3, -44, -1, 18, 24, -11, 11, 6, 7, 20, 13, 30, -3, -1, 0, 39, 8, -6, 2, 4, 1, 13, 3, 4, 1, -12, 0, -2, 8, -12, 29, -16, 36, 4, -5, 0, -28, 39, -24, -5, -49, -42, 2, -5, 7, 24, 25, -1, 6, -21, 9, -35, -35, 4, -10, 33, -5, 6, 16, 7, 5, -6, 0, -3, -2, -4, -19, -2, 2, -13, 2, -7, 4, -6, 41, -18, 13, 4, 5, 24, 12, 9, 4, -7, 21, 25, -8, 4, 22, -11, 4, -12, 0, -1, 25, -8, -23, 17, 30, -98, -36, -4, -4, -7, -4, 5, -3, 15, 28, 5, 21, -10, 0, -12, 9, -4, 10, -1, -1, -67, -7, -37, -2, -2, 48, 10, 6, 8, 3, -12, 3, 12, 11, -12, 41, -3, -9, 7, -1, 37, 0, -26, 1, 18, 6, 0, -2, 3, -7, 15, 5, 12, 18, 22, -5, -5, 32, -11, 6, 12, -24, 6, 2, 9, 14, -11, 1, -4, 0, 44, 0, 11, -11, 23, 5, -3, -20, -21, -10, -22, -37, -16, -3, -3, 28, -7, 8, -3, -4, -3, 0, 11, 8, -10, 10, -1, -4, -31, 12, 3, -15, -2, -4, 10, 5, 1, 28, 18, 15, -3, 15, -14, -19, -31, -4, 4, 15, -23, -7, -3, -4, 34, 9, -9, -42, 8, 23, -18, 5, 5, -12, -20, 0, 15, -3, -21, -10, -7, 0, 51, 26, -43, 6, 4, 9, -2, 23, -1, -47, 0, 1, 2, 21, -11, -12, -20, -9, -31, 2, -27, 12, -3, 13, 2, 5, -40, -4, -13, -2, -10, 0, -33, 18, -50, 4, -11, 5, 0, 6, 5, -6, 18, 6, 5, -11, -13, 19, 23, 6, -17, 0, 16, 27, -11, -40, -2, 8, 1, 0, -7, -9, -12, 10, 5, -8, 9, 0, 9, -8, -9, -6, -1, 47, -8, 1, -23, 0, 5, -6, -19, 8, 14, 37, 3, -5, -2, 20, -6, -23, -4, 7, 4, -1, 6, 22, 1, 4, -64, 16, -6, 2, 12, 35, 19, 16, 9, 3, -5, 3, -16, 3, -19, -84, 13, 13, 40, -44, -1, -10, -41, -1, 12, -14, -16, 16, -10, -17, -12, 16, 6, -52, -25, -46, 0, -27, 17, 21, -17, 1, -2, 2, -12, 18, -17, -43, 10, 2, -57, 5, -15, -29, -5, -28, -17, 14, -52, -3, -19, -5, -81, 4, 3, -7, 6, -3, 30, -3, 32, 0, 20, -3, -4, -81, -24, 2, 17, 8, 2, 22, -15, -5, 19, 13, -7, -29, -34, -2, 19, 28, -10, -29, 0, -39, 19, 29, -6, -19, -37, -12, -1, 105, -8, 24, -33, 4, 8, 7, 1, 22, -25, 0, -2, 4, -6, 2, -3, -35, 4, -6, 0, -8, 7, 17, -9, 0, -41, -27, -54, -43, -51, 39, 22, 21, 49, -3, -12, -3, -25, -9, -9, -53, 13, -13, 35, -34, 0, 17, 34, -9, -2, -5, -17, 4, 12, -22, 35, 34, -36, -40, -11, -51, 0, 20, 19, -19, -31, 11, 5, -5, -10, 5, 12, -8, -32, 6, -50, 5, 5, 9, -3, 6, -20, 0, -1, 2, -7, 7, -74, 0, 0, -11, 5, 0, -27, -6, -14, -8, 5, 4, -3, -91, -55, 8, 12, 55, 9, -43, 0, 2, 4, 13, -5, 4, -83, -9, 12, 23, 2, -1, 1, -6, 25, -17, -3, -71, -12, -19, 31, 44, 0, 19, -38, 7, -6, -5, -24, -8, -38, 59, 2, 3, 12, 1, 0, -31, 7, -17, 9, 3, 2, 8, 1, -31, -33, -21, -56, -43, -51, 47, -2, 32, 43, 8, -9, 5, -7, -26, 12, -40, 11, 15, 26, -24, 8, 5, 41, 9, -4, -9, 16, 19, 33, -11, 18, 33, -29, 9, -19, -13, 0, 10, 21, 23, 21, -23, -9, -33, -69, 23, 23, -13, -20, 3, -41, 3, -6, -29, -3, 40, -4, -2, 3, 4, 1, -1, -56, 11, 20, 17, 13, 0, 20, -2, -4, -12, -6, 5, -5, -21, -8, 0, -4, 52, 46, -23, 28, 30, -13, -13, -1, -20, -68, 29, -34, 43, 27, -7, 3, 15, 17, 1, -11, 0, 17, -12, -4, 0, 11, 0, 5, -6, 6, -5, -13, 0, 11, 17, 2, 1, -11, 0, -6, 0, -2, 0, 8, 43, -8, 8, 12, 11, -28, 5, -29, -64, -64, 19, -31, -2, -15, 28, -9, -1, -24, -15, 24, -12, 13, -6, 8, 26, 4, 4, 0, 23, 19, -9, 3, -22, 9, -10, -16, 24, -7, -20, 2, -30, 8, -16, 14, 2, 4, 9, 3, -28, -14, 2, 8, 6, -21, 12, -20, 23, -4, -2, 7, -2, 0, 35, -24, 3, -29, -6, 0, 3, 4, 3, 4, -5, 4, 2, 9, -12, -20, -6, 3, -43, 14, 2, 0, 3, 10, 12, -19, 9, -2, 14, 0, -17, -40, -10, -19, 16, -14, -8, 5, 13, -8, -15, 10, -45, 3, -21, 4, 15, 7, -13, 8, -3, 3, 3, 7, 12, 7, -39, 4, 5, 14, 4, -4, 16, -7, 0, 8, -3, 0, 3, 2, -9, 16, -32, -7, -25, -27, -28, 1, 15, -17, 0, -11, -5, 17, -20, -37, -10, 8, 8, -8, -16, -7, 0, 0, 5, 1, 0, -23, -32, 5, 6, -34, 10, -19, 0, -10, -10, -4, -17, 0, -9, -28, 13, 0, -36, -1, 7, 0, -43, -57, -6, 0, 25, -11, -4, 4, -7, -1, 4, -15, -1, -4, -6, 13, -8, 32, -23, -4, 2, -6, 0, 30, 7, -2, 4, 1, -11, -4, 10, 9, 8, -1, -13, -12, -9, -42, 7, 2, -29, -29, 36, 33, 33, 19, 30, -4, 20, -13, 34, -35, -32, 7, 9, -14, 22, -2, 6, 3, -2, 5, -4, 21, 13, 4, 7, -1, -3, -15, 3, -7, -4, -4, -9, 3, -15, -3, -31, 3, -21, -3, -16, 30, 1, -6, -3, -3, 25, 0, -5, -14, 5, 14, 53, -11, 0, 17, 5, -33, -3, -2, 6, -12, -5, 3, -2, 11, 17, 15, -9, 22, -9, -5, -24, -23, -25, -1, -40, 0, -39, -47, -12, 2, 21, -12, 8, 8, 0, -27, 0, 13, 1, 4, 9, -2, 31, -19, 5, 21, 2, -14, 4, 16, -5, 19, -9, -29, 3, -1, 1, -20, 7, 24, -4, 7, 41, -28, 4, 1, -24, 20, -14, -19, 8, 0, 17, 0, 1, 15, -8, -8, -39, 0, 6, 6, 29, 0, 28, -1, 6, -18, -4, 7, 49, 4, 5, 0, 10, 2, -3, 5, 15, -70, -33, 0, 4, -10, 17, -5, -15, 1, -13, 17, 2, -6, -25, -4, 0, -33, -22, -15, 0, 9, 34, 4, 21, -5, 16, -19, 0, -34, 12, -30, -31, -13, 22, -21, -37, -9, 5, -69, -11, 3, -5, -1, 31, 0, -44, 20, -11, -35, -39, -29, -43, 5, -17, 25, 18, -18, -14, 4, 5, 6, -6, -17, -41, 12, -2, -18, 30, -9, 23, -6, 18, 1, 12, 23, 0, -29, 1, -18, 7, -1, -1, -19, -1, -18, -2, 1, 21, -4, 0, 6, 11, -21, 22, -5, -38, 11, -41, 1, 10, 24, 62, 0, -4, -16, 6, 7, -41, -10, 17, 9, -9, 7, 4, 9, -14, -2, -15, 0, -17, -9, -11, -1, 7, 0, 0, 11, 22, -50, 14, -3, 6, 8, -6, -5, -14, 6, -19, 26, 5, 3, 9, 8, -12, -57, -3, 51, 12, -5, 7, 26, 12, 2, 16, -7, -3, -32, -43, 10, -21, 5, -3, 17, -15, 0, 13, 55, 5, -9, -4, 5, 2, -7, -34, 22, 29, 6, -21, -37, 5, -1, -19, 19, -19, -39, -47, 1, -11, -4, 5, 36, -10, 28, 0, -34, 2, 12, -56, -5, 38, -59, 21, 1, 4, 4, 0, -73, 7, 29, -3, -7, 5, 22, 7, -24, 0, -4, -4, 1, -63, 6, -16, 2, 7, 44, 0, -8, 9, 1, 3, 4, -24, 10, -4, -27, 11, -8, 18, -3, -36, 0, -21, 2, -17, -54, -11, 8, 29, 6, 10, -23, -6, -3, -3, 5, -27, -39, 6, -3, -7, -31, 2, 0, 3, -2, -17, 8, 0, -6, -8, 23, 2, -54, 10, 12, -5, -32, 8, 13, 27, 8, 15, -12, -1, -32, -11, 13, -14, 12, -1, 0, -35, -2, 6, 1, 1, 3, -8, 8, 23, 33, 5, -2, 13, 2, -51, -14, -14, 1, 27, 10, -11, 4, 43, -3, -8, -3, 30, 21, 9, -41, -9, -19, 27, -3, -40, -3, 35, -7, 0, 11, 6, -10, -9, -57, -6, 13, 14, 11, -6, -15, -6, -30, -10, -26, 0, 0, -54, -36, 16, -29, 35, 23, -57, -3, 11, -33, 5, 8, -11, -41, -12, -40, 19, 17, 20, -2, -19, 29, 15, -34, 4, -46, 0, 4, 6, -8, -2, 2, 0, 2, 7, 12, -2, -29, -5, -6, -9, -51, 13, 1, -11, 4, -41, -1, -9, -4, -27, -17, -14, -25, 17, -19, 0, -39, 27, -25, 11, 41, -1, -6, 6, -18, 2, -16, -3, 14, 26, -6, -15, 2, -17, -13, 22, 3, -11, -10, 46, 33, -25, 6, 11, 4, -55, -2, -14, 2, -4, -6, 5, -18, -17, -9, 9, 16, -19, 23, -23, -14, -18, -33, 23, 2, -35, 3, -11, -24, -8, 2, 4, -43, 0, -53, 10, -1, -10, -2, 6, 21, 3, -6, -4, -6, 0, 9, -86, -28, 49, -4, 11, 2, -10, 0, -8, -9, 36, 0, -9, -35, -40, -12, -11, 13, 3, 3, -31, 15, -9, -18, -3, -7, -16, 30, 27, -2, 4, 7, -8, 7, 6, -2, -2, -7, -23, -1, 1, -7, -1, 2, 0, -5, 13, -3, -24, -1, 18, 0, -34, -42, 6, -9, -23, -6, -8, 0, 23, -23, 7, -4, -1, -1, -37, 52, 10, 31, 8, 4, -23, -2, 19, 20, 4, 0, -6, -12, 10, -12, -27, -17, -4, 5, -35, 17, -43, 2, -17, -28, 6, -16, 13, -2, 12, 8, -3, -33, -21, -9, 27, 2, 13, 0, -81, 2, 11, -33, 16, 9, 1, -17, -8, 16, 10, 2, 35, -29, 6, -11, -4, -30, -1, -9, -1, -3, -13, -2, 22, 12, -7, 3, 9, -8, 9, 2, 27, 3, -20, -44, -7, 14, -2, -16, 1, 0, 2, 20, 18, -2, -23, -37, 0, -5, 45, -1, 17, 21, 1, -3, -4, -13, -16, 22, -5, -1, 0, -26, 3, 1, 23, -3, -1, -12, -5, 2, 5, 2, 13, 13, 22, 43, 0, 22, -26, 22, -23, -11, 14, -3, -1, -9, -34, -34, -41, 14, 2, -9, -32, 2, 22, -13, 13, 10, -8, -28, -21, 3, -14, -9, -11, -13, 7, 5, 0, 4, 9, -14, -30, -23, 0, -9, 15, -5, 10, 10, 0, -29, 17, -26, 20, -23, -55, 3, 15, 0, 25, 5, 4, -39, -4, 50, 4, 13, -7, -9, -1, -28, 0, -7, 11, -25, 0, 4, 10, -7, 15, 6, 32, 17, 0, -3, -10, 33, 32, -4, -3, -1, 21, -33, 1, -10, 29, -5, 34, -27, 7, -18, -35, 37, -9, -16, 53, -2, -41, 1, -3, 0, -4, -5, 41, -9, -18, -2, 6, -3, 3, -1, -11, 7, 20, -14, 33, 2, -18, -22, 40, 38, -3, 34, 4, 21, 32, 3, -4, 1, -8, -2, 2, -12, 10, -1, 2, 12, 0, 2, -21, -3, 23, -21, 17, 22, 1, -28, 32, -8, -29, 9, -11, -25, -18, -22, 1, 4, -15, -3, 43, 1, 43, -8, -27, -16, 12, -24, 15, 26, 9, 31, 3, -8, 20, -4, 20, 23, -8, -9, 0, -9, 3, 5, -1, 0, -22, 3, -7, -24, 7, 1, 7, 11, 0, 3, 44, -25, 27, 7, 7, 9, 8, -29, 1, 10, -15, -7, -18, 8, 4, -7, -3, 22, -4, -5, -4, -43, 2, -12, 14, 7, -15, -11, 29, -6, -3, -9, 4, -5, 3, -5, 6, -33, -30, -6, 2, 1, 18, -5, -4, 3, 12, -10, -34, 7, 0, 9, -4, -14, -17, 19, -2, 1, -7, -6, 40, 19, 4, -13, 1, -34, 14, 1, -26, 34, 41, 20, -8, -3, -7, 7, 26, 11, 3, -10, -6, 0, -38, 15, -4, -5, -21, 29, -24, -1, -21, 25, -7, -23, 2, -2, -6, 11, 12, 1, 14, 24, -2, -13, -3, -2, 0, -1, 9, 2, 18, -8, 4, 3, -6, -38, 1, 24, 26, -8, 3, -19, 4, 9, 19, -12, 2, -5, -6, -3, 2, 28, -17, 12, -14, 2, -4, -29, 11, 10, -12, -40, -1, 19, -8, -29, 6, 1, -37, -23, 17, -10, 3, -17, -22, -4, 0, -5, 9, -1, 15, 0, 5, 20, 30, -26, -10, -4, -3, -17, 8, -4, 10, -2, -6, 18, 47, 6, 10, 8, 23, 1, 2, 10, 16, 32, -25, -1, 44, -4, 6, -11, 1, 8, -6, -33, 25, 12, 21, 10, -2, 5, 24, 22, 7, 18, 10, 20, -14, 18, -35, 20, 30, -42, -3, 3, -8, 2, 12, 24, -9, -72, -6, -3, -11, -11, 24, 0, 31, 23, -1, -52, 0, 11, 35, 6, 25, 6, 8, 33, 1, 0, -1, -30, -3, 25, 2, 5, -1, 3, 0, -8, 23, -30, 2, 6, -4, -30, 32, 7, 41, 21, -31, 18, 18, -3, -42, 1, -32, -37, -29, 13, -7, 11, 39, 4, -14, -15, 22, 2, -19, -42, 4, 21, 55, 6, 0, 12, -3, -1, 0, 8, 28, -54, -4, 0, -3, -4, 0, 0, -10, 9, 1, 33, 0, 5, 1, 3, -20, -20, 4, -8, 3, 23, -9, 8, 29, 0, 0, -1, 5, -9, -3, -19, -17, 29, 1, 4, -25, -8, 16, -67, 21, -19, -2, 11, 50, 20, -25, 7, 24, 3, -22, 26, 1, -1, 22, 17, 16, -29, 6, -4, -54, 5, -26, -9, -26, -3, -9, -35, -49, 6, 9, -6, -3, -42, -16, 27, 6, -8, -4, -40, 6, 38, 2, 0, -3, 27, 0, -21, -2, -13, 1, 0, -24, -6, 27, 7, 48, 19, -33, 12, 20, 7, 17, -2, -3, -6, -12, 29, -2, 2, 25, 0, -18, 25, 3, -12, -25, -23, -16, 4, -34, 4, -19, 0, -6, -3, -1, 31, -26, -50, 20, 1, 4, -19, 9, 1, -15, -1, 17, 5, -3, 5, -1, 7, -15, -16, 24, -33, -14, -12, -30, 22, 29, 4, 0, -9, -3, -23, -4, -18, 25, 24, 18, -6, 1, 0, -2, 27, 24, -2, -7, -4, -11, 25, -31, 59, 9, 3, -26, 13, 2, -4, -12, -2, 24, 36, -27, -4, -14, -24, -26, 17, 10, 1, 0, -37, -7, -11, -1, -7, 38, -8, -15, 17, 1, -36, 0, -15, 5, 26, -10, 0, 0, -53, 5, -8, 0, -22, 3, -1, -8, 11, 18, 3, -23, 27, 7, 23, 3, -7, -21, 3, -11, -46, -10, -49, 6, -13, 13, 6, 2, 27, 13, -3, 6, 14, -14, 4, -22, -6, 19, -41, 7, -4, -4, 24, 18, -56, 12, -3, -1, -3, 0, -1, 2, -10, -17, -16, 16, 1, -10, -12, -20, -20, 3, -30, 0, -19, -22, -9, 34, -17, -3, 0, 8, -11, 8, 15, 18, 39, 1, -26, 26, -1, -8, 6, 7, 9, -10, -44, -7, 26, -19, 20, -3, -20, -9, 1, 21, 5, -6, -53, -15, 17, -4, -3, -38, 7, 4, 10, 11, 21, 15, 6, 3, -20, -29, -6, -14, -4, 1, -11, -5, -18, 0, -13, 8, 15, 8, -4, 2, 29, 0, -21, 0, -13, -5, 6, -1, -4, 33, 13, -26, -2, 5, 7, -2, 49, -48, 1, -24, 1, -37, -27, 21, 12, 14, -1, 1, 27, 21, -17, 27, 16, -13, -1, 7, 0, 0, 12, 2, -1, 4, 7, 11, -7, -7, -2, -6, -28, 0, -2, -1, 1, 29, 18, 3, 0, 5, 2, -7, 21, 8, 15, -19, 8, -29, 18, 29, -11, -2, -11, -8, 0, -33, -10, -1, 7, 13, -16, 0, 1, -16, -3, 4, 10, -11, -18, -3, -8, -28, 7, 11, 0, -29, 8, -2, 0, -1, -23, 46, 0, 1, -7, 14, 4, 1, 7, -4, 22, 17, 42, 9, -8, -38, 7, 34, -2, -2, -4, 5, -19, 7, 31, 5, 5, -6, -1, 3, -5, 2, -1, 11, -20, -5, -1, 23, -3, 0, -3, 43, 7, 11, -8, -15, 5, -15, 6, 10, -18, 7, -20, 26, -17, 25, 2, 28, -15, 15, -11, -13, 36, -7, -7, 40, -2, -17, 18, -8, 7, 3, 41, -18, 9, -27, -8, -6, -40, 12, -3, 10, 4, 44, -39, 8, 2, 14, -3, 0, 49, -3, -3, 12, 40, 14, -8, 7, 39, -7, 0, -1, -11, 20, -19, -21, -7, 42, -29, -29, -7, 15, -14, 13, 8, 0, 14, 16, -22, 1, -4, -21, 5, 32, -22, 49, -3, -5, 2, 1, 22, 6, 1, 33, -12, -8, -14, -8, -26, -14, 33, 4, -10, 30, 5, -9, 24, -14, 7, -5, -8, -6, 24, 10, -22, -27, 3, 3, 22, -2, 15, 8, -8, -6, -5, -13, -16, 36, 28, -42, 13, 4, 18, -26, 15, 20, -1, -9, -7, 21, 18, -7, 24, 19, -4, -9, 4, 11, 25, -27, 5, -15, -14, -16, 3, -7, 10, -6, 6, -6, 23, -19, 6, 0, 4, -4, -5, 14, -1, 16, -3, 27, 12, -12, -3, 9, 20, -21, -10, 11, -27, 0, 2, 4, 8, 45, -29, -22, -5, 0, 34, 10, -76, -8, 7, 36, -28, -11, -7, -24, -5, -2, -10, -2, 2, 6, -7, -21, 12, 2, 21, -4, -1, 26, -3, -32, 38, 18, 32, -20, -5, 40, 0, 22, -14, 35, 5, 11, 11, 11, 4, -19, 0, -24, -5, 1, 24, -5, -14, -5, 27, 14, -8, 19, 10, 4, -19, 6, -8, 31, 6, -5, 5, -40, -5, 43, 5, -4, 17, 2, -3, 7, 11, -1, 3, -17, -31, 0, 38, -16, 4, 0, 0, -10, -7, 26, -8, -7, -14, -7, 12, 23, 2, 20, -27, 1, -6, 5, 2, 11, -36, -18, 3, -4, -16, 14, 0, -7, -2, -10, 6, -1, -2, -10, 19, -18, 30, 6, -18, 23, -27, -16, 22, 20, -24, 4, -5, 6, -7, 21, -30, -15, 50, 24, -7, -19, -6, 10, -20, 14, 21, 9, -8, -22, 7, -27, 22, -7, 11, -43, -27, -26, 4, 5, 24, -6, -29, -28, -4, -47, -21, 32, -18, -51, 14, 13, 2, -40, -3, -27, -2, 28, 20, 16, 25, 0, -10, 3, 7, 1, -17, 8, 10, 1, -23, -3, -35, 27, 8, -1, -2, -26, -8, -21, -26, 1, -8, -15, 15, 3, 38, 21, 7, -19, -53, -8, 2, 22, -4, 16, -2, 8, 4, 6, 0, 11, 22, -7, 8, 34, -5, 29, -3, 7, -5, 0, 6, -6, 14, 53, -2, 0, -20, 19, -5, 25, -1, -16, 0, -2, 0, -4, -1, 2, 19, 7, -21, 2, 13, -7, -12, -8, -29, -14, -5, -4, -9, 9, 8, -2, -10, 0, -31, 9, -6, -7, -57, 4, 19, -9, 11, 60, -1, -5, 29, 12, -27, -24, 8, -15, -1, 4, 9, -2, -47, -11, 1, -61, 1, 20, 16, 17, -21, -15, 23, -7, 6, 14, 2, -7, 17, 2, 7, -5, 6, -3, -21, 5, -22, 1, 19, -1, 58, 2, 0, 13, -11, -5, -5, 3, 35, -16, -46, 24, 10, 6, -26, 14, 25, 5, 4, -7, -15, 22, -29, -4, -12, -8, 0, 8, 31, 38, 8, -18, 21, -6, 26, -5, 0, -14, -28, 6, 3, -1, 40, -4, -38, 22, 1, 3, 2, 9, 4, -1, 5, -5, -15, 13, 0, -10, -17, 9, -28, -3, -10, -21, -27, -14, 16, 15, 36, -16, 0, 4, -9, -24, 33, -34, 18, -20, 10, 7, 3, -25, 8, 11, -22, -12, 4, -5, 6, -43, 36, -2, -6, -6, -11, -6, 6, 15, -35, 26, 15, -35, -6, -21, -33, -35, -10, -10, 12, -7, 11, 8, 10, 16, -6, -6, -23, -4, 9, 4, -27, 5, -5, 15, -10, -11, -3, 1, -80, -2, -1, 0, -30, 1, -1, -17, 23, -5, -1, 20, 5, -11, 13, 27, 0, 24, 1, -18, -18, 5, 25, -27, -24, -1, 6, 18, 3, -12, -21, -7, -7, -6, 36, 27, -2, -14, -3, -9, -2, -1, -1, 11, -11, 31, 1, 0, -8, 16, 0, 2, -5, 11, 1, -18, 3, -9, -5, -13, 3, 13, -9, -19, 4, -10, 5, 30, 25, -37, -4, 9, -8, -38, 13, -5, 7, 17, 12, -7, -2, 8, -12, 16, -16, 2, -4, 4, 4, -9, -10, 4, 3, -2, 3, 13, -4, 4, -3, -19, -33, -13, -6, 19, -13, -28, 0, -10, 12, -2, 8, 4, 3, -11, -4, 17, -14, -34, -24, 6, -51, -2, -5, 1, 1, -25, -7, -6, 6, 6, -8, -2, -35, 5, 8, -33, 8, 2, -29, -68, 3, 1, 10, 7, -7, -14, 1, 0, 10, 37, -34, -31, -14, 4, 1, 10, 18, 13, 17, -34, 10, 2, -18, 17, -3, 5, 1, -2, -4, 0, 23, -53, 44, 45, -2, -7, -17, 14, -7, -7, -4, 30, -23, -27, -3, 23, -2, 10, 50, 18, 21, -23, 31, 5, -8, -4, -12, 4, -1, 5, -6, -10, -3, 22, 40, 20, 38, 18, -2, -18, -46, 44, -32, -8, 0, 28, -13, -11, 0, -24, 3, 56, 16, -6, 8, -31, 1, 8, 15, -9, 6, -9, -16, -62, 5, -26, -11, 0, 17, 4, 8, 1, -3, -6, 40, 0, -25, -7, 5, -5, -1, 12, -11, -3, 8, -7, -9, 7, 6, -13, -38, -3, 7, 10, -6, 17, -5, 29, 7, 24, 24, -25, 19, -18, 0, 14, 0, 3, 30, -14, -13,
    -- layer=2 filter=0 channel=4
    -32, 3, 5, -22, 10, -2, 5, -7, 8, 5, -43, 4, -24, 8, -4, -7, 4, 10, 22, 18, 12, 6, -6, -28, -8, -6, -18, -4, -69, 1, -11, -4, 15, 15, -14, 22, 0, 17, 16, 26, 23, -8, -29, 44, -15, 1, 1, -12, -2, 38, -20, -42, -9, -78, -39, 0, 22, -47, -36, 18, -1, 25, 1, -3, -2, -11, 16, -14, -14, 26, -2, 0, 3, -8, -25, -26, 15, -1, 0, 27, 15, -9, -4, 1, 15, -9, -19, -2, 11, 7, 4, -2, -40, -18, 1, -2, -6, -60, -1, -26, -25, 13, -5, -53, -7, 17, 1, 29, 7, -8, -57, -11, -26, -31, -29, -17, 14, 2, 0, 7, 13, 5, 0, 12, -7, -38, 18, 23, -6, 2, -8, -23, -14, 23, 1, -20, -1, -5, 22, -5, 16, -5, 0, 0, -4, 6, -11, 11, 31, 3, -3, 31, 3, 0, -4, 2, -80, 8, 18, -1, -4, -19, 1, 17, -35, 20, 5, 3, 36, -11, -25, 32, 6, -2, 4, 5, 35, 14, -36, -31, -41, -55, -20, -7, 16, -27, -33, 21, 5, 14, 16, 10, -13, -1, -2, -42, -47, 6, -11, -4, 19, 23, 5, -7, 3, -8, -10, 1, 3, -17, -1, -9, 3, 10, -21, -6, 21, -3, 33, 27, -3, -3, 6, -2, -1, -4, 5, -27, 9, 8, -1, -10, -6, -14, -15, 0, 3, -5, -25, -21, -20, 5, -12, -17, -4, -18, -13, -20, -3, 7, -3, -20, -25, -29, 15, 1, 6, 6, -18, 16, -44, -1, -14, -24, 11, -14, -24, -2, -16, -26, 12, 5, 0, 16, -11, -12, 26, -1, 1, 55, -13, 5, -2, -1, -87, -8, -19, 3, 6, 9, 13, -8, -20, -10, -6, -10, -1, -39, -21, 34, -4, -2, 5, -18, 44, -33, -8, -8, -28, -19, -36, -2, -8, -33, -20, 13, 1, -29, 9, 0, -17, -16, 11, 11, 6, 20, 9, -2, -28, -16, 14, -7, -30, 0, -19, -24, -11, 11, -16, -4, 8, 25, 10, -11, -18, -3, 7, 6, -11, 12, 4, 30, -4, 10, -1, -11, -15, 1, 4, -14, 5, -15, 1, 7, 6, -1, -27, -16, 4, 9, 20, -19, 12, 26, 1, -51, -10, 0, -41, -54, -1, -63, 1, -11, 4, -6, -33, -19, 0, -14, -17, -12, -3, -20, -9, -2, -11, -33, 1, 4, 1, -3, -40, 8, 60, -1, 0, 15, -21, 5, -26, 0, -70, -5, 26, -2, 23, -1, -11, 15, -43, 25, -3, -40, 20, 15, -14, 51, 0, -3, -2, -2, 39, -19, 0, -26, -23, 28, -9, -2, 10, -39, -21, 19, -3, -21, 23, -1, -19, 9, 23, -46, -16, 44, -35, 7, -1, -9, 18, -56, -28, -1, -65, -14, 13, -11, 33, -10, 25, 19, 56, -10, 2, 0, 22, -2, 6, 25, 3, 57, 2, 15, 0, 3, -26, 4, -3, 11, 1, -21, 0, 2, 1, 2, 8, -14, 9, 6, -9, -19, 18, -7, -5, -9, -30, 0, -32, -18, -8, 22, 12, -3, 15, -9, -2, 24, -54, -9, -17, -7, -2, -15, 36, -7, 17, 1, -5, 2, 1, 25, -6, -29, -28, 2, 3, 42, -13, -1, -35, 2, -53, -18, 18, -6, 4, -12, -13, 26, 8, 8, -8, 8, 18, -2, -76, 26, -17, -1, -9, -28, 13, -1, -22, -56, -52, -22, 2, 4, -28, -63, -34, 3, 5, 10, 27, -13, -14, -4, 21, -20, -9, 43, 6, -2, 27, -25, 8, -68, 27, 0, -25, 6, 1, -8, 13, 7, 5, 25, 10, -7, 16, -4, 15, -24, -19, -17, -1, 52, -1, -19, -3, 19, 4, 3, 0, 10, 0, -48, -19, 3, 0, -5, -30, 0, 32, -13, 19, -8, 22, 13, -6, -6, 7, -2, 23, 13, -5, -71, 1, -27, 3, 4, -8, 73, -30, 0, -15, -11, -8, 5, 21, -2, 2, -24, 5, 4, -1, -12, -59, -27, 32, -1, 0, 29, -21, 4, -11, 3, -39, 1, -7, 7, 30, -6, -10, -11, 1, 1, -18, 10, 29, -14, -32, 29, -30, 4, 0, -2, 11, -1, -21, -11, -37, 33, 9, -8, -27, -13, -8, -3, -3, 6, -10, -3, -27, -6, 14, -43, -30, 21, 5, 2, 5, -36, 14, -62, -7, 3, 13, -21, -10, -16, 13, 0, 4, 10, 18, 0, -5, 1, 13, 1, -27, 16, -2, 25, 0, -11, 5, -10, -26, 29, 2, -21, -6, -35, -4, 3, 0, -5, 1, -20, -3, 0, -12, -18, 18, 28, 27, -9, 4, 3, 30, -33, 3, -85, -9, -16, -15, 1, -23, 44, -51, -1, 31, -18, 1, 54, 52, -2, 11, -15, -1, 0, 0, 15, -9, 3, 30, -3, 0, 18, -25, -1, -43, 3, -79, -44, -8, -2, 5, 2, 11, -20, 24, -2, -9, 28, 46, 6, -29, 27, -6, 2, -3, -20, -11, -1, -1, -20, -27, -66, -20, 2, -79, -15, 3, 3, 1, 25, -30, 16, -3, -20, 36, 7, -18, 4, -14, 2, -25, -24, 20, 13, 29, -5, -45, 18, -2, -10, 41, -24, 10, 3, 12, -23, -8, -2, 24, -13, -31, 0, -6, 18, -2, -7, 0, 1, -11, 23, 7, 6, 7, 2, -9, 22, -4, -1, -2, -11, 17, 11, -48, -10, 2, -18, 45, -9, 21, 4, 18, 7, -14, -21, -4, -31, 6, 0, -10, 1, 1, 4, 26, 17, 10, 11, 10, -2, 10, 24, 4, 5, -4, 38, 45, 22, 15, 3, 1, 16, -23, -7, -12, 13, -72, 12, 11, 2, -4, -15, 38, 0, -25, 10, 3, -1, 30, -18, 29, 38, -1, 2, -4, 10, 11, -7, 18, -1, -9, -76, -23, 2, 13, -9, -30, 5, 5, 0, -5, -30, -25, -2, 16, 26, -5, 16, -23, -3, -7, 10, 9, 0, 3, 4, -25, 32, -23, 17, 13, -14, 14, -3, 50, -6, 14, 0, 6, -14, -2, -10, -5, 43, 0, -7, 0, 10, 3, 18, 4, 49, 4, -4, -11, 17, 0, 6, 12, -41, -19, -9, 9, -19, -3, -9, 6, 15, -15, 0, -13, 5, -12, -5, 9, -6, 1, 0, -20, -17, -15, 14, -1, -29, -2, 10, 40, -8, 21, -11, 3, -1, 4, 9, 20, -3, 9, -4, 4, -13, -18, 5, 0, 0, -79, -7, 0, -3, -4, 20, 36, -20, -22, 2, 7, -28, 7, -2, 4, 10, 2, -6, 0, -5, 25, -37, -20, -24, -5, -63, -19, 4, 11, 38, -22, 1, 0, -10, -14, -19, -27, -5, 4, -21, 13, 7, -15, -4, 18, 69, -6, -5, 22, 2, 15, -19, 1, 8, -23, -22, 5, -6, 24, -11, -9, 4, -4, -20, -8, 6, -9, 9, -1, 33, -5, -3, 39, -4, -7, -18, -3, -42, 0, -5, 5, 6, -18, -27, 7, -2, -39, 2, -18, -13, 37, -9, 9, 0, -24, -48, -10, -50, 17, -19, 2, 0, 1, 6, -34, 8, 1, -22, -7, 25, 18, 1, 0, 0, 3, -7, -4, -4, -10, -44, -39, -8, -2, 33, -15, 4, 14, 2, -69, 8, 4, 6, 15, 17, 14, -2, -39, 5, 4, -9, -26, -3, -46, -1, 19, 3, 1, 7, 15, -31, -29, -70, -61, -14, -13, -7, -4, 0, -43, 12, -5, -10, -30, 3, -34, -21, 25, 41, 13, -8, -22, 6, 5, 23, 25, -36, -6, 3, 31, 10, 7, 0, -14, -2, 18, -11, 29, 4, 5, -3, 22, 6, 19, 21, 3, 23, -3, 48, 2, 10, 42, -7, 3, -21, -5, -6, -20, 6, 4, 1, -9, -14, 21, 46, 14, -21, 14, 29, 14, -17, 24, -1, -4, -74, 18, -3, 28, -8, 41, 0, -20, 38, -57, 21, -18, -36, 6, 5, 9, -4, -17, -19, 5, 6, 2, 61, -23, -14, -58, 4, -3, 7, -31, -4, -13, -11, -47, 7, 11, -7, 21, 0, -20, 2, -9, 8, 0, -25, -6, -4, -44, 38, 9, 4, 4, -20, 18, 21, 0, -70, -56, -11, -6, 5, -37, 0, -29, -10, 8, -29, 6, -2, -32, -36, 12, 39, -10, 1, -7, 5, -17, -10, 13, -77, -25, 2, 2, -17, -18, -29, -5, 3, 12, -20, -29, 4, 20, 1, 11, -2, 45, -16, 5, 21, -4, 51, 14, -6, 9, 3, 6, -63, -5, 11, -31, 17, -4, 4, 1, 13, -29, 32, -31, 0, 31, 18, 16, -11, -23, 6, -6, -76, 23, -27, 36, 7, 32, 6, 6, 30, -49, -10, 14, 8, 0, -3, 40, -5, 39, -30, 0, -5, -5, 8, -15, -31, 33, -9, -2, 2, -2, -6, -6, 7, -41, -16, -10, -4, -9, -6, -32, -11, -22, 14, -16, -8, -12, 15, -28, -8, 8, 1, -3, -35, -5, 29, -14, -40, -6, 34, 9, 0, -34, -1, -46, -13, 8, 0, -22, 6, -9, -10, 10, -10, 15, 6, 0, 7, -44, 36, 8, -64, -26, 1, -23, -45, 4, 6, 35, 11, 23, -15, 16, -18, -55, -6, -11, -45, 28, 33, 3, 15, 4, 23, 16, 12, 7, -4, -6, -32, -1, -23, -10, 12, -6, -5, 6, -6, 23, 37, -10, 11, 23, 34, 0, -20, -15, 5, 20, -39, 6, -72, 25, -15, 40, 5, -7, 52, -20, -9, 2, 3, 6, 6, 70, -2, 24, -2, 5, -6, -3, 9, -53, -2, 6, -2, 2, -49, -10, -2, 23, 7, -14, -36, -24, -7, -3, 24, 6, -21, 3, 2, -6, 20, 5, 19, -50, 26, -19, 2, -4, -35, 19, 15, -38, -53, -21, -2, 36, 3, -34, -26, -1, -12, -9, 8, 20, -5, -2, -1, -14, 16, -15, 3, -22, -2, -2, -47, 1, -51, -39, -9, -50, -39, 50, -17, 11, -17, -9, -10, -1, -7, -22, 5, 3, 0, -24, 29, -5, 20, 4, -1, 7, -5, -2, -24, 5, 0, 1, 9, 7, 5, -1, 6, 14, -29, -17, 9, 17, -13, -8, 14, -6, -12, 31, 6, 19, -34, 13, -65, -11, -2, 1, -3, -22, 61, 38, 10, 23, -24, 7, 5, -8, -3, 31, 20, 8, -6, -4, 19, -1, -39, -1, 0, 4, 2, -4, 0, 20, -5, -27, 13, 12, 4, -18, -2, 13, 4, 4, -25, 7, 15, -10, -16, -32, -4, -24, 7, 2, -51, 12, -2, -36, 12, 0, -7, -17, -8, -30, 0, 4, 0, 6, -13, 4, -8, -18, -36, 12, 21, -36, -9, -22, 2, 28, -25, -2, -41, -9, 0, -18, -21, 21, 2, 22, -17, -8, -10, -27, -9, 20, 3, 47, 4, -7, -22, -4, 23, 1, 7, 10, -11, 18, -24, -6, 6, -5, -12, 16, -5, 2, 0, -17, -23, 0, -19, 60, -34, -11, -4, -19, 46, -7, -4, 7, -33, -1, -37, 0, 18, 14, 6, 19, -8, 29, -18, 19, 10, 11, -16, 21, 0, -6, 26, 9, 5, -5, 7, 43, -6, 24, -3, -4, 15, 12, -4, -3, -3, -74, 3, 11, 3, -18, 2, 15, 8, -5, 23, 26, -9, 42, -5, -4, 25, -5, -6, -4, -14, 21, -13, -3, 4, -52, 0, 0, 7, 8, -38, -10, 30, -5, -58, 18, -7, 6, 19, 3, -50, -16, 20, -16, -2, -15, 2, -15, 0, -26, 2, 17, -2, -20, 15, -9, 33, 2, 10, 3, -17, -9, 7, -17, -20, -11, -18, 3, 12, -7, -9, 5, -28, 22, 2, 0, -20, -1, -32, 0, 12, 5, -4, 34, -16, 23, -18, 6, -2, 5, -36, -3, 32, -3, -5, -49, 19, 18, -23, 3, -18, 15, -6, 2, -4, -5, 15, -5, 14, 17, 18, -2, -6, 7, 15, 2, 2, -8, -1, 39, 15, 11, 3, 3, 13, 0, -1, 12, 1, -80, -22, 3, 7, 6, 30, 4, 3, -12, -8, 38, 0, 40, -26, -2, -17, -8, -4, 0, -3, 40, 7, -10, -35, -6, 28, 5, 4, 26, -84, -23, 15, 10, -10, -4, 5, -16, 18, 0, -22, -7, -15, -15, -4, 26, 47, 11, -54, 0, 6, 17, -36, 4, -5, 4, 23, -1, -11, -13, -6, -7, 1, 36, 9, 1, -8, -5, 0, -9, 7, 4, 13, 9, 0, 1, -62, -1, 2, 29, -11, 1, -6, 20, -3, 8, -27, -9, -11, -5, -1, 15, -5, 10, 4, -33, 24, 28, 33, 0, 3, 34, -5, 5, 16, 0, 22, -6, -20, 8, -4, 16, 4, 4, 13, 0, -1, 7, -14, -1, 11, -45, 0, -6, 19, 8, 1, 11, -5, -83, -1, -34, 5, 23, 30, -20, 5, 4, -10, 20, -2, -32, 0, -10, -41, -9, 1, -7, 5, -27, 28, -43, -24, -32, -18, 30, 0, 22, -29, -4, -12, 8, 19, -3, 7, -3, 41, -2, -32, 1, -16, 25, -5, -5, 22, -54, -7, -9, 0, 7, -4, 17, -20, -24, 36, 12, -20, 25, -7, -45, 5, 1, -22, 11, 10, -3, -28, -4, -12, 1, 22, 11, -7, 2, -71, 6, -9, 15, 13, -5, 4, 32, 4, 8, -34, 0, 45, 0, -1, 22, 27, 25, 2, -3, 4, -8, -46, 29, -11, 21, 0, 17, 34, -18, 14, -31, 37, -1, 14, -5, 5, 3, -12, -3, 6, -3, 18, -3, 11, -50, -5, -7, -3, 0, -3, 6, 0, -34, 16, -19, -8, 4, 1, -19, 13, -5, -2, -6, 11, -16, -38, -41, -16, -8, 0, -5, 30, -19, 15, -6, -9, -6, 22, 50, 0, -14, -59, -13, 8, -4, 15, 14, 6, 26, -23, 8, 0, -6, -23, 16, 4, 0, 8, -14, -32, -32, 1, -21, -8, 20, -11, -55, 28, 6, -54, 0, 1, -18, -3, 32, 5, 29, 58, -5, -2, 7, 27, -2, 16, 13, -1, -1, -52, -3, 19, -1, 18, -4, 5, 39, 28, -25, -49, -20, 19, 19, 20, 18, -13, -5, 8, -14, -2, 11, -11, 14, 0, 27, 2, 18, 19, -34, -13, 4, 6, 3, 0, 20, -5, 12, 6, 0, -4, -4, -10, -18, -13, -29, -6, 7, 10, -28, 3, -16, -7, 25, 12, -11, -6, -2, 20, -19, 0, 10, -31, 6, 12, -43, 9, -43, 6, -37, -7, -11, -8, 2, -41, -7, -59, -14, -61, 45, -9, -8, -17, -25, -7, 2, -11, -21, -4, 17, -47, -4, -17, -6, -12, 33, 6, 22, -5, 1, -16, 3, 2, -27, -14, 11, 1, -26, 22, 8, -54, 10, 5, 24, 5, 17, 0, 5, 19, 4, 4, 3, 30, 16, 28, 28, -28, 3, 8, 0, -37, -14, -4, -6, 0, -7, 11, -39, -2, -58, 10, 14, 16, 15, -46, -23, -3, 54, 12, 14, -32, 6, 22, 15, -1, -4, 54, 2, -43, 7, 34, 8, 26, -1, 0, 10, 5, 0, 2, 5, -12, -20, -24, -3, 0, -7, -1, -16, -5, 24, 6, 25, 2, -41, -7, 17, 30, -2, -7, 1, -4, 33, -10, -22, 10, -35, -20, -17, -5, -9, 25, -12, -36, -18, -45, -40, 19, 23, 4, -16, -21, 16, -8, 6, -38, -15, 6, -2, 10, 16, 23, 30, -7, 5, 0, 2, -12, 1, -10, -28, 0, 31, 4, 25, -9, -25, 19, 4, 1, -4, -9, 0, -4, 36, 1, -6, -6, -2, -22, -7, 38, 5, -12, 22, -22, -1, -17, -1, -25, 18, 0, -2, 4, 17, 10, -18, 4, -19, -12, 9, 19, 4, 1, 34, -5, 40, -2, 50, 25, 20, 36, -4, 6, -13, 55, -9, -30, 39, 19, 10, -19, 22, 0, -25, -7, -2, 2, -3, 31, -30, -10, -5, 1, -9, -3, -12, 4, -52, -5, 15, 16, -29, -1, -19, 24, -12, 9, -7, -28, 2, 34, 49, -7, 4, 23, 8, 3, -3, -46, -2, 26, -3, -5, -8, 21, 10, 3, -23, -6, 17, -6, 5, -19, -19, -16, -32, 2, 17, -34, -13, -5, -16, -3, 6, -76, 22, 2, 2, 4, 8, 15, -7, 9, 8, 29, 7, 21, -9, 12, -2, -2, -37, 15, -4, -10, 6, -63, -2, -1, -7, 1, 2, -3, -1, 0, 0, 9, -6, 4, -3, 2, 37, -29, -12, 5, -3, -47, 20, -18, -19, -27, -3, 2, 0, 6, -7, -19, -18, 10, 29, -7, 13, -27, -1, -3, 3, 11, 4, -14, 55, -6, 0, -21, -7, 6, -8, 7, 17, -12, -10, -6, -1, -3, -8, -8, -9, -6, -29, -20, -23, 7, -8, -12, -15, 21, 6, 8, 31, 4, 11, 24, -7, 3, -10, 1, -4, -23, 23, 27, 27, 0, -20, 55, 6, -4, 1, 8, 10, 3, 4, -40, 5, 9, -46, 15, 0, 13, -31, -9, -60, 0, -1, -11, -2, 28, -22, -10, -15, -26, -18, 15, 13, 15, 0, 21, -12, -4, 3, 2, 50, 17, -20, 16, -5, 3, -8, 31, -3, -7, -9, 1, 7, -26, 2, -3, -12, 15, -3, -2, -8, -21, 9, 11, 33, 38, 0, -35, 0, 13, 3, -2, -10, 0, 60, -32, 16, -22, -4, -1, 7, 6, -7, -22, -1, 11, 9, 17, 43, -1, -21, -2, 4, 0, -4, -16, -11, 49, -20, 0, 4, 25, -15, 0, 12, -5, -41, -12, -11, 5, 26, 33, -6, 1, 10, 37, 29, 20, 37, -10, -38, -9, 9, -9, 6, -20, -22, 16, 1, 30, -33, 3, -10, 0, 7, -5, 20, 34, 7, -9, -2, 5, 0, 22, 1, -13, 4, 0, -20, 1, 6, 0, -19, -26, -61, -4, -12, 5, -2, 39, -3, 34, -1, -15, 20, 10, -7, 6, 46, 1, -8, 15, 2, -16, 3, -8, 2, 29, -14, -4, -3, -30, -6, -50, 32, -13, -4, 2, -32, -15, 22, -62, 21, 31, -4, 5, 6, 1, 20, -3, -27, -31, 12, 22, 16, -7, 11, 1, 8, -6, 18, 3, 0, 1, 9, 22, -39, 0, 0, 8, 2, 0, 0, 7, 0, 39, -70, -4, 2, 28, -30, 0, 1, -1, -19, 3, 0, 0, 36, 21, 19, 9, -9, -8, 41, 9, 4, -15, -1, -11, 4, -9, -4, 7, -15, -1, 25, 16, -25, -10, 28, -7, -10, -49, 13, 29, -8, -18, -30, 0, -4, 5, -14, -21, 35, 21, -1, -6, 21, 10, -46, -8, -14, 5, -10, 24, 11, 6, 15, 39, 13, -13, 21, -2, -18, -1, -2, 8, 30, 5, -7, 22, 5, -24, 8, -1, -10, -18, -1, -6, 4, 10, 3, -19, -5, 7, -3, 2, -21, -32, 59, 35, -3, 46, 10, 8, 44, -4, -22, 10, 7, 58, 31, 37, -17, -8, 10, 38, 7, -34, 0, 23, 2, 14, -2, -5, 2, -6, 3, -3, -6, -51, 0, 23, -95, -8, -1, 30, -24, -1, 8, -3, 1, 17, -7, -3, 24, 31, 12, -46, 21, -3, -20, 19, 2, -8, -22, -20, -32, -10, 2, 8, -32, -31, 31, -6, 5, 13, -7, -5, -6, 9, -3, 15, 4, -37, -59, -10, -6, -77, -17, 10, 1, 1, 14, -6, 11, -3, -77, -9, -47, -7, 33, -3, 14, -12, -16, 43, 14, -91, 17, 8, -59, 3, -64, -40, -34, -37, -1, 6, -9, -42, 10, 3, -15, -42, -3, -6, 3, -24, 35, -33, 3, 6, 7, 18, -76, -74, -13, 14, 1, 31, 12, 29, 25, -2, -14, 29, -40, 9, 7, 0, -11, 5, 48, 5, 48, 4, 32, 61, 17, 39, 68, -8, 9, 0, 0, -3, 0, -7, -8, -1, -64, 2, 6, 5, -13, 7, 37, -2, 12, 21, -6, 2, 26, 13, -9, -49, -17, 6, 3, 32, -7, 17, -26, -2, -30, -4, -4, 1, -20, -46, 28, 4, -19, -2, 7, 2, 18, -37, -3, -5, 7, -9, -25, 4, 6, -7, -12, -22, 5, -5, 16, -3, 27, 0, -33, -1, -9, 1, -50, 14, 24, -23, -32, 14, 0, -80, 31, -5, -45, -1, -9, -19, -26, 43, -6, 5, -5, -70, -2, 13, -25, -31, 4, 43, 0, -2, 38, -38, -5, -3, -21, 17, -24, -57, 6, -5, -7, 40, 31, 25, 8, -4, 9, 54, -4, 16, 16, 23, 10, 2, 26, -14, 1, -2, 5, 13, 7, 22, 11, -2, 2, -11, -1, 5, -4, 5, -6, -6, -28, 3, 0, 17, 9, 0, 20, -4, 4, 2, -4, 5, 8, 6, -8, -4, -1, 37, 38, 6, -14, 1, 0, 0, -16, 4, 1, -10, -22, 21, -32, 13, 1, 2, -1, -1, 5, -10, 17, -20, -2, 11, 5, 0, -7, -1, 17, -2, -22, 12, -21, -3, 0, -19, -51, -26, -18, -3, 7, 5, 4, -12, 9, 8, 1, -12, 5, -14, 12, -7, 3, 33, 14, 47, 1, -10, -5, 0, 14, -54, -3, -6, 2, 34, -3, 8, 28, -7, -6, 1, -29, -15, -7, -13, 9, 10, 0, 21, 10, 14, 35, -1, -1, 31, 14, 69, 5, 5, 20, -9, 0, 14, -34, -24, -15, 30, 14, -6, -35, 0, 13, -14, 5, 1, 5, 22, -19, -24, -45, -2, -1, 18, -21, -7, -5, -15, 29, -4, -24, -4, -26, -8, 15, 9, -63, -22, 45, -2, -15, 36, 28, 50, 0, -2, 0, -16, 42, 6, -11, -7, -1, 21, 29, -2, 4, -53, -24, -20, -10, -13, -10, -10, -47, 34, 2, -14, 17, -4, -14, -5, -6, -22, 14, 33, -47, 0, -61, 10, -55, 14, -12, 19, 9, 14, -5, -3, 47, 0, -13, 23, 1, 51, 2, 4, 2, 22, 2, -27, 13, -22, 6, 45, -2, -41, -11, 2, -1, 3, 17, -8, 27, -10, 43, -1, 13, 5, 8, 9, 11, -8, -38, 4, 15, 12, 5, 9, 24, 3, 9, 54, -11, -15, 5, -3, 0, -17, 2, -3, -6, -18, -3, 6, 0, -33, 15, -23, 44, 2, -4, 25, -4, -8, -14, -3, -48, 4, 0, 0, -18, -4, 4, 31, 17, -17, 68, 26, -4, 0, -28, -37, 0, 4, -2, -29, 0, 8, 11, 0, -63, -50, 0, -4, -11, -20, -5, -4, 7, -49, 36, 21, -38, 16, -17, -15, 3, 8, -21, 0, -10, -35, 6, 12, -79, 3, 11, 8, -24, 2, 25, 45, -4, -1, 9, 3, 23, 3, 2, 59, -3, 10, -4, 7, 3, -9, -11, -8, -25, 6, 5, 22, 0, -61, -3, 3, 7, -2, -15, -12, 50, -11, 23, 13, 4, -1, -27, 0, 67, 6, 16, -46, 19, 19, -7, -8, -1, 2, 11, 26, -6, -18, 15, 3, 0, -2, 39, -1, 17, -1, 7, 0, -7, 31, 0, 11, -14, -2, -7, -2, -17, 0, 22, 6, -36, 10, -3, -3, 22, 10, -18, 14, 27, 9, 1, 23, 18, 9, -17, -25, 6, -8, 0, 5, -50, -4, 36, -5, -33, -56, 2, 0, 10, -21, 12, 18, 0, 0, -3, 20, -43, 14, -15, 18, 25, 0, -23, -2, 16, 7, -4, 11, -37, 0, -53, -32, 3, 6, 38, 16, -13, -8, -3, 17, -2, -5, 3, 17, 5, -14, 7, 6, 2, 12, -3, 6, -11, -23, -5, 56, 0, -37, 18, -19, 3, -2, -5, -1, -22, 7, 14, 0, 18, 9, 13, 11, 25, 0, -16, -9, 80, 53, 6, -4, -19, -8, 3, 3, -21, -26, 3, -13, 16, 26, 41, -1, 8, 2, 0, 0, -1, 23, 13, 32, -41, 3, -5, 17, -20, -2, 36, 1, -4, -11, 0, -5, 1, 18, 22, -38, 5, -16, -16, -28, 1, -46, -12, -9, 34, -5, 0, 0, -21, 1, 45, -10, 22, -18, -6, 3, -4, 1, 7, 10, -1, 10, 1, -1, -15, -12, -25, 26, 2, 0, -9, -1, -6, -8, 9, 13, 1, 0, -23, 25, 23, -23, 10, -4, -4, -14, -3, 6, -18, 0, -7, 17, 9, 31, -3, 0, -1, 29, 2, -11, -30, -14, 6, -36, 0, -22, 22, -36, -3, 6, 8, -15, -56, 7, 22, -22, -26, 25, 25, -15, 28, 5, -38, 10, 6, 23, -15, 13, -17, -1, 14, -7, -89, -6, -33, 2, 6, 14, 10, -3, -18, -43, 8, -4, 0, 2, -58, 33, -66, 4, -6, 35, -12, -7, 15, -7, 31, 31, 49, -1, 2, 15, 22, -92, 31, -8, -75, -23, 20, -39, 37, 32, -21, 1, -7, -18, -55, -23, -7, 13, 68, 0, 0, 1, 8, 17, 41, 25, -2, -10, -45, 18, -25, -18, -2, -11, 0, 3, 3, -5, 34, 2, -43, -18, -66, -3, -12, -19, 15, 27, -27, -6, 14, -27, 17, -6, -73, 2, -37, -47, 60, -44, 6, 9, -7, 15, 16, 0, 8, -13, 2, -27, -7, -28, 16, -25, -10, 1, 8, -13, -118, 15, -35, 0, -7, 10, 29, -2, 15, -4, 0, -22, -32, 7, 4, 6, -34, -5, 12, -21, -18, 1, -10, 42, 10, -2, -10, -7, 13, -13, -4, 4, -7, -32, -2, 26, -58, 2, 0, 1, -8, -3, 20, 4, 37, 6, 30, 6, 12, 20, -2, -43, 2, -15, -23, 33, 11, -21, 0, 37, -4, -3, 6, 0, -41, -1, 3, 15, 7, -24, 36, -4, 37, -15, 11, 20, 11, 14, -54, -1, -18, -28, -10, -11, 44, 29, 15, 4, 47, 12, -18, 10, -1, -6, -19, -22, 4, 22, -6, -25, 10, -35, -5, -3, 0, -4, -40, -11, 33, -2, 0, 36, -5, -21, -3, 34, 5, -5, 5, 3, -5, -10, 19, -39, 4, -2, 35, 20, -79, 5, 28, -6, -15, 7, 7, -18, 22, 6, 10, 3, 18, 5, 12, 21, -27, -1, 21, -22, 8, -29, 7, -14, 8, -12, 13, -6, -15, -12, 4, 2, 2, -32, -19, 3, -14, 2, 0, -8, 6, 4, 0, -3, 1, 19, -2, 6, 16, 10, -1, -14, -13, 6, 33, 19, 11, 1, -24, 17, -7, -3, 2, -10, -7, 5, 18, -46, 10, 46, 20, 6, 0, 4, -10, -5, -5, -29, 17, 28, -15, -2, -9, 1, -14, 9, 23, -5, 14, -20, -21, 15, -7, 7, 20, -11, -7, 39, 23, 0, 4, -23, -6, 13, 20, -7, -12, 13, 5, 18, 1, 15, 6, 6, 2, 34, 1, -24, 5, -53, 1, -40, 12, -10, -1, -4, 8, 0, -31, 5, -13, 0, 2, 14, -8, -5, 35, -5, -18, 17, 32, -26, -1, 0, -1, 2, 27, 38, -5, 4, 17, 37, 10, -9, 7, -6, 13, -4, -1, 7, 6, 7, 1, -16, 10, -7, -9, 7, -12, -3, -6, 0, -8, 2, 1, -5, 10, -5, 16, 11, -12, -18, -2, -24, 9, 17, 24, -6, -15, -2, 2, -11, 29, -45, -16, -30, 18, 27, 21, 0, -6, -28, -12, -7, -7, 1, 9, 13, -35, 10, 17, -26, 2, 15, -20, -2, -6, -5, 23, -8, -41, 2, 26, -9, -2, -4, 45, 18, 17, 44, 6, 17, 25, 5, -1, 0, 14, -22, 1, 25, -2, 21, -1, -4, 28, 3, -2, 26, -3, -26, 7, 26, -4, 0, -8, -23, -6, 1, 22, 2, 30, -34, 3, -18, 58, -6, -18, -6, 6, 31, -7, -26, 3, 0, -2, 55, 27, -33, -3, 4, 7, -3, 47, 5, 0, 25, 10, 2, 3, -12, -7, -6, 6, 0, -5, 3, -1, -1, -13, 0, -49, 3, 6, 1, -2, 3, 23, 34, -43, 36, 42, 19, 19, 0, -69, 8, -14, -8, -5, -46, 6, -41, 45, 0, -74, -100, -4, 0, -8, 9, 3, -11, 8, -47, 6, -2, -15, -27, -18, 8, -16, 16, -16, 0, 14, -23, -9, -45, -39, 0, -51, 8, 26, -11, 16, 5, 0, 20, 23, 2, -31, 0, -30, 20, -18, -2, 6, 45, -1, -15, 6, 32, -6, 9, 2, 7, -6, -27, -5, 1, -1, -5, -10, -14, 11, -5, 10, -37, 15, -10, -17, -24, 33, -4, 2, 26, -22, -6, -2, 5, 36, 1, 25, 6, -11, -18, -13, 43, 5, 10, 12, 0, 13, 6, -4, 3, 3, -26, 3, 23, 0, 5, 4, 24, -6, 4, 7, 0, 8, -6, 0, -7, 5, -8, -15, 7, 10, 2, 1, 25, 0, 0, -61, 16, 0, -9, -11, -10, -14, -29, -16, -22, -15, -5, 8, 2, 22, -13, -32, 9, -12, 4, 37, -13, -29, -31, 2, 22, 0, 17, -16, 0, 14, -34, 31, -3, -31, 1, -10, -2, 40, 47, 19, -22, 0, -7, 15, -6, -20, -1, 27, 26, 20, -3, -3, 32, -3, -54, 1, 9, -25, -13, 5, 42, 1, -24, -8, 1, 0, 6, 16, 14, -11, 16, 41, -11, 8, -30, -20, -2, 39, 7, -1, -24, -8, 8, 18, 17, 19, 0, 34, -4, -21, -42, -4, 21, 3, -8, -8, 0, 0, 0, 0, 7, -4, 32, 12, 7, -35, -7, 0, 47, -7, -9, 5, -3, 19, 17, 18, 1, 2, -3, 8, 0, -8, 36, -20, -10, 9, 5, -37, 8, 36, -6, -1, -69, 10, -13, 17, -12, 5, -70, -16, 0, -14, -17, 23, 11, -8, -35, 33, 25, -39, -4, -11, 60, 0, 12, -13, 5, -4, -31, 54, -41, -5, 5, 3, 23, -4, 36, 21, -16, 5, 39, 40, -7, 48, 2, 0, 4, 12, 2, -4, 22, -3, 13, 12, 16, -19, -13, 0, -8, -7, -31, -6, -24, 6, 6, 13, -3, 26, 28, 25, -23, -9, -12, -8, 39, 56, -5, -32, -29, 1, 73, -5, 10, 12, 1, 42, 8, -45, -27, -12, 18, -17, 6, -8, 1, -9, -31, 11, 0, -3, -7, 34, 39, -20, 5, -5, 57, -19, 0, 12, -10, -38, -18, 4, -1, -3, -25, 13, -15, 30, -42, -55, -9, 7, 32, -24, 8, 1, -9, -15, -1, -10, -19, 23, 3, 8, 27, -13, -6, -3, 9, 14, 22, -6, 6, 10, 12, -8, -15, -8, 17, -9, -16, 26, 5, -12, -13, -9, -9, -56, 0, -42, -44, -8, 31, 2, -55, -9, 1, 19, -3, -16, 2, 5, -20, 48, -42, 5, 25, 3, 4, 15, 17, 1, -9, -2, -21, 1, -46, 4, -29, -6, -1, 37, 34, -33, 34, 12, 9, -25, 12, 1, 16, -18, 0, -51, -24, -30, 25, -8, 13, 24, 1, -2, -34, -1, -20, 21, 9, 8, 3, 31, 3, 31, -29, 7, 4, -9, 15, -12, -3, -20, -2, 1, 26, -1, -5, 33, -7, 5, -9, 7, 5, -15, -6, -17, -9, -4, 39, -50, -2, 6, 7, -4, 26, -1, 5, -1, -5, 19, 4, 18, 18, 30, 3, -13, -4, -9, -89, 24, -2, 12, 24, -16, -41, -8, -19, 0, 31, -9, -13, 31, 0, -4, 3, -11, 0, -27, -2, -5, 1, 7, -22, 1, -40, -3, 7, 14, -10, 21, -2, -33, -10, 63, 7, 0, 30, 0, -33, -1, -40, -13, 1, 5, 39, -6, -26, 33, -28, -6, 1, -8, -3, -71, 11, 1, -15, -14, 23, -2, 15, 63, -5, -16, -36, -5, -25, -6, 38, 8, 0, 11, -1, -44, -11, 0, 2, 10, 5, 0, -3, 0, -5, 5, 5, 4, 7, -12, -5, 16, -2, -8, 10, -4, -4, 22, -8, 11, 21, 10, -6, -7, -6, 17, -29, -28, 14, -11, -6, 8, -18, -7, 4, -19, -4, -6, -16, -34, 3, -29, 3, 21, 16, 4, 6, 2, -12, -4, 9, -3, -3, 12, 23, -41, -23, -9, 32, -11, 1, -22, 3, -5, 3, -25, 29, -32, -2, -32, 6, 14, 23, 30, -41, 6, 12, 28, -14, 15, -3, 0, -5, 13, 7, 0, 26, -3, -5, 4, 8, -16, 7, -7, -49, -3, -13, 5, -3, -2, -2, -18, 0, -23, 5, 3, -23, -3, -19, -18, -15, 40, -2, -26, -29, 49, 8, -16, 5, 23, 2, -15, -39, -14, 22, 27, -11, 2, 8, 15, -8, 9, 28, 3, 0, -6, 8, -5, -17, -13, -4, 2, 42, 0, 1, -14, 7, -15, 0, 21, -4, 38, 1, 17, -4, -12, 16, -15, -1, 0, -17, 0, -11, -1, -4, 4, -45, -1, 1, 0, -45, 13, 27, 8, 0, 17, 25, 3, -11, -1, 4, 23, -11, -34, -8, 42, -19, -6, 31, -41, -4, 0, 37, 0, 9, 17, -5, -73, -9, 13, -3, 45, -40, 11, 21, 15, 6, 57, 4, -13, 2, 16, 7, 0, 31, -3, -23, 15, 24, -12, 24, 6, -21, 0, -14, 4, 11, -4, -5, -6, -20, -27, -11, -2, -15, 9, -19, -3, 28, 17, 3, -104, 9, -7, 22, -1, -1, -25, 6, -22, 5, 27, -9, 9, -18, 12, 26, -5, 1, 12, 24, 14, -1, -5, -24, 10, -24, -21, -8, -8, 43, -8, 7, -26, 5, -38, 16, 35, -1, -12, 20, 9, 44, 36, -29, 31, 63, -7, 28, -46, -22, 8, -9, 3, -46, 37, -94, -24, -21, -70, -2, -29, 1, -11, -67, -8, 13, 1, -8, 4, 4, -8, -29, 11, -1, 26, 20, 17, 7, 24, -27, 40, -43, -40, 0, -37, 40, -1, 0, 0, 5, 30, 23, -3, -3, 15, 6, 33, 29, -41, -27, -2, 27, -4, -14, 2, 21, 17, -4, 3, 23, -4, -32, -27, 8, 3, -4, 0, -47, -8, -30, 30, -41, 12, 12, 2, 0, -30, -5, -5, 22, -14, -13, -8, 6, -4, -5, 14, 0, 7, -31, 19, 5, 14, -13, 42, -3, 16, 1, 0, -2, -1, 9, 27, -16, -41, -4, 0, 25, -23, -4, 18, -5, -29, 41, 35, -5, -6, 14, -9, 28, 11, 14, 4, 2, -13, 3, -50, -7, 5, 6, -7, -29, 15, -76, -18, 0, -49, -21, -24, 4, 29, -30, 0, 12, 0, -49, 9, 15, -30, -23, 25, -38, 14, -4, -38, 0, 23, -23, 1, -79, -86, -2, -58, 8, 15, 15, 22, -2, 28, 35, 3, 3, 0, 1, 21, 0, -5, -2, -2, 25, -3, -21, 0, 11, 0, 0, 6, 51, 3, -35, -9, 3, -2, 5, 0, -18, -51, -7, 34, -54, 5, 0, 1, -1, 15, 0, -9, -7, 8, 39, -5, 21, 23, -2, -5, -4, -2, -9, 22, -14, 8, -15, 41, 5, -11, -3, 1, 2, 2, -27, 22, -18, -13, -7, 1, 27, -5, -4, -6, 11, -41, 37, 43, -1, 0, -14, 9, 11, -18, 15, -38, -2, -4, 8, -51, -6, 13, 3, 1, -30, 26, 21, 22, -19, -24, -14, -35, -2, 5, -1, -17, 4, -10, -37, 16, 30, -49, 15, 19, -1, 11, -1, -38, -3, 19, -55, 51, 19, -14, 0, -67, 26, -16, -20, 27, -26, 15, 33, -12, 3, -12, 1, -4, -10, 0, -12, 5, 41, -9, -14, 4, -16, 18, 6, 0, 37, -6, -30, -33, 11, -2, -1, -25, -29, -21, 14, 23, -55, 7, 9, 6, 9, 31, 7, -32, -37, -16, -7, -14, 9, 3, -4, 3, -4, -30, -34, 0, -1, 0, -9, 17, -3, -6, -10, 1, 5, 7, -19, -31, -10, -75, 4, 0, 38, 2, 5, 0, -1, -72, 0, 26, 4, -2, 2, 14, -35, 4, -20, -51, 3, 3, 9, -28, 8, 40, 4, 0, -35, 8, -37, 1, -27, -46, -36, -15, 5, 8, -32, 2, 8, 5, -19, -13, 13, -26, 0, 14, 0, -30, 6, 16, 7, 21, -70, -2, -12, 1, -2, -78, -10, -17, 18, 6, -40, 16, 5, 4, 5, -57, 4, -30, -19, 62, -13, 3, 44, -3, -34, 6, 27, -9, 3, -9, -11, 2, -42, -31, -6, -1, 8, -10, 9, -35, 31, 32, -36, 15, -12, -5, -28, 0, -2, -46, -4, -37, 14, 2, 35, 21, -8, 0, -72, -32, -16, -11, 14, -5, -43, 3, -5, 15, 2, 12, 3, 1, -54, 10, -7, 0, 5, -6, 31, -5, -7, 11, -3, -36, 19, 28, 1, 0, -9, 22, -7, -25, 10, -23, 7, -14, 8, -20, -2, 34, -10, 1, -37, 16, -51, -10, -19, 1, -33, -30, 3, 12, -54, -12, 6, 0, 4, 18, -24, -48, -17, 5, -24, -3, 9, -2, 4, 10, -6, -1, -10, -40, -1, -64, -33, 13, -12, -29, -48, 9, 2, -13, -2, -27, 0, -6, -18, 38, -10, -7, 44, -10, -14, 3, 6, 11, 8, -1, -22, -3, -44, 7, 11, -7, -4, -6, -8, 6, 14, -14, -59, 10, 7, -23, -23, -8, -3, -47, -6, 47, 36, 5, 38, -16, 0, 1, -8, 12, -10, -2, -8, 12, -11, 28, -6, -22, 16, 3, -1, -1, 10, -12, -15, -41, -3, -2, 21, -18, 6, -1, 7, -58, 19, 8, 6, 21, -12, 45, -11, -18, -8, -14, -27, -23, 13, 8, -7, 21, -7, 0, -28, 40, -63, 19, -32, -8, -21, -17, -5, 16, 9, -15, 0, -5, -18, 22, 17, -52, -21, 5, -3, 14, 7, -34, 9, -16, -26, -10, -9, -62, -3, -21, -15, -10, 9, 20, -27, 31, 16, 23, 6, -5, 5, 2, -34, 25, -1, -7, 12, 1, -2, -6, 10, -6, -2, -5, -34, -3, -67, 2, 21, 6, 0, -19, 2, -39, -31, 48, -30, 22, -24, 0, -11, 32, -6, -24, 2, 30, -7, 11, 8, -20, -6, -9, -14, -15, 9, 19, -12, 5, -34, 59, 0, 25, 25, 12, 9, 4, -32, -29, 15, -63, 0, 6, 18, -13, 1, 7, 7, -63, -19, -8, 5, 24, 17, 21, -10, -7, 23, -6, -36, -11, -22, -31, -11, 2, -3, -1, -49, 0, 21, -40, -22, -36, 20, -7, 0, 12, -27, 10, -1, 3, -42, -6, 6, -17, -25, 32, 28, 19, 24, -21, -2, 15, -31, -29, -15, 5, -9, -24, 1, 22, 15, 1, -22, 30, -4, 26, -1, 0, 0, 0, 17, 1, -46, -2, 2, -5, -22, 2, 22, 23, 3, -6, 34, 2, -23, 0, 32, -4, -3, -46, -35, -23, -32, 15, -57, 28, 13, 2, -1, 9, 0, -58, 9, 18, -21, -10, 27,
    -- layer=2 filter=0 channel=5
    -12, 3, -27, 18, -83, -15, -61, 24, -13, 9, -77, -3, -1, -24, -1, -5, -1, 22, 32, -18, -12, -8, 1, -22, -1, 1, 13, -1, 47, -26, 2, -7, 0, -4, 0, 11, 1, 16, 12, 30, -3, -47, 21, -27, -19, -8, -9, 8, -21, 0, -24, 36, 42, 47, -12, 0, -66, -3, 36, -3, 8, 27, -7, -4, -26, -29, 30, -34, 14, 2, 23, 3, -26, -13, -3, 13, -47, -5, 13, -45, -1, -14, 17, 26, 8, -21, -8, 17, 42, 6, -33, -12, 0, -6, -5, 10, -1, 23, -6, -34, 0, 0, 1, 30, 3, -41, -21, -10, -4, 4, 3, 18, -36, 22, -22, -19, 17, -9, -3, -69, -43, 1, 4, -18, -15, -4, 0, 11, -15, -2, -3, 38, -13, -12, -2, 26, -10, 33, -7, 2, -7, 11, -1, -6, -5, -4, 19, 0, -30, -6, 0, -30, -17, 3, 0, -10, 60, -11, -11, 1, 12, -13, 3, 1, 6, 21, 9, 16, 0, -15, -20, -19, -52, 3, -4, 5, -32, 20, -46, -36, 44, -30, -12, 3, -31, 13, 9, -44, 7, 29, -2, -2, 21, -9, -4, 7, 37, 8, 24, -7, -18, -43, -26, -16, -14, -7, 51, -12, -10, -13, -8, 6, -14, -42, 26, 11, 15, -6, -27, -31, -41, 2, -1, -23, 0, 9, -11, -14, -30, -1, 3, -29, 4, -14, -20, 10, 3, 0, -22, 2, -27, -3, -3, -3, 16, 2, 13, -45, 17, 3, 38, 2, 11, 15, -14, 0, -10, 0, -13, -11, 17, -21, 19, -19, -19, 12, 12, 5, 5, 11, 4, -5, -4, -29, -50, 31, -64, -7, 0, -22, 3, -1, 0, -3, 36, 7, -9, -1, 12, 7, -7, -2, -15, 17, 16, 16, 10, -5, 0, -31, -13, 2, -8, 21, -11, -8, -27, 33, 34, -19, -1, -2, 14, 5, 22, -41, -1, 0, 5, -16, 0, 8, 11, 8, 22, 0, 41, -1, 28, -51, -21, 17, -5, -1, 7, -1, 19, -2, 15, -20, -9, -23, -8, 0, -41, 5, 8, 3, -14, 2, -4, -17, 1, 19, -10, 7, 12, 0, 3, 73, 5, 0, 28, 4, -7, -1, 38, -15, 0, 2, -8, -12, -16, -4, 1, 26, 16, -8, 19, 14, 33, 29, 20, 55, -18, 0, 17, -25, 11, -25, -34, 33, -9, -3, -14, 5, -25, 9, 2, -1, 3, -7, 18, 10, -56, 0, -7, -11, -6, 0, -22, 1, 34, 13, -10, -6, 42, 2, -4, 3, 15, -26, 36, 52, 27, 0, 18, -31, -21, 0, -1, 2, -13, -42, 5, 32, 27, -61, 17, -2, 9, 6, 6, -9, -5, 11, -7, 3, -15, 16, -10, 3, 5, 50, -1, 5, 6, 8, 2, -5, -13, -3, 0, -3, -3, 14, 13, 2, 11, 9, -17, 7, -32, -1, -23, 0, 8, -6, -7, -41, 4, -4, 16, 7, -13, -9, -6, -2, 6, -6, 7, -24, 0, -1, 3, 12, -7, -3, -4, 13, 3, -6, -9, 41, 0, -5, 0, 7, 15, 8, 0, -4, -31, -9, -40, -8, 43, 4, 3, 5, -24, -24, -16, 2, -3, -9, 10, 3, 6, -7, -8, 0, 3, -8, 4, 8, -15, 7, -15, -3, 26, 14, -2, 6, 16, -9, 6, 20, 11, -17, 0, -7, -29, 24, -5, -54, 9, 0, 0, -24, -3, 2, 7, 19, 5, -3, -7, 3, 23, 13, 7, 7, -8, -21, 2, 5, 0, 24, 26, -16, 2, 34, 3, -5, -6, 10, -1, 14, -18, 2, -26, -15, -16, -25, -19, -31, -3, 33, 16, 2, -8, 2, -19, -9, -18, -39, -6, -14, -3, 22, 1, -13, -23, 0, -5, 5, -2, -13, 21, -13, -6, -3, -21, 12, 3, 21, -21, 16, 5, -1, 1, 30, -10, 6, -57, -2, 15, 15, 20, 5, -9, 5, 10, -56, -4, 40, 5, 24, -9, -27, 2, 5, -10, 4, 9, -2, 5, 31, 12, 42, 8, 0, -9, 13, 2, 2, 21, -6, -4, 26, -2, -6, -4, -23, 41, 24, 6, 47, 22, -76, 14, -16, 12, -35, 22, 7, 6, 24, 10, 0, 17, 39, 0, 39, -8, 4, 22, 5, 32, -1, 0, -5, -8, -28, 5, 13, 2, -17, 22, 30, 14, -2, -18, 29, -17, 11, 0, -4, 39, 19, -12, -18, -31, -5, -6, 21, 7, 0, -9, 0, -5, -26, -1, -25, -4, -3, -8, -7, -6, -19, -8, 22, -2, -23, 0, -17, 25, -20, 3, -7, -38, 1, -45, -35, 2, -6, -10, 0, -5, -1, -20, -3, -60, 33, -15, 14, 2, 0, 3, 5, 10, -36, -39, 19, -43, 29, -22, -25, -6, 2, -1, 8, 5, 6, 6, 0, 14, -19, 2, -10, -6, 18, -17, -3, 4, 1, -5, 2, 17, 4, 9, -23, 59, 33, -26, 36, 35, -24, 7, -22, -34, -5, -3, 7, -2, 13, 21, 5, 1, 26, -24, 3, -12, 1, -19, -21, 27, 6, 3, 9, -30, -14, -31, -8, 4, -25, 51, 30, 17, -2, 24, 23, -7, -2, -19, 1, 9, -4, -17, -26, -42, 21, -7, 9, 4, 15, 28, -4, -43, -18, 27, 8, 2, 10, 5, 38, 0, -10, -14, -2, -6, -23, -7, -30, 6, 20, 0, 4, 1, 17, -35, -33, 0, -21, -4, -25, 18, -13, -20, 4, 4, -10, 0, 7, 2, 0, 1, -9, 4, 9, -3, -14, 22, 20, -9, -18, -29, -5, 13, -23, 1, -4, 4, 1, -35, -26, -14, 2, -7, 16, 9, -2, 20, 1, 12, -40, -32, -5, -17, -1, -10, 28, 29, -8, 14, -32, 10, -6, -20, -15, -33, 3, -4, -17, 33, -40, -28, 14, 24, -25, -24, -1, 13, 11, 0, -23, 3, 1, -7, -7, 27, -24, 0, -15, 9, -13, 11, 0, -55, -37, -21, -7, -42, 4, 33, -17, 12, -14, 2, 7, -21, 5, 29, 14, 4, -7, -20, 3, -15, 13, -3, -9, -1, 34, -4, -44, -33, -28, 0, -9, -7, -13, -3, 22, -5, -1, 3, -13, -23, -3, 25, 12, 0, 0, -20, -4, 3, 4, 8, -49, -13, -23, 0, 2, -22, 0, 23, 3, 18, 10, 4, 25, -10, 1, -31, -5, -5, -16, 10, 0, 1, -18, -34, 1, -74, 4, -2, -7, 4, -7, -6, 0, 21, 11, -25, 5, -24, 14, -19, 14, 23, -8, 15, 18, -28, 18, -18, 2, -35, -4, -4, 3, 11, -8, -30, 41, 11, -32, -22, 3, -2, -58, 23, -13, 0, 6, -11, 5, 17, -26, -4, 0, -19, -38, 14, -4, -3, -70, -20, 16, -16, 0, 25, -28, 18, -10, 21, 8, 0, 16, 7, 23, -18, 7, -15, 14, -43, 2, -1, -17, 3, -8, -15, -32, -15, 3, -7, 28, 0, -3, -19, -12, -7, 4, -10, -1, -7, -23, 14, -16, -22, -2, -24, 25, -1, -2, 20, -6, 37, 15, 4, 39, -4, 0, 20, -5, 69, 23, -31, 35, -7, -20, -36, 4, 28, 20, 7, 4, 4, -3, -30, 16, -57, -10, 2, -14, -6, -4, -4, -5, 25, -3, -28, 0, 16, 21, 43, -6, 44, -61, -25, 37, -1, 15, 17, 27, -22, 4, -4, 26, -2, -66, 19, 5, 44, -8, 3, -6, 12, -56, 26, -15, -7, 5, 3, 13, 45, -33, 13, 3, 3, -9, 43, 6, 26, -43, -13, 36, -37, 4, 7, -16, 14, 61, 5, -49, 17, -6, 31, 11, -76, 7, 5, -23, -29, -9, 0, -7, -5, 24, -12, 8, 5, 4, 5, 12, 0, -25, -13, -6, 0, 4, -4, 3, 2, -13, -5, 5, -15, 13, 12, 40, -2, 5, -4, 10, -18, -5, 23, 31, -15, 0, 38, 23, 0, 9, -8, 53, -3, 31, -37, 0, 57, 27, 8, 7, 6, -28, -5, -14, 8, -3, 6, 9, -13, 4, 14, 0, 9, 0, -28, 7, 25, 33, 0, 3, 33, -23, 22, 47, 34, 34, 20, 30, -18, 4, 7, 26, -2, -30, 15, 25, 54, -14, 19, 5, 24, -7, -14, -4, -1, 17, 4, -8, 11, -5, 5, 2, 26, 17, 15, -8, -12, 3, 12, 33, -24, -7, -24, 15, 3, 42, -5, -4, 24, -3, 19, 11, -93, 0, -7, -2, -51, -5, -5, -5, 2, 16, 6, 32, 40, 8, 3, -11, 1, -42, -14, -13, -5, 5, 19, 25, -6, 10, -32, 9, -14, 30, -4, 22, 55, -8, -10, -20, 26, 24, 10, 25, 2, 6, 5, -44, -16, 10, 13, 19, 5, -7, -42, 6, 18, 15, 5, -5, -5, -12, -31, 6, 21, -3, 3, -10, -8, -8, -17, 5, 9, -6, -28, 4, 41, 14, 27, -4, 29, -6, 2, 46, 39, 29, 3, 1, 14, 1, 0, 18, -15, -15, 29, 28, 18, 12, -8, 2, 44, -30, 8, -6, -6, 16, -10, -11, 8, -1, -10, -4, 4, 11, 18, -7, 6, 17, 9, -5, -21, 6, -15, 10, 17, 13, 7, -7, 13, 11, 12, 5, -65, 0, 21, -24, -12, -12, 4, -10, 1, -2, 3, 34, 22, 22, -6, 5, 2, -3, 6, -5, -1, -7, -13, 2, -4, -52, -44, 34, 14, -5, 4, 19, 38, -5, -17, 4, 22, -9, 9, 13, -8, -2, -9, -22, 0, 25, -20, 18, 2, 0, -16, -2, -21, -10, 11, 0, -5, -5, 8, 29, 15, -5, 1, 29, -5, -8, -15, -1, -31, 24, -7, -5, 16, -19, 16, 15, -36, 5, 14, 0, 49, 12, 14, 15, 30, -2, -3, -1, -19, 10, 21, 27, 19, -32, -65, -4, 1, -19, 3, -9, -14, 3, 4, -48, -6, -39, 0, -5, 1, 1, 3, 2, -10, 34, 6, -6, -8, -6, 49, 0, -9, -34, -17, -8, -4, 31, 45, -9, -22, -6, -39, -5, -2, -25, -2, -20, 0, 9, 0, 0, -9, 17, -2, 5, -4, -11, 0, 5, -6, -4, -16, -8, -3, -51, -38, 33, -8, -8, -4, 29, 31, -5, -13, -5, -13, 28, 22, -3, 0, -1, -1, -30, -28, 9, -16, 23, -21, -33, -30, -5, 6, 1, 9, 5, 5, 12, 15, -17, 1, -5, 7, -7, -5, -2, 6, -8, -31, 14, 9, 7, -35, -21, -26, 17, -8, 22, 6, -16, 23, -3, 14, 14, 5, -4, 3, 9, 14, -37, -8, 19, 1, -3, -18, -7, -33, -7, 2, -18, -7, 9, -11, -6, -23, -17, -26, -22, -5, -10, 16, 0, -7, 37, -2, -5, 1, 0, -9, -25, -14, -3, -5, 29, -13, 35, 26, 12, 21, -2, -6, 20, 20, -2, -1, 14, 0, 5, 5, -32, 13, -10, 0, -27, 4, -29, 6, 3, -4, 5, -26, -8, -35, 12, 2, -9, -26, -13, -23, -7, 1, 6, 13, -5, -31, 66, 5, 8, 6, 0, 3, -38, -31, -9, 1, 47, 12, -23, -8, -1, 2, -18, 1, -8, -6, -40, -6, -25, 6, -8, 4, -5, 2, 0, -3, 1, 23, 0, 2, -1, 0, -18, -23, 29, 4, 2, 34, 8, -19, -3, 13, -14, 0, -7, -8, -7, 18, -38, -56, 5, 18, -28, -4, -8, -1, -70, -8, 8, 0, 0, -8, 0, -13, -13, 22, -6, 34, 0, 29, -1, -26, -31, 44, 34, -19, -2, 54, -13, 10, -28, -5, 54, -13, -4, 25, 6, 57, -5, -5, 53, 17, 32, -1, -60, 7, 5, -2, -4, -14, -34, -4, 21, 7, -1, -11, 19, -3, 4, 11, -4, 20, 2, -11, -20, 22, -7, -5, -34, 15, 0, -44, 26, -13, 14, 7, -8, -16, -8, -5, -43, -2, -34, -12, 5, -2, 32, 40, -6, 0, -9, 0, 6, 5, -9, -13, -8, -17, -5, 9, 6, -7, -4, -6, -7, 28, 9, -20, -2, 1, 4, 7, -24, 8, -2, -18, 4, -15, 4, 21, 29, -12, 3, -7, -30, -28, -7, -16, 39, 16, 0, -23, 4, -23, -15, 6, -21, 2, -22, -28, -5, 15, -21, -17, -28, 5, -39, 23, 1, -6, -54, 15, 18, -56, 0, -17, -24, 2, 8, -5, 14, -11, -8, 3, 7, 4, -1, -8, -22, -8, 36, 3, 6, 9, -1, -5, -6, -15, -4, 1, 45, 4, -30, -16, -34, 0, 0, -12, 15, -9, 10, 10, -2, 11, 35, -18, -11, -46, -6, -1, -9, -4, 9, -6, 25, 9, -6, 15, -24, -1, 4, 29, 38, -19, 25, -56, -4, 13, 8, 3, -5, -2, -23, -18, -6, -10, -2, 2, 47, -4, 5, -3, 3, 10, 10, -3, -3, -6, 0, 13, -14, 10, -35, -20, 10, 2, 40, -5, 43, -24, -6, 1, 36, -14, -41, -4, 2, 11, 26, -50, 0, -15, -1, 8, -16, -1, -1, -5, -12, 11, -37, -10, 13, 0, -30, 8, 6, -1, 16, -6, 8, -38, 2, -26, -17, 3, 26, -1, -78, -3, -21, -8, 3, 12, 0, -29, 7, -29, 10, -5, 33, -1, -48, -7, -26, -39, 10, -2, 4, 4, -31, -34, -29, 4, -5, -22, -28, 15, -31, -8, -3, -29, 42, 0, 2, -35, 0, 20, -18, 18, -6, -4, 29, -33, -4, 13, 30, 13, 13, 26, 2, 6, 21, -44, -3, 3, -23, 6, 0, 6, -21, -15, 13, 27, -5, 7, 14, -17, 0, 7, -1, -7, -1, 9, 4, 19, 22, -10, 6, 20, -88, -30, 38, 16, -15, -11, 26, -3, -3, -1, 0, 3, -23, 24, 7, -13, -36, -41, -4, 7, 44, -43, -12, -3, -14, -11, -43, 8, 10, -29, 26, 0, -30, 15, -6, -22, 13, -60, -19, -21, 2, -45, -25, 7, 10, 17, -49, 21, -4, 33, -6, -15, -2, 14, -2, -41, -39, -1, 28, 9, -25, -5, -1, -18, 16, -1, 12, -1, -21, -11, -44, 2, -5, 4, 24, -1, -16, -52, 4, -26, 40, -8, 17, -44, 0, 19, -1, -44, 4, -4, 5, -7, 1, 3, 11, 33, 35, -7, 11, -7, -26, -14, 4, -8, -1, 16, 3, 6, 18, -74, -18, 23, -7, 0, 1, -15, -4, 0, 3, -18, 23, -23, 1, 21, 12, -38, -37, 14, -36, -14, 39, 87, 35, 11, 52, -10, -3, 0, 14, -33, 15, -3, -6, -10, 63, -42, 2, 36, -24, -10, 14, 0, -21, 21, -51, -8, -6, -17, 18, 6, -42, -24, -1, 31, 34, -29, 12, -18, -5, -66, -13, -7, 24, 19, -31, 5, -10, 17, 10, -46, -2, 29, -28, -22, -16, -7, -4, 3, -38, -5, -21, 28, -2, -4, 3, 0, -32, -20, -33, -3, 5, 10, -18, -6, -11, -43, -22, -20, 25, -3, 3, -16, -5, -33, -15, 22, 42, 10, 1, -6, 0, 3, -1, -39, 21, 40, 17, -6, -25, 18, -2, 2, 6, 0, 0, 3, -42, 6, 29, 28, 0, 6, 18, -9, 1, -2, 10, -43, 13, 2, 0, -12, 16, 3, -23, -13, 11, -15, 0, 34, 20, 20, 35, 16, -2, 5, 14, -10, -7, 2, 3, 30, -24, -32, 4, 21, -17, 7, 5, 1, 1, -40, -45, -25, -1, -10, -36, 1, -3, -5, 5, 8, 30, -2, 3, -37, -1, -47, 10, 15, -2, 6, 1, -1, -20, 19, -3, 4, 4, 15, 4, -3, -12, 3, 21, 0, -15, -8, 0, 6, 19, -5, -28, -3, 11, 4, -20, -6, 0, -23, -42, -16, -10, 7, 10, -1, 15, 0, 5, -31, -3, -55, -21, -7, 36, 21, -7, 7, -6, -12, -32, 16, -18, -16, 28, -3, -9, -16, -3, -5, 22, 5, -2, -6, -15, 18, 17, -55, -8, -2, -12, 8, 0, 21, -2, 19, -1, 34, -2, 9, -8, 7, 5, -23, 64, -11, -3, -23, -8, 19, 16, 7, -15, 0, -4, 17, -10, -29, 36, 13, -27, -14, -5, -49, 19, 12, 10, -17, -20, 3, 13, -29, -7, 5, 22, 17, 2, 28, 8, 29, -5, -11, 6, -53, -8, -24, -14, 3, -17, -4, 29, 4, -22, 4, -7, 42, 5, 3, 6, 38, -17, 2, 0, -10, 14, 5, 3, 13, -40, 0, -48, -1, -6, 13, -3, 6, 0, 9, 3, -26, 13, 4, 15, 7, 11, -11, 34, 5, -8, 18, 4, 7, 61, 27, 17, 13, -1, -21, -18, 10, 0, -22, 25, 5, -14, -3, -4, -8, 7, 2, 2, 0, 1, 18, 4, 15, -2, -5, 0, -12, -9, 3, 9, -18, -8, 8, -3, -33, -34, 3, -17, 1, 24, 26, -11, -15, 21, 8, -11, -10, 0, 2, -6, 37, -31, -29, -13, 3, 69, -13, -5, 11, 22, 1, 5, 1, 4, 3, 1, -7, 11, 24, -4, 31, -11, -1, -1, -40, 22, 8, -71, -35, -4, 9, -38, -7, -13, 4, 28, -12, 10, 25, 15, 3, 4, 11, 15, 30, -1, -6, 0, 2, -9, -3, -3, 8, -14, 6, 5, 5, -22, 1, 14, -5, 5, 10, -3, -25, 11, -9, -5, 11, 0, -3, -21, 2, -3, -28, -19, -26, 0, 0, -3, -16, 0, 17, -23, 44, 5, -6, 42, -9, 1, 52, 4, -6, -16, 5, -4, -3, -1, -19, -8, 13, 6, -1, 3, -15, 4, 6, 3, -7, -14, -13, -7, -27, -1, -11, -36, -7, -7, -46, 0, 23, 44, 18, 9, 1, -13, -1, -35, -17, -33, 10, -2, 4, 23, 6, 5, 45, -33, -16, 5, 2, -13, -18, 5, -19, 12, -25, 36, -13, -7, -4, -2, -32, -6, -54, 29, -54, -2, 30, -10, 31, 13, 26, 1, -22, -33, 18, 15, -18, -2, -46, -24, -2, 20, -6, -7, 0, -39, -1, -8, -14, -18, -3, 20, -6, 0, 14, -34, 4, -9, -4, -4, -5, 19, -20, 17, -10, -22, -10, 17, -20, -5, 32, 22, -36, -12, -4, 10, -10, 0, 21, -16, -39, -25, -12, -16, -2, 7, 1, -2, 15, 4, 4, 3, -3, -45, -2, -13, 0, 3, -6, 14, -11, -5, 15, 5, 1, 9, 23, 2, 19, 9, -3, -55, 22, -41, -48, 14, -4, 28, 26, 20, 15, -10, -4, 9, 4, -59, 2, 6, -17, 18, -10, -7, 14, -23, 13, 3, -8, 4, -59, 5, 4, 7, -1, 14, -18, 1, 10, -6, 12, -12, -14, -5, -50, 5, -59, -42, 29, 3, 8, -21, 8, -68, 20, -5, -9, -5, 13, -20, -15, 18, 7, 17, 1, 16, 2, -47, 0, -2, 2, -28, -3, -36, 1, -28, 3, -2, 19, 10, -41, -4, -8, 28, -17, 21, 13, -16, -41, 3, 31, -42, -3, -36, -3, 16, -8, -5, 23, -2, -28, 17, 21, -34, 0, 45, -49, -2, -6, -40, 3, 6, -5, 16, -9, -15, 47, -1, 7, 33, 0, -5, -2, 3, 11, -25, 4, 0, 14, 4, 20, -8, 34, -34, -60, 5, 84, 12, 29, 16, 2, -2, -2, -6, -22, -13, 8, 28, 19, 30, -73, 0, 23, 24, 2, 0, 10, -24, -57, 6, -3, 16, -1, 12, -4, -27, 3, -5, -8, -3, -45, -20, 13, 0, -35, -48, -21, -45, 7, -35, -16, -78, 3, -12, -21, -7, 0, -41, -1, 0, -1, -4, -2, -39, -1, -47, -22, 3, -6, -15, -1, -26, -17, -25, 3, -2, -3, 26, 6, -13, -25, 11, -59, 38, 17, 0, -68, -6, -2, 0, 7, -30, -35, 5, 1, -1, -21, 29, -31, 17, 46, 9, -1, 1, -11, 1, -9, -10, 9, 1, -7, -35, 1, 34, -6, -4, 2, 23, 0, -2, -4, -7, 10, -21, -27, 1, -6, -2, 34, -6, 12, -28, -25, 14, 33, 44, 23, 14, -24, 7, -5, -2, -24, -21, -16, 29, 20, -9, -20, 8, -36, -45, 8, 8, 12, 9, 5, -31, -24, 13, -25, 11, 15, -19, -4, 6, -2, 19, -22, 20, -25, -8, -28, -6, -13, 22, 17, -2, -5, -23, 31, 16, -12, 7, 5, -17, -9, -10, 6, -11, 5, 1, 15, -12, -38, 4, 0, -7, -4, -23, -32, -31, -5, 2, 0, -6, 9, -10, 22, -17, -47, -7, -13, 36, -66, -3, 21, 10, 8, 1, -11, -2, 0, -8, -6, 19, -16, 7, -21, 8, -18, 15, -81, 4, 5, -4, 9, 5, 3, -11, -7, -12, 12, 5, 5, 9, -23, 0, 4, -2, -6, 18, 6, -7, 13, 19, -3, -4, 0, -9, -44, 2, 20, 14, 10, 0, -9, 3, 0, -1, -59, -14, -39, 13, 7, 0, -17, 6, 48, -42, -21, 7, -10, -48, -23, 24, -29, 23, 1, 33, -7, -20, 18, 1, 38, 13, -14, -35, -69, 0, -24, -56, 12, 24, 23, -47, 15, -17, 38, 12, -7, 3, 24, -10, 2, -20, 2, 11, 6, -14, 10, 15, -9, -10, 0, 18, -4, -60, 20, -37, -6, 5, -15, 7, 5, -21, 40, 20, -30, 1, 0, 26, -16, 6, -51, -2, 41, 38, 16, 6, 15, -1, 1, -32, -11, -10, -24, 15, -7, -4, -8, -9, -17, 6, 0, -2, -3, -40, 5, 30, -4, 1, -8, 2, -11, -8, -18, 6, -9, 12, 21, -2, 3, -7, 20, 27, 19, 0, -7, -30, -8, -24, -8, 1, 36, -9, -3, -13, -26, 21, -52, 28, 2, 16, -41, 6, 29, -2, 14, 17, -2, 8, 3, -12, -12, -9, 17, 17, 13, 19, 0, -1, 11, 3, 1, -15, -18, -4, 22, -23, 25, 6, 0, 14, 15, 27, 6, 26, 36, 0, -11, 12, 44, -33, -7, 0, 0, 52, 2, -16, 6, -13, 6, 11, 6, -48, -18, 10, 5, 5, 27, 16, 17, -10, 24, -16, 10, -17, -13, 23, 0, -1, -3, 31, -9, -26, 1, -7, 28, 1, -7, -40, -12, -16, -38, 35, -13, -9, -11, 3, 1, 17, 9, -3, 0, 20, 47, -8, 21, -5, -1, -2, 2, -7, -6, 7, 6, 8, -1, -7, 16, -33, -14, 22, -7, 16, 12, -15, -7, 10, 14, -8, -3, 3, 0, -36, -8, -41, 24, -11, 46, 10, 21, -6, 0, -17, 2, 2, 3, -19, 20, 14, -12, -47, -3, 19, -13, 12, 8, 5, 15, -6, 2, -38, -6, -3, 45, 28, 4, 17, -6, 20, -10, -3, 30, 6, -9, 1, -4, -4, 14, 23, -7, -31, 2, 12, -3, 0, 3, -34, 2, -15, 5, -2, -22, 6, 5, -2, 3, 33, 12, 5, 23, 4, 22, -15, -23, -33, 12, 5, -35, -16, 15, -21, 15, 7, 21, -6, 6, 0, -23, -29, -36, 7, -4, -12, 27, -2, -2, -12, 10, 7, 1, -6, 28, 18, -9, 3, -2, 6, 13, -2, 3, -7, 17, -18, 28, 7, -7, -2, 10, -10, 7, -2, -21, -3, -2, 27, 11, 7, 14, -13, 0, 2, -30, -17, -19, 23, 14, 28, 0, 2, -18, -45, 23, 21, -4, -47, -16, 16, 0, 26, -6, 17, 6, 14, -7, -1, 2, -2, -40, -5, -55, 2, 25, 10, -4, 7, -25, -12, 3, -27, -15, 4, -13, -1, 23, -61, 39, 24, 7, 0, -5, 2, 6, -31, -10, -24, 7, 12, -7, -47, -6, -15, 2, 0, -15, 18, 0, 26, 4, 20, -10, -7, -13, 3, -8, -2, -35, 20, -34, -13, 1, -7, 26, 0, 9, -7, -46, -3, 18, 4, -1, 24, 65, -5, -3, 2, -2, 0, 7, 7, 19, -37, 18, -1, -4, 26, 11, 1, 25, 4, -27, 11, 7, 0, -7, 0, 19, 0, -5, -24, -17, -8, 6, 45, -5, 7, 6, 4, 0, -19, -46, -25, -21, 16, -11, -41, 1, -7, 37, -3, -2, 40, -10, -18, -1, 55, -24, -36, 3, 19, -10, 13, -13, 2, 3, -4, -35, 35, -10, 5, 11, 2, -15, 18, 39, -35, 0, -23, -14, 0, -10, 0, -30, -20, 18, 8, -5, 33, 1, 34, 0, -8, 23, -20, 4, 10, 3, -57, -3, -40, 1, 6, -19, 11, 28, -1, 22, 18, -53, 23, 21, 28, -9, -4, -18, -12, 24, 2, -2, -4, 10, -2, 3, -3, -1, 0, 25, 22, -7, 24, 18, 0, -18, -6, 7, -3, -6, 15, -14, -29, 56, 0, -9, 32, 14, 3, 0, 0, -21, -14, 0, -2, -8, -9, 32, 0, 15, -41, -31, -3, 38, 56, -2, -17, 18, 2, -5, -5, -35, -2, 0, 1, 5, -23, 25, -4, 33, 13, 7, 19, -9, -25, -15, 2, -20, 31, 13, 8, -4, -25, -19, 0, 14, 16, -19, -10, 5, -7, -50, -46, -1, 29, -2, -6, -9, -54, -15, -12, 63, -4, 10, -21, -14, 20, -1, -1, -2, 1, 2, -12, -24, -7, 1, -16, 2, -30, 30, -40, -3, 7, -10, 43, 23, -32, -57, 36, -74, 2, 14, -8, -10, -4, -6, 0, 17, 4, -28, -17, -13, -2, -14, -10, -8, -19, 10, -6, -5, 22, -17, -9, -8, -52, -6, -5, 10, 6, -43, -11, 17, 5, 4, 8, -3, 5, -3, -1, -1, -1, -7, 0, 5, 7, 11, -50, 0, 2, -27, 36, 14, 53, 19, -12, 5, -6, 3, -29, -19, 22, -13, 1, 28, 49, -28, 0, 11, -28, 1, 30, -5, 13, -19, 34, -20, 22, -17, 5, -43, -21, -13, -5, 33, 1, -37, 4, 9, -10, 3, -48, 19, -6, 24, -37, 20, -54, 9, -10, 2, -2, 24, -26, -13, 0, -6, -6, 0, -28, 4, -25, -27, -30, -6, -23, 3, -81, 15, -19, -1, -6, 23, 2, 4, -12, -22, 13, -16, 16, 11, -7, -19, 5, -20, -23, -20, 28, -18, 0, -1, 5, 17, 6, 1, -27, -31, 36, 2, 33, -13, 2, 3, 0, 11, 5, -6, 4, 3, 0, -28, 6, -4, 23, -2, -6, 9, 0, -36, -7, 6, 1, 8, 13, 25, 8, 0, 4, -29, -14, 1, 2, 32, 3, 73, 7, 5, -15, 6, -16, -18, 36, 23, -11, -8, -4, 4, -51, 12, 20, -11, -6, -6, 17, -30, 42, 10, 13, 8, 12, -20, -1, 24, -4, -16, -22, -19, 6, -10, -17, -8, 38, -22, -59, 2, -30, 22, -7, 4, 7, -4, -3, 58, 12, 3, -25, -4, -18, 6, 45, -3, -16, 1, 0, 0, -33, 8, -9, 8, 2, -1, -7, 8, -10, 28, 13, -12, -1, 10, 0, -11, -8, 21, -39, -7, 26, 9, -14, 35, 4, 11, -25, 15, -28, -42, 30, -16, -49, 41, -2, -13, 5, 9, -7, -6, 15, 54, -3, -46, -2, 4, -6, -18, 2, -13, -3, 5, 15, -31, 0, -21, -6, 16, 43, -3, -4, -5, -16, 3, -33, 3, -21, 24, -7, 0, 1, 35, 42, -4, 29, 26, 16, 6, 4, -7, -38, 21, -5, -1, -38, 29, 10, -13, 6, -7, 3, 15, -3, -22, 3, -8, 42, -1, -4, -27, -4, -36, -5, -40, 18, 10, 4, 5, 20, 15, 0, 61, 4, -13, 22, 28, 2, -7, 5, 0, 16, 4, 31, 28, -27, 3, -29, 3, 10, 0, 5, -1, 6, -10, 34, 33, -8, 1, -27, 6, -16, 7, -19, -14, -4, -8, -11, 1, 22, 6, -11, 25, 6, -5, 26, 40, -28, -8, 12, -8, -19, 3, 8, -10, -19, -5, 6, -5, 28, -7, 18, -31, -2, 4, 4, 2, -8, -21, 0, 48, -19, -15, 4, -5, -18, -68, -7, 58, 0, 13, -7, -30, -15, 25, -13, -20, -10, -7, -27, -22, -19, -20, 0, 29, 50, -30, -9, -7, 11, 1, -23, -1, -18, -3, 2, -14, -10, -1, -5, 7, -6, -18, 6, 15, -10, -25, -31, 1, 3, 21, 13, -30, 30, -9, 7, 11, -23, 12, 0, 21, -7, 0, 22, -2, -25, -3, -28, -4, -6, -6, -6, 42, -11, -5, -1, -5, 19, -33, 15, 2, 3, -4, 0, -13, 23, 27, -17, 23, -44, -14, -33, 23, 2, 3, 4, 3, 0, -1, -36, -18, 7, -12, 39, 24, -38, -43, 1, -6, 7, 34, -2, 0, -7, 7, -3, 0, 16, 28, 0, 14, 0, 3, -16, -5, -4, -17, 1, 23, 22, 10, -5, -6, 8, -11, 0, 33, -10, -15, -31, 8, 3, 40, -47, -13, -3, -1, -15, -11, -31, -22, 7, 23, -27, -13, 6, 21, -38, 8, 16, 3, -27, 12, 16, -30, 6, 13, -4, -13, -30, -1, -3, 28, 21, -4, 2, -75, 4, 20, -20, -11, 27, -18, -10, 6, -6, -13, 11, -46, -7, -25, -51, -42, -3, -2, -10, -1, 32, -1, -11, 8, -10, -6, -20, 0, 1, 29, -13, 2, 5, 21, -4, 5, 0, -1, -16, -7, 9, 6, 19, 32, -9, -1, -18, -27, 22, -21, 24, 25, -7, 10, 22, 12, -13, 18, -33, 2, 33, 27, 5, -1, 8, 3, 1, 2, -4, 1, 4, 37, 3, 5, 3, -3, -3, 7, 3, -35, 3, -12, 5, -7, 15, -24, -23, -18, -59, -41, -30, -12, 0, 27, 3, 3, 0, 0, 1, -1, 37, 8, 30, 15, 15, -32, 0, 24, -65, -2, 5, -9, -17, 13, -5, -23, -12, 20, 13, -8, -18, -18, 8, 3, -24, -9, 11, -39, 3, -34, -14, 0, -1, 2, -64, -10, -50, 16, 2, -56, 2, 0, -33, 5, 34, 6, 9, 2, 0, -1, -1, -7, -1, 0, -45, 0, -14, 37, -25, -5, -6, -3, -8, 19, -4, -15, -38, -40, 0, 6, 13, -34, 1, -7, -30, 7, -25, 1, 12, -17, -1, -5, -32, 13, -29, -2, -1, -8, 0, 42, -5, 0, -6, 15, 1, 0, 46, 0, -4, 19, 1, -4, 0, -18, 0, 14, -3, -17, -31, -30, -6, 2, 19, 8, 0, -15, 0, -26, 9, 13, 13, 9, 2, 15, 10, -9, -15, -32, -2, 7, -10, -7, 27, 0, -3, 2, 0, -7, -15, 0, -5, -28, -4, -26, 30, 8, 4, -30, -26, -17, -1, 18, -5, -40, 25, -32, -7, -24, 6, -5, -24, 0, -32, 2, -13, -5, -8, 30, 5, 19, -5, -19, 18, 4, 7, -4, -48, -7, -24, -12, -18, -2, -89, 5, -17, 33, -24, 7, 6, 8, -23, 12, -26, -41, -18, -42, -7, 1, 12, -21, -1, -12, -1, 16, -22, 2, -4, -6, -5, 34, 15, 10, -41, -30, 6, -8, 9, 4, 7, 0, -18, 0, -6, -7, 7, -11, -7, 20, 0, -3, 12, -21, 3, -6, -1, -9, 10, -14, 7, -27, -11, 27, -19, 6, -27, -7, 35, -33, -5, 2, -25, 20, 2, 0, -5, -69, 23, -31, -3, -32, 6, 6, 1, 23, -51, -3, -22, 4, -15, 6, 6, -23, 18, -11, -28, 7, -22, -9, 5, -1, 5, -16, -15, -7, 0, -53, 4, -2, 8, 14, 7, -5, -31, -35, 4, -25, 0, -4, -40, 3, -27, 2, 18, -4, -58, 5, 12, -9, -16, 0, -8, -6, -37, 6, -29, -5, -2, -62, -12, 22, -41, 23, -1, -40, -5, 15, 3, 19, -4, 0, 25, -30, 3, 11, -20, 8, 3, 2, -32, 56, -25, -41, -20, -8, 4, 6, 2, 20, -5, 10, -6, -6, 4, 5, -16, 9, 6, 0, 9, 4, 0, 6, -5, 8, -4, -6, 2, 0, 10, -14, -44, 10, -10, -28, -7, 22, 34, 18, 7, 18, 2, 0, -6, -36, 6, -19, 32, 21, 8, -27, -6, 39, -19, 20, -12, -15, 15, -1, -13, -31, 23, 1, 1, -29, 14, -19, -2, 2, 12, 8, -30, 0, -6, -35, -23, 0, 18, -2, -13, 3, -17, -20, 17, -59, 2, -39, -48, 12, -23, -1, 13, -1, -44, 1, 14, 5, -7, 2, 6, -2, -65, 15, -15, 0, -5, 16, -3, 21, -25, 31, 0, -26, 3, 15, -5, 16, -2, -6, -32, -43, 4, -10, -5, 5, 0, 11, -30, 36, 3, -13, 2, -13, 11, 32, -11, -26, -7, -1, 2, -3, 5, 12, -3, -27, 0, -2, -26, 11, 4, -14, -8, 3, -10, -25, -7, -2, -8, -10, -3, 6, -2, -9, -45, 8, -20, 1, -41, 21, -8, 4, -2, 2, 0, 6, 46, 20, 6, -13, -8, 7, -28, 2, -4, 3, -20, -2, -21, -4, 9, 2, 3, 5, -6, -11, 3, 6, 32, 0, -24, 0, -6, -31, -6, -41, -2, 5, -7, 4, 12, -2, 3, 15, 4, 0, 0, 26, -3, 1, 2, -4, -4, -1, 12, 19, 3, 3, -2, 0, -39, 7, 7, -4, -4, 17, -13, 15, -33, -39, -17, -14, 3, -3, 18, 62, -8, -5, 0, -5, 28, -3, -15, 15, -4, 12, 0, 11, -29, -23, 19, -2, -29, 16, -3, -17, -8, 3, -6, 5, 6, 40, -28, -22, -9, 6, -16, -22, -1, -17, 0, 14, -3, -13, -3, -21, -46, -28, -7, -4, 24, 49, 25, -50, -12, 22, -58, -41, -1, -3, 8, -24, -19, 7, 20, 39, -50, 2, 4, -30, 6, 0, -1, 6, 54, 26, 20, 22, 15, -7, -7, -39, -7, -9, -7, -28, -32, -31, -9, -2, 1, 27, -8, -19, -31, 17, 32, -22, 14, 8, 0, 50, -7, 16, 25, 13, 41, -5, -20, -4, 38, -1, -2, -17, -5, 1, 30, -6, 26, -10, 27, 0, -4, 26, 16, -18, 32, -7, -1, 25, -28, -26, -34, 11, 6, 22, -7, 28, -23, -13, -6, 17, -4, 21, -2, 18, -44, -9, 17, -2, 9, 21, 0, -4, 8, 0, 4, -6, 40, 1, -30, 0, 6, 2, -10, -1, -5, 13, 3, 28, 1, -1, 0, -19, -3, 11, -25, -22, 3, 7, 2, -11, -27, 12, 23, 0, -8, 4, -25, 31, 21, 30, 17, 46, 10, -22, -7, 13, -14, 2, -6, 5, 10, 42, -12, -22, -7, 6, 21, -37, 18, -14, -1, 23, -17, -10, -7, -37, -6, 45, -37, -15, -9, -18, -1, -23, 10, -2, 3, -7, 0, 9, 9, 4, 7, -6, -19, -7, -7, -4, 21, -10, -3, 4, -18, 3, 6, 0, 25, -1, -1, 25, -3, -11, 5, -23, -15, 21, -13, 24, 12, 32, -2, -15, -18, 0, -37, -3, 6, 5, 0, 23, -13, 17, -14, -63, 28, 8, -8, 37, 6, -9, 12, -7, 0, 1, 17, -4, -7, 16, 1, 0, 8, 10, 4, 4, 3, 56, -15, 11, 1, -19, -5, 16, -20, 2, -7, -42, -18, -37, 22, -26, -26, 0, -2, -2, 2, 4, -2, 15, 21, -2, 27, 0, -5, 3, 36, 3, -10, -6, -41, -19, -4, -27, 7, 12, -17, -2, -2, -18, -3, 24, -33, -14, 1, -17, 0, 30, -38, 10, -9, 26, -14, 3, 37, 0, 0, 44, -4, -4, -45, 6, 2, 0, 3, -6, 0, -10, 11, -13, -6, 7, -33, 4, -29, 26, -12, -2, -3, 19, 23, 25, -17, 0, 3, 10, 9, -18, -3, -17, 3, -24, 6, -20, -1, 6, -3, -2, 5, 3, -32, 49, -24, -20, -16, 0, 4, 36, -5, 23, 8, 0, 1, -2, 6, 29, -16, -23, -8, 4, 3, -5, 2, 1, 9, 24, -23, -13, -8, -19, 18, 27, 9, 12, 32, 6, -14, -83, 27, 31, -30, 1, 2, 4, -35, -30, -10, 18, 36, 41, 41, -1, -6, 36, 10, 23, -11, 1, 10, -28, -9, -36, -19, 24, 24, 0, -37, -16, -6, 15, -3, 15, -18, -10, 2, -14, -15, -34, 13, 7, 28, 0, 46, 25, -3, 19, 4, 2, 0, -14, -6, 0, -6, 1, 32, 2, 7, 29, -27, 0, -49, -1, -62, 5, 23, -3, -2, -7, 2, -2, -20, 15, -6, -11, 0, 1, 6, 29, -1, -4, 17, -37, -9, -23, -25, 11, 3, 4, 5, 29, 0, -17, 20, -13, -12, 3, -4, 0, -12, -5, -6, 0, 32, 28, -40, 12, 2, 3, 4, -8, 3, -6, 0, -6, -20, -16, -3, -18, 5, 0, 14, 22, 2, -14, 6, -42, -6, 15, -43, 4, -5, -2, 6, -6, -32, 6, 0, 0, -46, 0, 4, 22, -23, -5, 5, 8, -30, 25, -25, -7, 16, -4, -13, -2, -20, -24, -1, -12, 19, 32, -30, -82, -1, -35, -4, -8, 9, 49, 13, -17, 29, 11, -5, 13, -4, 24, 19, -27, -7, 0, 6, -3, -36, -11, -6, 11, -2, -3, 9, 4, -41, -5, 7, -1, -1, 36, -16, 19, -38, -8, -10, -7, -23, -1, 13, -10, 6, 5, -23, -54, 18, 8, 16, 16, 0, -9, -30, 28, 8, -17, 8, -11, -16, -24, -1, 9, 16, 13, 1, -1, 7, -7, -2, 38, -6, -4, 23, -3, -2, 6, 1, 49, -11, 16, 4, 2, 28, -27, -8, 3, 2, -5, -13, -62, -45, 17, -54, 17, -5, -9, -20, -11, 3, -46, 40, 32, -56, 3, 0, 8, -77, 13, 24, -8, -14, 33, 2, -18, 24, -1, -5, -12, -27, -40, 0, 7, 33, 37, -11, -47, -4, -77, -9, -1, -17, 30, 9, -9, 58, -8, -2, 34, 4, -25, -10, 4, 45, 6, 10, -4, -5, 0, -3, 8, 8, 6, -4, 5, -15, 0, 0, -6, -5, 27, -19, 20, -16, 54, -32, 0, -34, 6, 34, 19, 3, -3, -37, -19, -2, -6, -3, 11, -2, -4, -43, 33, -39, -42, -8, -19, 9, 11, 2, -10, 19, 9, -6, -5, 18, 49, -17, -34, -5, -4, -7, -8, 5, 16, 0, 8, 0, 18, -6, -17, 7, -28, -8, 16, 6, -5, -33, -34, -38, -13, -8, -1, 5, 5, -20, -2, -6, -14, 18, 1, -5, -3, -4, 0, -9, -16, 20, -5, -12, -7, -4, -19, 57, -9, -44, -19, -36, -17, 1, -5, -1, 3, -2, -23, 3, 5, -21, -8, 0, 13, 42, -12, 60, -23, 6, 12, -3, 20, -38, -6, 48, 3, -32, -4, 30, -7, -9, -9, -18, 2, -21, 1, -21, 12, 20, -2, 6, 22, -1, 12, 3, 22, -8, -10, -38, -17, 9, 31, 5, -25, 24, 28, -49, 10, -4,
    -- layer=2 filter=0 channel=6
    -15, -9, -4, 59, -36, -48, -38, -5, 5, 28, 9, -1, 55, -4, -1, -4, -5, -28, -9, -16, -35, -7, 2, 0, 1, -1, 28, 9, 22, -1, -19, 2, -7, 26, 7, -8, 13, -13, -17, -8, 20, -8, -33, -2, -4, 2, -1, 0, -33, -45, -55, -21, -15, -30, -11, 0, -6, -20, -3, 26, 0, 8, 5, 20, 39, -58, -1, -7, -26, -17, 26, 0, -4, 0, -27, -27, 12, -3, -56, -28, 10, -20, -43, 19, 21, 37, -38, -9, -44, -7, -39, -11, 5, -61, -7, 18, 7, -18, 9, -7, 9, 18, 0, -43, 5, -1, 18, 33, -4, 2, -11, -1, -28, 8, -76, -17, 23, 8, 13, 10, -43, -5, 31, -31, -27, 23, -7, -18, -10, -6, -10, 45, -52, -39, 4, -8, -3, 21, 16, 1, 0, 2, -14, -5, -7, -5, -19, 2, 27, 2, -4, 39, 0, 6, 18, -3, 0, -11, 5, 3, -10, 22, -34, -15, -30, 6, 9, 10, 13, 13, -23, 1, 40, 6, -4, 13, -54, -78, -36, -54, -49, -17, 11, 0, -15, -27, -18, 22, 2, 35, -30, -21, 11, -49, 12, 21, 3, -8, 2, 8, -15, 34, -20, -19, 7, -4, -36, -27, 8, -28, -3, 22, 12, 9, -1, 14, -7, 5, -12, 20, 20, -40, 1, 50, -1, 0, -4, 17, 3, -6, 3, -65, -4, 0, 6, 25, 2, -6, 7, 5, -33, 36, -49, 8, 20, 30, 8, -14, -32, 0, 15, 24, -30, 3, 1, 11, 5, 1, 7, 34, -23, 19, 4, 1, -10, -25, 29, 8, 0, -3, -3, 6, -3, 33, 19, 4, 8, 3, -6, 13, 10, 1, 43, 0, 3, -9, -1, -4, 0, -5, 15, -4, 7, 11, -20, -24, 32, 40, -8, -6, 9, 2, 3, -20, -15, -22, -32, -50, -25, 7, 6, 3, -27, -13, 3, 22, -8, -22, -19, -24, 5, -26, -7, -21, -2, -2, -17, 1, 23, 17, -3, -5, -19, -9, 1, 9, -6, -7, -28, 0, -1, -17, -32, 3, 17, -5, -41, -20, 27, -34, 0, -9, 3, -14, 2, -11, 13, -3, 0, 0, 0, 14, -2, -7, 3, 0, 10, 20, -53, -11, 9, -13, 5, -3, -1, 0, -39, -4, 27, 38, -53, 23, -22, -19, 11, 6, -12, 42, 2, 7, -11, -10, -11, 22, 17, -8, 0, -6, -11, 2, 6, 29, 19, -18, 7, -6, 1, 14, 9, -1, 33, 7, -4, -11, 6, 1, -16, -3, 18, 5, 1, 5, 2, -22, 14, -20, -17, 10, 11, -3, 5, 11, 0, -137, -15, 6, -35, -21, -2, 2, -18, -6, -32, 10, -10, -28, -16, 19, -10, 14, 18, -17, 1, -20, 25, -1, 60, 25, -7, 32, -49, -1, 4, -19, -16, 6, -66, 17, 8, -15, -87, 2, 23, -7, -6, -20, 26, -23, 3, -22, 0, -12, 9, -12, -17, -2, -3, -46, 4, -8, 8, 2, 4, -7, 30, 19, 4, -9, 25, -5, 3, 18, 17, 0, 0, -8, 30, 0, -24, 18, -7, 13, 1, 6, -5, 53, -14, -29, 3, -12, -11, -2, 49, 2, 34, 23, -15, 0, 0, -7, 0, 6, 73, -8, 3, 7, -15, 0, 24, 4, -45, 7, 15, 5, -13, 12, -8, 10, 43, -23, -4, 2, 29, -5, -21, 8, 2, 1, -3, 32, -24, -8, -13, -2, -5, 29, -7, 2, -16, -53, 8, 6, 2, -7, -1, -8, -18, -17, -10, 0, -5, -24, 10, 6, 55, 25, 1, 3, -22, -9, 14, 1, 7, 7, -65, -22, 3, -45, -62, -9, 25, -2, -5, 21, 6, -17, -6, 37, 0, -5, 3, -3, 3, -18, 0, -49, 1, -5, 13, 0, 1, -6, 14, -14, -15, -15, -23, -23, 16, 7, 0, 1, 0, 3, 53, 0, -24, -8, -23, 16, 0, 0, 6, -7, -49, 15, 11, -7, -13, 7, 35, -8, -7, 12, -8, 1, -7, 2, 17, -27, -11, -7, 0, -9, -9, -6, 16, -5, -71, 7, -4, 7, -6, 18, -10, 2, -26, 0, -5, -38, 4, -11, -23, 2, 6, 6, -5, -13, -23, -8, -24, -57, -27, 4, -2, 1, 15, -12, -43, -12, 2, -10, 20, 6, 2, -17, 15, -7, 45, -22, 2, -1, -8, 85, 2, 37, 9, -1, -5, 0, -25, 11, -6, -16, 19, 13, -40, -6, 1, -4, -16, -6, 14, -5, 0, 33, 3, -2, 4, 13, 20, -10, 4, -51, -3, 6, 18, 16, 2, -5, 18, -3, -6, -10, -8, -7, 1, 13, 17, -34, -35, 2, 21, -7, 27, -57, -10, -8, 0, 0, 1, -1, -41, 15, -5, 1, 5, 8, -28, 2, 35, -24, -10, -5, -5, 24, 32, 6, 53, 4, -2, 2, 1, -3, 17, 9, -52, -16, -14, 1, 2, 4, -57, 1, -27, 37, 22, -1, 25, -8, 0, 19, 36, -7, -3, 4, 8, -66, -15, -9, -17, -16, 11, -1, 18, -9, -8, 5, -7, 18, -24, -36, 3, -18, 6, -5, 16, -15, 6, 4, -39, 67, -4, -2, 16, 0, -49, -9, -2, -7, -4, 6, 18, 22, -18, -3, -21, 6, -41, 31, 54, -40, -5, 12, 1, -8, 5, -11, 24, 22, 5, -19, 7, 12, 24, 14, 7, 0, -14, 19, -38, 18, 10, -3, -3, 18, 25, 6, -35, 1, -16, -19, -40, -6, -4, -4, -3, -5, 1, 44, -5, -8, -32, -3, 11, -1, 11, -8, -2, 18, -1, 1, -6, 5, -8, 0, -29, 6, -9, -15, -1, -2, 15, 1, 49, -18, 3, -1, 3, 13, -49, -8, 37, 8, -17, 23, 9, 7, -25, 16, 13, 3, 0, 0, -31, 7, -24, -16, 11, 38, 16, -4, 1, -44, 21, 12, 1, 4, -15, 23, 30, 1, 9, -10, -30, 0, 30, -4, 1, 20, 7, 22, -13, -7, 5, -19, 0, -21, -8, 17, 5, -5, -9, 6, 9, -1, 0, -42, 22, -5, -4, 6, 0, -32, 0, 3, -3, -2, -6, -18, 4, -21, 23, -2, 3, 3, 17, 21, -30, -4, -47, 20, 9, 20, 3, 4, -19, 5, 36, 23, -3, -26, 6, 19, 21, -3, 0, 28, 15, 12, -10, -13, 10, 12, 3, -2, -12, -7, -11, 7, 4, 15, -16, 17, 22, 2, -9, -23, 15, -7, -12, -4, -11, -13, 1, -3, 19, 18, -13, -13, 4, -19, -15, -12, 0, -4, -21, 27, -9, 1, 3, -2, -20, 0, -54, -12, -14, 28, -6, 5, -22, -34, 5, -10, -2, 12, 16, -43, 10, 18, -6, -55, -26, 3, 0, 5, -1, -22, 25, -26, 14, -11, 14, 5, -15, -50, -12, 0, 11, 22, -15, 10, 27, -4, 13, 1, 0, 20, 4, -5, -7, 17, 7, -21, -24, 16, 6, -17, 0, -6, -5, -12, 0, 5, 14, -15, -28, 0, 3, -9, -1, -9, 7, -27, 13, 5, -6, 47, 54, 17, 0, -9, -1, 4, -41, 25, -28, 1, -11, -27, 0, 6, -5, 0, -40, 5, -16, 4, 1, -1, -47, 17, 24, 5, 2, -10, 21, 3, -15, 2, -50, -19, 17, 0, -21, -12, -35, 7, 17, -16, 5, -13, 38, 2, -68, 1, -34, 1, 2, -16, 6, 27, -49, -58, -66, -47, -18, 0, 15, -17, -25, -10, 3, -1, 3, -32, -7, 15, -11, -43, -5, 19, -32, 5, 4, -39, -1, 4, -17, -9, -2, -10, -15, -25, 0, 1, -13, 6, -38, 8, 37, 3, 1, 14, -38, 0, -3, 26, -6, -42, -3, -23, -31, 13, 5, -20, 7, -13, -5, 1, -6, -3, 22, -7, 10, -21, -11, 7, -8, -39, 9, -29, -14, 3, 30, 22, -12, -42, -13, -19, -16, -2, -8, -11, 2, 20, -13, -9, 3, 5, -10, -8, -38, 14, -15, -4, -3, -10, -8, 19, -33, -4, 4, -39, -2, -6, -41, 2, -1, 40, 0, 7, -2, 4, 9, 9, -11, 3, 34, -36, -19, -12, -47, -36, -4, 2, 4, -5, -32, -16, -54, -14, -82, 40, 6, 3, -19, -47, 21, 3, 3, 12, 24, 31, 35, -9, 27, -47, -14, 39, 12, -5, 33, 1, -5, -26, -10, -9, -48, 13, 42, -10, -35, 47, 16, 18, -85, 0, 19, -1, -46, -25, -17, -9, 1, -18, 0, -13, -5, 4, -23, 7, -2, -59, -2, -1, -18, 5, 2, -3, 30, 10, 22, -42, 41, -31, 15, -16, 4, -40, -2, -5, 41, 33, -4, 32, -8, 24, -32, 4, -53, 15, 11, -4, 6, -59, -3, 8, 5, 1, -36, 47, -15, 3, 1, -18, 17, -1, -103, 2, -1, -8, -2, 4, -6, -4, -65, 16, 1, -3, 12, 19, -7, -15, -85, -31, -17, -58, -16, -28, -36, 5, -8, -11, -4, -18, -25, -96, -44, -41, -100, -45, 9, 2, -2, -10, -47, 16, -6, -5, 18, 16, -13, 5, 22, -49, -14, 13, -63, -3, 28, 22, 20, -15, -4, -10, -5, 0, 2, 20, -77, -1, 6, -16, -87, -8, 4, -4, -26, -17, -41, -24, -1, -4, -3, -32, -1, 26, -12, 2, 4, -75, -1, 13, 5, -4, 1, -6, 24, -2, -24, -33, 64, -38, 0, -28, 13, -6, 5, -7, 14, 8, -58, 19, -4, 16, -12, 0, -13, -21, -35, 11, 0, -55, -1, -5, -16, -1, 3, 25, -14, -4, 4, -9, 34, 6, -29, -10, -4, -10, 5, 5, -4, -4, -15, 9, 13, -6, 20, -1, -3, 6, -39, 16, -30, -52, 10, -30, -4, 0, -1, -9, 2, 8, -30, -11, 12, -15, -52, 58, -21, -6, -38, -77, -33, -4, 0, -18, -3, -16, 14, 17, -2, -47, 12, -7, 0, 0, 25, 34, 6, 13, 16, 0, -79, 12, -32, 28, -36, -30, 13, -33, -5, 0, 15, -1, 11, -10, 3, -13, -2, 8, 3, -4, -2, 17, -16, 3, 6, -41, 0, 2, -5, 21, 6, 3, -16, -11, 4, -35, 44, -32, 3, -9, -10, 1, -5, 0, 54, -14, 44, 11, 12, -31, 29, -4, 21, 0, -12, -12, -12, 0, 3, -15, 0, -7, -23, -17, -16, 3, -2, 26, 34, -12, -66, 1, -3, -15, 11, 3, -14, 2, -29, -28, -12, 6, 3, 5, -2, 4, -24, -46, -11, -13, 8, -24, 6, -6, -2, 0, -5, -29, 2, -43, 9, -16, -10, 17, 12, 5, 14, -4, -2, 6, 5, 7, -6, -15, -31, -5, 20, -41, 3, 3, -7, -2, -51, 50, 3, 0, -29, -10, -6, -32, -19, 13, -28, 9, 6, 14, 0, -18, -27, -5, -9, -13, 25, -8, 4, -25, -4, 13, -2, 9, 14, -9, 2, -27, 1, -50, 33, 19, -4, 0, 23, 24, 0, -8, -3, 1, 6, -11, -21, -7, -7, -2, -18, -32, -25, -19, -12, -19, 4, 0, -26, 37, 34, -30, -68, -22, 1, -29, -24, 10, -6, -17, -14, 0, 5, 9, -49, 15, -1, 7, -5, -24, 8, 5, 43, 6, 4, -15, -18, -6, 2, 3, 30, -3, -1, -15, -19, -36, 46, 38, -1, -10, 18, 8, 0, -9, -45, -3, 7, -1, -7, 30, 34, 0, -7, -25, 2, -16, -6, 9, -20, 11, 8, 6, -15, 4, -18, -11, 33, 9, 2, 60, -14, -39, 13, -11, 30, -61, -14, -23, -7, 9, -6, 27, 0, 6, -39, -6, -34, -15, 14, -7, 4, 25, 7, 49, -7, 14, -20, 10, 2, -46, 2, -28, 10, -24, 6, -2, -1, 17, -11, -9, -59, 19, -6, 6, -7, 10, -47, -3, 44, -33, 3, -29, -16, -19, -6, 4, -60, -5, -16, 6, -49, -58, -1, -1, -35, -8, 8, -24, -2, 7, 3, 11, -55, -10, -63, 0, 1, -13, 0, 2, -8, -4, 18, -8, 13, -2, 2, -9, -57, 19, 0, -8, -46, -13, 21, 3, -23, 17, -1, -2, -4, 7, -14, -52, -39, -7, -11, 19, -11, 3, 2, 11, 28, -4, -14, 10, -8, -67, 15, -32, 2, 0, -9, 5, 2, 7, 2, 75, -26, -34, -25, -9, -16, -10, 14, -55, -81, -54, 12, -28, -30, 6, 48, -4, -6, -28, 2, -15, 0, -42, -4, -20, -6, -43, 12, 13, -2, -96, -4, -1, -16, -10, -5, 7, 28, -26, 22, -11, 3, 8, 2, -4, 10, -25, -114, -6, 25, -38, 33, -53, 8, -6, -16, 0, -38, -36, -53, 28, 3, -47, -7, -4, 53, 4, -5, 31, 0, 4, 1, 1, -1, 12, 12, 6, -5, -18, -14, -5, 4, 1, -16, 17, 36, -6, 16, -11, -28, 0, 1, 44, -37, -23, 17, -10, -56, -14, -32, 0, -4, 9, -4, 51, -83, -12, -26, -33, 13, -6, -34, -23, -30, 12, -9, 20, 13, 21, 2, -49, 28, -75, -14, 22, -11, -4, 48, 62, -14, 4, -9, -3, 9, -5, 18, -35, -48, -28, 2, -3, -54, 13, 76, 0, 0, -31, -8, 5, -7, 11, 1, -25, -2, 34, -11, 16, -2, -22, 3, 14, 0, 14, -1, 0, 9, -7, 5, 4, 11, -29, 8, -30, 0, -53, -43, -6, 29, -8, 11, -8, 14, 20, 13, 1, 2, -64, -57, 13, -5, 15, -1, 17, 2, 0, -13, 51, -4, 6, -4, -25, 4, -40, -109, 8, 0, -20, -12, 2, -28, 11, -48, 34, 56, -6, 24, -3, -2, 47, -39, 43, 9, -59, -48, -33, -12, -42, -22, -2, -8, 1, -1, -19, -47, -22, -13, -56, 34, -10, -36, 2, -12, -4, 9, 23, 3, 52, -7, 16, 43, -112, 14, 69, -30, 6, 31, 9, -22, 1, -17, -6, 42, -3, -5, -15, -68, 34, 14, 15, -95, -2, 28, 7, -21, -16, 11, -32, -5, -42, -1, -38, -5, 18, 0, 30, 6, -3, 1, -25, 7, 54, -6, 4, 19, -4, -34, -38, 37, -6, 52, -32, 24, -45, 2, -1, 33, -46, -49, 1, 1, 3, -8, 0, -91, -65, -54, 11, -38, -58, -11, 4, 44, -8, 11, 52, -11, -1, 1, 3, 18, -17, -86, -2, -7, -9, -5, 2, 11, 7, -1, 4, 23, 0, 39, 15, 18, -21, 14, -25, -24, -109, -79, -12, -19, -48, 3, -10, 2, -34, -24, -56, -75, 3, 8, -10, -81, -1, -79, -55, 22, 11, 0, -12, -5, 3, 14, -40, 29, -101, 0, 45, -3, 9, 42, 11, 13, 26, -55, -11, 46, -23, 10, 10, -10, -25, 28, -33, -64, 9, 20, -1, -26, -34, -7, -25, -1, -14, -7, -37, -19, 36, -5, 18, -7, -31, 7, 9, 12, 39, 0, -3, 11, -17, -23, -5, 61, -17, 30, -29, 23, -14, -33, 5, 34, -31, -83, -28, 17, 4, -2, -4, -39, 6, -13, 20, -69, -104, -9, -5, -7, -5, 28, -13, -12, -3, 6, 8, 27, -20, -69, -1, -7, -23, -17, -7, -7, -8, -3, 12, 13, -5, -3, -2, 29, 19, -11, -16, -14, 3, -11, -66, 17, -17, -4, -2, 3, -5, 13, -47, -11, 21, 4, 28, -62, -9, -19, -64, 16, 19, -2, 22, -1, -44, 19, 3, 14, -70, -17, 1, 23, 0, 43, 22, 7, 13, 7, 0, -22, -47, 8, 22, -55, -47, 14, -28, -1, 3, 0, -1, -18, -32, -5, 14, -6, -41, 1, 5, 0, -6, 0, 11, -4, -52, -1, -56, -14, 19, -7, 0, 15, -33, 23, -27, 54, 10, 3, 8, 18, -13, 18, 3, 29, -2, 35, -13, 19, 10, 43, -1, -8, 20, -13, 8, -25, -26, 6, 4, -26, 1, -3, -1, -19, 1, -4, 6, 22, 4, 12, 1, -2, 15, 1, -3, -9, -5, 14, -22, -26, -1, 12, 11, -37, 4, -7, -42, -14, 9, -10, 3, 3, -11, -19, 6, 0, 15, -23, 14, -28, -47, 22, 8, 0, -9, -47, -12, -18, -8, 4, 18, 11, -2, 38, 53, -7, -13, 3, -3, 15, 9, -42, 44, 8, -13, -11, -6, -47, -85, -34, 3, -23, -35, -6, 9, 5, -24, 7, -6, 20, -37, 11, -10, 5, -19, -1, -11, 4, -18, -21, -11, 3, -50, -7, -47, 20, -9, -2, -3, 17, 14, -14, 0, 0, 27, -19, 24, 6, -22, 30, -1, 29, -8, 40, -13, -10, -32, 16, -1, 16, 76, 0, -10, -29, -3, -10, -25, 0, 1, -23, -3, -5, 2, 8, 10, -23, 17, 23, 3, -1, -23, -17, -5, -1, -1, -12, -28, -40, 3, -9, -4, 0, 15, 23, -22, -15, -39, 46, 39, -28, 15, 11, 7, -4, 40, -54, -10, 23, 4, -10, -25, 47, 4, -26, -59, 32, -18, -2, 23, 8, 6, 6, 38, -13, -35, -13, -17, 51, 4, 9, 22, 10, -32, -19, -4, 47, -48, -21, -21, -54, -19, -3, 43, -29, 11, 0, -5, 9, -33, 15, -10, -1, -17, -1, -16, 13, -16, -16, -6, 2, -34, 7, -49, 1, -37, 1, 0, 17, 15, -5, -1, -20, 3, -26, 26, -25, -6, -26, 0, 46, 32, 7, -22, -22, -17, 38, 1, -28, 31, 2, 32, -26, -46, 0, 4, -29, -11, 15, -35, -8, -6, 3, 0, -28, -1, -55, 3, -1, -13, -28, 5, -33, -5, 1, 5, 5, 0, -10, 0, -28, 0, -14, -37, -32, -76, 42, -29, 33, 34, -17, 6, 4, 26, 17, -33, -44, 25, -1, 48, -64, 6, -2, -15, 26, -9, 0, 9, 10, -30, -18, -49, 4, -62, -11, -10, -12, 0, 11, 53, -38, -29, -16, -11, -62, -47, -3, -61, -36, -49, 32, -10, -44, 5, 16, -6, -48, -47, 13, 17, 3, -35, -3, 16, -4, -40, 18, 13, 0, -66, -7, 20, -20, 17, -1, -3, 52, -32, -23, -7, 19, -20, -3, 5, 17, -16, -57, -3, 15, 10, 34, -43, 16, 16, 16, 4, -28, -39, -38, -11, -25, -8, 1, 15, 33, 1, 15, -24, -15, -3, 6, 2, 19, -35, -67, -4, -2, -17, -1, 4, -36, -7, -49, 20, 43, -3, 3, -8, -52, 15, -19, 10, -34, -48, -23, -44, 4, 27, -23, 2, 0, -8, -13, 11, -34, 22, 9, -29, -27, -8, -11, 24, 13, 7, -8, 6, 30, 25, 3, -25, 36, -110, -11, 24, -6, 6, 1, 36, 38, 15, -2, -10, -69, -66, 4, 0, -73, 9, 35, 18, -61, 3, 18, -3, -18, -16, 5, -21, -2, -15, -9, -5, -8, 16, 19, 24, -2, -25, 0, -25, -21, 39, 1, 2, 4, -2, -24, 22, -29, -26, 30, -7, -1, -94, -16, -2, 7, -36, 7, -52, 12, -7, 13, 1, -39, -56, -50, -21, -61, -7, -8, 1, 45, 2, -14, -2, -4, 2, 8, -20, 22, -53, -65, -7, -9, -70, -8, -8, -46, 7, -32, 4, 52, -4, 51, 21, -50, 4, -14, -20, -10, -99, -81, -26, -28, -16, 19, 8, -4, -38, -2, 62, -83, -9, -27, 5, -25, 4, -21, -46, 30, 57, -12, -7, -3, 19, 16, 10, 57, -110, -34, 49, -12, -3, -36, 1, 6, -47, -12, -2, -1, -70, 14, -28, -29, 43, 44, 35, -126, 6, 32, -6, -39, -28, 36, 16, 0, -46, 5, 2, 8, 23, 27, 24, -5, -59, 0, -14, -9, 66, -1, 7, 25, 12, -18, -2, -20, 1, 70, -33, 39, -48, -29, 7, 15, -58, 68, -104, 30, -4, -8, 2, -20, -44, -41, -10, -51, -5, -2, 17, 27, 5, 21, 2, -5, 6, 6, 24, 2, -46, -50, -1, -8, -43, -10, 4, 0, 0, -16, 28, 40, -3, 45, 8, -39, -16, 19, -14, -31, -95, -26, -65, 0, -3, 20, -4, -8, -3, 48, 14, -87, 28, -3, 16, 11, -3, -36, 0, 36, 26, -8, 31, -2, 0, 3, -6, 44, -82, -36, 53, 5, 1, -6, -17, 6, -65, -11, -6, 9, -9, 3, -30, -70, -2, 47, 4, -41, 14, -12, -4, -30, 12, 59, -71, 4, -21, -6, -22, -13, -14, 44, 26, -6, -112, -6, -5, -23, 59, -4, 2, -10, 15, 7, -18, -9, 8, 45, 20, 32, -53, -2, 6, 22, -53, -85, -32, 14, 2, -21, 3, -40, 7, -12, 37, -44, -92, 5, 17, -33, -6, 8, -37, -13, -6, -2, 4, 12, 4, -36, 5, 7, 7, 8, 1, -27, 5, -2, -24, -3, -1, 15, -9, -10, 24, -9, -28, -53, -18, 5, 6, 31, 34, 19, 2, -4, 14, -22, -24, -43, 24, 0, -67, -72, -6, -50, 39, 16, 7, 0, 17, -10, -26, 5, 37, 8, -109, -1, -2, 5, 1, -15, 22, -6, -16, 3, -9, -58, -62, 14, -16, -57, -54, 7, -38, -27, -7, 20, 7, 15, -77, 5, 3, -5, -4, -3, -40, 13, -22, 4, 23, 1, -64, -6, -24, -39, 31, -4, -4, -19, 1, 13, -9, 5, 14, 0, 18, -1, -33, -17, 0, 58, 3, -25, -22, 23, 13, 51, -2, -8, 37, 34, 5, -1, -38, -6, -5, -29, -3, 0, -1, -1, 1, -3, 5, -2, -17, -27, 2, 0, -26, 8, -5, 4, 4, -27, 3, -16, 5, -12, 13, 4, -11, 29, 3, -29, 22, 60, 13, 6, -12, -1, 0, 4, 34, -35, -39, -41, -21, -6, -75, -21, -9, -11, -48, 10, -21, 13, 9, 35, 7, 22, 40, 20, -14, 15, -27, 13, 0, -1, 6, 39, -2, 4, -8, 5, -16, -24, -11, -45, -46, -9, -12, 0, -11, -55, -4, 4, -46, 0, 47, -3, -6, -2, 5, 3, -13, 1, 21, -2, -13, 2, -8, 8, 13, 4, -1, 54, -31, 4, -23, 0, 58, -18, 17, 4, -1, -11, 0, 73, 8, 66, 6, -9, -24, 32, 0, 0, 7, 15, 4, -29, 27, 1, -6, -19, 0, 2, 15, -6, 2, -4, 18, -26, -13, 25, 0, 9, 17, 0, -6, 37, -3, -7, -15, -8, -4, -20, 10, 13, 4, 13, 23, -55, -48, 37, 26, 8, 56, 29, -4, 2, 5, -72, -31, -20, 4, -10, 16, 31, 6, 29, 37, 16, 6, -6, 23, -33, 9, -7, 17, 5, -45, -26, -28, 9, 7, -7, 31, -44, -30, -10, 2, -37, -46, -9, -18, 5, 1, -1, 21, -14, 4, -26, 4, 13, -27, 13, 26, -6, 5, -4, -19, 2, -24, 20, 12, 0, 0, 4, -49, 21, -6, 0, 7, 8, -3, -6, 29, -13, 12, -1, 18, 0, 19, -73, 5, 0, -30, -22, -65, -10, 8, 17, -8, -43, 29, -5, 3, -28, -26, -19, 15, -59, 1, 31, 9, -3, -2, 7, -43, -20, 11, -14, 0, -1, 11, 13, 1, 23, -1, -1, -12, 3, 0, -5, 23, -18, -17, 13, 9, 22, 3, -3, 1, 4, 28, -22, 1, -8, 7, 31, -66, -40, 16, 27, 29, -35, -10, 0, 7, 5, 14, -1, -26, -21, 13, -18, -3, 3, -21, 18, -13, -19, 8, 14, 44, -62, -56, -44, -5, -9, -13, 4, -30, -38, -4, 5, -11, -40, -2, -2, -3, 7, 21, -4, 8, 5, 3, 2, 11, 1, -24, 6, -4, 5, -37, -7, 46, 5, 8, -7, -3, -9, -14, 21, 10, -33, -17, -18, 2, 22, 5, -26, 5, 34, -26, 27, -2, 2, 34, -31, 5, -27, -39, 0, 24, -15, -47, 9, -9, 6, -5, 31, -29, 0, 0, -6, -39, -15, 0, 4, 2, 3, -6, 11, 2, -27, 6, 12, 21, 42, -1, -10, 11, -31, 21, -13, -19, -5, -38, 10, -40, 33, -11, -9, -2, -3, 48, 31, 0, 13, 16, 15, -2, -57, -10, -31, 18, 18, 20, -14, -5, -5, 38, 31, 27, 10, -33, 22, 7, 24, -3, -17, 64, 23, -11, -46, -5, -21, -43, 13, -51, 0, 30, 25, -26, -63, 4, 21, -6, 58, -10, -9, -25, 4, 17, 1, 19, -5, 0, 31, 35, 3, -55, 1, 2, -27, 19, -5, -7, -61, -14, -7, 12, -5, -21, 22, 14, 6, -31, -33, -7, -9, -61, 41, -64, 19, 6, 9, 0, -16, -25, -55, 0, -28, -24, 5, -7, 8, 2, 29, -8, 1, -3, 6, 10, 24, -27, -31, -7, -5, -51, 11, -9, -16, -7, -59, 6, 21, -4, 29, 11, -86, -34, -5, -25, -5, -16, -1, -6, 19, -25, 27, 0, -3, 0, 55, -57, -43, -10, -11, -44, -23, -5, -36, -25, -5, 1, -9, -37, 41, -17, 6, -20, 26, -72, 6, 6, 10, -3, -54, 37, 47, -27, -16, -8, 0, -58, 16, -29, 4, -13, 33, -30, -17, 18, -30, 5, -42, -18, 11, 35, 2, -14, -3, 4, 9, -10, 17, 2, -4, -11, 0, 8, -3, 16, 0, 8, 27, -24, 37, 13, -74, 19, 31, 8, 12, -10, 17, 5, 34, -35, 13, -19, 21, 10, 29, 0, -3, -8, -4, -2, 9, -30, -4, 40, 60, -4, 25, -8, -2, -4, -1, -7, 29, -29, 11, -7, -7, -22, 5, 4, -11, -3, 6, 22, -6, 0, 28, 14, -47, -14, 30, -8, -43, -3, 17, 52, 31, 3, 20, -8, 5, 4, -22, -38, -18, 5, -15, -31, -37, -3, -18, -5, 32, 9, -8, 44, 8, -10, 15, 42, 21, 5, -17, 43, 17, 3, -13, -30, 19, -73, -25, -4, -1, -23, 38, -16, 19, -4, 22, -15, -83, -2, -30, -6, -31, -18, 5, -14, -5, -8, -7, -40, -11, 12, 49, 43, -6, -81, 5, 21, -22, 37, -6, 7, -10, 4, -1, -22, -40, 27, 46, 16, 15, 15, -8, -1, 52, -13, 9, -27, 15, 20, -14, -6, -17, 12, -38, -12, 6, -48, -7, -8, 16, 8, 22, -30, -13, 0, -3, 24, 18, -47, -11, -5, -8, -11, 4, 5, -4, -8, 26, 13, 15, 4, -7, 24, -14, 4, 34, 10, -9, -20, 5, 5, 32, 38, -12, 6, -10, 34, -24, -55, -80, 2, -6, -53, -76, -8, -35, 23, -10, 4, -5, 35, -44, 18, 24, 17, 31, -35, 12, -3, 10, 6, 43, 29, -17, -5, -10, 3, -57, -35, 9, -5, 1, -18, 14, -8, -46, -1, 9, 6, 17, -43, -5, -26, 4, 0, -2, -35, 0, -40, 13, 27, -6, -38, -4, 0, 19, 37, 7, -5, 12, -18, -24, -6, 26, 37, 20, -11, 20, -21, -12, -2, 67, -44, -19, -78, 6, 37, 42, -7, -6, 1, -29, -22, -10, -26, 12, 45, -23, -8, -4, -6, -9, 7, 0, 39, 5, -29, 1, -7, 1, 0, 9, -3, 34, -6, -34, 8, 4, -7, -9, 23, -50, -2, 0, -22, -52, -40, 23, 18, 6, 27, 12, -2, -5, 3, 28, -58, 10, -6, -11, -25, -36, 2, 6, -25, 25, 5, -11, -10, -14, 42, -12, -10, 19, -28, -17, -20, 18, -2, 12, 2, 24, -18, -48, -9, -20, -50, 6, 5, -5, -41, -7, -13, 2, 13, -42, 4, 10, -61, 12, 31, -4, 32, 1, -39, 9, -18, -5, 8, -7, -67, -2, -56, 34, -9, -7, -6, 15, -7, 7, 15, 1, 28, -28, 32, -6, 0, -43, -5, 10, -27, 6, -16, 11, 16, 12, -8, -4, -29, -6, 8, -16, 8, -5, 0, -8, -7, 3, -1, 0, 7, -1, -2, 6, 0, -1, 0, -1, -4, -16, 6, 26, -9, -28, 5, 7, 2, -11, 1, -21, 22, -14, 0, -44, -78, 10, 13, 15, 18, 23, 1, -10, 40, -22, 11, -40, 5, 0, 18, -1, -1, -8, -21, -13, 10, -3, 4, -55, 14, -13, 4, 0, -17, -36, -4, -12, -3, -6, 53, 7, 27, -53, -6, 21, -50, 2, -1, -37, -21, -6, -1, -7, -9, -39, -2, 1, 2, 22, 22, -6, -6, 7, -13, -4, -30, -1, 5, 5, -19, 0, -5, 37, 14, 6, -1, 12, -1, 7, -17, -20, -2, -2, 2, -1, 5, -18, -7, -8, -64, 0, -12, 18, 7, 3, -6, -37, -4, -6, 16, 1, -21, -8, 3, -12, 10, 15, 9, -21, -6, -1, 29, -8, 8, 9, 4, -5, -10, -32, 0, 13, -3, -22, 29, 5, 0, 1, 21, -14, 2, 5, 5, -22, -46, -22, -9, 11, 21, 1, 0, 0, 22, -4, -131, -12, -5, -12, -37, 7, -6, -25, 10, 17, -3, -2, 19, 12, 33, 2, 39, -5, -24, -12, -7, -3, 2, 19, 77, 26, -10, -41, 2, -46, -25, 24, -54, -9, 24, 13, 21, -13, 5, -48, -1, -3, -36, -2, 34, -2, -8, -2, 11, 4, 9, -28, 12, 3, -67, 6, -29, 21, 14, -3, -3, 24, 30, -1, -42, -39, -8, -4, -15, 9, 0, -19, -7, 10, -19, 0, -25, 6, 27, -36, -7, -8, 9, 7, 34, -11, -6, -4, 18, -3, -1, 12, 12, -14, 0, -4, -4, -20, -31, 17, -2, 3, -18, -23, -8, 22, -7, 4, -6, -30, -2, -7, 16, -23, -35, 8, -8, 43, 27, 12, -11, 5, -14, -8, 1, 6, 37, 1, -62, -20, -7, -4, -6, 7, 5, -34, 23, -25, -21, -5, 5, 6, -2, 2, -6, -23, 8, 8, -23, 1, 5, 4, 52, 9, 9, -24, 0, -31, -25, 17, -18, 16, 20, 0, 3, -20, 20, -54, -1, -33, -5, -16, 38, -5, -3, -7, 34, 0, -20, 0, 20, 1, -44, -5, -17, -6, -9, -2, -4, 6, 19, -107, -29, -29, -25, -13, 21, 5, -55, -6, -1, -21, -12, 46, -54, 2, -7, -13, -8, -28, 10, 20, 13, 4, -21, -4, -12, -35, 4, 26, 16, -19, -6, 0, -26, -41, 12, 21, -8, 2, 0, -28, 4, 12, -2, 22, 5, -46, 5, 0, 13, -13, -21, 10, 13, 20, -23, 7, -19, 32, -1, -13, -2, 3, 54, -22, 9, -50, 32, 18, 19, 8, -5, 12, -11, 1, -21, 3, 15, 11, -35, 8, 4, 2, -4, 43, -16, 39, -5, -18, 43, 22, 4, -32, -8, 22, 5, 15, -29, 7, 15, 14, -5, -5, 11, -2, 4, -49, 11, -25, 40, 4, 1, -4, 25, 0, -43, 10, 29, 4, -62, 1, -13, 5, -17, 5, -2, 12, -49, 8, -42, -31, -30, -16, 15, 5, -20, -31, 6, 28, -42, 21, 4, 2, 20, -14, 6, -24, 22, 3, 13, 33, -20, -2, 10, -14, 0, 10, 42, -6, 0, 0, 24, -35, -26, -6, -5, -1, 6, 4, -2, 32, 2, 15, 20, -27, -4, 20, 5, -15, -3, 49, 1, -4, 1, -5, -5, 27, 22, -22, -7, -9, 13, -16, 19, -11, 24, -7, -6, -13, 0, 1, -29, -9, -3, -1, 43, 34, -2, 41, 7, -23, -13, 41, 9, 25, -4, -18, 36, -17, -36, -26, 4, 13, 11, 0, 27, 22, 1, 4, 21, 29, 11, -37, 7, 12, 2, -38, -22, 0, -13, -9, -15, 10, 22, 19, 16, -8, -86, -7, -3, -12, -10, 0, 5, -21, -8, 12, -21, -24, -29, 2, 11, 8, 8, -13, -4, 23, -53, 13, -25, -7, 17, 0, -1, 26, 32, -6, 8, -3, -12, 13, 13, 24, 6, -2, 36, -11, -5, 7, 16, -2, -3, 3, -5, -3, -18, -20, -6, 20, -3, 26, 9, -4, 6, -3, 19, -5, 5, 16, -26, 0, 14, 30, 9, 0, 0, -13, 5, -7, -8, -22, 33, -38, -2, 10, 3, -14, -9, -25, 6, 15, 7, 0, 7, -25, -4, 13, 24, -14, -42, 43, 3, 26, 3, 52, 31, 10, -4, -22, 1, -2, -20, 18, 9, 10, 13, 22, 20, -12, 1, -49, 0, 43, -41, -44, 44, -1, 0, 0, 39, 2, -1, -10, -3, 6, -58, 5, -25, 0, 0, -4, 7, 19, -21, 7, -23, -12, -2, 7, 31, 0, 13, -17, -7, 27, -42, 37, -38, 12, 20, 34, -4, 12, 36, -12, -16, -18, 11, -1, 28, -42, -3, 27, 20, -15, -1, 0, 3, -28, -42, -76, -5, -2, -7, -6, -7, 23, 2, 15, 4, -13, 1, 2, 6, -14, 16, 3, -12, 25, 0, -5, -6, -33, -7, 4, -1, 0, 4, 10, -29, -6, 17, -17, 11, -32, -2, -24, -56, 12, 2, -6, 20, 7, 10, -39, 20, 13, -3, -2, -36, 27, 6, 23, 8, 4, -1, -45, 0, 19, -8, -21, -31, -33, -12, 0, 5, -30, 1, -73, 6, -3, 9, -3, 33, -2, -19, 3, 26, 0, -31, -1, 2, 0, -44, -6, -41, 14, 11, -2, 5, 5, -23, -12, 18, -22, 22, 13, 37, 23, -3, -53, 5, 22, 5, 54, -28, -6, 39, 37, 4, 6, 12, -40, 28, 0, -26, -11, -6, 18, -8, -11, -8, -4, 2, 2, 37, -1, -31, -32, -8, 0, -15, 10, 2, 30, -4, 3, 12, -7, -7, -6, 14, -8, 47, -34, -18, -45, -45, -29, -8, 3, 67, 18, 0, 1, 67, -13, 17, 21, -15, -10, -9, -14, -5, -7, 46, -18, 3, 0, -17, 17, -3, -24, 25, 18, 5, -13, -28, -15, -2, -14, 30, 23, -22, -1, -7, -77, -22, 5, -12, 58, -52, 22, -1, -21, 1, -37, -5, 37, -6, 18, 1, 4, 33, 5, 11, 2, -20, 16, 50, -5, 23, 3, -22, 30, 16, 2, 8, 37, -23, -25, 27, -7, 19, 0, 13, 15, -35, 9, 5, -13, -60, 21, -20, 31, -29, 10, 5, 19, -25, 14, 17, -37, -1, -2, 0, -18, 2, 15, 0, -9, 2, 5, 25, 17, -12, -20, 4, 5, 11, -8, 2, 11, -1, -56, 0, -10, -2, -16, 17, 5, -1, -14, -51, -17, -31, -5, 4, 30, 29, -13, -1, 3, 16, -30, 14, -1, -9, -11, -5, 6, -10, 22, -16, -24, 4, -13, -4, 12, -2, 1, 43, -16, -36, 26, -38, -18, 5, -42, 37, 0, 24, -19, -3, -92, -17, 2, -2, -21, -22, -1, 4, -57, 10, -19, 0, 18, -9, 3, 17, 6, 33, -3, 26, 2, 16, -13, 19, 4, -19, 0, -36, 25, 12, 1, -6, 34, -10, 11, -20, -82, 39, -8, 17, -5, 18, 9, -2, -62, -26, 44, -35, 13, -32, 12, -4, 28, -30, 43, 30, 3, 2, -8, 4, -25, -12, -12, -1, -8, 6, 6, 42, -21, -12, 13, 0, 4, -39, -17, 1, 14, 0, 27, -25, -7, -2, 3, 10, -10, -3, 11, -22, 5, -15, 3, -18, 16, 10, -25, -6, 1, 6, -18, -7, -35, 18, -7, 5, 5, 3, 31, 0, 26, -6, -7, 31, 21, -25, 0, 29, -22, -14, 5, -8, 12, 0, -36, 48, -12, -14, -24, 1, -35, 12, 25, -9, -32, -17, -4, 9, -18, -5, -1, 2, 22, -14, -20, 49, -7, -21, -3, -32, 1, -3, -32, 26, 7, -38, 0, -4, 28, -8, 0, -5, 23, -2, 3, -46, -84, 38, -25, -14, 1, 22, 18, 3, 6, -14, 30, 10, 2, 3, 9, -6, -6, 19, -20, 18, -18, 6, -5, 0, 21, -7, 3, 35, -6, -1, 3, 15, -21, 7, 0, 7, -5, -33, -18, 3, 20, -3, 34, -17, -49, -3, 9, -9, -19, -3, -12, 19, -9, -14, -14, 21, 4, -7, -19, 1, 0, 60, 1, -61, -47, 22, -33, -5, -25, -7, -29, -16, -11, -26, -11, -15, 3, 1, -13, 34, -17, -28, -3, -26, -11, 0, -4, 47, -3, -21, -38, -5, -52, -6, 29, -35, -15, -5, 0, -4, -56, 13, -49, -1, 39, 0, -51, -24, 1, -18, -5, 3, 5, -14, -44, 8, 3, -27, -5, 16, 24, 0, -6, -4, -1, -17, 11, -53, -18, 21, -4, 7, -11, -7, -2, 4, 18, 6, 35, 21, 8, 0, 10, 1, -25, -3, 27, 12, 4, -31, 0, 16, -13, -4, 9, 41, -16, 7, -2, 7, -73, 5, -93, 0, 3, -55, 2, -1, 24, 0, 35, 4, -16, 5, 6, 6, -38, 10, 4, -25, 9, 12, -44, 25, -27, -36, 26, -3, -6, 3, -7, -105, -15, 3, -1, -16, 3, -8, -21, -19, 11, -7, -11, 19, 7, 21, 26, 7, -12, 20, -10, -4, 13, 2, -15, 18, -3, -44, -7, 2, -1, 5, 30, 8, -51, -20, 5, -5, -34, 8, -16, 2, -16, -24, -8, -17, -3, 9, -3, 11, 8, 3, -26, 14, 7, -23, -2, -12, 25, -3, -5, -7, 3, -15, -5, -53, 22, 59, -9, 4, -3, 6, 10, 5, -33, -11, 21, 18, 5, 7, 26, -4, 6, 58, -18, -10, -2, -1, -3, 5, -48, -1, 8, -3, -8, 1, -6, 9, -44, -22, -39, 1, -3, -12, 8, -2, 17, -11, 47, -19, -29, 0, 16, 7, -32, 7, 6, 0, 6, -8, 9, 30, -29, 15, 1, 9, 2, 54, -17, 13, -23, 35, 7, -9, -13, -3, 2, 20, 38, -1, -14, 33, 1, 4, -12, 22, 16, -12, -5, -15, 13, -2, 11, 14, 6, -47, -18, -4, -62, -6, 11, -17, -49, -47, 23, -8, -35, 12, -32, 6, -11, -9, 0, 23, -2, 14, -5, -5, 8, -26, 23, 1, 1, -81, 1, -36, 32, 18, 1, -3, 53, -25, -3, 21, -58, 31, 6, 8, 4, -13, 46, -8, 35, -32, 3, 11, 9, 11, 44, 4, -6, 31, 3, -17, -32, 5, -4, 25, 0, 4, 3, -8, -15, 8, 5, 2, -28, -30, -42, 5, 2, -10, 8, 3, 50, -6, 17, 0, 10, -6, -7, 19, -40, 30, -5, 5, -2, 16, -13, 23, -12, 24, 4, 7, 3, 20, 8, 1, -38, -3, -15, -58, -63, 2, 4, 21, 1, 19, -1, 7, 11, 0, -14, 21, 20, 11, -22, 2, 11, -5, 46, 38, 10, -65, -41, -9, -68, -30, -20, -47, -8, -23, 23, 3, -79, 0, -23, 3, -16, -11, -4, -1, -5, 21, 3, -42, 0, -61, -8, 14, 6, -89, 5, -48, 17, 27, -3, -2, 5, -32, 34, 12, -55, 30, 11, 31, 21, -11, 3, 2, 19, -54, -5, 4, 22, 41,
    -- layer=2 filter=0 channel=7
    11, -4, -3, -13, 59, 24, 23, -23, 12, -9, 7, 2, -30, 9, -16, -6, -6, 17, -33, 6, -15, 8, 0, 23, -3, 4, 14, -1, -4, -32, -8, -4, 7, -27, 7, 3, 4, -19, -6, 33, 10, 3, 7, -6, -26, 2, -1, -5, -19, 6, 31, 21, 15, -6, 16, 2, 34, -30, -6, -40, 1, 1, -1, -12, -28, 15, -8, 13, 19, -1, -42, 5, 18, -37, -20, 15, -10, -1, -50, 27, 3, -21, 0, -18, -12, 0, 32, -4, 2, 0, -11, -18, -13, -1, 2, 20, 5, -15, -16, 1, -6, -3, -2, 15, 5, -23, -25, -10, 3, 6, 13, -29, 45, -24, 36, 13, -20, -30, -22, 14, 37, -10, -25, 10, 6, -34, -2, -23, 13, -3, 17, -2, 28, 32, 46, 16, 6, -34, -41, 1, -32, -1, -1, 2, 5, 20, -11, 8, -33, 4, 1, 32, -5, -5, 6, -6, -26, 3, -6, -2, -10, -17, 4, 12, 4, -4, -5, 16, -31, 7, -27, -31, -29, 3, -8, 19, 20, 5, 19, 23, -28, -1, 27, 0, 20, 5, -32, -44, -8, -17, 24, 2, 3, -7, 32, 2, 13, 0, -13, -4, -14, 20, 19, -4, -10, -1, -51, 37, -19, 4, -19, -5, -2, -6, -23, 3, 0, -4, 0, -18, -4, 2, 1, -13, -6, -23, -20, 21, 8, 7, 7, -94, 1, 20, -7, -5, 2, -4, -14, -5, 29, -66, 41, 16, -15, -37, 3, 16, 19, 1, -30, -5, 8, 11, -15, -41, 3, 8, -30, -18, 18, 32, 9, 13, -6, -4, -5, -2, -53, -17, -4, 6, -7, 19, 18, -12, 13, -5, -6, 56, -2, -6, 8, 0, 5, -19, -2, 6, -9, -18, 10, 12, 28, -6, -26, 5, -30, -1, -18, -12, -22, 4, 10, 22, -6, -30, 5, 5, -17, 24, -4, -10, -21, 28, -27, -20, 0, 31, 11, 30, 9, -7, 43, -13, -12, -6, 10, -1, -38, 63, 16, 10, -2, -2, -23, -31, 10, -1, -5, -20, -10, 29, 9, 0, -11, -2, 18, -17, -20, -23, -7, 10, 0, 1, -16, 20, -8, 28, -2, -66, 0, -27, -20, 42, 7, -5, -22, -8, 17, -18, 7, 24, 0, -29, 2, 2, 13, 5, 12, -9, 7, -29, 25, -30, -9, -4, -12, -7, 12, 11, -12, -27, -8, -3, -25, 2, 3, -10, -15, 0, 0, 13, -42, -2, -1, 0, -9, 32, -12, -2, -2, 2, -30, -30, 2, -6, -43, -15, 14, -3, 23, 0, -15, 7, -3, -13, -2, -52, -25, 0, -3, 25, -19, -10, 7, -6, -11, 55, -49, -5, -16, 25, -18, -9, -1, 18, 13, 25, 14, -3, 16, -6, 10, -37, 16, -6, -14, 26, 9, -33, -28, 5, -6, -10, -27, -36, 37, -19, -9, -11, 49, 4, 13, -4, 26, -30, -59, -6, -6, 58, -4, 11, -17, 1, -14, 8, 2, -76, 0, -25, -15, 34, 0, 0, 14, -14, -28, -37, 5, 10, -29, 10, 5, -4, 8, -1, -56, -42, 9, -13, 9, -13, 27, 8, -5, -14, 10, -37, 0, -4, -8, 7, -12, 6, -18, -13, -16, -2, -3, 18, -36, -5, 8, 4, -7, 0, -26, 5, -24, 6, 22, -50, -10, -5, 0, -31, 34, -17, 31, -17, -9, 16, -38, -16, -12, 20, -18, 2, 2, 14, 4, -10, -41, -12, -16, 17, -16, 4, -7, -32, -35, -34, -5, 23, 26, -1, 26, 8, 7, 30, 3, -15, 5, 1, -43, 13, -3, -9, -24, -4, 27, -14, -8, 7, 40, 18, -17, -19, 5, -6, -3, -4, 34, -16, -7, 11, 3, 24, 0, 9, -16, 29, -26, 6, 2, -68, -5, 0, -45, 23, 1, 0, 16, -13, 14, -20, 12, 30, -10, -9, -17, -11, 25, 2, 14, -12, 32, -10, -3, -25, 5, 3, 4, 1, 17, 5, 0, 25, 11, 7, -5, 4, -44, 6, -16, -2, 6, -17, -11, 16, -26, 1, 0, -6, -2, 5, 10, 0, 50, -18, -10, 6, 8, -20, 12, -3, 32, -15, 12, 16, 7, -13, -31, -35, -35, -4, 1, -19, 2, -18, 1, -33, 11, -27, 17, -6, 11, 21, -19, -24, 1, -18, 0, 1, 32, -5, 16, -18, 2, -12, -9, 8, -28, -41, 16, 10, -10, -8, 28, -6, -6, -15, -20, 5, 0, -5, 24, -12, 23, -3, 20, 14, -24, 31, -5, 12, 7, -32, -32, 34, -43, -2, -7, 0, -7, 56, -35, 31, 4, 0, 35, -12, 19, -49, -24, 33, -7, -54, 25, 7, 1, -3, 23, 18, 32, 20, -12, -47, 15, -3, 6, -3, 47, -27, 35, -7, 1, -12, 38, 0, -42, 6, -17, 1, 9, -16, -22, 14, -2, -1, 0, 15, 7, 5, 13, 2, 2, 7, 29, -4, 0, 17, -19, 20, -1, -12, 9, -25, -27, 16, -2, 1, -54, -12, 3, -67, -10, -18, 60, -40, 24, -13, 16, 0, 11, -10, -54, -15, 0, -60, -3, 14, -5, 10, 19, -25, -41, 17, -44, 0, 11, 0, -3, 31, -32, 0, 45, 17, 29, -19, -24, 14, -4, 15, -8, -1, 31, -1, 31, 4, -40, 26, 1, -25, -9, -33, -25, -8, -12, -5, 0, -55, -4, 15, 4, -8, 7, -6, 25, -34, 4, -52, 15, 19, -6, -49, -5, 4, 12, -3, -37, -31, 30, -62, -2, -5, -6, 1, -14, 27, -8, -20, 10, -6, -4, 24, -36, 1, 22, 3, 5, -6, -7, -48, -38, -13, 10, 1, -2, -15, 5, 1, 26, 13, 35, -34, -43, -1, -12, 10, -9, -13, 0, -18, -20, -3, -14, -18, 9, -19, -9, 3, 0, 3, -34, -18, 0, 12, 0, 40, 24, 1, -22, 21, 11, -14, -1, 17, 6, 4, -2, 16, 9, 26, 4, 10, -8, -1, 57, -108, -6, 0, 36, 1, -61, -15, -11, -23, 10, -14, -5, 24, -17, 15, -13, -4, 0, -7, -12, 7, -6, 9, 6, -33, -27, -3, -30, 1, -7, -20, 4, 14, -26, 11, 3, -4, 22, -10, 15, 5, -22, 8, 8, 1, 5, -48, -3, -5, 25, 13, 24, -31, -13, -14, -3, 6, 7, 32, 25, -19, 12, 22, -16, 3, 2, -9, -4, 20, -11, -3, 0, 48, 11, 17, -20, -4, 0, 1, 19, 4, 23, -5, -12, -42, -11, -4, 4, -11, 1, 12, 1, 0, 16, 23, -2, -6, 6, -27, -21, 5, 2, -4, -18, -18, 19, -13, -12, 15, 46, 5, 0, -21, -18, 0, -1, 23, 26, 8, 10, 18, 8, 7, 20, 9, 4, 3, -1, -3, -39, 5, -14, 5, -35, 0, -40, 17, 13, 23, -12, -38, -11, 0, 0, 4, -2, -24, 0, 30, 1, 7, -2, -51, -9, 0, -19, -11, 1, -3, 5, -1, 24, 4, 7, -3, 4, 24, 11, -21, 36, 12, 17, 35, -3, 1, 23, 8, 28, -23, -8, -6, -7, 8, 18, 5, 27, 3, -1, 7, 14, 27, 4, 0, -2, 7, 7, -6, -3, 8, 9, 0, 61, -25, -17, 0, 0, 22, 26, 4, 16, 3, -23, 4, -27, -5, -24, 6, 0, 12, -31, 3, -8, -25, -9, -19, 42, -8, -12, 5, 3, -6, 29, -20, 35, 6, 32, 16, -8, -1, 20, -37, -1, 29, -11, -21, 28, -24, -7, -16, 4, -7, -4, 9, -29, 7, -53, 52, 13, 33, -36, -3, 9, 12, -21, -11, -11, -11, -20, 9, -28, -1, -22, 1, 22, -13, -5, 11, 6, -38, -1, -29, -4, -9, -37, 9, 2, -56, 2, 12, 46, 14, -9, 0, 23, -14, 13, -44, 28, -10, 22, -31, 24, 14, 15, -1, 2, -23, -37, 8, -26, -29, -1, -2, 10, -25, -2, -14, -32, 48, 3, 4, -6, -3, 8, 9, 3, 4, 1, 34, 26, 0, 30, 0, 6, 11, 12, -1, 24, 3, 15, -34, -22, -6, -16, 11, 14, 4, 12, 35, -31, 0, 0, -3, 9, 16, -1, -2, -5, -16, 24, -46, -15, 27, 12, 16, -14, 3, -12, -54, 23, -7, -8, 12, 4, -46, -6, 1, -18, -23, -22, -34, 35, 4, -10, 34, -13, 19, -16, 2, -3, -6, 4, -44, 16, -28, -32, 14, 56, -2, -12, -5, 23, -33, -18, 9, 0, -25, -2, 26, -13, -24, -46, -4, 1, -70, -2, -43, 27, 0, 3, 2, 12, -25, -24, -25, 11, -19, 0, 16, -24, 17, 0, -1, -6, 1, 6, 16, -4, 3, -40, -1, 48, 42, 48, -71, -23, 42, 12, 0, -17, 3, -18, -57, -10, -6, 3, 10, -7, -12, -25, -7, 5, -3, -9, 2, 16, 0, 78, -7, -20, 0, -38, -2, -9, -27, 36, 32, -27, 36, -7, 13, -16, 17, -47, 0, 1, -23, -10, 8, -15, 21, 15, 0, -21, 4, 16, -28, 57, -12, -5, 8, 7, -13, -3, -30, -8, 8, -30, 6, 41, -2, 3, 3, -47, 3, -37, -10, 42, -1, -6, -24, -13, -12, -17, -62, 31, -20, 18, 6, 9, -25, -15, 10, 3, 10, 8, 7, -16, -24, -20, -25, 3, -4, -7, -7, 15, -33, 3, -6, -15, -9, -1, 36, -20, -40, -5, -11, -19, 3, 16, -6, 43, 4, 16, 26, -22, -1, -13, 6, 32, -3, 33, -20, -7, 53, 5, -20, 12, -1, -27, 34, -4, 2, 0, 7, 9, -14, -22, -4, -2, -5, -6, 8, 26, 7, -23, 16, -16, 7, -5, 18, 12, -9, 24, 56, 0, -5, -9, 8, -24, -14, -34, 4, 7, 8, 2, -15, 10, -15, -16, -1, 14, 8, 30, -16, -9, -10, -6, 8, 5, 29, -17, 4, 20, -3, -30, 13, -2, -5, -3, 9, 6, -2, -41, 3, -1, 4, -17, 14, -35, 9, -12, -23, -13, 0, 13, 4, 9, -12, -12, -9, 0, -46, 2, -3, -26, 21, -4, -14, 5, -27, 3, 8, 25, 18, 7, -6, -8, 17, 28, -22, -4, 0, 6, -13, 18, -2, -14, 0, 1, 21, -11, -17, -5, -7, -26, -3, -37, -19, -20, 46, 29, 8, 7, 15, -4, 1, 9, 5, -4, 5, 1, -11, 13, 33, 71, 4, -2, 19, -13, 2, 4, 5, -36, 17, 16, -4, 15, 15, 36, 9, -17, -2, -5, -8, -45, -43, 23, -5, -31, 1, 2, 38, -4, 2, 43, 0, -12, -45, -3, -6, 13, -24, -52, 12, -7, 9, -6, -29, -5, 0, 52, 34, 4, 12, -28, 3, -3, 38, 41, 47, -1, -10, -32, 52, 11, -10, 15, -44, 7, 7, 4, -8, -18, -7, 8, -20, -53, 6, 2, 14, -1, 0, -12, 8, -36, 40, 0, -2, 3, 28, -10, 41, -6, -1, 13, -35, -16, -20, 25, -4, 6, -14, 65, -7, -6, 6, -64, 58, -25, -15, 5, -6, -26, 7, -30, 52, -5, -4, 51, -9, -16, 52, -51, -2, 16, -27, -15, 1, -4, 8, -28, -32, -21, -5, -3, 11, -2, 1, -8, 8, 37, -34, -6, 4, 14, 9, 0, 9, 44, -36, -11, 27, -10, -47, -10, 24, -58, -3, 2, -9, -33, 58, -32, -5, -4, -35, 7, -6, -4, -23, 15, -30, -2, 17, 13, -58, -13, -14, 33, 58, 14, -4, 3, 0, 2, -87, -4, -22, 3, 0, -72, 50, -2, -21, 22, -34, 22, 12, 17, -14, -20, 4, -4, 5, -72, -30, -5, 8, -4, 10, -18, -19, -17, 23, 5, 2, -4, 42, -34, 10, -1, 3, 1, -20, -20, -21, 21, -25, 0, 18, 18, 16, -24, 0, 76, 28, 4, -1, -26, -9, -30, 0, 59, 58, -22, -28, 6, 29, 14, 0, 4, 0, 3, -12, -18, -1, -6, -3, -17, 29, -23, 3, -1, 6, 9, -5, 16, -1, 34, -29, 7, 0, 15, 3, 11, -4, 13, -18, -16, -1, -32, -1, -7, 0, -2, 3, 8, -3, -37, -15, -22, 5, 22, 2, 14, 0, -50, -8, 15, 0, 0, 13, 6, 18, -3, -29, -3, 33, 7, 15, -14, -1, -13, -50, -10, 5, -14, 2, -8, 29, 2, 34, 2, -38, 0, 3, 5, -1, -12, 5, 2, -10, -55, -8, -2, 2, -2, -22, -15, 13, -15, -17, -4, 30, -6, 8, 11, -8, 5, 0, 11, -3, -15, -1, -8, -14, -14, 10, -8, -7, 68, 0, 38, 17, -28, 11, -20, 1, -2, -5, -9, 29, 8, -20, -24, 6, 1, 21, -5, -8, 0, 5, 0, -6, -7, 45, -11, 36, 21, -5, 6, -28, -4, 1, 20, 1, -4, -19, -28, 0, 15, 24, 47, -40, 1, 40, -17, -7, 7, 5, 5, -17, 23, 0, 0, -32, -4, -58, 36, -9, -10, 22, -51, -7, 22, 29, -1, -8, -10, -13, 18, -22, 14, -11, -21, 15, 6, -26, 7, 4, -12, 15, 2, 2, -52, -10, -36, -14, 36, 16, 20, -31, -23, -33, 17, -3, -109, -6, 20, -37, -17, -5, 0, -41, 3, -7, -9, 9, 0, -28, -3, 52, -3, -10, 47, -63, 6, 0, 16, 1, 8, 2, 0, 0, -58, 20, 20, 18, 37, 3, 15, 9, 11, 38, -19, -9, 15, 7, -19, -22, -5, -4, -25, -30, 8, 3, -4, 1, 10, 27, -14, 0, -7, -2, -1, 16, 15, -2, 0, 13, 12, -4, 25, 6, 23, -27, -52, -1, -3, 20, 6, -55, -12, 61, -56, -24, -28, 64, 34, -32, 22, 1, -7, -3, -36, -94, 5, 5, 15, 16, -29, -2, 11, 26, 20, -57, -2, 2, 25, -5, 10, 16, -39, 20, 40, -30, 53, -6, 20, 30, 32, 4, -41, -2, -9, -14, 8, 7, 18, -47, -35, -16, 4, 5, -110, -2, 26, -76, 0, -24, -6, -14, -6, -27, -4, 27, -18, -40, -1, 15, 3, -34, 60, -114, -1, 1, -28, 14, 41, 14, 4, 46, -81, 52, -17, 16, -4, 0, -15, 5, 34, -4, -27, 13, -11, 0, 31, 62, -8, -26, -11, 22, 8, -9, -23, 7, 18, 2, -8, -5, 0, -22, -36, 10, 37, -3, -5, 5, 11, 6, 15, 3, 13, -27, -16, -2, -18, -3, -2, -43, 23, 60, -27, 14, -9, 54, 6, 11, 10, 2, 0, 2, 16, -31, 4, 11, 14, 10, -20, -9, 64, -6, 35, -34, -10, 29, -18, 8, -3, 26, -32, 29, 11, -4, 48, -1, -24, -2, 35, -45, -29, -9, -6, 13, 23, -40, 2, -64, -35, -21, 12, -6, -57, 1, 42, -31, -10, 12, 3, -23, 0, -2, -21, -10, -76, -9, -2, -17, 6, -38, 41, -95, 0, 2, 13, -6, 28, -14, -19, 26, -47, 7, -14, 16, 75, 5, 26, -27, -31, 63, -37, 23, -4, -2, 21, 8, 10, -15, 3, 12, -7, -4, 24, 8, 6, 47, -1, -3, -5, 1, 0, -20, 3, 3, 4, 44, -6, 2, 19, -9, -9, 14, -3, -8, -11, -2, -5, -24, -13, 54, -23, -48, -20, -8, 0, 44, -9, -2, 0, -19, -11, 25, 6, 10, 9, -21, -20, -2, 17, 9, 3, -9, -12, -13, 5, 1, -7, -47, -3, 16, 14, -10, -3, -5, 25, -11, -44, 24, -39, 2, -27, 3, -46, 12, 0, -29, -9, -56, 16, -5, -42, 1, 22, 18, -35, 23, 3, -3, 2, -40, -24, 16, 5, -15, 3, 10, -7, -10, 20, -12, 4, 4, -11, -32, 4, -26, -27, 0, -32, -5, 13, 14, 48, 1, -39, -43, -6, 15, -25, -6, -30, 0, 12, -32, 8, 72, 34, 16, -6, 9, -1, 8, 0, 16, 0, -6, -1, -3, 37, 5, 12, 3, 8, 36, -5, 1, -2, -3, -49, 10, 13, 0, 3, -16, 51, 25, -14, 21, 14, -37, -43, -48, -14, -3, -40, 7, -4, 21, 29, -50, 64, -1, -13, -19, -5, 5, -2, 7, -19, 12, -8, 3, -23, -15, -10, -26, 39, -45, -3, -13, -63, -9, -20, 49, 13, 4, 34, 5, 15, 21, 20, 33, -2, -1, -11, -12, 16, -7, -43, 2, 19, 3, -44, 0, 7, 4, -4, 4, -22, 23, -19, 40, 2, -16, 5, 30, -26, 34, -4, -6, -38, -21, 3, -34, 26, -23, -13, -19, 56, -26, 21, 5, -64, -12, 29, -13, 24, -2, -1, -3, 20, 21, 25, 12, 27, 26, -5, 18, -13, -9, -3, -33, 0, -2, 6, -45, -1, 1, -4, -3, 1, 21, -9, 2, 0, 5, -14, 23, 28, 0, 17, -4, 6, 26, 10, -33, 54, 22, -20, -38, -13, -7, -32, -7, -12, -14, -6, -20, 18, -1, -30, -5, 20, -2, 1, -33, -13, 10, -16, -17, 0, -23, 23, -6, 28, -21, 3, 41, 36, -4, 11, -60, 10, 5, 11, 8, -22, 18, -28, 0, 32, 33, 37, 7, 35, 4, -26, 1, -35, 4, -26, -1, -1, 16, 4, -33, -9, 40, 0, 20, 0, 19, 3, -10, -23, 13, 2, 5, 48, 29, -6, -15, 1, -14, 19, 0, 31, 39, 8, 4, 21, 45, 24, 23, 5, -11, 1, 1, 4, 51, -45, -52, 32, 29, 0, 5, -9, 7, 11, -17, -12, -6, 0, -45, -6, -21, 0, 2, 0, 39, -15, 5, -4, 6, 53, 2, 8, -3, 11, -2, 6, -45, 35, -13, -28, 38, -3, 4, 1, 25, 24, -5, 5, -14, -34, 8, -3, 14, 22, -1, -33, 1, 1, 18, 17, -22, 3, 12, -7, -38, 0, -45, 32, 21, -9, 1, 0, 1, 29, -65, -11, -36, -27, -4, -29, 13, 0, 14, -12, -58, 33, -7, -9, -16, -67, -5, 15, -32, -2, -77, -6, 37, 8, 6, -22, 25, 5, -6, -4, 3, -1, -22, -17, -5, -5, 7, -12, -22, -33, 2, 13, -18, -3, 16, -15, -34, -2, -5, 16, -32, -29, 33, -4, 14, -28, 0, 6, -12, 29, -6, 4, -4, -5, -8, 17, 1, 1, 38, -8, -4, 7, 15, -59, 3, 13, -4, -2, 2, 11, 1, 26, 2, -16, -2, -3, -6, -39, -11, 10, -42, 6, 22, -69, -4, -39, 47, 18, 4, -6, -4, -3, -1, -46, -27, -3, 27, 2, -47, 30, 5, 17, 17, -13, -3, 7, -19, 27, 7, -31, -9, -18, 30, 43, -20, -17, -1, 32, 0, -34, 16, -78, 0, 1, 61, -3, 45, 16, -71, -9, -42, 48, 3, -88, -1, 9, -49, 3, 19, -2, 10, 0, -1, -19, 9, 3, -14, 2, -8, 6, -13, 33, -75, -7, 0, -38, 17, 33, -10, 40, 20, -49, 3, 0, 35, 26, 0, -7, -26, -23, 68, -5, -5, 7, 4, 45, -18, -12, -2, 0, 60, -15, -19, -36, -12, 16, 58, -14, 0, 4, 5, -41, 37, 0, 1, -3, -5, 4, 0, 55, -10, 3, 0, -29, 5, -27, 0, -12, -52, -49, -15, -35, 12, -61, 83, -6, 30, 17, -13, 0, 26, -73, -75, 20, -52, 30, -8, 98, 3, 1, -24, -34, -36, -1, 22, 23, 10, -4, 32, -58, 19, 18, 7, 6, 3, 24, 29, 5, 40, -57, 0, -57, 50, -15, 78, 34, -69, -14, -86, 44, -11, -127, 6, 58, -46, -31, 23, 6, 13, 4, -47, -12, 34, -18, -18, -7, 10, 2, 4, 9, -82, -5, -6, -66, -9, 2, -10, 6, 49, -43, 11, -36, 33, -52, -8, -23, -20, -23, 72, -19, 8, 5, 4, 45, 8, 17, -27, -9, 22, 7, -22, 13, -5, 0, 4, -11, -9, -10, 18, -4, -1, -1, -7, -2, 17, 19, -6, -3, 7, 1, -6, -25, 4, -54, -22, -33, -42, 26, -6, -43, 31, 2, 55, -19, 12, -8, -14, 9, 0, -7, 16, 6, -37, 5, 10, 42, 2, 66, -25, -18, -17, -3, -11, -20, 13, 6, -21, -42, -2, 4, -15, -14, -5, 22, -43, -15, -26, -59, -2, -6, 39, 13, 3, 52, -47, -28, -48, 22, 4, -60, 0, -1, -59, -45, 8, 3, 11, -3, -20, -19, 25, -5, -57, 0, 54, -3, -58, 12, -45, 7, 1, -49, -41, 44, 12, 0, 16, -55, -13, -34, 3, 66, 8, -2, -31, -6, 35, 0, 4, 20, 3, -18, -14, 0, -12, -27, -1, -6, -13, -2, -11, -18, 30, -9, 6, 6, 17, 28, 1, 18, -4, -3, 19, 3, 5, 7, 9, 8, 4, 8, 8, -11, -4, 24, -23, -13, -26, -46, -16, -15, -11, 6, 12, -29, -9, -5, 29, 3, -22, 19, -23, 11, 25, -45, -4, -39, -19, -1, 3, -9, 3, 8, 38, 23, 2, -5, 15, 25, -15, 14, 7, 12, 7, 5, 39, -54, 5, 24, 23, -14, -3, 15, -1, -8, -38, 5, -22, -73, -6, 11, -45, -36, 51, 4, 11, 5, -33, -18, 16, 6, 1, -7, -47, -4, -53, 2, 0, 7, 3, 28, 15, 5, -33, -30, -36, -35, 20, -7, -30, 20, -9, -84, -63, -14, -69, 6, 8, -5, 1, 10, -44, -15, 25, 25, 34, -12, -5, -9, -1, 16, -8, -6, 6, 5, 17, 53, -16, -1, 0, 0, 9, 2, 7, 15, -1, -53, 6, 5, 3, 7, -16, 26, 21, -3, 39, 43, -19, 6, -46, 3, -1, -31, 6, 12, 8, 36, -9, 28, 15, 12, -49, -4, -1, -1, 12, -3, 11, -1, 14, -28, 0, -13, 1, -9, -10, -16, 8, -32, -1, 0, 21, -7, 8, 19, -7, 21, 13, 8, 11, 9, 51, 2, -3, 50, -7, -29, 3, -6, 39, 7, 5, 3, 44, -6, -31, -24, 17, 10, 13, -4, -29, 7, -18, -11, 11, 0, 0, -8, 14, -20, -12, -26, -12, -3, 10, 18, -8, 17, 0, -57, -61, -35, -25, 26, 20, -24, 5, 9, 5, -24, -44, 13, 18, -5, 10, 0, -5, -8, -35, -16, -6, 6, -77, -29, -49, -25, -2, 6, 37, -10, 8, 0, -5, 44, -6, 28, 4, 42, 33, 6, 3, -10, -33, 44, 30, 1, 31, -37, 15, 5, 5, 0, -41, 28, 19, 0, -7, 13, -3, 38, 3, 17, -33, 1, 9, -7, -14, -46, -24, 4, -25, 11, 30, -19, 56, 24, -3, 19, -89, 2, -4, 18, 1, 2, 32, -16, 25, 22, 1, 45, 18, 16, -3, 36, 4, -16, 67, 6, -20, -7, 4, 9, -33, -18, 48, 31, -1, 0, -8, -1, 33, 0, 6, -6, 2, 43, -13, -22, -7, 16, -15, 29, 2, -13, 2, 18, -3, -8, 11, -15, 87, 17, 13, 3, 7, 11, 32, -31, -17, -34, 22, -5, -17, -72, -7, -4, -22, -3, 2, 4, 23, -27, -35, 9, 1, 3, 31, 1, 6, -28, -1, 37, 16, 9, 4, -2, -18, -53, -20, 54, 53, -40, 4, -4, 2, -31, 37, -6, -1, 5, -46, -4, 10, 9, 14, 28, 31, 13, 4, 26, 45, 23, 0, -3, 5, -13, -12, 6, -36, 15, 8, -59, 8, 15, 3, 10, -78, -6, -55, -4, -3, -10, -20, 11, 29, 17, -61, 24, -2, 42, -3, -21, 5, -9, -12, -1, -54, 0, 14, -3, -18, -22, 12, 34, -10, -7, 14, 2, -66, -9, 21, -5, 2, 29, -21, -10, 23, -36, -18, 32, -8, -22, -43, 5, -1, 29, -12, -86, 13, 4, 36, -13, 9, 0, 23, -8, -20, -26, 19, -3, -25, -33, -10, -26, -22, -13, -5, 6, -19, -34, 5, -11, 0, 0, 39, -11, 4, -17, 3, 29, 10, 15, 1, 5, -14, -3, 1, 0, 2, -38, -2, -48, 0, -16, 20, -7, 3, 6, 0, 4, -49, -36, 3, 3, 15, 17, 0, 14, -18, -10, -4, -14, 20, 3, -24, -5, -50, -17, 16, -13, 16, -32, 5, 8, -40, -11, -30, -9, -8, -27, 17, -9, 27, 38, -23, 1, -13, 36, 7, -24, -6, 20, -30, 6, 26, -7, 8, -3, -28, -9, 14, 4, 17, 3, -2, 0, -42, -10, -17, 3, -4, 14, 53, 8, -23, 23, -5, 22, -16, -23, -47, -3, -1, -35, -43, 3, 99, 4, -3, -29, -4, 11, 7, 12, -11, 53, 32, 1, -26, -2, -6, -34, 17, 0, 3, 11, -26, 21, -7, -11, 7, -5, 63, -17, -2, -5, 4, -2, 18, -7, -1, -2, -27, 7, 19, 7, 8, -30, -4, -61, -31, -35, -13, -28, -3, 9, 22, -25, -20, 22, 18, -24, 25, 3, 0, 15, -25, -21, 2, 0, -6, 23, -25, 2, -68, -24, 66, -29, -10, 0, 5, -19, 1, 0, 7, 33, -7, 29, 101, -26, -6, 0, 0, 8, -10, 18, -4, -1, 4, -13, -5, -27, -3, -5, 20, 11, -31, -12, 12, -8, 22, 0, -33, 0, -3, -26, 27, 8, -5, -31, 12, -11, -4, 55, -26, 44, 2, -19, 26, 13, -1, -15, -11, -10, 51, 15, 2, -10, 4, 48, -6, 5, -39, 6, 32, -5, -25, 0, -1, -9, 11, -3, -6, -3, 7, 21, -17, -18, 4, 1, 58, 0, -2, -18, 6, -20, 37, -11, -1, -21, -49, 21, 0, -20, -27, -13, -11, -45, 13, -27, 6, -10, 3, 4, 3, -14, -17, 38, -23, -3, -33, 27, -4, 39, -12, -53, 8, -5, -30, -35, -4, 3, -13, -11, 28, 9, -20, 21, 0, -7, -20, 17, -3, 1, 4, 0, 30, -7, 0, 43, 19, 12, 0, 56, -10, 22, -8, -9, -9, 22, 10, 0, 18, 0, 15, -13, 36, 0, -2, -7, 20, 2, -39, -14, 16, 6, 1, -16, 24, 1, 14, -4, -14, 6, -5, -32, 16, -40, 6, -18, -32, -33, 34, 6, -2, 29, 3, 19, -30, -30, -10, -16, 30, -2, -11, -24, -1, 7, 14, -5, -2, -4, -7, 46, -13, -33, 1, 8, 36, 8, 8, -8, -1, -30, 33, 25, 1, -1, -14, 20, 4, -41, -20, -75, -76, -7, -7, 23, 37, -12, 0, -7, 2, -23, -50, 36, -18, 20, -1, 17, 5, -26, 10, 9, 12, 6, -18, -1, -1, -18, -29, -5, -25, 1, -28, -2, 2, -27, 27, 34, 15, -43, 2, -19, -5, 20, 19, 23, -43, -7, 9, 69, -21, -61, 6, 23, -16, 7, -23, 0, 24, -3, -50, -4, 12, -3, 27, -6, 25, -4, -44, -15, 5, 2, 2, 16, 21, -1, 16, -21, -6, -16, 4, -28, 14, 38, 3, -65, -7, 11, 30, 23, 11, 2, 5, 14, -46, -18, 3, 23, 12, -7, -2, -30, 5, -23, 36, -2, 7, 4, -2, 35, -37, 28, -1, -5, 35, 0, 5, -4, 5, -76, 19, 20, 0, 7, 14, 16, -1, -57, 4, 68, -58, -23, -6, -3, 23, -14, -4, 2, 0, 17, 25, 49, -4, -22, -17, 7, 4, 0, -12, -49, 31, 7, -11, -19, -16, -29, -4, 2, 1, 20, 9, -7, 5, 6, 35, 42, -1, 3, 1, 10, 22, 21, 32, -20, 56, -10, 9, 37, -6, -29, 1, -9, 37, -5, 18, 6, 38, 2, -15, -31, 10, 3, 6, 3, -11, -3, -11, 8, -24, -1, 3, 20, 0, 9, -7, -5, -26, 6, 20, 1, -4, 65, -7, -80, -45, -22, 10, 4, 7, -15, -1, 7, 5, -26, -23, 30, 32, -20, 23, 24, 0, 29, 9, -8, 3, 0, -36, -48, -21, 39, -3, -6, 38, -5, -3, 29, 0, 13, -3, -18, -7, 13, 47, -16, -23, -17, -15, 46, 34, 7, 49, -57, -4, 19, -1, -1, -28, 50, -16, 11, 0, 5, -75, 57, 1, 27, 31, 9, 13, -2, 9, 12, 1, -12, 9, 11, 47, 8, 39, 48, 4, 42, -69, -11, -45, 60, -1, -12, 63, 19, 30, 24, -14, 14, 13, 13, 7, 52, -3, -9, 68, 12, 22, 7, 6, 5, -9, -12, 25, 16, -3, 1, 47, 0, 21, 15, -14, -2, 9, 9, 12, -37, 8, 0, 17, 6, 17, 7, 53, 14, -3, 14, 9, -2, 31, -5, 41, 4, -2, 16, 28, -13, -16, 17, -3, 7, -47, -20, -5, 15, -28, -4, -2, -6, -33, -49, -41, -1, -2, -3, 20, 9, 3, -32, -1, -9, 14, 43, 5, 14, 0, -27, 12, 5, 0, 19, 38, -5, 21, -53, 31, 34, 10, -2, -30, 3, -7, -25, -10, -31, 2, -7, 1, -10, -11, 3, 17, -16, 0, 3, -26, -46, -25, 3, -13, -12, -17, -8, -6, 28, -72, 15, -88, 31, -4, -8, 10, -8, -19, -7, -19, 14, 27, 5, 0, 8, -7, 9, 68, 15, 6, -7, 3, 1, -41, -18, 34, 8, -12, -7, 34, -4, -19, -8, -1, -4, -1, 39, -30, -25, 24, -26, -22, -14, -15, -7, -1, 24, -6, 6, -4, -33, 3, -6, -4, 0, 6, -5, -19, -26, -42, -7, 28, -4, -30, -9, -9, 13, -49, 2, -4, 1, -32, -52, -10, -39, 3, 0, 36, 16, 9, -13, 2, 2, -4, 7, 0, 22, 0, -27, 2, 1, 44, -28, -17, -47, -1, -90, -1, -3, 2, -3, -17, 26, -70, -18, -27, -38, -2, 29, -5, 3, 38, -13, 17, -6, -18, -6, 14, -34, -52, -15, 2, -23, -11, 0, -5, 28, -11, -6, -60, -19, 3, -1, 3, 16, 6, 7, -3, 6, 38, 3, 1, 35, -5, 2, 14, 26, 51, -3, 3, -4, -38, -16, -3, 24, -2, -4, 10, 7, -9, -10, 19, 2, -5, 39, 6, -33, 15, -25, -6, 18, -39, -31, -37, 36, -6, -8, -25, 10, 38, 28, -1, 16, -3, 20, -18, 2, -2, 4, 27, -6, -17, 22, 0, 15, -36, -14, 6, 0, -23, 3, -37, -63, 2, 4, 16, -9, 3, -32, 7, -19, 39, 54, 3, 3, -21, -13, 9, 21, 0, 0, 6, -53, -37, -42, -13, 15, -9, 3, -17, 38, -23, 10, 7, 0, -24, -3, 3, 15, 29, 0, 27, -2, -19, -10, 24, -27, -8, 15, -6, -47, 25, -49, 8, 41, -8, 41, -6, 0, -1, 42, 16, 2, 15, 0, 0, 20, 26, 25, 2, -18, -3, -75, 31, 29, 16, -2, 32, -4, -19, -6, -26, 26, -2, -3, 61, 1, -8, -10, 37, -4, 0, 38, 5, -13, 24, -23, 7, 18, -46, 1, -24, 11, 0, -22, -26, -59, -10, 25, -27, 4, -5, 43, -48, -33, 10, 0, 25, 0, -18, 49, 3, -6, -28, -9, 2, -1, -55, 35, -6, -34, 1, -2, 65, 3, 8, -12, 10, -22, 12, 14, 4, 3, 5, 10, 9, -49, -10, -14, -27, -29, 16, -45, 6, 23, -3, 5, 5, 35, 21, -4, -12, -5, -27, -9, 1, 0, 23, -30, -1, 2, -38, -17, 17, -37, -41, 15, -2, -8, 15, -34, -4, 22, 11, 4, -9, -11, -3, 21, -36, 12, 41, 4, -45, 7, 37, 46, -2, -30, -6, -26, 24, 14, 38, 3, 46, 3, 52, -20, 4, 12, 15, 0, 6, 5, -16, 7, 35, -7, -6, 46, -6, -10, 8, 22, 13, 28, -31, -2, 4, -70, 8, -21, -28, 5, -14, 0, 0, 7, 8, 21, -83, -22, -31, 8, -18, -18, -2, -18, 0, -17, -14, -13, 5, 1, 8, -19, -18, -37, 4, -4, 65, 0, 6, -5, 7, -17, 14, 27, -4, -8, -24, 3, 9, 0, -4, -28, -23, -40, 16, 1, 6, 3, -3, -2, -31, -5, -57, 35, -26, -5, 0, -5, -5, 37, -13, -16, 7, -7, -33, 4, -25, -47, -33, 37, -26, -1, 0, 4, -6, -16, 8, -54, 40, -35, 1, 27, -23, 3, 5, -1, -49, -19, 2, 76, 1, 35, 0, -16, 25, 33, 18, 2, 34, 1, -7, -16, 9, 36, 21, 7, 4, -5, -46, -1, -2, 3, 5, 12, 5, -31, 1, -28, 17, -10, -24, -10, -11, -22, 6, -93, -5, 18, 7, -4, -7, -18, 6, 25, -58, -9, 8, 1, 7, -18, 12, 12, -4, 3, 10, -9, 2, -5, -26, -6, -23, -24, 1, 2, 37, -3, 4, 9, 4, -74, 34, 14, 7, 3, 18, 30, 2, -16, 4, 17, -3, -22, 33, -12, 10, -18, -3, 0, 18, -7, -15, 5, -19, -19, -38, 2, -4, 24, -17, -52, 9, -5, -7, -5, 8, -9, 5, -22, 12, 26, 26, 24, -5, 14, -11, -18, 15, 7, 1, 27, 20, 7, 38, -3, 29, -5, -26, 27, 0, -8, -1, -36, 31, -23, 2, -5, 21, 8, 12, -14, 15, 12, 8, 1, 7, -1, -24, -1, -20, -3, 2, 7, 16, 24, 7, 7, -18, -10, 15, -1, 0, 21, 7, -55, -35, -14, 26, -5, -5, -34, 7, -16, -28, 15, 12, 36, 11, -6, -12, 16, -6, 33, 50, -7, 7, -3, -44, -24, -8, 27, -3, 4, 23, -22, -5, 32, -5, -44, 6, -16, 5, 0, 33, 9, -23, -34, 45, 71, -28, 34, 11, -22, 11, 46, -11, 2, -4, 31, 33, 0, -44, -29, -29, 50, -7, 51, -6, -8, 2, -5, -54, -27, -15, -12, 14, -3, 8, 15, 27, 14, -3, 46, -42, -34, -48, 33, -8, -2, 34, 25, 54, -20, 24, 10, -39, 25, -12, -45, -6, -51, 63, 14, -35, 0, 20, 6, -63, -22, 71, 3, -22, 0, 3, 3, 2, 34, 2, 3, 7, 6, 16, 6, -27, 22, 5, 5, 1, 11, 42, 20, -3, -42, 6, -29, 2, -10, 31, -23, -1, -50, 9, -19, -11, 14, -2, -18, 6, 9, 2, -3, -28, 0, 1, -5, -52, -22, -23, 0, 8, -2, 32, -13, -1, -14, 4, -43, -27, 0, 3, -1, -5, -12, -22, -8, 49, 11, 18, -12, -14, -70, -4, 38, -4, 7, -33, 0, -4, -27, -49, -45, 13, -18, 5, -55, 12, -1, 16, -2, -4, -54, -27, -48, 0, 24, 12, -17, 12, 8, 5, 10, -39, 26, -101, 8, -11, 23, 19, 0, -1, -16, 8, -3, -37, 28, 0, -32, 1, -5, 23, 2, -62, -1, 46, -5, -24, -27, 10, 12, -23, -1, -66, 0, 3, 15, -17, 7, -4, -19, -12, 5, 5, -9, -36, 14, -5, 3, 9, 14, 2, -21, -13, -24, 50, 8, 28, -12, -5, -17, -4, -43, -19, 16, 39, -6, 15, 48, 0, 18, -35, -11, -4, 0, 7, -12, -29, -10, 7, 4, 23, -8, -4, -2, -1, -29, -8, -26, -6, 2, -12, -38, -13, -9, 16, 8, 66, -14, -31, -66, 4, 21, -6, 4, -4, -23, 9, 7, -21, -14, -2, 14, -5, -41, -42, -18, 11, -8, -10, -19, -53, -54, -29, 13, 17, -49, -5, -15, 8, -41, -16, 17, -69, -24, -10, 22, 16, 8, -3, 0, -27, 2, -33, 39, 7, -80, 1, 20, 16, 9, -33, -5, 9, -3, 0, -22, 40, 18, -10, 5, 10, 5, 27, 3, 7, 1, 5, 41, -17, -31, 3, -22, -33, 1, -12, 16, -41, -2, 4, 3, -20, -15, -17, 4, 11, -19, 2, -3, -21, 13, -2, -12, 16, 0, 8, -10, -6, 1, -40, -9, 2, 6, -8, -5, -30, -78, 0, -5, 38, -2, -1, -14, 3, 8, -8, 20, 4, 13, -26, -47, 5, -5, 8, -5, -15, -35, -16, -44, 27, 9, 6, 6, -4, -20, 34, 23, 4, 8, 32, 14, -4, 2, 19, 3, 21, -1, -22, -14, -44, -59, -15, 16, -22, -34, 23, 7, 7, -34, 0, 1, -32, -17, -9, 42, 4, 7, -5, 29, -21, -5, -44, 15, 3, -63, -6, -25, -27, 13, -30, -5, 39, 0, -56, -17, 11, 35, 5, 1, 21, 0, 16, 0, 1, 0, 4, 28, -33, -8, 15, -30, -21, 14, 2, 29, -37, -33, -5, -3, -13, -35, 11, 22, 24, 3, -3, 20, -40, -2, -18, 55, 20, -12, -9, 16, 1, -6, 6, -12, 6, 8, 3, 7, 11, -43, 4, -4, 14, -11, -5, 34, -2, -33, 27, 10, -6, -1, 2, -2, -17, 3, 9, 26, -16, -55, -1, -37, -16, -7, -8, 1, 6, 7, 42, 40, -18, -5, -19, 22, -3, 4, 9, -16, 27, -8, -27, 23, 8, -35, -2, 39, -25, -23, -3, -4, 7, -7, -16, -2, 7, -11, 0, 0, 15, 11, 30, 22, 4, 4, -21, 26, -4, -24, -3, -53, 11, 8, 8, -5, 42, -3, -16, -11, 9, 3, 1, 2, 27, 1, 1, 19, 17, 6, 0, 14, 0, -32, 16, 8, 30, 5, -29, 22, -5, -19, -1, -28, -14, -6, -25, -5, 2, -4, -2, 21, -59, 13, 21, 20, 16, -17, -11, 17, -6, -4, -19, -6, -3, -4, -52, 13, -6, -27, 0, 5, 19, -35, -2, -15, -4, -82, 19, 0, 1, -12, 0, 16, -5, -36, -48, 7, 0, -57, -4, -5, -34, -2, -5, -2, -8, 13, -16, 0, -57, -36, 27, -8, -4, -1, -30, -39, 15, -2, -19, -7, -51, -58, 12, 27, -46, 0, 14, -6, 2, -16, -28, -3, -7, -49, -3, 77, -12, -2, 26, 6, -17, -9, -12, 49, 0, -61, -2, 12, -12, 1, -45, 0, 31, -6, -11, -17, 31, -26, 12, -5, 38, 4, 19, -13, 2, 5, 5, 23, 1, -14, 9, -21, -5, -3, -20, 2, 17, -72, 7, -72, -43, -48, 16, -1, -15, -28, -3, 4, -50, 14, 26, 33, -2, -1, -5, -24, 1, -13, 12, -7, 7, -4, 5, 16, -15, -4, -3, -3, 12, -13, 9, -22, -4, -73, 34, 0, -3, 6, 6, 33, -2, -18, -26, 6, -13, -28, 16, -17, -10, -6, 1, -2, 30, 1, 12, 33, -7, -12, -67, 42, 5, 18, -23, -35, 3, 7, 8, -1, 5, -26, 10, 10, -14, -7, 41, -2, 7, 18, -26, -27, 19, 44, -5, -12, 38, 15, 38, 18, 15, 13, -72, 37, -14, -18, 3, -15, 13, -4, -57, 0, 22, 6, -22, -19, 38, 6, 18, 0, 22, 1, 20, 14, -6, 0, 0, 9, 7, -17, 29, 44, -11, 0, -2, 21, 0, -11, 6, -36, -24, -49, 22, 1, 11,
    -- layer=2 filter=0 channel=8
    -11, 0, 10, -49, 9, -27, 28, -4, -29, 47, 1, -6, -29, 5, 2, 4, 5, -14, -26, 27, -20, 0, 1, -45, 12, 0, -30, -1, -9, 16, 39, 3, -11, -6, 22, -23, -72, -55, -3, 33, -6, 22, -18, -8, -4, 3, 0, 24, 13, -6, 17, -73, -26, -66, 20, 0, 21, 16, -60, -20, 1, -6, 11, 4, -1, 16, 4, 28, 18, -14, -42, 5, 19, -15, 13, -3, -32, 4, -17, 7, -13, 15, -53, 9, -42, 7, -21, 13, 13, -3, 10, 17, -9, 31, -4, -16, 3, -10, 1, 7, -26, -15, 0, -4, -6, 20, 4, -11, 4, 3, -14, -8, 19, -36, 27, 23, -55, -8, -20, 0, -10, 4, -5, 8, 24, 29, 16, 8, 17, -5, 1, 36, 17, -26, 9, 9, -14, -5, 39, -6, 15, -18, 2, -5, 8, 2, -2, 1, -110, -6, 1, -12, 11, 6, -19, 3, -63, 19, 8, -5, -12, -11, 33, -20, 2, -47, -3, 34, 2, 11, -1, -5, 8, 2, 1, 13, 31, 22, 48, -31, -30, 11, 13, -3, 0, -8, -17, -5, -16, -35, 5, 4, 19, 7, -2, 42, 8, -26, 31, -7, 20, -31, 15, -5, -19, 4, 31, 5, 13, 38, 36, 8, -34, 11, 7, 7, 3, 0, 6, 7, -2, 32, 0, 0, -10, 2, -2, 7, 16, -8, -6, 47, 4, 7, -3, -6, 6, 5, 1, -6, 22, 8, 15, 25, -35, 9, -40, 32, -24, 0, -39, -8, 1, 37, 16, 20, 10, -1, 2, 12, -4, -15, 0, -9, -6, -45, 1, -5, 20, -20, 5, 0, 3, -21, 7, -27, -37, -9, -3, 7, 20, -5, -42, -6, -47, 31, 14, 0, 0, -33, -8, -23, -53, -26, -11, 11, -17, 16, -6, -12, 4, 2, -4, -7, -1, -57, 7, -39, -11, -7, 6, 1, -23, -28, -52, -4, -18, 3, 12, 3, -12, 21, -39, 3, -14, -22, -3, 1, 9, -33, -3, -2, -12, -1, -8, -29, 11, 12, 4, 23, -31, 10, 10, 0, 4, 1, 15, -20, 13, 19, 0, 21, -3, -3, 3, -1, -6, -35, 5, -96, 6, -5, -9, -12, -7, 2, 3, 3, 15, 8, 11, 12, -14, -14, -18, 23, -33, 2, -24, -10, -1, -19, 4, -11, 0, 0, 3, 4, -30, -16, 9, 3, 0, -7, -40, -3, 15, -22, 5, -1, 0, 14, -17, -27, -35, -7, -7, 15, 20, -2, -50, -2, -24, -9, 24, 4, 11, -13, -15, -26, -10, 10, -26, -22, 2, 4, -28, -54, 5, 1, -6, -11, 3, 18, 13, -25, -42, -2, -22, -4, 2, 17, -27, -14, -8, -33, -2, -9, -16, -10, -30, 23, -10, -16, -28, 0, -11, -3, 3, -37, -3, -7, -30, 14, -10, -5, -10, 0, -31, -19, 26, 0, -23, 6, 11, -14, 10, -4, 7, 12, 0, -7, 8, -8, 27, -18, 2, 9, 3, -2, -9, -9, -2, 0, 0, 0, 8, 17, -3, -4, -25, -23, 3, -17, -20, -5, 0, -23, 14, 10, 11, 4, 5, -6, -5, -12, -25, -37, 16, -1, -3, -32, -11, -1, 27, -19, -1, 6, 6, 0, 2, -6, -31, -7, 1, 3, 12, 5, -18, -4, 5, 13, -9, -7, -8, -2, -34, -36, 0, -38, -24, 6, 11, 17, -51, -11, 2, -7, -3, -10, -22, 22, -24, -42, -26, -17, -10, -6, 3, 24, -20, 2, 0, -30, 2, 0, 17, -9, -38, 26, 0, 10, 28, -3, -2, -17, 7, -5, 13, 2, -53, 13, -2, 25, 0, 12, -14, -36, -1, 11, -9, 6, -2, -12, -2, 9, -1, 37, 4, -6, 2, 18, 39, -39, 4, -73, -2, 6, -10, -4, -2, -1, -11, 6, 25, 26, -5, 12, -4, 9, -39, 3, -18, 2, -40, -20, 7, 32, -3, 13, -1, -8, 3, -55, -34, -18, 23, -6, -2, 28, -5, 3, 42, -24, -6, -5, 0, 2, -24, 14, -19, 1, -2, 9, 22, 0, 4, 2, 23, 4, 2, 4, 3, 25, 0, -23, -6, 6, 2, 15, 4, 36, -65, -46, 12, 1, 5, 11, -12, 43, -42, -54, -54, -4, 26, 1, 9, -7, -49, 1, -5, -21, 3, 18, 7, 0, -8, 57, -2, 12, 0, -7, 34, -25, -1, -29, 2, 4, -30, 16, 23, 39, 19, 9, -21, -12, -4, -1, -10, 1, 11, -1, 6, -10, -3, 33, 2, 7, -8, 7, 21, -39, 7, -42, -2, 3, 0, -5, 0, -2, -19, 14, -7, 10, 29, 11, -6, 25, -11, 22, 0, 0, 36, -5, 25, -11, 31, 6, 10, -1, 2, -37, -21, -7, 3, 7, -2, 42, 5, -6, 27, 8, -1, 2, 3, 15, -5, 26, -90, -2, 1, -35, 0, -7, 12, 7, 23, 19, 36, 3, 7, 18, 47, -36, -38, 13, 8, -6, -22, 35, -20, -41, 9, -2, 1, 14, -11, 14, -3, -24, -34, 66, 27, -3, -2, 2, -37, 27, -12, -41, 12, 13, 24, 20, -33, 39, 27, 4, -6, 0, 27, -74, 19, -20, -1, -2, 23, 23, 14, 46, -8, -1, -24, -14, -6, 5, 17, -3, -8, 1, -2, 6, -6, -8, 1, -1, -2, 22, -3, -41, 0, 36, 0, 24, -2, -22, 6, 5, -7, 3, 15, 6, 32, 20, -32, -5, 8, 24, -3, 7, 17, 25, 2, 13, 0, -8, -2, 1, 7, 8, -16, 2, -9, 15, -14, 0, 54, -5, 19, -18, -3, -1, 4, -1, 14, -21, 2, -7, -5, 15, 31, 0, -29, 4, -9, 23, 26, -1, 17, -4, 0, 5, -48, 0, -6, -36, 18, 23, -15, 18, 6, 6, 0, -15, -4, 34, -7, -13, -32, -22, 7, -8, 13, -12, -36, -7, -7, -2, 6, 16, -5, -7, -33, 20, 33, -33, 0, -6, 22, 31, -7, 30, -43, 1, -28, -8, 51, 46, -37, -10, -1, -9, -64, 2, 6, 3, 12, -4, 12, 6, -2, -23, -8, -9, 6, 44, 0, -2, 0, -10, -1, -25, -8, -8, -5, 0, -17, 14, 11, -10, 60, 8, -19, 11, -63, 11, 4, 2, 25, -16, 6, 3, 34, 18, 0, -4, 11, 5, 0, -6, -4, 23, -4, 64, -14, 0, 10, -20, -3, 3, 2, -21, 3, -16, 0, 1, -8, 8, 33, -4, -21, 0, 4, 22, 7, -5, 6, 11, 14, 6, -31, 2, -7, -3, -3, 17, -16, 11, 2, 2, -4, -14, 3, 9, -6, 6, -27, 17, 18, 0, 17, 38, -15, 1, -10, -11, 10, 21, -9, 16, 27, 14, -5, 0, -5, -6, 31, -34, 19, -1, 4, -1, -34, 10, -6, 29, -46, 3, 14, -9, 13, 14, -20, -3, 14, 15, 16, 27, -5, 23, 5, -2, 14, 46, 62, -13, 0, -73, 3, 0, -4, 19, -3, 6, -4, 25, 20, 12, 0, 12, 5, -15, -10, 16, 10, -4, 1, -8, -1, -12, 29, -8, -6, -4, 0, -10, -40, -19, 12, -6, -16, 4, -22, -8, -9, -13, -3, 6, -1, 37, 23, -25, -80, -3, 4, 16, 17, -2, 0, 0, -3, 9, 12, 1, -13, -11, -5, 3, -36, 1, 2, -12, -42, 10, -51, -40, 18, -7, 8, -18, 13, 5, 32, -16, -27, -16, -10, -9, 15, 14, -36, 13, -16, 28, 18, 2, 11, -12, 0, 11, -42, 6, -15, 0, -67, 9, -10, -15, 22, -9, -85, 9, -15, -16, 19, 7, -13, 0, -13, 15, 5, 7, 10, -12, 9, -2, 0, 47, 3, -6, -9, 38, 22, -2, 5, -17, 6, 16, -12, 2, -7, -4, -22, 19, -16, 38, 2, 9, -6, 6, -20, -47, -10, 0, -34, 1, -9, -20, -45, -54, 3, -6, -20, -14, -5, -3, 34, 2, -14, -27, -23, 0, 6, -67, -1, 5, 3, -4, 11, -34, -11, 2, -9, 15, 2, 3, 15, -3, 23, -19, 3, 1, -4, -11, 24, -7, -27, -19, -10, -26, -9, 11, -14, -48, 19, 3, 3, 6, 33, -16, 34, -27, -9, 20, -38, 1, 0, -4, -51, 22, -5, 6, -1, -12, -9, -16, 8, 18, -36, -18, -67, 0, -10, -8, -4, -9, 29, -6, 1, 41, 9, -16, -40, -27, 9, 4, -2, 2, 2, 6, -4, 0, 23, 8, 1, 16, -4, -14, -1, -14, 50, 18, 4, -44, 1, 5, 5, 20, 4, 3, -18, -14, 0, 28, -23, -1, -12, 18, 3, -16, -19, 2, -37, 1, -19, -42, 0, -33, 7, -4, 9, -29, -44, -1, 11, 33, -8, -9, 16, 0, 21, -45, -6, 0, -2, 21, -14, -37, 16, -3, -2, 24, 8, 4, -6, -6, -47, 20, 23, -3, 9, 1, 12, 0, -53, 0, -14, -12, -50, 4, -19, -20, 23, 3, 0, 10, 12, -15, 3, -10, -21, -26, -10, 0, -11, 42, -25, 1, 1, -6, 10, 0, -18, -9, 25, 19, -20, -14, -55, -5, -13, -25, 0, 3, 43, -1, -42, 43, -6, 5, 6, -3, 18, -2, -12, -7, -10, 4, -11, -18, 33, 3, -7, 39, 4, -5, 2, 12, 43, 24, 7, -39, -4, 1, 18, 23, 4, -5, -4, 6, -7, 33, 2, 10, 16, 29, 17, -21, -1, 0, -16, -12, -28, -108, -18, -23, -9, -4, 2, -22, 2, -7, 14, 32, -13, 19, -39, 0, 26, -63, 1, 0, 6, 36, -44, 5, -4, 2, -5, -6, 13, -3, -7, 2, -12, -9, -1, -3, -12, 26, -22, -9, -31, -43, 17, 33, 14, 19, -74, -33, 2, 2, 4, 25, -10, -29, 12, -54, -86, 31, 26, 6, -26, -15, -55, 16, -7, 1, -1, 10, 7, -23, 8, 44, -25, -13, -9, 1, -29, -14, -2, -34, 23, 3, -34, 21, -7, -1, 46, 14, 12, 10, -7, 5, 33, 6, 13, 7, 4, -1, -6, 36, 0, 6, -9, 25, 13, 10, 7, -64, 5, 19, 0, 10, 3, -1, -4, 26, -3, 25, -26, 9, -4, 38, 16, -11, -8, 0, -25, 25, 2, -7, -2, -45, -2, 1, 6, 13, -8, -11, 22, 19, -18, 1, 26, 1, -12, -64, -1, -6, 9, 34, 13, 16, 15, 2, 0, -18, 13, -4, -32, -2, 19, 32, 21, 7, -7, -16, 9, -19, 4, -59, 10, 18, -4, 15, -27, -18, 0, 1, 6, -33, -4, 8, -3, -42, -34, 32, 25, -6, -22, -6, -14, 16, -1, -52, 0, 18, 33, 23, -9, 12, -2, -16, -5, -6, -59, -25, 1, 12, 13, -8, 20, 16, 34, 31, 4, 36, -39, -10, -16, 8, 14, 0, -8, -1, 18, 11, 4, -4, 0, 0, 0, 53, -6, -18, 2, -8, 1, 18, 7, 6, 3, 5, -12, 31, 14, 12, 5, 10, -8, -4, -8, -29, 1, -3, -21, 54, 23, -52, 9, -11, 4, -1, 13, 13, -25, -35, -18, 3, -15, -12, -8, -5, -8, -34, 5, 1, 6, -4, 26, -20, -28, -1, -7, -13, 26, 0, -4, 0, -2, 0, -2, -2, -6, 0, 51, -16, -60, 24, 19, 21, -2, 11, -35, -35, 4, 6, -8, -2, -5, 36, -15, -4, -37, 27, 0, -7, -12, 20, -30, -15, -3, -46, 2, 23, 9, 11, -35, 8, -17, -23, -14, 6, -6, 27, 2, 23, -17, 0, -11, 30, 14, 26, -8, 20, -2, -11, -30, 3, -5, 6, -14, -11, 17, 7, -3, -15, -6, 27, 10, 3, -12, -11, -7, -35, -4, -31, 0, -3, 1, 5, -13, 3, 2, -22, 37, 23, -31, -4, -26, 0, 49, 1, 0, -12, 27, -94, 48, -31, -1, -9, -5, 50, -10, 8, 3, -5, -15, 10, 26, -2, 16, -34, -3, 6, 1, 1, 12, -33, -16, 0, 4, -28, -1, 1, -18, 0, -32, -4, -17, -7, 40, 24, -18, 21, -89, -21, 17, 4, 14, 15, -47, -24, 1, -3, 1, -14, 11, 0, -2, -66, -48, -7, 4, 5, -11, -8, -59, -2, -5, -7, -5, 20, -13, -7, 29, 16, -31, -10, -18, -5, -13, 8, 9, 6, 3, -6, -50, 28, -2, 2, 11, -4, 37, -14, -35, -3, -29, -4, -8, -16, 24, -7, -4, 27, -7, 30, 2, -12, 56, 2, -5, -22, 0, -23, -7, 22, 5, -3, 18, 15, -16, 20, 12, 9, -24, -11, 31, -16, 9, -2, 8, -23, 12, -16, 46, -16, -10, -4, 16, 7, -2, -5, 23, 8, -22, 16, 42, -6, 10, -24, -1, 3, 4, 6, 9, -48, -92, 3, 0, 10, -2, 5, -11, -3, 17, -14, -18, 0, -48, -8, -8, 5, -55, 30, -3, -19, 1, -15, -13, 4, 2, 9, -2, -4, -28, 26, 15, -3, -31, 7, -15, 0, 0, -6, -10, -23, -4, 20, -4, 15, -20, -3, 15, 31, -23, -50, -9, 5, 2, -24, 4, -6, 12, -6, 13, 26, -21, 23, 7, -24, -26, -2, -32, 4, -6, -4, -9, 4, -3, -22, 1, 37, -5, 6, -3, 23, 42, 16, 1, -9, 0, 5, -4, 3, 2, 3, -21, 10, -49, -10, 29, -1, -80, -22, 12, -10, -5, -1, 26, -6, 5, -54, 3, 0, -23, 0, -23, 11, -4, -2, 35, -19, -5, 30, 29, -5, -12, 17, 2, -2, 6, 8, 55, -34, -54, 6, -8, 15, -17, -7, 19, -5, -24, -33, -63, -6, 13, 2, 2, -9, -45, 37, -16, -38, 6, -12, -30, -18, 17, 0, 0, -14, 0, 49, -2, -27, -11, -1, -13, 4, 5, 37, -14, -22, -1, 18, 15, -3, -38, -4, 10, 37, -20, -1, -38, -1, -48, -32, -12, -49, 37, -4, 11, 53, -32, 14, 28, -34, -19, -3, 1, -11, -14, 2, 1, 8, 16, -30, -7, 35, 1, -5, -9, 28, 23, 51, -5, 2, 1, 14, -3, 18, 5, 1, -34, 12, -25, 35, 9, 0, -76, -20, 5, -13, -33, 7, 2, -60, 16, 3, -24, -32, 1, -7, 12, -68, -13, 14, 4, 14, -17, 1, -17, -5, 16, -30, 4, -1, 6, 19, 4, 27, 24, 4, -6, 57, -2, 0, 3, 9, 8, 12, 27, 0, -54, -8, 34, 0, 8, 16, -6, -36, -63, -4, -37, -32, 28, -1, 1, -30, -12, -26, 10, -6, 2, 9, 13, -8, -32, 66, -22, 21, -10, 17, 5, 35, -16, 5, 24, 9, -17, -46, -25, -3, -42, -11, 3, 9, 35, -3, -34, 33, -13, -1, 2, -20, 0, 6, 5, 8, 11, -2, -35, -8, 4, -15, 3, 21, 4, -23, 9, 33, 28, 25, -8, -39, -7, 34, 0, -5, 3, 0, 4, 21, -6, 61, -25, 20, -32, 35, 22, -11, -32, -5, -13, -9, -38, -30, -34, -5, -2, 1, -2, -21, 26, -5, -2, 21, -5, 57, 32, -6, -11, -55, 4, -1, 0, -7, -38, 10, 9, -8, -3, -23, -12, 3, 10, 1, -52, -11, -20, 2, -53, -20, 38, -11, -15, -21, -7, 4, -57, 5, -44, -69, 11, -3, -2, -26, 5, -64, -14, -39, -66, -6, 24, -5, 18, 49, -36, 32, -13, -7, 0, 19, 3, 14, -14, -27, -1, -29, -28, -5, -26, -23, 13, 23, 22, -11, -13, -13, 15, 7, -14, 25, -36, 17, -50, 9, -20, 5, 3, -11, 12, -3, 1, 32, -7, -10, -10, 45, 0, 20, 5, -27, 2, -14, 16, 0, 3, 4, 7, 37, 18, 21, 5, 16, -9, 2, 3, 0, -13, 3, -11, 22, -21, -67, -18, -16, 8, 0, 8, 30, 10, -16, 15, 14, 6, 0, 21, 4, 13, -57, 7, 6, -2, -15, -13, 8, -33, -3, 2, -24, 2, 5, -79, 4, -15, 5, 8, 0, -8, -25, 28, 0, -50, -85, 12, 6, -13, 9, -36, 25, 8, -6, 4, -20, -23, -26, 5, -37, -22, 1, 41, -3, 15, -42, -45, -22, -9, -25, 16, 6, -15, 36, -13, 4, -4, 18, -22, -1, -59, -50, 35, 0, -38, -9, 27, 22, -73, 18, -4, 47, -20, -4, 0, 1, -4, -5, 39, -5, -27, 24, 0, -5, 3, 5, 6, 20, -11, -36, -4, -33, -4, 11, -26, 8, -3, 6, 8, 52, 15, 15, 31, 15, -11, -17, -22, -4, 45, -1, -7, 9, -2, 0, -21, -55, -3, -6, 6, 33, 14, -6, -22, -24, 0, -8, 33, 1, -13, -25, -1, -1, -2, -4, -18, 18, 1, 2, -2, -10, -3, -1, -11, 0, -19, -8, -33, 0, -25, -34, 11, -7, -29, 35, 12, 43, 53, 33, 7, 7, 4, 0, -6, 0, 9, 12, 7, -2, -4, -25, -2, 0, -6, -78, 4, -24, -14, 20, 16, -24, 1, -15, -12, 7, -44, -47, 6, 5, 3, 45, 0, 21, 16, 4, -53, 16, -32, -18, -2, 15, -34, 0, -62, -13, 28, -4, 16, 5, 12, 1, -3, 10, -8, -9, 11, 18, 15, 1, -6, -20, -1, 4, -2, -30, 6, 7, -21, -5, 23, -9, -9, 11, -38, -30, -12, -17, 29, 5, -12, -9, 11, 15, -12, -5, 1, -9, 12, -24, 18, 4, 5, -29, -7, 14, -21, 3, 17, -10, 11, -4, -6, 18, -12, 13, -5, 0, 2, 12, 10, -1, 23, 7, -17, -15, 46, 4, -8, -17, 42, -14, -19, 26, 5, 24, 2, 24, -13, 31, -11, -4, -9, 7, 23, 41, 23, 5, -37, -65, -7, -4, -10, -21, -16, -14, -7, -6, -11, -3, -19, -13, 33, -5, 2, 9, -9, -7, -5, 45, -14, 0, -1, 0, -32, 22, -34, -21, 0, 43, 2, 9, -16, -12, 0, -2, -22, 3, 0, -2, 6, 27, -7, -29, 8, -18, 26, 9, 0, -8, 2, -11, 0, 0, 3, -7, -7, 8, 1, 4, 12, -11, -32, 9, 13, -34, 29, 0, -37, 9, 28, 26, 23, -10, -8, 1, 0, -16, -17, 25, 6, 22, -8, -7, 34, -4, 28, -24, 13, 7, -1, -1, -13, -1, 0, -4, -4, -13, 6, -8, 7, 3, -20, -20, 22, -2, 0, 0, -1, 0, -56, 32, 6, -7, -26, -14, -66, 7, 15, 8, -7, 23, 8, 53, -21, -23, -46, 30, 22, 0, 2, -9, -29, 28, -8, -5, -2, -31, -2, -42, 16, -3, -5, -13, 1, -1, 8, 7, -33, -34, 31, 4, -25, 21, 22, -13, 31, 19, -10, -11, -16, -3, -18, 0, -1, -2, -1, -17, -4, 7, 3, -31, 0, 33, 34, 14, 0, -42, 3, 5, 14, 1, 2, 0, 11, 13, -11, 37, -30, 4, -53, 11, 13, -35, -53, 3, -24, 28, 21, 2, -5, -16, 11, 5, -9, -15, 25, 32, 30, 14, 2, 14, -6, 0, 10, -24, 15, -5, 0, 7, -68, 4, -48, 1, 5, 11, 13, 1, 13, 0, -66, -20, -30, -6, 7, 6, 16, 12, -1, 45, 35, 10, -23, -17, -81, -62, -16, -4, -8, 0, 5, 52, -26, 0, -69, -15, -4, -1, 33, -1, -2, -28, -11, 3, 9, -75, -20, -56, 11, -11, -8, -16, -12, 2, -2, -53, -12, -27, 33, 1, -29, 44, -16, -22, -28, 32, -29, -11, -32, -20, 6, 5, -26, 44, -10, -7, 4, 62, 0, -30, -3, 13, 21, 12, 0, 42, 1, 40, 8, -16, -7, 0, 12, -55, -17, 63, -65, -13, -40, 1, 30, -10, -44, 0, -20, 30, -32, -34, -14, -12, -3, -4, -16, -24, 5, 1, 19, 1, 7, 19, -25, 0, 37, -7, 1, -7, 3, -7, 13, -20, -10, -7, 2, -10, 7, -2, -1, -5, -38, 3, -12, -8, -24, 0, 29, -2, -43, -19, 33, -4, -76, -39, -31, 11, -5, -5, 0, -2, 3, 83, -8, -26, -36, -81, 13, 2, -8, -3, -41, -1, -17, 4, -14, -14, -17, -3, -10, -12, 6, -52, -3, 0, 23, -38, -6, -25, 56, -3, 10, 32, 11, 26, 35, -4, -22, 10, -26, -12, 1, 3, -9, 27, -19, -10, 6, 20, -5, 9, 9, 33, 42, 26, 1, -73, -5, 32, 26, 0, 0, 0, 32, -56, -31, 52, -15, -30, 0, 12, 7, -22, -21, 2, 3, 17, 18, -8, -56, -1, 5, 6, 4, 16, 13, -10, 3, 25, -3, 7, 8, 1, 44, -44, 1, 2, -5, -31, -14, 5, -35, 3, 0, -18, 12, 0, 6, 3, -38, -25, -31, -2, -44, -4, 49, -22, -19, -34, -1, -16, -21, 8, -15, -43, 8, 4, -5, 0, 16, 14, 10, -38, -19, 38, 16, 1, -9, 14, -40, -8, -6, -6, -9, 0, -25, -20, 5, 0, -13, -10, -12, 0, -13, -15, -25, 3, 30, 1, 27, 48, 7, 6, -12, -11, -13, -3, -59, 0, -9, 0, -27, 17, -20, 0, 1, 25, -4, 29, 3, 41, 37, 15, 1, -38, -4, 18, 9, 2, 1, -6, -18, -30, 0, 46, -15, -9, -13, -14, -4, -9, -1, 3, 20, 54, -13, -15, -27, 0, 13, -3, -2, 37, -39, -39, 7, 5, -13, 5, 26, -5, 28, -64, 5, 3, -8, -14, -15, -21, -31, 0, -2, 10, 6, -3, -35, 3, -9, -35, -12, -3, -46, -12, 33, -7, 26, -81, -20, 25, 6, -7, -15, 21, 1, 3, -5, -55, -8, 9, -5, 35, -6, 10, 47, -5, -8, 13, -12, -20, 1, 6, 0, 11, 5, 46, -2, -18, -34, 8, 20, 5, -27, -19, 14, -4, 8, -1, 14, -5, 8, 17, 22, 33, -15, 0, -31, 0, -33, -7, 8, 21, -27, 16, -4, -3, 6, 0, 10, 18, 18, -10, -5, -49, 7, 16, -20, -16, 6, -7, 7, -1, -11, 31, -2, -4, -24, -17, -48, -2, -11, -6, 26, 49, 12, 20, -47, 0, 3, -5, 1, -13, -10, 24, -4, -42, -10, -41, -32, -4, -2, -30, 8, -5, 3, 3, -20, 38, -8, -6, 0, -10, 14, -2, 3, 1, 2, -50, 20, -3, -39, -37, -4, 19, 3, 19, 22, 64, -17, 2, 7, -22, -16, 3, 0, 43, 30, 8, 29, 10, -11, 41, -30, 5, -19, -2, 7, -10, 1, 30, -4, 2, 20, -21, -30, 31, -10, -69, 24, 4, -70, 45, 9, 7, -12, -3, -59, 6, -38, -46, -29, 20, -42, 19, -46, -5, 6, 3, 2, -12, -7, -7, 6, 15, -7, 10, 18, -62, -25, 59, -5, 3, 2, 7, -42, -43, -6, 2, 4, 0, -49, -8, 12, -32, -89, 0, -15, -7, -21, 8, -7, 2, 8, -59, -6, 8, -18, -5, -22, -51, 36, 25, -6, -4, -11, -19, 16, 3, 48, -22, 8, -2, -4, -42, -2, 13, 31, 4, 0, 2, 0, 6, -25, 1, -50, -53, -25, 4, -22, -10, 0, 20, -42, 11, 15, 13, 9, -2, -9, -26, -13, -1, 11, 22, 37, 68, -22, 16, -14, -70, -2, -6, 5, -56, -2, -5, 5, 16, -32, -11, -7, 0, 36, -15, 0, -3, 24, -1, -14, 0, -4, 40, 44, -1, -88, 22, -15, -24, -3, 47, 1, -27, -21, -16, -10, 3, -39, 1, 2, -7, -5, 0, 3, -6, 0, 2, 33, 8, 7, -4, 7, 18, 0, -4, -1, 6, -6, 8, 20, 12, 26, -27, -2, -15, 29, -12, -5, 6, -39, 39, -26, -21, -50, -54, -35, 1, -20, -40, 18, 23, 4, 8, -8, 0, -31, -6, 39, 4, 5, -5, 5, -11, 26, -5, -63, -5, -6, -26, 2, 1, -5, 0, -56, -5, -42, 1, -32, -27, -20, 18, -21, 37, 45, 20, 31, -37, 12, -49, 12, -3, 2, 8, 7, 58, 0, 8, 0, -11, 7, -8, -5, -43, -5, -6, -2, -20, -10, -29, -1, 3, 12, -9, 0, -6, -4, 8, -22, 6, -15, 20, 37, 0, -18, 32, -34, 1, -65, 68, -28, -25, -33, -7, -5, 0, 24, 43, -20, -6, 5, -34, 0, 5, -9, 39, 52, 6, -3, 44, 3, 38, 18, -17, 10, 0, -4, -48, 2, 76, 10, -47, 4, -15, 13, -1, -39, -6, -14, 0, -27, -11, -32, -12, -27, -4, 6, -25, 32, 20, 11, 38, -23, 23, -38, -6, 38, 0, 4, -1, 7, 17, 27, -16, -16, -6, -7, -30, 3, 5, -5, 0, -66, -4, -5, 0, -33, -19, -14, 7, -90, -19, 29, -15, 45, -38, 3, -5, -29, -4, 0, -10, 51, 20, -3, -79, -38, -31, 29, -1, -1, 24, -21, 9, -7, 30, 6, -49, 8, 30, -20, -43, 16, 2, -10, 4, -51, -32, 8, -11, 30, -1, -25, 43, -39, 5, -80, 46, -21, 0, -35, -14, -18, 2, 50, 1, -32, 5, 1, -23, 1, -10, -2, -4, 34, -6, 6, 60, 3, 32, 28, -37, -1, 4, 35, -22, 5, 57, 15, -62, -7, 19, 14, -7, -34, 4, -16, 38, -31, -36, -52, -24, 9, -6, -11, -19, 26, 38, -30, 13, -19, -4, -34, 4, 10, 11, 4, -7, -2, 15, 34, -1, 6, -3, 2, -70, 8, -6, 23, -4, -16, -6, 14, 2, -6, -16, 15, -8, 0, -41, 48, -37, -8, -28, -17, 17, -18, -10, -3, -19, 5, 76, 9, -29, -1, 40, 25, -3, -21, -3, 0, -9, -10, 5, -3, -51, -3, 1, -13, -30, 1, 8, 5, -3, -4, -46, 17, -19, 60, 3, -60, 8, -33, 10, 14, 29, 3, 10, -45, -9, 48, -5, 15, 21, -22, 0, 4, -30, 5, 17, -5, 10, 27, 1, -3, -51, -2, 34, 23, -33, 0, -1, 13, -2, 5, 46, -15, -40, -1, 39, 2, -10, -55, -1, -11, 40, 9, -3, -31, -9, -10, 6, -8, 9, 0, 34, 24, -25, -19, -1, 15, -4, 11, 6, 4, 0, -2, 4, 4, 20, 2, 3, 5, -39, 0, 2, -1, 0, -31, 16, 27, -7, -19, 28, 55, -6, 23, -70, 0, -57, 13, -8, -10, 24, -20, -5, -4, 22, -1, 6, 11, 33, 27, -31, 1, 1, 32, 3, 15, 4, -9, -4, -13, -16, 1, 2, 16, -11, -11, -2, -6, 2, 9, -31, -12, 40, 23, -1, 20, 10, -5, 17, -7, 26, -3, -6, -29, -1, -21, 2, 39, 4, -40, -24, 2, -21, -4, -20, 3, 17, 28, 21, 7, -12, -4, 20, 11, -8, -4, 1, -7, -7, -22, 38, 7, -19, -34, 24, 6, -6, -25, -2, 8, 19, -29, -7, -21, -3, -3, 3, 3, 17, -4, -26, 8, -61, -23, -13, 51, -5, 8, -62, 4, 1, -4, 6, -12, 15, -9, 1, 2, -3, -7, -9, -12, 3, 38, -28, -45, -3, -32, 5, 90, 2, 24, -63, -11, -2, 32, -4, 11, 6, -4, -1, -4, -23, 0, -6, 29, -6, 19, -3, -12, -2, 0, -6, 28, -19, -8, 5, 9, -74, 0, 21, 10, -12, -2, 0, 11, 4, -79, -30, 1, 26, 3, -7, 26, -14, -22, 1, 30, 9, -19, -7, 19, -4, -40, 5, 4, 35, -17, -24, -6, -27, 5, -15, 13, 5, -42, -15, 4, -15, 3, 26, -31, -36, 0, 1, 0, -24, 9, -18, -10, -32, -57, 38, 24, 4, 0, -1, 28, 6, -21, -2, -38, -23, -4, 1, 12, -11, -27, 28, 2, -9, 6, -32, -77, 0, -37, -10, -5, -4, -1, 25, 32, 16, -34, 4, -2, -32, 24, 6, -3, -4, 49, 8, -21, 6, -7, -25, -10, 34, -9, 6, -27, 37, -26, -39, 34, -22, -3, 1, 7, 29, 25, 34, 0, 31, 49, -27, 7, -4, -14, -42, 20, -4, -11, 18, 5, -22, 7, -21, -56, 17, 27, -75, -9, 5, -40, 34, 8, 11, 16, 4, -38, -12, -22, -16, 7, -42, -31, 36, -31, 2, 42, 6, -2, 0, 15, -15, 0, 27, -7, 11, -6, -14, -33, 30, -7, -27, 0, 31, 0, -42, 1, 5, 13, 0, 3, 9, -26, -29, -86, 19, 15, -66, -1, -4, -9, -3, -2, -13, -4, 10, -19, -3, 28, -100, 35, 30, -6, -9, 11, -11, -16, 7, -14, -2, 10, -2, -4, 7, 27, 27, 54, -2, -6, -31, 9, -8, -1, -4, -22, 2, -23, 0, 27, 35, -14, -5, -8, 18, 9, 33, 38, -17, 52, -61, 11, 4, -6, -3, 12, 59, 14, 48, 36, -38, 5, -1, 15, 18, 52, 25, 3, 29, -7, -10, 10, -3, -26, -17, 16, 1, -10, -6, -7, -9, -10, 14, 22, -9, -67, 1, -13, -2, -35, 17, 1, -19, 0, 14, -18, 6, -32, -15, 14, 2, 1, -40, 0, -14, 2, 17, 0, 18, 6, -59, -1, 23, 34, -14, 5, 4, 18, -2, -30, 1, -7, -29, 16, -5, 15, 15, 22, 1, -62, 39, 3, -9, 8, -40, -24, 2, -1, -26, 32, 19, -7, 8, 7, -17, -21, 4, 12, 30, 5, 3, 7, 0, 54, 29, 8, -5, 3, -118, -18, 0, -9, -5, -35, -58, -21, -7, 27, -5, -13, 0, 7, 8, 37, 22, 41, -18, 14, -55, 23, -5, 0, 0, -1, 100, -29, 48, 10, 50, 19, 0, 2, -18, 67, 1, 3, -5, 24, -18, 45, 29, -38, -17, -10, 41, 20, -2, 21, -64, -9, 59, 19, 2, -22, 6, 15, -28, -60, 45, 2, -22, -18, 7, -8, -3, 20, 33, 53, -20, 1, -68, 0, -10, -4, -18, -1, -12, 0, 50, 1, 38, 18, 0, -4, -3, -18, 20, -23, -11, 17, -2, 8, -37, 10, -10, 27, -1, 1, 38, -13, -39, 9, -34, 0, 0, 2, -13, 27, 22, 1, 48, -7, -5, -26, 3, -21, 48, -4, -5, 0, -3, 55, 12, -19, -1, 3, -103, -4, -7, -30, 1, -33, -32, 8, -4, 30, 26, -6, 14, -18, 25, 18, -17, 44, -20, -15, -46, -11, 5, -5, 1, 6, -15, -10, -24, -9, -1, 61, 0, 7, -20, 7, -4, -8, 12, 22, -27, 13, 25, -42, -20, 9, 24, 13, -2, 14, -43, 29, 12, 22, 0, -8, 3, -10, -46, -84, 30, 20, -3, -106, -3, -2, -5, 65, 14, -17, 38, -5, -127, -1, -17, 13, -3, 13, -12, -1, -35, 2, 39, 16, 0, -1, 0, 1, 28, -2, -30, 21, -17, 33, -25, 6, 6, 1, -6, -7, 44, 5, 15, -27, -12, -8, 3, -9, 18, 53, 48, 4, 19, 0, 16, -19, -3, 13, 42, 0, -9, -3, 17, -14, 31, -26, -2, -3, -101, 15, 0, 7, 0, 2, -43, -18, 1, 17, 5, -28, 8, 5, 13, 5, -3, 61, -33, 8, -32, -15, 0, -7, -9, 20, 37, -5, -14, 22, -30, 20, -3, 14, -37, 29, 5, -8, -16, 4, -42, -2, 0, -4, 15, 3, -10, -8, 5, 3, -78, 3, -21, 21, -7, -37, 30, -41, -16, -73, 13, -9, 9, -52, -4, 16, -4, 13, 8, -12, 3, -1, -130, 0, -13, -3, 26, 21, -2, -8, 14, -3, 41, 40, -9, -1, -8, 21, 0, -7, -22, -39, -53, -2, -13, 15, 37, -29, -3, 6, 39, -31, 29, -62, -6, -11, 1, 22, 37, 75, 23, 10, 6, -20, 41, 33, 6, -24, 17, 12, -5, 3, -4, 20, 0, -3, 3, -3, -25, 21, -7, 5, 0, -48, 8, -6, -6, 3, 11, 8, 17, 27, 24, 20, -38, 65, -38, 0, 0, 2, -4, 0, -16, -2, -25, 9, 33, 4, -81, 17, 0, 19, 18, 59, 17, -4, -14, -1, 0, 11, 29, -15, -16, 7, 25, 0, -8, -8, -42, -20, 1, 37, 0, 15, 24, 10, 14, -61, 50, 7, -5, -43, -15, -3, -2, 4, 28, -17, 4, 7, -87, -2, -36, 15, 11, -13, -7, -2, 39, -4, 29, 18, -12, 1, -8, 14, 4, -30, 32, -11, -46, -19, -1, 19, 13, 14, -5, -3, 46, -21, 36, -37, 33, 36, 2, -12, -3, 25, -82, 25, -8, -13, -10, 25, 3, -79, -24, -2, -3, -6, -12, 31, 5, 34, -3, 2, -16, 11, -5, 0, -3, 38, -26, -12, 0, -27, 4, 38, -3, 23, -19, -19, -10, -2, -23, -28, 2, 13, 8, 5, -24, -21, 22, 32, 26, 15, -20, -16, 2, 66, 10, 80, -33, 5, 2, 31, -33, 23, -5, -21, 47, -21, -57, 16, 7, 11, -59, 36, 64, 4, -3, -32, -20, -26, 21, 27, -45, -11, 14, -15, 8, -2, 2, -3, 16, 0, -9, -4, 15, 1, -10, 14, 0, -9, -29, 7, 48, -4, 42, -48, -35, -6, -1, -7, 0, 3, -16, -36, -7, -60, 3, -11, -72, -29, -6, 34, 45, 0, 35, -83, 15, 36, -2, -17, -6, 10, 1, -9, -33, -1, -35, 22, -6, -14, -55, -4, -8, 5, -20, 22, 43, 27, 0, 0, -36, 14, 3, -55, -1, 69, -22, 7, 3, -38, -30, -31, 42, -3, 17, -32, -24, 24, -15, 84, 22, -17, 0, -3, 16, 47, 76, -29, 66, 44, 0, 5, 8, -47, -6, 24, -23, 3, -3, 64, -51, 15, -3, -50, 7, -42, -91, -27, -5, -4, -36, 15, 9, -24, 3, -74, -43, 33, -36, 52, -33, -37, 98, -6, 4, 1, -2, -15, -14, 9, 53, 4, -9, 3, 40, -1, -78, -36, 32, 4, -67, 0, 21, -38, -44, 0, -1, 38, 0, 11, 13, 0, -21, -122, -27, -43, -90, -7, 2, -27, 17, -10, 87, -3, 21, 15, 2, 5, 9, 27, 0, -7, -1, -6, -36, 8, -2, 1, 40, -1, -3, 4, -22, 26, -1, -40, -5, 1, -7, 0, -2, -13, -6, -23, -27, 10, 2, 16, 12, -6, 8, 21, 27, -11, -14, -31, -40, 89, 9, -11, 0, -2, -23, 8, 5, -19, 31, 59, -34, -15, -2, -4, -11, 58, -11, -1, 6, 27, -23, 25, -17, -11, -3, 6, 11, 0, 0, 25, -41, 19, 21, 5, 0, -42, 29, 46, -27, -36, 12, 20, 17, 20, -9, 7, 3, -26, 12, 24, 3, 2, -64, 0, -35, 8, -36, -2, -18, 2, 1, -1, 18, -24, -18, 0, -7, 7, -8, 20, -37, 32, -24, -10, -15, -16, -7, 1, -2, -5, 37, -34, -45, -6, -3, 0, 4, 6, 14, 70, 35, -8, -6, -4, 1, -25, 4, -13, 51, 5, -4, 5, -30, 44, -3, -27, 0, -3, -89, 10, -1, -18, 1, -63, 45, 30, 5, 25, 42, -6, 16, -4, 37, 9, -19, 27, -24, 85, 21, -16, 4, -8, -26, -5, 21, -4, 41, 31, -37, 0, -1, -28, -8, 76, -20, -1, -5, 23, -13, 35, -5, 0, -41, 49, 26, 11, 2, 5, -44, -3, 24, 22, 4, -38, 7, 30, 7, -65, 23, 16, 20, -37, -12, 8, 2, 15, 10, 25, 11, 0, -127, 5, -29, 13, 25, 9, -3, -7, -52, 0, 9, -9, 0, 3, -1, -8, -6, 42, -21, 67, -20, 14, -13, -7, 1, -7, 1, -9, 6, -7, 37, 23, -1, 2, 2, 13, 11, 24, 24, -3, 16, -7, 6, -48, -1, -42, 55, 0, -2, -1, -6, 53, 3, -33, -3, -1, -103, -17, -4, -29, 6, -18, 47, 1, -3, 25, 31, -23, 32, 3, 2, 7, -16, 15, -34, 41, 16, -26, 1, -7, 22, 10, -48, 23, 10, 33, -22, 15, -8, -43, -7, 90, -6, 7, 0, -5, -5, 30, -1, 7, -4, 11, 46, -12, 4, 3, -23, 32, 46, 20, 0, 2, 27, 50, -41, -76, 9, 41, 1, -70, -9, 6, -1, -22, 10, 5, 31, 0, -140, -3, -13, 0, 1, 15, 14, -9, -53, 0, 44, -6, 18, -7, -4, 17, 0, -10, -9, 0, -27, 7, 16, 2, 2, 27, 7, -17, 14, -26, 4, 2, -18, 2, 1, -8, 3, 21, 30, -31, -14, -3, -1, 1, -4, 7, 40, 11, -1, -2, -11, 53, 23, -11, 5, -4, -152, -27, 5, -21, -6, -21, 0, 14, 0, -5, 15, -15, 15, -18, -9, -11, -23, 46, -11, 49, 6, -1, -4, 1, 5, -13, 53, 20, 37, 51, -33, -6, 0, -12, 0, 45, 9, 12, 1, -22, 12, 28, 20, 5, -14, -15, 34, -16, 6, -6, -66, -19, 54, 32, 2, 3, 14, 27, -15, -77, 6, 25, 11, -48, -10, 26, -4, 23, 3, 18, 19, 1, -167, -8, -33, 4, 15, 9, 2, 5, 29, 5, 36, -20, 11, -7, 5, 1, 18, 6, 8, -14, -21, 8, 17, -24, 0, 16, -5, 17, 30, -15, 0, -11, -13, 11, 0, -22, -30, -1, 13, -6, -12, -7, -1, -2, 3, 5, 13, 0, -1, 0, 8, 45, 50, -60, 3, -8, -72, -5, -6, -26, -7, -23, -4, 12, -7, -26, 0, 0, 20, 35, 21, -12, -26, 15, 18, -9, 29, 27, 2, -7, 17, -16, -21, 34, 64, 24, -25, 8, -4, -19, 4, 62, -2, -2, -9, -4, 1, 64, 9, -33, -20, 1, -19, 24, 0, 10, -39, -20, 78, 55, 6, -15, 23, 58, 0, -20, 22, -9, 29, 5, -1, 23, 6, 43, 7, 34, -6, -1, -49, 4, -23, 10, -11, 22, 0, -5, 48, -5, 35, -20, -14, -6, -8, 0, 27, -18, 24, -18, -1, -23, -14, -18, -4, -18, -3, 2, 62, -35, 0, -2, -23, 59, 5, 1, 5, -39, -91, 0, -16, -3, -57, 43, -7, -59, -36, 2, -6, -2, 9, 112, 19, -48, -2, 3, 17, 16, 3, -34, 0, 40, -80, -39, 1, -77, -20, 15, 12, 44, -18, -10, -54, -27, 35, 0, -9, -13, 3, -8, -66, 38, -11, 42, 28, 66, -57, -10, -6, -21, 11, 84, -48, 0, -26, 34, -26, -7, -14, -12, 39, -33, -58, 26, -1, -8, -53, 54, 19, 6, 5, 78, -17, -71, 14, 7, -37, -61, 32, 27, -2, 27, -4, 19, 22, -7, 37, 0, 11, -7, 15, 9, -25, -32, -50, 6, -23, -3, -15, -66, -75, -3, 0, 45, 6, 64, -15, -16, 16, -124, -33, -69, 12, -3, -1, 20, 62, -20, -23, -96, -36,
    -- layer=2 filter=0 channel=9
    33, 2, 9, 5, 20, 1, 4, -11, -1, -65, 33, 1, -1, -53, -5, 9, 3, 8, -15, 11, -54, 3, -1, -6, 4, -6, -30, 0, 6, -1, 8, -5, -19, 0, 0, 2, 22, -23, -2, -21, -43, 27, 32, -38, 4, -1, 2, 1, 19, 34, 11, 28, -30, 51, 12, 3, 45, -1, 42, -27, -10, -39, 23, 0, -21, 31, -7, -1, 27, -41, -54, -1, -35, 11, 11, -31, -17, 1, 40, -12, -17, 31, -35, 1, -22, -11, 13, -20, 27, -5, 56, 10, 19, 13, 4, -16, 3, 34, -13, 30, 28, -50, 5, 29, 2, 35, 10, -27, 3, -1, 57, 5, 53, -3, 34, 11, -34, -10, 15, 32, 18, -5, 23, -38, 29, 24, -6, -39, 6, -4, 10, -5, 30, 0, -23, -24, -5, -26, -36, 4, -1, -56, -2, 7, 6, -3, 0, 8, 4, 0, 1, -35, 0, 7, -19, -4, 41, 18, 3, -4, -14, -1, -31, -16, 32, -22, -10, 7, -56, 2, 10, 0, -4, -2, -2, -46, -8, 58, -4, 58, 30, 15, 22, -4, 12, -12, 42, 16, -4, 0, 16, 4, -15, 28, 15, -21, -15, -4, -59, -5, -45, -5, 0, 0, 12, 3, -3, -28, 36, 18, -35, 6, 0, -11, -16, -15, -4, 0, 22, -15, 4, -8, 0, -4, 6, 16, 0, 16, -36, -20, 7, 4, 2, 2, 3, -31, 4, 7, 19, 7, 5, 22, -42, 9, 27, -10, 0, 8, 18, 0, -4, 0, 13, -36, 20, -22, -6, -7, 1, 5, 28, 14, -9, -19, -11, 16, -36, 0, 26, -12, 3, 3, -1, 19, 12, 33, -15, 7, -3, -34, -17, -4, 12, -1, 0, 11, 14, -3, -8, 15, -10, -11, -10, 14, 4, 5, 12, 17, 29, -8, -25, 0, -1, -11, 18, 22, 28, 10, 9, 33, 7, 4, 0, -80, 37, -11, -12, -8, -12, -16, -3, 10, -40, -11, 26, -16, -32, 2, -48, -15, 7, -42, 1, 2, -19, 32, -13, 0, 5, -4, -17, -11, 13, 1, 2, -6, 31, 10, -43, 13, 2, -8, 0, 22, 7, 7, -12, -1, -1, -61, 2, 7, 9, -27, 1, 8, 9, -21, 5, -34, 7, -16, 28, -11, -6, 26, 25, 0, 10, 19, 4, 7, 10, -36, -13, -4, 17, 6, 44, 29, 19, -7, 6, 19, -31, -2, -17, 18, -5, -5, 5, 6, -4, 19, -21, 4, -6, -17, 0, -9, 23, -8, -42, 19, 36, 5, -10, -13, -32, -14, -9, -6, 20, 17, -13, 5, 40, -20, -26, -3, 1, 39, 2, 49, 16, 52, 5, -8, 31, 3, 5, -20, 25, -21, 0, 21, 29, -37, 12, 12, -6, 22, 15, 4, -16, 7, 15, -6, 10, -11, 27, 3, -7, 33, 9, -1, 0, -21, -12, -21, -48, -10, 8, 5, -2, 37, -44, 2, -2, -9, -4, 12, -24, -8, -5, 8, 6, 14, 2, 35, 15, 5, 4, 7, 3, -19, 1, -31, -4, -20, 15, 14, 8, 58, -2, 0, -23, 56, 0, 57, 10, 29, -4, 4, 3, -11, 37, 13, 34, -37, 5, 0, -13, 2, -24, -43, -9, 1, 3, -28, 9, 22, 5, -5, -4, 3, 8, -7, 15, -3, 6, 40, 24, 4, -5, -7, -33, -14, -21, 31, 1, -13, -62, -3, 56, 10, -20, 6, -6, 18, 8, 13, 19, 35, 17, -39, 0, 0, -9, 1, 54, -11, -18, 36, 3, -47, 26, 13, 15, -23, -16, 5, -6, 2, -20, 3, -8, -28, 37, 0, 38, -17, 41, 13, 0, -42, -16, -3, -57, -8, -5, -2, -3, 18, -2, 8, -7, -18, 6, -8, -15, -3, -35, 26, 2, 6, 5, 25, 35, -15, -7, 5, 11, -11, -4, -43, 0, -19, -2, 5, 3, 19, 3, 1, -15, 21, 1, 10, 38, -19, 8, 2, 7, -25, 39, -7, 19, -16, -10, 22, -29, -5, 11, -43, 3, 0, -3, 30, 19, 25, -9, -5, 0, 2, 5, -2, -9, 5, 23, 13, 45, -5, 5, -28, 9, 0, -10, -7, -14, 26, -59, -14, 71, 9, 0, 2, 4, -20, 9, 0, 16, 56, 40, -70, -13, -7, 38, -11, 30, 5, -10, 26, 16, -18, -1, -6, 31, -23, -15, 0, -36, 0, -26, 6, 5, -24, -10, 4, 0, 2, -14, 0, -12, 1, -11, -16, 15, -13, -15, 0, -8, -13, -14, 25, 0, -53, -6, -3, -7, -3, 10, 3, -7, -49, -1, -4, 0, -9, 0, 3, 31, -21, 42, 11, -7, -1, 13, -7, -3, 20, 33, 6, -56, -9, 14, 12, 21, -9, 31, 4, 7, -8, 38, -15, 2, -23, -1, -15, -15, -8, -16, -51, 4, -1, -4, 20, 14, 5, -34, -1, 5, -12, 19, 6, -11, 8, -21, 19, 54, -4, -15, -33, -29, 11, -7, -26, -9, 26, -21, 16, 62, -20, 7, -4, 7, 13, 0, 0, 5, 23, 30, -31, -26, -2, 30, -1, 22, 13, -11, 28, 34, -2, -1, 27, 43, -39, -21, -31, -37, 5, -35, 24, -6, -13, -13, 0, 21, -23, -49, -13, 29, -20, -15, -7, 29, -12, 0, 1, 8, -19, 0, -5, 7, 16, 3, 32, -5, -18, -3, -12, 0, -12, -7, -8, 3, 14, 6, 7, 32, -1, 33, 5, 16, 29, 4, 12, 1, -21, 21, 7, -36, -11, 37, 44, 28, -49, 9, -5, 2, 8, 6, 23, 28, -25, -9, 17, 16, 6, -5, -31, -1, -4, -3, 4, 4, 12, 1, 3, -2, 17, -6, -2, -30, 7, -4, 17, 0, 4, 31, -10, -11, 0, -3, -35, -54, 11, 5, 18, 6, 14, -10, 1, -1, 2, -10, 31, 33, -14, -5, -30, 2, -1, -2, -48, 6, 1, -10, -24, 19, -2, 5, -8, 8, 2, -25, -13, -56, 6, -26, 4, 21, -7, -24, 2, -25, -13, -27, 2, 17, -48, 3, -8, -5, -13, -3, 2, 24, -25, -5, 4, -6, -8, 0, -28, 0, -22, 20, 8, -4, -73, -7, 27, 14, 1, -4, 4, -29, 1, 14, 5, 8, -5, 9, 1, 29, -2, 51, 4, -70, 0, -2, 50, 20, -3, -10, 2, 20, 7, 15, 0, -9, -32, -14, -35, 5, 3, 2, -16, 0, 3, 0, -18, 12, 7, 26, 0, 3, 26, -16, -2, -9, 9, 0, 50, 64, 7, -13, -10, -5, 5, -3, 0, 0, -19, -7, 14, -4, -2, 19, 0, -1, -16, -26, 9, 7, 6, -5, -23, -4, -2, 14, -9, -6, 5, -2, 10, 21, 1, -7, 9, -24, -56, 13, 21, -34, 9, -37, -12, -16, -44, -15, -3, -17, -22, 28, -47, 14, 16, 16, 34, -15, 8, 19, 4, 3, 7, 12, -31, -5, 13, 2, 4, -7, 19, 8, -13, -2, 36, 2, 18, -19, 1, -1, -1, 0, 3, 1, 4, 6, -16, 32, -6, -14, 0, 6, 2, -19, 36, 3, 29, 8, -9, -12, -1, 0, -43, 29, 31, 48, -23, 1, -54, -34, 8, 11, 11, 0, 5, 1, 0, 0, 18, -3, -4, -5, 12, -9, 6, 13, 0, 4, 7, 19, 4, -25, -11, 0, -2, 5, 51, 26, 4, -20, 0, -6, 41, -18, 6, 3, -7, 6, 34, 23, -25, 3, -71, 2, -6, -6, 12, -8, 5, -9, -26, 10, 0, -14, 13, -4, -11, 20, 2, -13, -4, 0, -56, -17, -17, -17, 5, 14, 14, -6, 14, -9, 15, -2, -24, 0, -16, 39, -2, -4, 24, -38, -31, 6, 8, 2, -9, -6, -28, -10, -3, 5, -4, 6, 0, -13, -22, 0, -2, -24, -3, -9, 28, -9, -2, 41, 12, -28, 10, 8, -2, 0, 57, 22, 19, 5, -2, 2, 7, -1, -34, 33, 13, 20, 23, 1, 10, -42, -2, -36, 6, -14, 6, 5, -2, -23, 30, 0, 6, 0, -7, 3, -5, -11, -6, -7, -6, 13, 4, -3, -13, 16, -1, -18, 2, 16, -7, -29, 7, 7, 43, 5, -1, 0, -3, 12, 40, -8, -16, 3, -45, 3, -4, 38, 7, -19, 14, -2, 7, 4, -2, 9, 26, -12, -34, 24, 10, 0, 6, 9, -29, 3, -48, 24, -2, 70, 8, 8, 5, 21, -15, -4, 7, -12, -3, 24, 1, 5, 37, 11, -37, -1, 32, -1, -20, -12, -24, -23, 8, -6, 14, -5, 30, 0, -26, 5, 1, -45, 14, -5, -7, 28, 5, 24, -36, -12, 2, 4, 2, -42, 63, -6, 16, -7, -4, 6, -5, -10, -67, -22, 24, 5, -28, -5, -9, -30, 6, -38, 3, 0, -5, 2, -17, -5, 31, 26, -6, -8, -1, 8, -2, -15, 1, -18, 14, 44, -5, -25, -23, 0, 10, 1, -19, -2, 19, -20, -16, 1, 0, -7, -4, -1, -12, -7, 53, -6, 1, 5, -62, -15, -6, 31, 40, 17, -3, 5, 8, 16, 0, 10, 12, -63, -4, 2, 3, -16, 0, 14, -43, -6, -11, 62, -3, 41, -1, 8, -8, 29, -8, -21, 27, -48, 2, 4, 0, 9, 24, -13, -19, 2, 30, -2, -35, -12, -33, 0, -1, -3, -35, -5, 23, -26, -35, -4, -1, -12, -3, -28, 2, 1, -51, 10, -39, -1, -16, 37, 2, -75, 45, -34, -4, -29, -9, 19, 5, 10, -61, 21, -14, 3, -11, -12, 19, -49, 8, -2, -13, -3, 7, 0, -19, 9, 22, -63, -6, 3, 23, -8, -7, -42, -5, 6, 9, 5, -7, 16, 2, -8, -2, 26, -20, 5, -18, 0, -23, 10, 41, 2, -2, 8, 4, 19, 24, 39, 30, 9, -31, 18, 1, 34, 58, -1, 1, 5, -25, 9, 3, 1, 7, -7, -42, -9, 8, -22, -3, -18, -9, -5, 23, 11, -6, 31, 9, -8, -1, 5, 20, -18, -14, -5, -12, -2, 1, -12, 30, -34, 39, -2, 23, -7, -8, -2, -28, 25, 26, 0, -46, 2, 19, -10, 1, -6, 2, 13, -14, 29, 23, -18, -10, -3, -3, -2, 0, 37, 5, -47, 16, -5, -8, -13, -43, 18, 0, -6, -30, 16, -21, -34, -27, -7, 12, -19, 4, -25, 3, -1, 6, 0, -19, 5, 17, -21, 2, 2, -7, -11, -5, -34, 0, 6, -47, 32, 4, 1, -4, 26, 15, -15, -18, -1, 17, -7, 14, -4, 34, 7, 3, 1, -20, -49, 40, -8, 16, -26, -51, 1, 0, 20, -22, -15, 8, -4, 14, 20, 6, -4, 2, 32, 5, 12, 13, -15, 2, 3, -24, 0, 11, -3, -7, 43, -12, 23, 7, 20, 21, 16, 2, -4, -13, 28, 0, 11, 1, 8, 7, 4, 7, -7, 13, -23, 28, -24, -13, 0, -11, -3, 0, 6, 3, -2, 4, 41, -5, 21, -1, -2, 5, 45, 12, 13, 37, 93, -6, -33, 0, 13, -9, 23, -21, -11, 0, 0, 8, 13, 16, 42, -41, -6, 0, 38, 0, 1, 0, -7, 3, 2, -5, -14, 6, -17, -5, 3, 32, -2, 5, -7, 0, 9, 0, 24, 1, -18, -24, 15, -13, -15, -16, -58, 15, 24, 15, -1, 7, -7, -7, 6, -8, -1, 0, -16, 0, 22, -27, -35, -1, 10, 11, -3, 0, -6, -11, -33, 5, 12, -25, 18, -1, 27, -28, -44, 7, 24, -12, -24, 27, 12, -5, -38, -9, 0, 30, 7, -70, -1, -24, 11, -13, 4, -4, 1, 3, -36, -1, 0, 19, 4, -56, -14, -39, 25, -2, 0, -4, -6, 27, -6, 44, -3, 7, -31, -44, -2, 12, -15, -7, 17, -18, -9, 18, 3, 0, -31, 13, -38, 55, -12, -28, 20, 5, 8, -11, 8, 10, 3, -21, -15, -48, 25, 1, 5, -1, -8, 4, -7, -21, -26, 2, 47, 4, 5, 23, 6, -2, -26, -5, 15, -42, -27, -5, -19, -16, -10, 10, -2, 13, 9, -14, 18, 7, 8, -8, 41, -4, -4, 31, -3, 5, 9, 30, -10, -38, -12, -3, 26, 8, 22, -19, 3, -5, -7, -13, -1, 4, -12, 14, 4, -27, -11, 2, -9, -55, 0, -3, 17, 1, -7, 20, -5, -27, 30, 0, -37, 27, 11, -21, 17, 4, -44, 29, 5, -19, -4, 28, -1, -3, -8, -33, 24, 6, 3, -40, -7, 33, -28, 9, -1, 5, -2, -23, 38, -37, 13, 12, -13, -3, -14, 6, 18, -4, -26, 24, -55, 55, -1, -12, -1, -2, -14, -11, 6, 4, 5, -21, -18, -46, -50, 2, -7, 4, -2, -6, -2, -12, 27, 0, -13, -5, 5, 27, -5, -2, -24, 0, -48, 3, 0, -1, -28, -28, -7, 20, -17, 38, 45, 31, -16, 7, 16, 1, 8, -4, -4, 13, 19, -9, 2, -22, 0, 0, -18, -9, -7, 15, -2, 0, -17, -13, 8, -2, 0, 0, -38, 25, 11, -10, -8, 4, -25, -52, 27, -15, 28, -3, 8, 12, -16, 7, 44, 15, -18, 32, 5, -7, 7, 0, 3, 30, 13, -2, 3, 31, 3, 2, -27, -35, 22, 16, -7, 4, 4, -5, -16, 19, -5, 2, 10, 6, -3, 18, -14, -14, 22, -29, -34, 9, 12, 6, -48, 8, -33, -6, 10, -18, 24, 0, -24, -49, 16, -12, -11, 16, -2, -35, -50, -2, 45, -14, -8, -7, -4, -34, 20, 1, -1, 0, -4, 41, 0, -7, -16, -7, -29, -6, 13, -3, -21, 2, -4, 14, -2, 47, 18, -20, -50, 20, -21, 21, 0, -4, 0, 4, -22, 22, 3, 0, -16, -12, 0, -9, 23, -25, 13, 6, -6, -24, 9, -21, -4, -13, 8, 10, -6, 14, 12, 3, -25, -54, 3, -5, 17, -1, 45, -10, -18, 24, 43, 0, -2, 0, 8, -21, 18, -7, -60, 23, 23, -4, -1, 61, 0, -3, -17, 36, 22, 6, 1, 30, 2, -7, -19, 13, 7, -4, 3, -26, 7, 28, -16, -2, 41, -41, -27, 64, -10, -5, -39, 16, -40, -55, -17, 12, 32, -5, 15, -21, -4, 4, 7, 1, 5, -11, 3, -1, -2, -16, -11, -5, 2, 2, -26, 14, 16, 0, -2, 31, -24, -1, -20, 0, -30, -19, 2, 0, -8, 2, -6, 14, -44, 23, -24, -25, -41, -18, -14, -18, 3, 5, -6, 4, -22, 46, 5, -26, 3, -19, 13, 0, 24, 26, -23, -23, 9, -2, 0, 7, -21, 44, -13, 30, 8, -8, -5, -3, -47, -38, 3, 20, 43, 6, 16, -13, -37, -11, 50, -21, -38, 25, 26, 0, 10, 1, 9, 31, 20, -18, -5, 69, 4, 15, 0, 17, -18, -11, 0, 62, 4, 22, -7, 37, -2, 1, 0, 30, -19, 38, -28, -21, 30, -29, -14, 19, 1, 0, -68, 18, 7, -52, -2, -11, 13, -6, 17, -31, -16, 0, 3, -10, 4, -13, -8, -8, -19, -6, -4, 1, -9, 34, 39, 10, -21, -2, -8, 8, 0, -7, -14, 1, -44, -4, -40, -3, 0, -21, -3, 0, -24, 9, 4, -71, -21, -18, -4, -15, -9, -3, -2, -31, 9, 39, 52, 9, -3, -50, 22, -10, -11, 21, -10, -16, 2, -29, 4, 0, -11, -1, -53, 2, -23, -19, -8, -6, -72, -51, 5, 0, 11, -3, -25, 0, -11, 0, 44, 31, -35, 28, 14, -22, 9, 7, 13, 11, 5, 29, 4, 14, -8, 0, -20, -16, -31, 0, 1, 5, 5, 17, -9, -5, -7, 7, 3, 34, 0, 13, -7, -33, -7, -18, -22, -3, 69, -3, -59, 13, 5, -9, -6, -19, 17, 0, 33, -19, 4, -29, 29, -10, -4, -22, 4, -5, 21, 24, -7, -5, 4, -27, 12, 5, -31, 7, 7, -4, 9, -6, 24, -1, 4, -33, -26, 2, 22, 17, 1, 7, -8, 5, -14, -36, -11, -19, 2, -22, -18, 0, 1, -41, -3, 26, 24, 4, -16, 14, -23, -5, 25, -5, -1, 1, 4, -25, -15, 2, -22, -30, -6, 22, -21, -62, -31, 1, -7, -9, -7, 0, -29, -6, -15, 7, 16, 25, 28, -39, -15, 14, -21, -13, 9, 0, -10, 2, -12, -28, -4, 40, 0, -34, -11, 0, 0, -13, -6, 48, -4, 22, 1, -10, 6, 6, -18, -48, 4, -11, 9, -42, 5, -11, -6, 5, 24, -4, -19, 57, -36, 17, 10, -9, -32, -4, -42, -20, 10, -14, 38, -91, 4, 21, -11, -2, -39, 15, -7, -8, 0, -8, -33, 8, -39, -1, -7, 21, 6, -5, -12, -6, -12, 23, 8, -6, 0, 5, -9, -3, -33, -20, -59, 16, -5, -17, -7, 29, -7, -4, 5, -15, -25, 12, -20, -2, 8, -48, -35, 0, 13, 68, -12, -17, 4, -4, 4, -7, -2, -68, -26, 18, 13, -38, -1, -1, -2, -18, 4, -18, 16, 7, -14, 32, 58, 9, 28, -107, 6, -25, -28, -8, -3, 3, -75, -8, -65, 2, -8, 17, 7, -30, -18, -11, -31, 11, -4, 20, -5, 18, 0, -37, 0, -2, -26, -56, 25, -21, -5, -53, -45, -5, 6, 34, -8, -5, -19, -6, -39, 1, -12, 5, 11, -8, 23, -42, 2, -17, 1, 10, 3, -48, -39, 4, -16, 16, -8, -5, -4, -12, 15, -1, -24, -4, -6, 29, 26, 0, 7, -8, -30, -21, -35, 0, -8, -4, 24, 28, -18, -2, 18, -9, -18, -4, -25, -45, -4, -2, 4, 21, -2, 6, -4, -30, -2, -64, 13, 1, -36, 54, 0, -6, 6, 21, 3, 39, 17, 11, -58, 18, 17, 21, -10, -2, -24, -27, 15, -56, 1, 6, -20, 24, 16, -9, 21, 17, -25, 39, 11, 0, 0, -7, -18, 19, -11, 19, -5, 51, 3, 49, -2, -4, 20, -9, -3, -27, 6, -2, -16, 27, 4, -6, 37, 49, 2, 35, -39, 9, 40, -42, -30, -5, 0, -4, -40, 3, 19, -55, -19, -13, 53, 2, 25, -17, 0, -2, -24, 44, 1, -37, -26, -1, 1, 13, 0, -3, 0, 14, -13, -20, -57, -3, -3, 38, 5, 1, 11, 4, 7, 20, -63, -6, 6, -16, -32, 28, -13, 18, -19, 12, 7, -2, -26, 4, 37, 4, 7, -8, -10, 39, 0, -55, -4, -57, -11, 5, -5, 53, -1, -20, -7, -10, -21, 28, 9, -4, -86, 7, 18, 17, 7, 3, -27, -76, -10, -95, 4, 4, 26, 9, 0, -49, 34, 21, -27, 14, -10, -11, 7, 4, -15, 13, 53, 38, 7, 49, 3, 17, -10, -58, 18, -18, 7, -34, -6, 18, 2, 16, 2, -5, 19, 34, 37, 42, -25, -16, 55, -24, -49, -29, -23, 4, -53, -4, -1, -30, -18, 19, 27, -3, 8, -70, -6, 6, -19, 55, -12, -12, -7, 0, 36, 15, -3, 6, 6, -24, 12, -21, -28, 6, 3, 21, -2, 4, 10, 1, 0, 18, -20, 0, 27, 0, -8, 4, -3, 12, 0, 24, -69, 5, -13, 29, 18, 5, -2, 5, -8, 43, 46, -29, 9, -49, 33, 4, 27, 40, -52, 1, 4, -24, 1, -20, -1, -14, 0, -1, 32, -26, 13, 3, -37, -54, -4, -15, -15, -6, -37, 7, 29, -3, 32, 25, 14, 1, 13, 0, 12, -1, -13, 18, 55, 0, -1, 67, -1, 16, -32, -18, 51, -5, 6, 30, -6, 30, 16, 10, 0, 2, 55, 22, -17, 74, -30, 15, 54, -7, -23, 1, -92, -7, -67, 36, 0, -67, 28, 31, 25, 1, -13, -33, -44, -21, -9, -4, -7, -31, -39, 3, 3, 23, 3, 6, 0, 9, 55, -5, -94, -5, -8, 54, -17, -8, -10, -1, -19, -3, -30, -4, -21, 12, -13, 6, -14, 26, -5, -29, -61, -1, -38, 6, 21, 6, 7, -11, -1, 41, 6, 0, 11, -56, 33, -4, 21, 43, -7, -8, -11, -39, -13, 11, -2, 2, -19, 11, -13, -20, 5, 8, -40, -44, 21, 13, 8, -7, -36, -24, 50, 3, 24, 10, -5, 13, 17, -13, 12, 3, -18, 9, 33, 11, 3, 62, -3, 8, 3, -10, 48, -21, 4, -43, 7, 5, 14, 17, -3, -1, 28, 40, -27, 65, -46, 0, 24, -16, -26, -16, -3, 4, -106, 8, 21, 2, -3, 0, 12, -2, -15, -65, -24, 6, 10, 11, 4, -54, 36, -4, -3, 8, -10, 3, 2, 23, 8, 5, -21, 2, 6, 32, 5, 3, 6, -2, -65, -25, -44, 5, -11, 3, -10, 23, -22, 19, 38, 23, -31, 2, -17, 41, 32, 7, -4, -15, 12, 14, 50, -22, -17, -43, 21, -6, -16, 45, -29, 16, -4, -18, -25, 0, -9, 48, -38, 33, 13, 25, 8, 0, -43, -58, 19, -14, 27, -3, -57, 34, 5, -16, 28, 41, -13, 22, 8, -8, 21, 7, 11, 15, 57, -1, -7, 63, 5, 11, -13, -20, 0, -10, -7, 7, 1, 22, 23, 9, -3, -4, -3, 32, -5, 19, -12, 7, 51, -2, -41, 3, 22, 5, -54, 10, 26, -45, 2, -15, -38, 8, -11, -7, 4, 9, 33, -8, -5, 9, 5, -4, -19, 4, -10, 4, 4, -21, 2, 10, 10, 1, -1, 25, 0, 3, -23, -1, -26, -16, -50, -5, -3, 15, -26, -5, -23, 1, -27, -9, -5, -8, -23, 0, -34, 5, -12, -26, -7, 11, 28, -15, -34, 33, -35, 0, 0, -43, -2, -40, -7, -21, 4, -3, -34, -35, -23, 23, 6, -45, 12, -5, 13, -12, 1, 16, -8, -3, -28, -18, 27, 8, 41, -22, -13, 12, -42, -9, 11, -3, -21, -47, -9, -65, -1, 18, 3, -23, -10, -14, 4, 17, -3, 0, 6, 15, 6, -27, -5, -5, -51, -23, -39, -17, 24, -62, -19, 8, -12, 34, -27, 7, -8, 21, -1, 10, -11, -8, -71, -4, -38, 16, 0, 10, 30, -52, -16, 31, 32, -7, -7, 34, -6, 3, -2, 15, -64, 19, -27, -7, 5, -31, -11, 4, 8, 0, -26, 21, 29, 1, -16, -15, 15, -18, 4, -3, -21, 23, 2, -52, -8, 22, -3, 10, 4, 17, -17, -44, -2, 14, 8, -76, -84, -4, 0, -14, 18, -29, 6, 28, -13, -47, 7, -19, -16, -6, 38, -29, 11, 0, 32, -7, 0, 32, -7, -2, 7, 35, 15, 13, -25, -47, -18, -65, 1, -4, -4, -3, -59, -11, -35, -55, 7, 5, -1, -62, -20, -7, -38, 6, -4, -55, 4, -1, 8, -24, 2, 5, -16, -56, 4, -25, 20, -67, -29, 14, 0, 12, -30, 2, 11, 31, -42, 20, 7, 30, -25, -3, 6, -1, 29, 2, -1, 20, -1, -24, 2, 2, -18, 27, 0, -7, 6, 10, -43, 11, 33, 6, 5, 26, 13, -9, 13, -5, -1, -51, -35, 4, 9, -4, 10, 1, -15, 7, 22, 22, 9, -1, -20, -10, 5, -1, -1, 7, -33, 38, -8, -9, 11, 15, -25, 3, -22, 50, -17, -59, -4, -4, -27, -33, 27, -3, -24, 21, 16, -1, 21, 5, -6, -49, -14, -27, -10, -5, 15, 11, 12, 2, 23, -9, -4, 23, -15, -2, -1, -2, -4, 7, -51, -40, 6, 24, 6, 37, -11, -38, -43, -7, -2, -52, 3, -14, -8, 3, -4, 2, 43, 23, 6, -21, 4, 42, 6, -3, -27, 6, -4, 7, -12, 12, -38, -53, -10, 7, -1, -5, -5, -7, -2, -2, 8, 10, -5, -39, 49, 2, 1, 35, 2, -6, -6, 19, -20, 2, -24, -1, -3, 11, 10, -6, 1, 0, -21, -57, -55, -7, -18, -2, -5, 28, -4, 1, 0, 27, 41, 38, -2, 14, 10, 9, -3, 39, -4, 7, -32, -51, -12, -38, -63, 4, -104, -4, -11, -31, 7, 9, 17, -29, 32, 36, -4, -15, 36, -8, 39, -3, -24, -63, 13, -77, -12, -7, -5, 18, 16, -31, 13, 36, -11, -22, 20, -7, 9, -2, -75, -20, 14, -34, -4, 25, -2, -9, 0, -101, -19, -22, 5, 3, 6, 9, -19, 10, -4, 3, 43, 16, -13, 17, -17, 10, 22, 1, -44, -7, 40, 10, 9, 34, -54, -34, -35, 18, 35, -5, 32, -58, 10, -21, 1, 38, -20, -3, 53, 8, 21, 40, -3, 4, 1, 0, 12, 3, -68, 0, 7, -4, 19, -2, 22, 7, -65, -24, -30, -2, 34, 5, -42, 16, -7, 18, 4, -1, -17, 29, -41, -30, 11, 3, -7, -13, -12, 4, -34, -25, -17, 3, -28, -7, -9, 14, -10, -30, -1, -9, -22, -4, 16, -5, -17, -37, 18, -17, 27, 8, -17, -52, 3, -53, -4, -10, -34, -20, 26, -61, 26, 48, -5, 20, 11, -5, 14, -4, -17, 4, -24, 41, 3, 35, -4, 27, -29, -83, 7, -5, 3, 0, 0, 0, 11, 23, 1, -3, 68, 34, -14, -13, -5, 11, 17, -6, -20, -6, -24, 2, 6, 7, 5, -74, 11, 39, 15, -6, 22, -42, -15, -9, 7, 32, -14, -29, 12, -5, 2, 9, -2, 3, -6, -26, 0, 10, -67, -9, -8, 29, 13, 1, 7, -4, -60, -19, -23, -6, 5, 3, 28, 29, -35, 10, -4, -56, -56, -32, -34, -52, 6, -2, -5, -5, -6, 5, -55, -17, -33, -17, -4, 0, -11, 16, -40, -18, -3, -15, 0, 26, 14, 2, -34, 15, 34, -40, 23, 4, -41, -11, -11, 33, -5, -5, -31, 12, 5, -27, 16, -3, -12, 40, 18, -9, 0, 0, -12, 4, 18, 2, -5, 47, -3, 59, -11, -53, 12, -4, -4, -8, -7, 4, 6, 15, 4, -1, 44, 47, 8, -23, 5, 13, 6, -24, -43, 27, -55, 4, -13, 11, 41, -73, 13, -38, 16, 0, -48, -18, -28, 0, 19, -11, -1, -15, 17, 3, 25, 4, 4, 2, -7, 6, -2, 6, 7, -3, 4, 10, -8, 6, 0, 2, -27, -22, 0, 2, 12, -16, 18, 1, -20, 33, -23, 31, 20, 15, -10, -17, 17, 2, 5, 1, -37, -36, -19, -17, -36, -20, -42, -2, 5, -17, -22, -36, 8, 10, 16, -17, 8, 12, -20, 19, 17, -60, 5, 2, -29, -11, 7, 14, 6, -4, -39, 31, 8, -60, 25, 1, -28, 16, 11, -2, 13, -5, -2, -3, 33, -4, 0, 37, -8, 40, -23, -62, -5, 14, -3, -24, -1, 1, -10, 3, 3, 3, -7, -18, 0, -9, 20, -2, 0, 7, -28, 11, -27, 4, -3, 25, 48, -68, 16, -30, -24, -7, -53, -26, 21, 32, 12, 3, -7, 16, 32, -2, 49, 20, 0, 1, 0, -47, -61, 25, -13, -5, 0, 9, 0, 4, 18, 5, 3, 8, 4, 1, 13, 9, 12, -28, 1, 19, -37, 58, 43, 12, -12, -8, -42, 4, 5, -8, -81, 9, -29, -20, 2, -11, -81, 2, -13, 38, -8, -37, 0, 5, -32, -31, -1, -41, -16, 3, 13, -24, -4, -3, 12, -60, 4, -24, -19, -4, -74, 28, 36, 0, -17, -53, -21, -13, -15, 4, 9, -1, -59, -2, -74, -25, -4, 5, 3, -51, -22, -85, 7, -2, -6, 4, 5, 16, -2, 15, -4, -1, 18, -25, -98, 4, 26, 0, -11, -7, 20, 39, 7, -5, 5, 45, -37, -25, 21, 19, -87, 2, -29, -9, 12, -20, 46, -63, -13, 32, 21, -8, 11, -6, -16, -5, 6, -39, -61, 19, 21, 1, 6, 16, -4, -6, 13, -3, -49, -16, 22, 5, 7, -2, 36, -46, 9, -38, -34, -11, -7, -34, 17, -24, -9, -1, 8, 20, -33, -6, -12, 10, -10, -3, -3, -2, -2, -30, -11, 6, -15, 6, -13, 4, 11, -31, 22, 4, 26, -8, -17, -4, 1, 9, -5, 21, -19, -3, 22, 0, 12, -52, 3, 1, 3, -54, -4, -4, -29, -3, -2, -28, -19, -27, -7, -13, -8, -30, -14, -19, -30, 16, -4, -17, -7, -34, 6, 10, 0, -2, -63, 15, -13, -48, 2, -36, 2, 13, 30, 3, 0, -6, -12, 2, -56, -47, 9, -11, -13, -8, -41, 5, -13, 10, 11, -26, -5, 10, 40, 4, -35, -7, -10, -3, -2, -19, -38, 28, -25, 2, 7, 9, -3, -2, 23, 13, -66, -46, -27, -1, 3, -26, 54, -20, 2, -30, -11, 2, 12, -27, -10, -1, -28, 5, -10, 14, -41, -28, -1, -11, -19, 30, -34, 4, -37, 9, -18, -47, 1, 1, -17, -7, 30, -19, -20, -8, 18, -27, 33, 0, 30, 14, -12, 2, 10, -4, -52, -12, 1, -43, 38, -17, -24, 4, -14, -18, 11, 0, -1, -5, -29, -41, 3, 0, -2, 15, -17, -60, -39, 20, -4, 40, -7, 11, -14, -8, -1, -9, -25, 30, 4, -28, 31, -3, -35, 12, -4, 40, -61, -4, -4, 37, -2, -10, -22, 6, 0, 2, -22, 41, -29, 7, 3, -53, -8, -2, 62, 0, -34, -18, -3, -1, 8, 5, -17, 14, -31, -1, -5, 20, -7, -4, -1, 6, -31, -26, -16, -2, -22, 0, 12, 8, 9, -14, -9, 36, 6, -15, -18, 42, -45, 0, 2, 8, 15, -22, 8, -24, -20, 16, -129, -3, -17, 3, -3, -17, -6, 4, -17, 22, 23, -21, 0, -3, -9, -17, 23, 0, -14, -9, 8, -44, 16, -9, -10, -14, -2, -37, -9, 37, -22, 17, -14, -5, 3, -5, 2, -18, -51, -45, 4, -9, -4, 5, 4, -50, -11, 6, -5, 7, -6, -5, -33, 8, 1, -7, -39, 44, -2, -33, 5, 22, -59, 42, 15, -20, -20, -6, 0, 48, 12, 12, -4, -8, 3, -6, 12, 5, -27, -4, -1, 6, 1, -4, 26, 7, 8, -17, 0, 4, 2, -11, -11, 19, -26, -5, 4, -3, 8, -7, 9, -3, -22, -23, -3, 3, -18, 16, 17, -17, -4, -1, -10, -17, 11, -2, 31, 37, -21, 1, 0, 15, 17, -58, -10, 8, -11, 0, -91, -3, 36, 6, 3, 12, -6, -2, -20, 28, 13, -18, -26, 12, 16, -10, 20, -3, 4, -13, 17, -24, 0, -2, 24, 4, 28, -31, -15, 41, -18, -2, -4, 5, -9, 3, -3, -26, -5, -6, -4, -11, 4, 36, 0, -74, 21, 0, 0, 7, -9, 8, 2, 5, 4, 4, -35, 73, 1, 0, -10, 2, -25, 15, -12, -30, 21, 4, 16, 8, -16, -20, 10, -6, -2, 4, -2, 17, 7, -28, 6, -29, 0, 10, -1, -9, -14, -2, -13, 6, -4, -20, -10, 28, 0, 0, 5, -10, -1, 1, 15, -7, -40, -1, -1, -3, 2, 17, 14, -26, -13, -7, -11, -1, -8, 26, -11, -12, 32, 8, -3, 5, -5, 3, -24, -27, -26, -7, -69, 3, 25, 28, -37, 18, -3, 7, -27, 36, 35, -2, -11, 5, -25, -2, -8, -5, -23, 11, -14, 0, 3, -5, 34, -6, 16, -76, -13, 34, -24, -10, 23, -3, -8, -5, -6, -34, -29, 7, 1, -5, 4, 21, -16, -102, -8, -16, -5, 0, -4, -13, -16, 31, 7, -7, -7, 65, -20, -39, 25, 34, -11, 18, -7, -1, 16, 1, -35, -2, 3, 1, 8, 4, -8, -8, -69, 12, -12, 14, 20, -61, 2, -21, -6, -4, -19, -23, -21, -9, 1, -36, -42, 39, -13, -3, -6, 12, 18, -8, -7, 0, -48, -10, -22, 5, 10, -15, 22, 2, 8, -6, -1, 12, 0, -6, -27, 31, 14, -3, -4, 25, 8, 19, -4, -25, -11, -5, -67, 4, -42, -8, -16, 13, 8, 7, -8, 38, 38, -41, -14, 2, 16, -12, 13, 0, -3, 22, 12, -39, 25, 4, -29, 0, 6, -28, 3, 56, -12, -11, -9, 0, 27, 6, 25, -31, 0, -28, 4, 0, -3, 27, 2, -24, -17, 7, -1, 21, 0, 36, -33, -17, 3, 4, 23, 39, -15, -35, 37, 22, -24, 14, 1, -13, -19, -4, 9, 42, 30, -62, -2, -15, -37, 0, -34, 0, -29, 16, 8, -25, 9, 14, 46, 7, 25, -9, 0, 0, 0, -29, -39, 26, -12, -7, -6, 4, 13, 3, 15, -8, -23, 16, 28, -1, 15, -20, 46, -24, 52, -17, -21, 10, 12, 5, -21, 23, -49, 0, 2, 28, -3, -1, -34, -11, -12, 28, -40, -2, 16, 22, 22, 6, 0, 26, -40, 25, 25, -73, 7, -22, 25, -17, 13, -5, 18, -2, -40, -72, -11, 1, -28, 13, 51, -21, 6, 34, -24, -31, -27, 6, 10, 0, -12, -61, -50, -50, 3, -2, 2, -13, -17, -47, -7, 0, 3, -15, -7, 0, -30, 33, -7, -6, -9, 13, -39, -5, 25, -11, -13, 16, 35, 4, -8, -6, 22, 11, -2, -35, 19, 9, -55, 1, 44, 8, -32, 7, 11, 31, -24, 37, -23, 7, -29, -9, -8, -1, -6, -15, 26, 15, -15, -6, -2, 2, -11, 1, 29, 0, -43, 10, 26, 6, 49, 16, 33, -73, -14, -13, -2, -54, -6, 0, -29, -72, 6, 3, 0, 8, -3, -19, 1, 19, -17, 59, 44, 2, -25, 14, 10, 24, -2, -26, -46, 60, 6, -26, 37, 3, -38, 43, -8, 1, -3, 30, 26, 21, -7, 2, 18, -7, -31, 0, -58, 53, 5, -45, 4, 15, -54, -6, 17, -39, 10, -6, 6, -10, -2, -21, -10, 6, -1, 5, -5, -67, 6, -20, 8, -6, 0, -4, -107, 67, -45, -75, 35, -2, -14, 2, 39, 16, -23, 0, -23, 12, 15, -32, -4, -34, -38, 4, 30, -20, -34, 28, 40, -7, -9, 7, -13, 8, -36, -35, 0, -4, 0, 7, -8, 68, -7, 0, 4, 29, -26, 5, -2, 6, -19, -27, -4, -6, -9, -33, 36, 1, 5, -26, -17, 3, 0, 33, -13, -8, -7, 3, -4, 23, -6, -43, 8, 5, -82, 13, 0, -2, -19, -20, -36, 0, 7, 2, -34, 62, 55, -5, 0, 21, 46, -10, 18, 2, 0, 20, -28, 19, 25, -7, -48, -5, -13, 9, 23, 34, -9, -16, -3, -2, 12, 2, 7, -48, 7, -6, -3, 41, 6, 7, -19, -42, -42, 4, 3, -80, 1, -16, -21, 1, -1, -6, -25, 89, 9, -48, 34, 36, 2, 30, -9, -8, -36, -6, 26, 29, 15, -3, 27, -22, -11, -4, 0, 17, -31, -4, 20, -28, -4, 16, -36, -4, -28, -24, 0, -6, 3, -16, -40, 21, 3, 3, 1, -15, -13, 4, 10, -3, 10, -11, 14, 0, -54, -31, 25, -26, -16, -38, 6, 23, 26, 31, -29, 27, -14, -1, -6, 12, 35, -13, 21, -39, -59, -17, -35, -6, 0, -4, -48, -7, 0, 29, 22, 47, 54, -47, -4, 20, 34, -22, 39, 5, -16, 28, -10, -22, 5, 0, 57, -10, -19, 19, 43, 48, -51, -5, -13, -4, 6, 6, -45, -22, -11, -24, 3, 11, 5, -16, 1, -66, -2, 0, -1, 10, -7, -12, -31, -2, 0, 6, -28, 65, -13, -37, 0, 46, -49, 38, 0, 14, -40, -1, 39, 21, 11, -10, -11, 4, -20, 4, 25, -8, -57, 0, 22, 2, -2, 19, -73, -8, -37, -23, 0, -4, -2, 11, -13, 11, 35, -1, 3, 9, -11, 5, -6, 7, -5, 14, 21, 3, -53, -35, 29, -15, -6, -77, -7, 13, 11, 46, -26, 4, -6, -2, -2, 3, 30, 45, -6, 34, 5, 28, 9, -6, 19, 2, -24, -4, 4, 15, -1, 46, 43, -13, 4, 19, -6, 0, 1, -5, -13, 23, 1, 1, 1, -8, 10, 2, -38, 10, -18, 42, -9, 4, -21, -17, -32, -2, 2, -34, 7, -2, -6, -29, -8, 0, -3, -36, -4, -13, 0, -53, 7, -15, -20, -3, -6, -1, -20, 54, -39, -6, -37, 52, -14, 37, 4, 11, -15, 6, 27, 15, 6, -49, 1, -26, -29, -3, -17, 30, 3, -19, -1, 20, -1, 13, -17, -3, -49, -11, 0, 1, -6, 2, -4, 31, 10, 6, 9, 23, 4, -3, -14, 3, -18, -45, -8, 3, -3, -11, 27, -25, 7, -22, 0, 19, 13, 61, -5, 24, 2, 5, 0, 29, 9, 21, 0, 34, 3, 15, 13, -4, 7, 28, -40, -4, -1, 32, -34, 69, 50, 26, 9, 5, 47, 15, 38, -4, 13, 22, -3, 28, 25, -7, 25, -13, -49, 1, -1, 53, -14, -15, -2, 15, -30, -7, 5, -14, 22, -15, 5, 0, 0, 0, 1, -52, -8, -17, -2, -33, 1, -6, -28, -6, -3, -7, 1, 73, -2, -11, 2, 65, -10, 32, 9, -1, -67, 1, 43, 36, 30, -32, -1, 0, -37, 6, 4, 5, -11, -13, 23, 17, 4, 18, 1, -14, -27, -14, -4, -2, 3, -2, -5, 36, 57, -7, 0, 2, 7, -5, -16, -6, -15, -8, -5, 4, -9, -22, 23, -28, 10, -44, 16, 14, 69, 60, 4, 9, 24, -8, 0, 20, 15, 69, -16, -23, -35, -35, 30, 0, -37, 12, -46, -21, 2, 24, -27, 51, 43, -32, -26, 20, 44, -11, 47, -5, 13, 19, -25, -42, 20, -8, -24, -4, -22, -38, 11, 44, -41, -35, 36, 0, -9, -4, -9, -9, 4, 9, 7, 0, -5, 26, -14, -42, -14, -2, -6, -16, -2, -17, -17, -18, 0, 6, -8, 58, 7, -17, -3, 53, -38, 50, -15, 1, -13, -5, 22, 60, 29, -1, -1, 6, -50, 0, 24, 22, -12, 5, 35, 31, -2, 37, -47, -5, 3, 12, -3, -4, 0, -32, -1, -22, 6, -2, 8, -50, 0, 5, 2, 0, 0, 2, -31, 2, 6, 6, 28, -30, -6, -45, 15, 8, 26, 17, 6, -20, 3, 0, -5, 11, 11, -13, -46, -50, 8, -9, 3, -9, -4, 14, 6, 3, 6, 36, -30, 30, 24, -23, 8, 5, 0, 11, 12, 6, -15, -17, -18, -85, 12, -1, 40, 9, 40, 0, 3, 61, -22, -34, -8, 6, -39, -1, -13, -52, -4, -11, 0, -18, -4, -37, -16, -37, -18, -23, 3, 14, 2, -11, -21, 12, -4, -3, -104, 44, -49, 6, -40, 34, -9, 11, 30, -40, -29, -4, 24, 30, 0, -22, 11, 36,

    others => 0);
end iwght_package;
