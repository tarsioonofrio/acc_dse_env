library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 13, 
    53, 0, 0, 0, 0, 13, 0, 
    39, 0, 0, 0, 0, 39, 0, 
    0, 14, 76, 12, 19, 70, 1, 
    101, 5, 230, 164, 194, 193, 206, 
    244, 99, 255, 206, 215, 242, 257, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 
    81, 0, 0, 0, 0, 0, 0, 
    0, 16, 0, 0, 0, 12, 0, 
    0, 82, 0, 0, 0, 0, 0, 
    0, 0, 131, 0, 0, 0, 0, 
    0, 0, 65, 0, 0, 0, 0, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    0, 0, 0, 0, 0, 0, 0, 
    75, 0, 42, 0, 0, 0, 0, 
    116, 0, 0, 49, 51, 21, 0, 
    174, 74, 0, 0, 0, 0, 0, 
    118, 166, 143, 48, 23, 0, 0, 
    68, 117, 0, 0, 0, 3, 70, 
    124, 35, 13, 13, 11, 24, 63, 
    
    -- channel=6
    63, 22, 56, 104, 14, 45, 63, 
    103, 30, 64, 51, 0, 27, 62, 
    136, 43, 0, 55, 10, 58, 0, 
    180, 80, 63, 42, 0, 82, 1, 
    49, 99, 135, 75, 150, 98, 76, 
    95, 116, 235, 103, 0, 0, 42, 
    84, 213, 85, 0, 0, 0, 17, 
    
    -- channel=7
    14, 22, 0, 0, 0, 0, 0, 
    8, 66, 45, 0, 0, 0, 0, 
    50, 40, 36, 20, 0, 22, 0, 
    67, 0, 0, 25, 4, 0, 0, 
    54, 78, 108, 36, 4, 38, 48, 
    107, 45, 55, 40, 54, 32, 75, 
    80, 37, 32, 22, 22, 43, 32, 
    
    -- channel=8
    71, 52, 67, 89, 14, 0, 60, 
    0, 0, 0, 0, 0, 0, 39, 
    1, 129, 35, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 48, 0, 
    0, 0, 0, 0, 63, 28, 0, 
    0, 0, 210, 62, 0, 0, 0, 
    36, 84, 51, 0, 0, 0, 11, 
    
    -- channel=9
    97, 188, 95, 45, 99, 132, 99, 
    159, 210, 119, 71, 104, 98, 79, 
    113, 17, 52, 132, 130, 94, 121, 
    152, 139, 8, 18, 52, 0, 90, 
    118, 152, 122, 83, 0, 0, 94, 
    0, 0, 0, 0, 67, 121, 80, 
    59, 0, 0, 85, 108, 100, 85, 
    
    -- channel=10
    186, 168, 104, 126, 111, 61, 190, 
    50, 120, 55, 14, 88, 0, 90, 
    0, 153, 89, 0, 30, 0, 16, 
    0, 51, 63, 3, 54, 15, 103, 
    0, 0, 0, 0, 4, 134, 130, 
    130, 0, 0, 79, 59, 20, 36, 
    113, 30, 91, 26, 25, 45, 0, 
    
    -- channel=11
    150, 170, 179, 132, 64, 72, 97, 
    50, 112, 116, 108, 40, 98, 56, 
    0, 83, 29, 107, 0, 65, 78, 
    0, 62, 51, 103, 19, 81, 104, 
    0, 0, 0, 0, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=12
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 38, 0, 
    24, 0, 0, 0, 0, 33, 0, 
    108, 0, 0, 55, 17, 17, 19, 
    133, 125, 47, 0, 0, 14, 0, 
    181, 34, 21, 75, 33, 38, 97, 
    110, 141, 126, 112, 102, 133, 116, 
    
    -- channel=13
    326, 294, 325, 235, 157, 72, 164, 
    0, 247, 156, 0, 19, 0, 0, 
    0, 199, 176, 0, 0, 0, 0, 
    0, 0, 163, 0, 26, 2, 3, 
    0, 0, 0, 89, 59, 0, 146, 
    2, 95, 0, 0, 0, 0, 0, 
    0, 33, 0, 0, 0, 0, 0, 
    
    -- channel=14
    0, 39, 0, 0, 0, 0, 0, 
    0, 55, 0, 0, 33, 22, 0, 
    0, 0, 0, 35, 28, 0, 78, 
    76, 0, 0, 0, 0, 0, 45, 
    134, 60, 0, 115, 0, 0, 36, 
    2, 6, 0, 0, 80, 226, 202, 
    86, 0, 0, 170, 209, 204, 222, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 37, 
    0, 0, 0, 0, 0, 12, 0, 
    77, 0, 0, 92, 122, 194, 190, 
    253, 73, 161, 215, 235, 262, 272, 
    
    -- channel=16
    0, 0, 0, 6, 1, 0, 28, 
    0, 0, 0, 0, 0, 0, 36, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 37, 0, 0, 0, 
    0, 0, 0, 0, 0, 44, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=17
    0, 9, 0, 52, 38, 62, 32, 
    88, 57, 38, 111, 90, 86, 92, 
    79, 131, 33, 106, 117, 126, 43, 
    94, 147, 66, 50, 91, 83, 28, 
    5, 104, 101, 9, 45, 0, 1, 
    0, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 11, 0, 
    109, 0, 8, 193, 289, 393, 370, 
    351, 143, 328, 393, 433, 459, 488, 
    
    -- channel=19
    16, 29, 107, 37, 112, 89, 46, 
    109, 87, 126, 104, 36, 28, 19, 
    131, 45, 190, 115, 92, 61, 89, 
    141, 94, 3, 8, 0, 41, 21, 
    41, 185, 169, 130, 75, 122, 107, 
    146, 178, 296, 141, 193, 166, 145, 
    54, 121, 92, 40, 54, 48, 55, 
    
    -- channel=20
    64, 25, 50, 58, 0, 0, 11, 
    0, 0, 0, 3, 0, 0, 4, 
    27, 109, 0, 0, 0, 9, 0, 
    0, 16, 102, 23, 40, 78, 0, 
    0, 0, 0, 0, 51, 0, 0, 
    0, 37, 117, 0, 0, 0, 0, 
    13, 91, 9, 0, 0, 0, 0, 
    
    -- channel=21
    51, 68, 63, 5, 74, 49, 32, 
    14, 45, 42, 86, 55, 49, 61, 
    0, 0, 0, 34, 6, 40, 107, 
    0, 31, 52, 20, 0, 52, 48, 
    0, 0, 77, 93, 90, 167, 88, 
    25, 2, 1, 47, 163, 191, 190, 
    106, 44, 129, 137, 170, 164, 170, 
    
    -- channel=22
    51, 89, 72, 106, 96, 86, 73, 
    64, 82, 57, 100, 23, 58, 87, 
    0, 79, 0, 16, 0, 46, 64, 
    0, 38, 7, 15, 6, 25, 30, 
    0, 0, 63, 0, 72, 70, 24, 
    0, 0, 64, 0, 13, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=23
    0, 0, 0, 0, 101, 29, 0, 
    137, 73, 33, 0, 121, 0, 0, 
    0, 65, 0, 0, 219, 0, 8, 
    0, 105, 48, 0, 35, 0, 0, 
    0, 126, 53, 30, 0, 76, 52, 
    0, 135, 0, 0, 96, 136, 78, 
    3, 0, 4, 0, 55, 10, 49, 
    
    -- channel=24
    73, 61, 17, 0, 19, 0, 43, 
    12, 60, 0, 0, 55, 0, 7, 
    0, 26, 120, 0, 88, 0, 5, 
    0, 26, 3, 0, 35, 0, 71, 
    0, 24, 0, 0, 0, 7, 0, 
    20, 0, 0, 0, 15, 10, 0, 
    37, 0, 40, 27, 40, 36, 4, 
    
    -- channel=25
    270, 254, 279, 297, 192, 164, 266, 
    277, 255, 168, 90, 27, 25, 147, 
    135, 210, 111, 11, 69, 0, 14, 
    0, 128, 95, 54, 85, 14, 41, 
    0, 49, 22, 0, 0, 0, 71, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    98, 85, 109, 85, 50, 59, 15, 
    54, 105, 153, 98, 14, 34, 55, 
    4, 159, 18, 59, 22, 19, 24, 
    0, 0, 0, 0, 30, 77, 7, 
    0, 92, 140, 78, 19, 111, 59, 
    0, 128, 94, 77, 131, 135, 139, 
    94, 50, 131, 98, 103, 94, 109, 
    
    -- channel=27
    21, 41, 91, 17, 58, 2, 36, 
    29, 66, 29, 0, 135, 0, 12, 
    86, 100, 146, 0, 174, 0, 31, 
    20, 29, 234, 0, 151, 0, 69, 
    122, 48, 0, 99, 21, 6, 83, 
    131, 341, 0, 69, 36, 89, 62, 
    38, 189, 74, 36, 87, 75, 121, 
    
    -- channel=28
    0, 0, 0, 25, 0, 70, 19, 
    152, 0, 2, 143, 0, 107, 134, 
    88, 68, 0, 159, 0, 279, 38, 
    105, 203, 0, 142, 0, 188, 0, 
    0, 105, 193, 0, 16, 149, 0, 
    0, 0, 319, 0, 87, 0, 0, 
    69, 0, 96, 25, 0, 0, 0, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 9, 0, 0, 
    27, 19, 4, 0, 0, 0, 0, 
    24, 44, 75, 12, 55, 94, 84, 
    135, 43, 118, 127, 150, 160, 171, 
    
    -- channel=30
    298, 341, 278, 176, 209, 80, 145, 
    30, 285, 177, 0, 0, 0, 0, 
    0, 41, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 48, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    0, 23, 31, 17, 22, 30, 22, 
    46, 0, 41, 97, 52, 85, 62, 
    110, 98, 89, 94, 75, 93, 38, 
    56, 90, 82, 115, 157, 90, 56, 
    60, 20, 36, 40, 0, 0, 21, 
    0, 112, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end ifmap_package;
