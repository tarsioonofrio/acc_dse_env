library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    500, 500, 497, 498, 503, 503, 502, 507, 507, 497, 485, 495, 516, 532, 536, 537, 522, 507, 489, 477, 472, 473, 479, 482, 481, 491, 502, 516, 517, 510, 
    515, 516, 509, 502, 505, 502, 504, 507, 502, 464, 445, 469, 505, 527, 527, 517, 505, 473, 439, 412, 407, 426, 448, 464, 473, 483, 494, 510, 514, 509, 
    516, 518, 519, 515, 511, 507, 508, 510, 497, 409, 381, 402, 465, 494, 495, 497, 475, 414, 369, 320, 310, 322, 364, 395, 421, 456, 479, 492, 503, 505, 
    497, 497, 505, 514, 514, 515, 514, 517, 508, 434, 397, 370, 439, 479, 469, 449, 418, 369, 298, 235, 221, 244, 282, 313, 374, 415, 453, 466, 480, 490, 
    469, 476, 496, 507, 516, 519, 520, 523, 518, 457, 398, 378, 403, 411, 400, 407, 381, 313, 231, 187, 193, 215, 234, 275, 311, 368, 424, 448, 466, 480, 
    402, 409, 466, 497, 515, 526, 525, 520, 515, 492, 435, 379, 362, 355, 347, 345, 327, 280, 219, 183, 200, 235, 259, 273, 300, 354, 397, 429, 455, 470, 
    322, 334, 388, 443, 496, 520, 508, 480, 475, 451, 396, 332, 295, 293, 303, 304, 301, 293, 251, 215, 219, 263, 293, 295, 308, 334, 390, 424, 447, 464, 
    209, 228, 294, 358, 459, 506, 443, 348, 301, 293, 293, 262, 231, 255, 279, 295, 312, 319, 270, 240, 222, 249, 285, 306, 313, 321, 361, 416, 448, 464, 
    134, 135, 185, 295, 421, 491, 380, 247, 150, 168, 175, 191, 190, 233, 278, 296, 324, 328, 278, 226, 181, 227, 273, 290, 299, 306, 342, 393, 430, 459, 
    82, 98, 108, 245, 389, 475, 384, 218, 74, 82, 124, 148, 168, 217, 270, 279, 339, 312, 242, 182, 139, 211, 253, 286, 286, 280, 305, 354, 396, 437, 
    71, 74, 87, 221, 377, 471, 418, 231, 140, 124, 150, 132, 145, 184, 243, 259, 310, 272, 210, 133, 117, 203, 253, 286, 282, 285, 283, 312, 344, 409, 
    61, 66, 96, 214, 377, 467, 468, 320, 235, 166, 167, 121, 108, 145, 213, 241, 286, 231, 173, 98, 127, 212, 269, 297, 293, 282, 267, 278, 304, 379, 
    56, 68, 85, 193, 368, 457, 483, 382, 296, 195, 175, 107, 104, 126, 179, 215, 263, 214, 152, 101, 129, 201, 252, 276, 280, 268, 253, 255, 294, 369, 
    43, 58, 65, 176, 312, 408, 448, 383, 309, 173, 95, 50, 72, 138, 194, 223, 252, 225, 171, 113, 144, 222, 267, 278, 279, 257, 245, 270, 314, 384, 
    25, 36, 33, 140, 225, 324, 365, 387, 318, 190, 113, 84, 110, 189, 214, 239, 282, 256, 215, 162, 165, 195, 253, 279, 276, 262, 270, 312, 361, 424, 
    0, 6, 5, 96, 167, 237, 264, 324, 295, 250, 146, 148, 209, 234, 259, 257, 272, 296, 326, 256, 226, 245, 292, 318, 310, 290, 300, 344, 403, 442, 
    0, 0, 0, 51, 128, 169, 200, 242, 282, 291, 232, 240, 255, 248, 262, 245, 261, 295, 298, 291, 302, 290, 319, 347, 345, 333, 352, 385, 431, 451, 
    0, 0, 0, 23, 116, 150, 176, 184, 217, 274, 275, 306, 257, 219, 208, 211, 241, 275, 282, 305, 304, 326, 368, 346, 354, 350, 387, 410, 437, 459, 
    0, 0, 0, 16, 97, 122, 115, 128, 194, 279, 279, 287, 202, 157, 136, 161, 227, 293, 308, 318, 325, 362, 372, 340, 342, 352, 400, 424, 444, 460, 
    33, 0, 5, 35, 107, 116, 60, 14, 42, 153, 197, 167, 115, 64, 41, 100, 179, 262, 309, 314, 316, 313, 290, 266, 251, 281, 320, 343, 356, 365, 
    28, 0, 10, 41, 93, 72, 11, 0, 0, 31, 115, 113, 71, 33, 37, 91, 160, 236, 263, 270, 253, 234, 206, 175, 162, 168, 177, 199, 203, 204, 
    11, 0, 0, 16, 56, 27, 0, 0, 0, 8, 59, 92, 77, 69, 77, 93, 120, 173, 197, 185, 158, 136, 113, 91, 73, 64, 64, 71, 70, 72, 
    7, 0, 0, 17, 35, 0, 0, 0, 0, 0, 75, 103, 100, 105, 105, 110, 117, 128, 124, 106, 91, 80, 63, 43, 30, 21, 18, 23, 26, 22, 
    0, 14, 13, 24, 0, 0, 0, 0, 0, 64, 101, 110, 111, 117, 120, 113, 106, 102, 91, 74, 59, 50, 35, 16, 10, 8, 9, 7, 0, 0, 
    0, 29, 43, 50, 0, 0, 0, 0, 32, 88, 79, 84, 88, 94, 101, 104, 99, 92, 81, 60, 38, 21, 11, 9, 7, 12, 0, 0, 0, 0, 
    0, 21, 49, 60, 0, 0, 0, 0, 73, 84, 70, 71, 79, 94, 98, 97, 89, 79, 62, 45, 27, 9, 0, 0, 3, 1, 0, 0, 0, 0, 
    0, 3, 33, 52, 11, 0, 0, 16, 89, 76, 57, 62, 65, 81, 92, 92, 80, 63, 47, 32, 13, 2, 2, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 32, 33, 6, 38, 53, 109, 94, 73, 61, 55, 66, 70, 70, 59, 48, 35, 25, 23, 20, 17, 4, 0, 0, 0, 0, 0, 24, 
    0, 0, 3, 15, 43, 44, 73, 103, 116, 108, 98, 86, 77, 75, 73, 70, 52, 26, 13, 16, 26, 33, 28, 4, 0, 0, 0, 0, 3, 55, 
    0, 3, 15, 18, 45, 75, 94, 119, 126, 124, 117, 102, 103, 110, 111, 95, 62, 29, 14, 16, 29, 50, 41, 7, 0, 0, 0, 0, 6, 64, 
    
    
    others => 0);
end gold_package;
