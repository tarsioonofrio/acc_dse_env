library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 5, 0, 0, 2, 84, 0, 0, 0, 27, 2, 0, 2, 5, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 7, 74, 0, 0, 0, 0, 28, 
    0, 117, 0, 9, 1, 12, 13, 0, 0, 49, 0, 0, 0, 0, 54, 
    0, 84, 0, 40, 52, 0, 0, 0, 0, 88, 0, 0, 10, 0, 6, 
    0, 31, 0, 0, 66, 0, 0, 0, 0, 217, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 68, 77, 0, 0, 0, 168, 0, 0, 4, 27, 0, 
    0, 0, 0, 0, 22, 81, 0, 0, 0, 98, 0, 0, 17, 0, 0, 
    0, 0, 0, 56, 0, 0, 0, 18, 23, 0, 18, 0, 6, 29, 18, 
    0, 0, 0, 71, 0, 0, 26, 14, 0, 0, 0, 0, 52, 55, 0, 
    97, 0, 0, 203, 0, 0, 43, 0, 0, 0, 23, 36, 16, 5, 0, 
    29, 14, 0, 146, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 31, 56, 0, 0, 0, 0, 0, 0, 4, 9, 13, 0, 0, 21, 
    0, 0, 79, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 5, 0, 0, 56, 0, 0, 
    
    -- channel=1
    164, 171, 171, 172, 168, 172, 174, 171, 163, 149, 131, 139, 147, 138, 122, 
    164, 171, 176, 175, 183, 273, 179, 158, 112, 149, 148, 116, 111, 132, 134, 
    120, 154, 173, 172, 174, 238, 142, 94, 84, 228, 205, 174, 116, 83, 147, 
    107, 170, 180, 185, 174, 181, 204, 122, 124, 223, 209, 146, 103, 40, 133, 
    224, 305, 191, 252, 381, 291, 242, 136, 92, 191, 264, 143, 137, 76, 57, 
    244, 351, 208, 149, 348, 287, 302, 188, 102, 299, 285, 140, 155, 128, 72, 
    256, 324, 187, 128, 238, 321, 359, 247, 145, 342, 256, 146, 140, 174, 133, 
    308, 353, 196, 190, 205, 387, 271, 216, 146, 291, 248, 144, 150, 173, 147, 
    365, 394, 193, 267, 180, 210, 191, 184, 201, 199, 173, 86, 89, 158, 173, 
    386, 388, 239, 296, 207, 145, 249, 299, 177, 156, 87, 41, 125, 206, 179, 
    399, 378, 250, 432, 405, 253, 327, 332, 186, 112, 97, 126, 167, 205, 169, 
    293, 373, 328, 549, 375, 174, 178, 169, 141, 139, 156, 171, 187, 201, 185, 
    182, 252, 377, 481, 186, 166, 155, 150, 147, 154, 181, 201, 206, 205, 246, 
    185, 173, 308, 363, 165, 185, 168, 151, 157, 175, 185, 193, 185, 224, 210, 
    189, 177, 178, 206, 129, 146, 163, 168, 188, 207, 176, 178, 259, 270, 156, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 51, 0, 0, 0, 35, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 71, 0, 9, 0, 0, 19, 
    0, 30, 0, 18, 5, 0, 6, 0, 0, 39, 11, 0, 0, 0, 0, 
    17, 71, 0, 4, 156, 58, 10, 0, 0, 98, 18, 0, 12, 0, 0, 
    8, 44, 12, 0, 72, 56, 63, 0, 0, 115, 5, 0, 0, 4, 0, 
    31, 42, 0, 0, 16, 122, 24, 38, 0, 87, 15, 0, 17, 23, 0, 
    48, 89, 0, 43, 0, 57, 7, 0, 14, 0, 52, 0, 12, 4, 0, 
    82, 86, 0, 66, 9, 0, 28, 6, 8, 25, 0, 0, 0, 0, 0, 
    117, 77, 0, 128, 0, 0, 80, 78, 0, 0, 0, 0, 9, 26, 1, 
    141, 114, 34, 148, 80, 41, 59, 56, 21, 16, 19, 29, 30, 32, 26, 
    14, 115, 109, 122, 9, 20, 18, 16, 11, 14, 22, 30, 38, 41, 40, 
    20, 27, 158, 77, 7, 28, 9, 18, 23, 28, 34, 47, 28, 52, 59, 
    17, 35, 39, 67, 13, 41, 40, 21, 24, 24, 21, 27, 48, 37, 0, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 6, 13, 23, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 11, 3, 6, 3, 17, 10, 0, 
    36, 0, 0, 0, 0, 0, 5, 14, 8, 21, 6, 10, 10, 15, 0, 
    45, 5, 0, 0, 0, 15, 0, 8, 6, 4, 6, 23, 11, 20, 21, 
    58, 0, 0, 0, 0, 0, 0, 14, 11, 0, 20, 19, 15, 17, 8, 
    45, 28, 17, 0, 0, 0, 12, 4, 13, 0, 6, 16, 17, 3, 0, 
    38, 29, 37, 9, 0, 7, 8, 0, 14, 0, 0, 17, 11, 0, 0, 
    21, 24, 31, 24, 20, 17, 24, 5, 8, 1, 13, 28, 5, 0, 0, 
    19, 24, 28, 29, 30, 27, 16, 31, 40, 35, 51, 53, 48, 36, 38, 
    52, 49, 42, 0, 11, 77, 63, 67, 72, 69, 73, 77, 83, 78, 83, 
    87, 57, 59, 0, 80, 76, 73, 72, 73, 77, 83, 84, 79, 87, 96, 
    100, 88, 56, 29, 70, 75, 76, 74, 78, 81, 84, 87, 93, 95, 80, 
    97, 94, 75, 62, 68, 72, 74, 78, 74, 79, 81, 88, 90, 85, 97, 
    
    -- channel=4
    129, 134, 133, 134, 132, 128, 139, 146, 134, 114, 100, 105, 108, 117, 114, 
    128, 139, 141, 136, 136, 120, 120, 120, 89, 54, 28, 44, 70, 95, 110, 
    98, 113, 136, 138, 140, 148, 65, 53, 39, 54, 32, 30, 25, 57, 97, 
    21, 73, 124, 140, 114, 87, 57, 31, 24, 72, 32, 41, 14, 17, 92, 
    0, 63, 102, 133, 81, 73, 47, 26, 25, 51, 46, 25, 33, 15, 57, 
    3, 45, 89, 99, 84, 60, 42, 40, 16, 81, 39, 16, 41, 23, 16, 
    0, 31, 72, 101, 103, 64, 65, 32, 23, 85, 17, 15, 25, 27, 30, 
    6, 24, 32, 64, 85, 97, 46, 48, 26, 98, 27, 17, 35, 46, 65, 
    11, 31, 0, 40, 43, 55, 34, 33, 46, 62, 53, 26, 34, 65, 108, 
    32, 33, 0, 36, 25, 48, 49, 32, 39, 54, 24, 15, 41, 105, 107, 
    34, 34, 0, 68, 0, 14, 45, 32, 0, 0, 0, 0, 0, 0, 0, 
    9, 15, 16, 89, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 22, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    42, 36, 37, 37, 39, 35, 42, 42, 35, 33, 32, 38, 31, 37, 33, 
    42, 39, 38, 37, 35, 32, 27, 34, 9, 15, 10, 33, 49, 43, 38, 
    39, 49, 44, 37, 44, 58, 1, 17, 18, 33, 11, 7, 14, 54, 45, 
    0, 87, 48, 39, 32, 16, 10, 6, 21, 53, 0, 22, 2, 30, 67, 
    0, 61, 27, 17, 0, 0, 0, 1, 26, 40, 4, 0, 24, 7, 67, 
    0, 39, 16, 25, 39, 0, 0, 0, 9, 79, 0, 0, 31, 5, 14, 
    0, 25, 35, 2, 59, 18, 4, 0, 0, 81, 0, 2, 28, 19, 21, 
    0, 0, 14, 12, 28, 44, 0, 17, 1, 74, 0, 4, 30, 36, 28, 
    0, 2, 0, 27, 15, 19, 7, 19, 32, 28, 41, 2, 40, 39, 43, 
    0, 6, 0, 33, 0, 19, 12, 0, 40, 14, 0, 14, 49, 63, 33, 
    35, 4, 0, 55, 0, 0, 25, 0, 0, 0, 17, 9, 29, 29, 6, 
    72, 12, 0, 57, 0, 0, 23, 17, 4, 9, 15, 15, 10, 19, 8, 
    17, 68, 19, 23, 0, 8, 9, 14, 15, 16, 14, 17, 16, 4, 9, 
    2, 19, 82, 0, 0, 16, 5, 15, 10, 13, 15, 17, 5, 21, 22, 
    0, 12, 25, 32, 17, 29, 17, 8, 9, 9, 10, 13, 13, 6, 0, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 18, 18, 5, 0, 0, 
    0, 0, 0, 0, 0, 12, 0, 1, 5, 59, 63, 46, 28, 11, 0, 
    6, 21, 0, 0, 0, 0, 16, 20, 38, 66, 43, 41, 33, 19, 4, 
    33, 68, 0, 0, 20, 18, 44, 30, 43, 41, 49, 21, 39, 19, 15, 
    70, 104, 0, 0, 110, 38, 49, 31, 32, 78, 65, 33, 49, 34, 13, 
    57, 111, 2, 0, 51, 51, 81, 42, 35, 108, 59, 40, 47, 49, 31, 
    72, 98, 30, 0, 11, 97, 72, 68, 32, 86, 56, 48, 53, 54, 4, 
    99, 124, 59, 66, 21, 61, 41, 49, 41, 32, 57, 34, 42, 21, 0, 
    111, 122, 72, 99, 54, 27, 45, 64, 58, 38, 31, 22, 30, 0, 0, 
    137, 107, 79, 122, 64, 56, 104, 114, 58, 43, 60, 69, 94, 99, 78, 
    197, 143, 78, 153, 147, 124, 139, 135, 119, 118, 133, 142, 150, 157, 150, 
    167, 177, 119, 165, 108, 128, 127, 127, 127, 135, 147, 156, 160, 157, 169, 
    172, 156, 177, 166, 110, 138, 130, 130, 132, 145, 161, 172, 163, 183, 194, 
    170, 167, 155, 165, 130, 145, 143, 131, 134, 149, 151, 153, 164, 189, 153, 
    
    -- channel=7
    120, 123, 123, 127, 126, 118, 124, 139, 130, 101, 83, 86, 97, 110, 115, 
    122, 129, 126, 129, 127, 97, 111, 99, 80, 50, 29, 32, 47, 80, 105, 
    71, 80, 129, 133, 131, 103, 78, 57, 42, 19, 29, 30, 29, 41, 77, 
    49, 33, 115, 127, 103, 83, 50, 41, 26, 26, 41, 35, 34, 31, 49, 
    40, 12, 103, 105, 43, 49, 41, 37, 24, 29, 40, 42, 28, 32, 34, 
    34, 6, 102, 104, 21, 54, 39, 47, 30, 4, 36, 41, 25, 30, 29, 
    43, 0, 62, 109, 40, 39, 28, 40, 37, 0, 39, 34, 25, 26, 38, 
    29, 12, 34, 59, 67, 14, 38, 30, 45, 34, 43, 38, 22, 30, 79, 
    18, 0, 28, 12, 49, 41, 50, 31, 29, 52, 41, 40, 28, 59, 92, 
    22, 12, 22, 0, 24, 35, 33, 24, 29, 37, 27, 20, 12, 64, 94, 
    0, 15, 22, 0, 20, 10, 0, 0, 1, 4, 0, 0, 0, 0, 0, 
    0, 0, 22, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=8
    5, 0, 4, 0, 0, 1, 3, 0, 0, 0, 2, 17, 4, 0, 0, 
    2, 0, 5, 0, 8, 0, 0, 0, 0, 21, 0, 0, 22, 28, 0, 
    0, 68, 4, 0, 8, 28, 0, 0, 9, 61, 0, 0, 0, 36, 34, 
    0, 95, 0, 8, 0, 22, 0, 0, 0, 109, 0, 2, 0, 0, 95, 
    0, 28, 0, 82, 0, 0, 0, 0, 0, 134, 0, 0, 0, 0, 51, 
    0, 24, 0, 25, 118, 9, 0, 0, 0, 210, 0, 0, 19, 0, 0, 
    0, 0, 15, 0, 95, 64, 0, 0, 0, 177, 0, 0, 11, 16, 0, 
    0, 0, 0, 0, 61, 84, 0, 5, 0, 116, 0, 0, 37, 15, 0, 
    0, 7, 0, 49, 0, 46, 0, 0, 39, 0, 32, 0, 43, 37, 11, 
    0, 13, 0, 85, 0, 12, 52, 0, 0, 3, 0, 4, 47, 41, 0, 
    90, 5, 0, 170, 0, 0, 62, 0, 0, 0, 0, 6, 22, 31, 0, 
    117, 76, 0, 122, 0, 0, 31, 26, 0, 8, 12, 16, 12, 13, 0, 
    0, 113, 132, 0, 0, 2, 0, 6, 2, 9, 13, 8, 6, 15, 14, 
    0, 17, 189, 0, 0, 12, 0, 1, 14, 11, 11, 16, 4, 32, 0, 
    0, 12, 35, 7, 0, 37, 24, 6, 11, 0, 0, 15, 45, 0, 0, 
    
    -- channel=9
    4, 0, 0, 0, 0, 0, 0, 0, 0, 22, 37, 28, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 69, 12, 0, 0, 29, 24, 0, 
    39, 67, 0, 0, 0, 78, 37, 43, 1, 0, 0, 0, 0, 30, 6, 
    0, 0, 0, 0, 0, 12, 0, 0, 0, 39, 0, 16, 10, 0, 31, 
    0, 0, 0, 14, 0, 0, 0, 0, 9, 7, 0, 0, 0, 0, 20, 
    10, 0, 0, 41, 100, 34, 0, 0, 0, 0, 0, 13, 5, 0, 0, 
    0, 0, 26, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 6, 32, 43, 0, 5, 1, 0, 11, 7, 0, 
    0, 0, 0, 0, 0, 84, 6, 0, 0, 0, 49, 58, 31, 0, 0, 
    8, 0, 0, 0, 0, 14, 0, 0, 0, 63, 55, 26, 0, 0, 5, 
    16, 0, 0, 0, 0, 0, 0, 47, 8, 0, 0, 0, 0, 39, 43, 
    101, 50, 0, 0, 80, 104, 70, 67, 30, 19, 5, 9, 0, 0, 0, 
    0, 73, 25, 0, 86, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 
    0, 0, 81, 65, 23, 0, 0, 0, 2, 0, 6, 19, 8, 0, 38, 
    0, 0, 11, 78, 31, 36, 36, 1, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=10
    168, 166, 175, 173, 173, 164, 184, 183, 170, 145, 123, 134, 143, 150, 138, 
    171, 179, 181, 178, 180, 196, 179, 160, 100, 87, 79, 82, 93, 128, 146, 
    114, 141, 182, 177, 182, 139, 84, 53, 65, 101, 70, 59, 53, 81, 133, 
    42, 148, 185, 183, 162, 127, 113, 63, 52, 105, 67, 61, 20, 30, 118, 
    47, 163, 173, 191, 198, 172, 90, 54, 28, 99, 105, 64, 59, 31, 79, 
    57, 119, 164, 132, 87, 103, 104, 73, 33, 172, 98, 31, 62, 44, 47, 
    68, 90, 124, 119, 110, 149, 123, 93, 36, 158, 61, 46, 53, 67, 66, 
    92, 84, 105, 124, 128, 174, 71, 65, 42, 143, 62, 34, 56, 75, 88, 
    90, 109, 43, 101, 116, 54, 59, 72, 95, 100, 68, 4, 34, 94, 163, 
    90, 105, 34, 94, 75, 83, 99, 106, 89, 64, 8, 8, 76, 167, 148, 
    109, 116, 31, 179, 124, 119, 133, 77, 31, 21, 17, 32, 41, 60, 45, 
    36, 79, 89, 222, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 33, 111, 141, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 90, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    
    -- channel=11
    12, 17, 11, 17, 14, 9, 13, 17, 13, 13, 14, 3, 9, 15, 19, 
    6, 9, 8, 20, 7, 0, 33, 9, 39, 0, 6, 0, 0, 0, 11, 
    19, 0, 9, 18, 7, 14, 58, 16, 0, 0, 49, 38, 46, 0, 0, 
    94, 0, 10, 1, 15, 0, 20, 39, 21, 0, 84, 26, 53, 19, 0, 
    125, 0, 55, 0, 24, 40, 82, 57, 34, 0, 35, 73, 7, 45, 0, 
    108, 9, 78, 27, 0, 76, 81, 59, 64, 0, 107, 95, 0, 39, 20, 
    104, 63, 19, 71, 0, 0, 65, 74, 89, 0, 121, 57, 2, 0, 40, 
    87, 78, 35, 33, 0, 0, 144, 50, 66, 0, 90, 69, 0, 19, 44, 
    101, 36, 125, 0, 29, 38, 49, 15, 0, 40, 0, 91, 0, 0, 0, 
    70, 48, 143, 0, 68, 21, 0, 47, 21, 45, 84, 7, 0, 0, 23, 
    0, 44, 137, 0, 141, 35, 0, 78, 105, 40, 0, 0, 0, 0, 0, 
    0, 12, 84, 0, 194, 100, 16, 17, 28, 9, 8, 8, 12, 15, 27, 
    33, 0, 0, 65, 182, 20, 26, 17, 17, 8, 4, 3, 21, 23, 3, 
    49, 6, 0, 145, 65, 11, 32, 16, 14, 12, 18, 20, 31, 0, 55, 
    64, 17, 7, 29, 31, 0, 21, 26, 11, 17, 34, 16, 0, 47, 80, 
    
    -- channel=12
    77, 83, 75, 83, 79, 74, 84, 85, 78, 74, 71, 64, 72, 75, 73, 
    74, 79, 74, 88, 73, 76, 104, 79, 84, 44, 65, 52, 38, 58, 72, 
    79, 50, 82, 87, 75, 73, 124, 64, 31, 9, 98, 80, 83, 23, 54, 
    142, 0, 91, 71, 89, 47, 86, 69, 58, 0, 142, 67, 92, 54, 0, 
    178, 37, 130, 4, 122, 83, 143, 101, 69, 0, 106, 117, 50, 80, 0, 
    148, 104, 161, 59, 68, 137, 170, 109, 108, 0, 169, 139, 41, 74, 54, 
    149, 149, 111, 134, 0, 56, 151, 137, 138, 0, 190, 107, 43, 47, 86, 
    149, 164, 86, 119, 9, 42, 190, 103, 123, 0, 153, 119, 28, 65, 90, 
    173, 121, 178, 66, 86, 80, 116, 77, 41, 92, 62, 119, 22, 50, 59, 
    151, 122, 214, 14, 141, 44, 43, 128, 63, 93, 109, 33, 3, 38, 95, 
    66, 127, 206, 0, 236, 96, 35, 146, 157, 74, 21, 13, 15, 40, 67, 
    6, 96, 157, 22, 273, 158, 63, 67, 74, 42, 41, 39, 48, 48, 64, 
    67, 1, 39, 172, 225, 54, 54, 47, 46, 37, 35, 40, 55, 54, 48, 
    84, 42, 0, 243, 102, 43, 66, 47, 40, 41, 45, 55, 62, 24, 87, 
    94, 47, 43, 85, 58, 30, 50, 56, 41, 54, 65, 43, 20, 87, 111, 
    
    -- channel=13
    58, 52, 59, 56, 57, 52, 66, 70, 57, 47, 47, 52, 50, 50, 44, 
    64, 59, 58, 59, 55, 31, 57, 55, 39, 12, 0, 8, 35, 55, 48, 
    36, 79, 65, 64, 60, 17, 37, 19, 1, 0, 0, 0, 0, 26, 46, 
    0, 28, 68, 61, 46, 31, 0, 0, 0, 0, 0, 0, 0, 0, 37, 
    0, 0, 56, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 61, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 71, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 49, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=14
    36, 36, 32, 30, 31, 28, 39, 41, 32, 36, 45, 41, 30, 33, 30, 
    31, 29, 33, 33, 23, 0, 29, 40, 61, 0, 0, 7, 35, 29, 25, 
    59, 49, 31, 35, 36, 66, 51, 34, 0, 0, 0, 0, 0, 30, 20, 
    0, 0, 25, 26, 27, 0, 0, 0, 0, 0, 10, 21, 13, 17, 20, 
    0, 0, 26, 0, 0, 0, 9, 6, 24, 0, 0, 0, 0, 0, 34, 
    8, 0, 30, 68, 43, 31, 0, 0, 0, 0, 16, 27, 0, 0, 0, 
    0, 2, 43, 32, 15, 0, 0, 0, 1, 0, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 50, 37, 10, 0, 13, 13, 0, 16, 19, 
    0, 0, 12, 0, 8, 56, 13, 0, 0, 30, 21, 61, 24, 0, 4, 
    0, 0, 0, 0, 0, 22, 0, 0, 14, 40, 51, 7, 0, 0, 30, 
    0, 0, 10, 0, 0, 0, 0, 10, 7, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 71, 46, 18, 13, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 23, 18, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 28, 0, 0, 0, 13, 12, 0, 
    34, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 21, 9, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 18, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 29, 20, 6, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 5, 12, 0, 0, 0, 
    0, 0, 0, 0, 4, 20, 0, 0, 0, 39, 22, 0, 7, 0, 0, 
    9, 0, 0, 0, 0, 0, 47, 46, 35, 0, 0, 0, 5, 25, 27, 
    45, 33, 0, 0, 21, 14, 0, 0, 0, 2, 1, 0, 0, 0, 0, 
    0, 28, 11, 11, 3, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 49, 31, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 0, 0, 0, 3, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 17, 61, 0, 0, 0, 
    0, 0, 51, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 8, 0, 
    12, 39, 2, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 104, 0, 
    0, 0, 0, 15, 0, 0, 22, 92, 112, 0, 0, 0, 0, 0, 0, 
    27, 115, 0, 60, 1, 11, 66, 0, 0, 0, 0, 17, 34, 46, 32, 
    260, 0, 23, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 20, 17, 
    0, 38, 0, 0, 0, 8, 142, 22, 35, 46, 68, 58, 0, 0, 39, 
    0, 7, 0, 0, 0, 1, 122, 0, 0, 0, 0, 0, 29, 26, 50, 
    0, 0, 3, 0, 0, 2, 59, 12, 0, 0, 54, 46, 1, 26, 33, 
    0, 0, 7, 5, 10, 12, 30, 22, 51, 67, 9, 0, 16, 21, 32, 
    
    -- channel=17
    527, 527, 527, 527, 528, 529, 529, 527, 527, 526, 528, 528, 528, 527, 530, 
    529, 530, 530, 529, 528, 528, 529, 530, 520, 459, 480, 522, 529, 529, 532, 
    524, 526, 532, 531, 532, 528, 527, 494, 438, 389, 413, 513, 531, 532, 535, 
    525, 529, 535, 535, 535, 497, 507, 483, 452, 441, 434, 511, 537, 537, 540, 
    325, 368, 513, 525, 530, 515, 523, 521, 523, 501, 451, 409, 376, 465, 542, 
    416, 451, 505, 441, 471, 379, 394, 423, 483, 505, 459, 443, 395, 472, 539, 
    254, 308, 382, 442, 448, 192, 218, 325, 446, 491, 444, 395, 394, 396, 436, 
    149, 306, 271, 384, 451, 413, 458, 422, 375, 345, 301, 296, 327, 372, 400, 
    274, 463, 419, 462, 498, 488, 478, 402, 390, 366, 383, 347, 327, 328, 321, 
    300, 296, 314, 318, 329, 340, 328, 296, 298, 243, 244, 206, 205, 220, 269, 
    10, 55, 39, 32, 47, 79, 111, 125, 135, 114, 108, 128, 184, 215, 260, 
    0, 26, 44, 0, 0, 0, 142, 121, 106, 113, 158, 196, 209, 232, 292, 
    0, 0, 0, 0, 0, 0, 145, 202, 186, 162, 136, 157, 190, 265, 356, 
    0, 0, 0, 0, 0, 0, 0, 58, 7, 51, 124, 203, 244, 291, 385, 
    20, 0, 0, 0, 0, 0, 0, 37, 64, 174, 223, 235, 270, 325, 403, 
    
    -- channel=18
    120, 122, 122, 122, 123, 123, 123, 123, 122, 122, 125, 122, 122, 122, 124, 
    122, 124, 124, 123, 124, 123, 124, 122, 120, 110, 141, 135, 123, 123, 125, 
    125, 126, 125, 123, 125, 123, 127, 115, 121, 91, 129, 149, 124, 125, 126, 
    126, 121, 127, 125, 127, 109, 138, 90, 75, 58, 55, 127, 124, 125, 126, 
    136, 154, 158, 128, 127, 101, 119, 112, 116, 116, 122, 128, 136, 164, 132, 
    36, 52, 113, 123, 136, 133, 160, 158, 152, 103, 63, 47, 20, 110, 131, 
    126, 155, 141, 97, 73, 0, 29, 51, 114, 128, 134, 133, 136, 130, 156, 
    46, 37, 45, 133, 103, 22, 50, 79, 114, 89, 48, 38, 43, 49, 81, 
    85, 84, 42, 84, 122, 120, 140, 82, 75, 88, 98, 91, 107, 113, 97, 
    123, 129, 138, 139, 134, 120, 97, 79, 91, 54, 74, 49, 45, 48, 66, 
    13, 40, 42, 59, 76, 93, 102, 97, 80, 63, 49, 43, 42, 31, 53, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 38, 39, 49, 
    0, 0, 0, 0, 0, 0, 129, 74, 46, 43, 51, 45, 20, 36, 69, 
    0, 0, 0, 0, 0, 0, 7, 62, 36, 11, 0, 9, 24, 50, 85, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 15, 21, 35, 52, 83, 
    
    -- channel=19
    20, 20, 20, 20, 20, 19, 20, 19, 18, 20, 22, 19, 19, 20, 19, 
    20, 20, 20, 19, 20, 20, 20, 19, 18, 16, 26, 23, 20, 20, 20, 
    20, 20, 19, 19, 20, 18, 22, 15, 29, 41, 24, 26, 20, 19, 20, 
    27, 24, 19, 19, 20, 11, 21, 28, 39, 42, 41, 22, 22, 20, 20, 
    38, 40, 23, 19, 19, 23, 13, 23, 24, 27, 24, 28, 29, 37, 21, 
    43, 35, 8, 18, 16, 18, 24, 25, 31, 31, 43, 40, 36, 19, 22, 
    45, 46, 38, 40, 16, 61, 53, 52, 30, 19, 21, 25, 29, 20, 33, 
    63, 21, 32, 14, 37, 45, 26, 9, 29, 44, 49, 48, 42, 42, 27, 
    49, 25, 37, 22, 24, 24, 24, 47, 43, 40, 45, 38, 39, 39, 48, 
    17, 59, 61, 67, 68, 68, 69, 70, 60, 70, 59, 69, 59, 51, 43, 
    42, 46, 51, 52, 48, 55, 69, 71, 70, 72, 69, 66, 66, 48, 30, 
    28, 26, 33, 28, 27, 34, 57, 63, 66, 68, 63, 45, 23, 29, 20, 
    15, 16, 20, 24, 25, 21, 17, 34, 22, 8, 4, 20, 19, 12, 13, 
    18, 18, 19, 22, 21, 20, 17, 0, 0, 11, 12, 0, 7, 12, 13, 
    20, 9, 11, 16, 17, 18, 10, 10, 16, 0, 0, 7, 9, 12, 14, 
    
    -- channel=20
    42, 44, 44, 44, 44, 44, 44, 44, 46, 42, 41, 43, 44, 44, 44, 
    42, 43, 43, 43, 43, 43, 44, 43, 42, 25, 34, 42, 43, 43, 43, 
    44, 45, 44, 43, 44, 44, 43, 33, 23, 8, 41, 47, 43, 44, 43, 
    32, 34, 41, 46, 45, 33, 45, 25, 11, 4, 2, 40, 35, 38, 41, 
    4, 20, 40, 47, 45, 35, 48, 37, 37, 28, 23, 18, 20, 39, 38, 
    17, 24, 52, 44, 44, 40, 43, 44, 40, 15, 3, 11, 1, 38, 39, 
    1, 18, 23, 27, 19, 0, 0, 0, 31, 43, 39, 36, 40, 39, 37, 
    9, 10, 19, 50, 22, 0, 31, 32, 20, 0, 0, 0, 1, 5, 22, 
    45, 42, 21, 46, 42, 27, 30, 5, 20, 19, 15, 14, 14, 11, 0, 
    48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 26, 
    4, 36, 13, 9, 9, 15, 0, 0, 0, 0, 0, 18, 39, 33, 34, 
    8, 16, 31, 16, 11, 14, 101, 90, 101, 96, 76, 51, 36, 42, 39, 
    0, 16, 22, 16, 16, 17, 81, 167, 141, 80, 55, 55, 40, 37, 39, 
    0, 19, 16, 14, 16, 14, 39, 78, 54, 70, 54, 35, 38, 37, 37, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 32, 0, 0, 0, 
    29, 31, 21, 0, 0, 0, 8, 0, 0, 0, 0, 9, 17, 18, 1, 
    0, 0, 23, 1, 8, 3, 14, 8, 0, 0, 0, 0, 0, 33, 3, 
    25, 23, 17, 0, 0, 0, 20, 28, 37, 5, 0, 1, 2, 10, 13, 
    13, 36, 21, 42, 0, 0, 0, 8, 9, 0, 0, 4, 12, 4, 22, 
    71, 3, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 7, 16, 8, 
    48, 0, 7, 0, 0, 0, 0, 0, 5, 0, 11, 0, 9, 13, 16, 
    35, 34, 28, 32, 37, 28, 16, 12, 11, 5, 8, 10, 12, 15, 21, 
    16, 50, 3, 12, 25, 31, 4, 0, 6, 4, 7, 12, 7, 7, 19, 
    21, 46, 37, 18, 27, 33, 99, 0, 0, 0, 0, 1, 10, 21, 28, 
    0, 34, 34, 28, 33, 34, 59, 0, 0, 0, 5, 29, 21, 27, 27, 
    0, 33, 36, 36, 34, 33, 46, 5, 1, 36, 24, 22, 26, 25, 25, 
    
    -- channel=22
    143, 144, 144, 144, 145, 145, 145, 144, 142, 146, 148, 145, 144, 144, 145, 
    145, 146, 146, 146, 146, 146, 146, 144, 146, 150, 157, 151, 145, 146, 147, 
    145, 144, 146, 146, 145, 146, 148, 151, 155, 144, 152, 156, 147, 147, 148, 
    155, 152, 152, 146, 145, 146, 149, 139, 133, 135, 131, 163, 157, 153, 153, 
    173, 169, 168, 144, 146, 140, 145, 142, 149, 157, 164, 168, 165, 163, 160, 
    106, 113, 155, 136, 153, 146, 159, 158, 158, 158, 136, 121, 108, 144, 161, 
    159, 158, 154, 124, 144, 86, 111, 125, 145, 157, 154, 149, 144, 154, 158, 
    77, 112, 108, 139, 144, 97, 113, 143, 150, 137, 121, 109, 113, 116, 136, 
    89, 139, 96, 117, 148, 159, 170, 131, 130, 137, 146, 145, 148, 158, 148, 
    149, 160, 176, 176, 175, 172, 166, 150, 153, 129, 145, 125, 116, 112, 117, 
    78, 93, 99, 104, 110, 121, 139, 136, 133, 119, 110, 105, 107, 97, 97, 
    9, 37, 20, 6, 3, 14, 53, 61, 73, 69, 66, 69, 70, 76, 83, 
    0, 11, 18, 0, 0, 0, 76, 8, 0, 0, 20, 39, 42, 72, 106, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 68, 89, 123, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 17, 49, 67, 79, 97, 126, 
    
    -- channel=23
    12, 11, 11, 11, 11, 11, 11, 12, 14, 10, 7, 10, 12, 11, 11, 
    12, 11, 11, 11, 11, 11, 11, 12, 10, 2, 0, 7, 11, 11, 11, 
    12, 12, 12, 13, 12, 11, 9, 6, 0, 0, 0, 0, 11, 12, 11, 
    0, 1, 8, 13, 11, 9, 10, 16, 6, 2, 0, 0, 4, 6, 9, 
    0, 0, 0, 14, 11, 13, 6, 11, 4, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 13, 1, 2, 0, 0, 0, 1, 8, 5, 3, 0, 1, 
    0, 0, 0, 3, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 6, 12, 17, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    25, 14, 20, 20, 21, 15, 0, 0, 0, 0, 5, 4, 5, 12, 13, 
    36, 21, 25, 29, 27, 24, 13, 73, 68, 55, 33, 32, 27, 17, 9, 
    40, 27, 23, 24, 26, 25, 25, 57, 49, 32, 34, 25, 25, 19, 9, 
    47, 40, 33, 31, 31, 29, 19, 28, 40, 42, 33, 29, 25, 18, 9, 
    
    -- channel=24
    0, 2, 2, 2, 3, 3, 3, 0, 3, 0, 4, 3, 2, 2, 4, 
    0, 3, 3, 2, 4, 2, 5, 1, 0, 0, 59, 31, 1, 3, 4, 
    5, 7, 5, 1, 5, 0, 11, 0, 1, 0, 63, 74, 1, 4, 4, 
    15, 0, 7, 5, 3, 0, 51, 0, 0, 0, 0, 57, 3, 3, 5, 
    63, 95, 86, 12, 5, 0, 22, 0, 5, 0, 0, 22, 37, 115, 19, 
    0, 0, 10, 13, 25, 4, 68, 64, 68, 0, 0, 0, 0, 79, 23, 
    63, 117, 61, 37, 0, 0, 40, 56, 78, 4, 7, 17, 37, 28, 91, 
    105, 28, 2, 108, 11, 0, 0, 0, 25, 5, 0, 0, 11, 0, 22, 
    214, 0, 0, 6, 22, 0, 22, 0, 0, 0, 14, 0, 34, 43, 29, 
    112, 51, 63, 57, 53, 38, 7, 14, 21, 0, 20, 0, 17, 26, 40, 
    20, 65, 29, 55, 73, 88, 70, 64, 47, 32, 31, 36, 44, 10, 35, 
    0, 74, 0, 0, 0, 26, 76, 0, 0, 0, 8, 0, 14, 12, 40, 
    0, 38, 36, 0, 0, 9, 233, 23, 6, 0, 15, 30, 13, 29, 51, 
    0, 0, 10, 0, 3, 4, 125, 34, 0, 14, 9, 23, 11, 39, 52, 
    0, 0, 0, 0, 0, 0, 43, 27, 4, 40, 7, 7, 23, 30, 44, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 38, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 58, 32, 40, 29, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    138, 132, 28, 0, 0, 0, 0, 0, 0, 0, 41, 94, 115, 91, 0, 
    0, 0, 0, 44, 42, 124, 154, 129, 83, 0, 0, 0, 0, 0, 0, 
    156, 165, 83, 0, 0, 0, 0, 0, 0, 3, 65, 103, 98, 95, 95, 
    44, 0, 6, 36, 0, 0, 0, 0, 78, 50, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 21, 48, 25, 0, 20, 21, 40, 84, 105, 72, 
    63, 133, 129, 122, 106, 81, 51, 26, 32, 20, 43, 35, 10, 13, 10, 
    82, 84, 92, 127, 150, 168, 156, 147, 120, 103, 78, 48, 3, 0, 0, 
    17, 32, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 27, 59, 39, 13, 8, 88, 13, 0, 0, 70, 65, 0, 0, 0, 
    0, 2, 12, 12, 6, 5, 15, 24, 90, 55, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    152, 153, 153, 153, 154, 153, 153, 153, 154, 151, 149, 155, 153, 153, 154, 
    152, 153, 153, 152, 152, 152, 152, 153, 149, 105, 113, 148, 153, 152, 153, 
    149, 151, 153, 153, 155, 152, 149, 130, 86, 62, 114, 139, 153, 153, 154, 
    146, 149, 154, 156, 155, 129, 143, 118, 118, 112, 123, 169, 150, 152, 154, 
    16, 47, 132, 151, 151, 134, 169, 146, 153, 132, 98, 65, 53, 102, 152, 
    145, 166, 164, 118, 119, 76, 70, 85, 108, 111, 118, 138, 114, 176, 152, 
    0, 15, 67, 122, 113, 0, 25, 80, 161, 137, 102, 74, 76, 75, 91, 
    8, 115, 60, 108, 95, 125, 180, 122, 56, 36, 38, 60, 88, 107, 134, 
    151, 134, 152, 173, 151, 120, 112, 78, 109, 90, 84, 69, 51, 35, 29, 
    86, 7, 8, 7, 11, 19, 13, 20, 25, 7, 8, 0, 16, 35, 55, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 50, 75, 
    0, 21, 15, 0, 0, 0, 24, 28, 7, 14, 48, 83, 76, 56, 100, 
    0, 0, 0, 0, 0, 0, 90, 82, 101, 84, 43, 24, 74, 100, 125, 
    0, 0, 0, 0, 0, 0, 73, 119, 59, 39, 88, 115, 88, 102, 120, 
    0, 11, 4, 0, 1, 1, 37, 56, 79, 127, 102, 82, 98, 112, 128, 
    
    -- channel=27
    71, 67, 67, 67, 66, 67, 67, 69, 67, 67, 65, 66, 67, 67, 65, 
    71, 67, 67, 67, 66, 67, 65, 68, 67, 103, 35, 42, 68, 66, 65, 
    72, 68, 66, 68, 65, 70, 64, 89, 82, 88, 16, 26, 68, 67, 66, 
    46, 61, 60, 67, 68, 99, 32, 101, 58, 63, 33, 0, 64, 63, 64, 
    47, 22, 8, 67, 66, 88, 32, 73, 55, 79, 96, 89, 73, 9, 56, 
    45, 26, 37, 73, 57, 109, 72, 71, 60, 88, 60, 46, 75, 0, 50, 
    53, 21, 30, 32, 87, 132, 0, 0, 0, 70, 95, 101, 78, 84, 29, 
    0, 0, 49, 0, 50, 64, 6, 87, 67, 61, 47, 12, 0, 2, 0, 
    0, 50, 33, 21, 43, 80, 59, 111, 54, 71, 60, 83, 67, 65, 58, 
    0, 69, 52, 56, 54, 51, 63, 42, 33, 60, 37, 54, 19, 21, 14, 
    25, 0, 29, 28, 26, 28, 40, 42, 48, 50, 33, 18, 0, 9, 6, 
    31, 0, 40, 32, 7, 0, 0, 12, 0, 0, 0, 0, 39, 34, 0, 
    34, 0, 0, 20, 0, 0, 0, 108, 99, 95, 79, 34, 0, 0, 0, 
    99, 0, 0, 0, 0, 0, 0, 15, 55, 1, 0, 0, 14, 0, 0, 
    95, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 18, 5, 4, 3, 
    
    -- channel=28
    177, 172, 172, 172, 171, 173, 173, 175, 171, 173, 171, 173, 173, 172, 172, 
    177, 173, 173, 174, 173, 173, 172, 175, 175, 202, 137, 153, 174, 173, 173, 
    175, 172, 173, 175, 171, 177, 168, 191, 173, 177, 92, 124, 177, 173, 174, 
    158, 171, 171, 174, 175, 208, 136, 202, 146, 149, 123, 80, 176, 173, 174, 
    125, 104, 125, 172, 173, 198, 135, 181, 155, 179, 179, 166, 152, 99, 168, 
    116, 99, 127, 162, 157, 176, 142, 146, 143, 193, 160, 135, 156, 44, 156, 
    112, 83, 124, 122, 181, 181, 42, 32, 42, 162, 174, 172, 152, 150, 111, 
    0, 33, 100, 47, 150, 156, 87, 155, 145, 149, 131, 96, 74, 91, 78, 
    0, 133, 119, 104, 128, 176, 157, 196, 116, 123, 124, 138, 119, 121, 129, 
    0, 120, 106, 118, 117, 123, 132, 108, 100, 115, 84, 100, 63, 66, 65, 
    40, 16, 47, 38, 35, 35, 54, 62, 72, 72, 57, 45, 35, 58, 55, 
    37, 0, 52, 32, 3, 0, 0, 40, 17, 14, 10, 24, 61, 79, 54, 
    41, 0, 3, 27, 1, 0, 0, 126, 95, 97, 90, 76, 56, 49, 57, 
    127, 0, 0, 0, 0, 0, 0, 58, 77, 39, 16, 23, 69, 59, 74, 
    129, 5, 0, 0, 0, 0, 0, 4, 1, 0, 59, 77, 68, 71, 83, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 19, 59, 49, 31, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 22, 4, 0, 0, 0, 0, 0, 0, 
    
    -- channel=30
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    65, 42, 0, 0, 0, 0, 0, 0, 0, 0, 7, 39, 55, 0, 0, 
    0, 0, 0, 14, 3, 64, 63, 44, 4, 0, 0, 0, 0, 0, 0, 
    87, 70, 16, 0, 0, 4, 0, 0, 0, 0, 26, 54, 32, 48, 15, 
    0, 0, 8, 0, 0, 0, 0, 0, 38, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 26, 44, 19, 
    15, 60, 54, 50, 39, 20, 8, 0, 0, 0, 10, 4, 0, 0, 0, 
    68, 52, 74, 94, 103, 101, 91, 83, 67, 62, 39, 17, 0, 0, 0, 
    24, 0, 0, 4, 17, 15, 0, 0, 0, 0, 0, 0, 2, 6, 0, 
    8, 32, 56, 46, 23, 19, 49, 86, 81, 91, 116, 64, 0, 0, 0, 
    9, 14, 21, 22, 16, 15, 57, 151, 173, 72, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 12, 39, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 4, 23, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 12, 2, 0, 0, 0, 0, 0, 0, 0, 29, 30, 29, 11, 0, 
    0, 0, 0, 13, 18, 67, 88, 75, 36, 0, 0, 0, 0, 0, 0, 
    43, 29, 19, 0, 0, 0, 0, 0, 0, 7, 43, 56, 54, 42, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 19, 17, 28, 36, 26, 47, 49, 55, 60, 34, 0, 
    55, 51, 38, 38, 26, 11, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 16, 29, 36, 48, 54, 41, 31, 21, 6, 0, 0, 0, 
    4, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    0, 2, 5, 0, 0, 0, 23, 3, 0, 16, 33, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 30, 59, 69, 17, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=32
    0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 65, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 1, 0, 0, 
    39, 7, 0, 10, 34, 5, 5, 0, 0, 0, 49, 58, 0, 55, 0, 
    11, 0, 0, 36, 22, 0, 10, 2, 27, 23, 55, 0, 0, 0, 0, 
    3, 18, 40, 35, 14, 0, 0, 0, 0, 0, 0, 7, 0, 0, 75, 
    0, 0, 20, 8, 0, 0, 0, 0, 4, 0, 41, 0, 0, 0, 0, 
    0, 56, 3, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 
    53, 0, 0, 0, 10, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 
    0, 4, 4, 6, 6, 2, 0, 0, 31, 0, 0, 0, 0, 3, 0, 
    
    -- channel=33
    418, 397, 495, 500, 521, 511, 535, 529, 534, 549, 527, 552, 534, 552, 541, 
    426, 396, 498, 488, 521, 492, 508, 527, 526, 470, 452, 549, 530, 548, 539, 
    423, 375, 481, 479, 507, 476, 471, 447, 474, 371, 384, 505, 501, 514, 522, 
    383, 334, 415, 440, 455, 451, 442, 386, 291, 221, 218, 212, 361, 429, 427, 
    216, 202, 230, 256, 274, 290, 304, 289, 218, 203, 195, 211, 279, 309, 233, 
    179, 189, 202, 205, 262, 245, 267, 232, 217, 219, 267, 382, 282, 341, 177, 
    208, 178, 170, 224, 298, 301, 310, 292, 297, 303, 351, 399, 347, 255, 106, 
    253, 268, 295, 341, 378, 393, 394, 362, 358, 291, 294, 343, 344, 215, 220, 
    249, 252, 303, 371, 368, 355, 349, 339, 338, 317, 328, 342, 333, 290, 303, 
    233, 273, 328, 323, 331, 346, 349, 315, 303, 352, 349, 316, 257, 189, 157, 
    295, 311, 303, 267, 271, 327, 290, 181, 209, 287, 254, 203, 142, 107, 79, 
    265, 287, 251, 183, 200, 270, 234, 175, 183, 183, 140, 121, 82, 55, 21, 
    198, 203, 178, 147, 151, 151, 135, 133, 117, 113, 80, 80, 50, 28, 20, 
    52, 50, 56, 68, 79, 81, 87, 78, 104, 85, 54, 35, 23, 26, 23, 
    15, 20, 35, 46, 57, 63, 65, 44, 94, 51, 28, 16, 18, 31, 0, 
    
    -- channel=34
    83, 99, 127, 125, 131, 126, 131, 118, 134, 139, 128, 133, 121, 129, 131, 
    85, 97, 132, 115, 128, 117, 130, 131, 130, 105, 140, 142, 122, 135, 135, 
    83, 92, 125, 104, 118, 107, 107, 131, 138, 49, 144, 153, 118, 130, 138, 
    83, 83, 119, 122, 110, 109, 93, 70, 73, 59, 62, 106, 166, 125, 132, 
    84, 67, 82, 107, 104, 110, 101, 75, 36, 27, 34, 18, 53, 52, 73, 
    19, 16, 8, 20, 23, 26, 49, 36, 29, 17, 35, 43, 0, 76, 0, 
    38, 19, 22, 48, 73, 42, 47, 22, 15, 28, 72, 97, 45, 62, 0, 
    31, 18, 29, 50, 73, 79, 81, 77, 92, 57, 89, 87, 68, 0, 0, 
    69, 72, 100, 105, 101, 100, 88, 65, 69, 22, 46, 62, 66, 49, 74, 
    25, 51, 70, 82, 74, 64, 69, 75, 80, 78, 75, 69, 61, 42, 36, 
    76, 67, 72, 65, 92, 95, 48, 24, 55, 84, 70, 46, 15, 0, 0, 
    84, 68, 39, 28, 25, 81, 52, 17, 27, 30, 15, 1, 0, 0, 0, 
    66, 63, 51, 33, 36, 38, 18, 10, 13, 9, 0, 0, 0, 0, 0, 
    6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 
    
    -- channel=35
    57, 60, 49, 48, 42, 39, 29, 25, 24, 24, 25, 22, 28, 21, 28, 
    45, 49, 35, 34, 24, 26, 20, 21, 23, 11, 39, 20, 24, 16, 25, 
    34, 42, 24, 22, 7, 18, 10, 15, 22, 21, 26, 21, 17, 9, 15, 
    25, 38, 10, 14, 2, 10, 11, 8, 22, 54, 36, 31, 23, 3, 8, 
    32, 30, 26, 16, 17, 15, 29, 34, 54, 45, 48, 50, 13, 2, 11, 
    46, 46, 33, 47, 37, 45, 48, 57, 47, 44, 52, 21, 6, 2, 25, 
    45, 49, 53, 50, 55, 61, 62, 67, 55, 46, 27, 12, 22, 3, 38, 
    64, 59, 60, 57, 59, 57, 57, 51, 48, 31, 26, 17, 21, 40, 27, 
    62, 57, 64, 63, 59, 57, 53, 51, 42, 40, 23, 22, 29, 27, 12, 
    77, 63, 54, 56, 65, 54, 42, 33, 42, 35, 33, 26, 23, 27, 30, 
    68, 64, 59, 55, 45, 52, 40, 53, 45, 25, 30, 36, 33, 36, 22, 
    49, 60, 52, 63, 57, 38, 44, 44, 36, 36, 31, 38, 36, 33, 36, 
    45, 47, 50, 47, 40, 41, 46, 36, 33, 37, 39, 34, 36, 37, 37, 
    38, 42, 39, 38, 32, 32, 36, 36, 43, 30, 38, 34, 38, 35, 32, 
    30, 30, 31, 33, 35, 33, 32, 31, 29, 43, 33, 37, 35, 35, 23, 
    
    -- channel=36
    0, 0, 7, 10, 18, 25, 34, 31, 39, 39, 39, 43, 35, 38, 41, 
    0, 10, 27, 23, 36, 34, 40, 40, 42, 21, 39, 49, 39, 46, 46, 
    11, 23, 42, 37, 51, 40, 40, 51, 50, 0, 46, 55, 40, 53, 54, 
    28, 34, 58, 61, 64, 57, 51, 30, 6, 0, 0, 12, 50, 62, 73, 
    20, 15, 25, 42, 44, 46, 30, 9, 0, 0, 0, 12, 52, 36, 36, 
    0, 4, 1, 6, 0, 0, 0, 0, 0, 0, 12, 34, 13, 57, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 50, 33, 67, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 32, 44, 37, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 32, 33, 24, 23, 54, 
    0, 0, 0, 0, 0, 0, 1, 10, 12, 16, 21, 21, 19, 13, 16, 
    0, 0, 0, 0, 3, 0, 0, 0, 5, 19, 12, 3, 0, 2, 8, 
    0, 0, 0, 0, 0, 10, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    3, 3, 0, 0, 0, 0, 0, 0, 17, 0, 1, 0, 0, 1, 3, 
    
    -- channel=37
    0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 9, 0, 2, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 2, 11, 0, 8, 0, 0, 11, 8, 0, 41, 7, 0, 2, 0, 
    0, 3, 11, 0, 0, 0, 0, 0, 4, 2, 38, 54, 36, 13, 11, 
    17, 14, 26, 35, 22, 20, 8, 1, 0, 7, 11, 13, 30, 22, 25, 
    24, 17, 8, 15, 7, 10, 5, 1, 13, 11, 22, 6, 0, 19, 0, 
    25, 11, 10, 21, 19, 0, 2, 0, 5, 13, 32, 17, 0, 31, 0, 
    2, 0, 0, 0, 0, 0, 0, 1, 3, 7, 29, 13, 0, 0, 8, 
    8, 6, 21, 1, 0, 1, 10, 7, 15, 0, 19, 7, 2, 0, 20, 
    0, 9, 5, 8, 3, 9, 11, 12, 5, 10, 7, 2, 7, 11, 21, 
    8, 5, 9, 1, 22, 14, 3, 5, 38, 25, 11, 13, 15, 18, 26, 
    40, 8, 3, 10, 13, 43, 0, 1, 23, 24, 21, 21, 24, 25, 22, 
    34, 16, 11, 14, 27, 30, 15, 25, 25, 26, 23, 32, 15, 26, 23, 
    33, 30, 29, 32, 32, 31, 29, 32, 23, 24, 25, 24, 23, 28, 30, 
    27, 31, 33, 33, 30, 30, 32, 32, 39, 8, 27, 22, 29, 29, 26, 
    
    -- channel=38
    171, 156, 185, 178, 177, 162, 162, 158, 161, 163, 150, 155, 150, 160, 149, 
    163, 141, 170, 156, 163, 147, 154, 157, 153, 157, 141, 152, 145, 157, 147, 
    146, 122, 149, 135, 145, 132, 142, 144, 145, 132, 140, 154, 142, 145, 142, 
    122, 98, 121, 113, 113, 115, 118, 113, 127, 123, 126, 135, 138, 127, 113, 
    109, 93, 109, 112, 107, 108, 115, 125, 103, 107, 104, 75, 84, 103, 87, 
    92, 81, 91, 85, 96, 99, 121, 122, 108, 102, 92, 92, 72, 90, 52, 
    115, 95, 98, 111, 139, 129, 140, 122, 120, 121, 117, 119, 83, 81, 38, 
    117, 107, 104, 129, 147, 156, 161, 156, 152, 131, 114, 99, 93, 45, 50, 
    142, 140, 155, 166, 171, 171, 168, 146, 129, 100, 94, 102, 108, 90, 100, 
    127, 126, 147, 159, 154, 147, 142, 137, 123, 131, 122, 115, 106, 92, 80, 
    154, 156, 154, 138, 149, 152, 140, 106, 108, 129, 120, 108, 83, 68, 61, 
    151, 149, 143, 117, 111, 139, 118, 88, 97, 101, 89, 84, 68, 58, 41, 
    125, 128, 120, 103, 110, 109, 87, 85, 86, 86, 68, 66, 55, 47, 40, 
    79, 75, 71, 71, 71, 72, 78, 74, 62, 67, 57, 48, 45, 45, 44, 
    37, 39, 49, 52, 55, 57, 63, 56, 66, 55, 46, 40, 44, 45, 31, 
    
    -- channel=39
    0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 11, 11, 11, 3, 10, 
    0, 0, 0, 2, 0, 10, 4, 3, 7, 0, 12, 7, 15, 7, 12, 
    0, 10, 6, 19, 14, 18, 9, 11, 11, 12, 0, 2, 16, 18, 16, 
    9, 19, 11, 22, 27, 29, 25, 11, 0, 2, 0, 6, 5, 14, 34, 
    0, 2, 1, 1, 9, 8, 4, 0, 0, 0, 0, 7, 10, 16, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 24, 19, 33, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 30, 22, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 18, 18, 31, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 6, 7, 15, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 9, 10, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 2, 5, 8, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 5, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 4, 6, 6, 5, 
    2, 5, 2, 1, 0, 1, 1, 4, 7, 0, 6, 6, 7, 6, 7, 
    11, 10, 8, 8, 6, 4, 1, 8, 4, 12, 5, 7, 5, 5, 15, 
    
    -- channel=40
    0, 41, 31, 10, 10, 10, 12, 0, 24, 8, 4, 15, 0, 0, 17, 
    0, 42, 41, 0, 13, 4, 10, 11, 20, 0, 82, 33, 0, 1, 26, 
    0, 40, 46, 0, 9, 0, 0, 32, 48, 0, 132, 65, 0, 13, 34, 
    0, 42, 37, 38, 6, 18, 0, 0, 0, 0, 56, 80, 140, 32, 60, 
    37, 48, 35, 72, 50, 57, 43, 0, 0, 0, 21, 12, 48, 0, 45, 
    30, 22, 0, 30, 0, 0, 9, 0, 4, 0, 52, 12, 0, 37, 0, 
    24, 7, 0, 64, 37, 0, 0, 0, 0, 0, 57, 29, 0, 0, 0, 
    0, 0, 0, 6, 7, 0, 0, 0, 14, 0, 69, 42, 0, 0, 0, 
    9, 26, 65, 35, 4, 13, 15, 0, 14, 0, 23, 3, 1, 0, 12, 
    0, 28, 19, 9, 14, 4, 0, 0, 40, 17, 10, 0, 0, 0, 26, 
    47, 6, 5, 0, 41, 57, 0, 0, 70, 33, 10, 0, 0, 0, 0, 
    83, 17, 0, 1, 11, 61, 0, 0, 25, 5, 0, 4, 0, 3, 0, 
    61, 22, 0, 18, 28, 25, 6, 5, 11, 12, 0, 20, 0, 3, 0, 
    24, 24, 14, 22, 15, 19, 18, 3, 30, 0, 5, 2, 0, 6, 0, 
    1, 11, 9, 11, 6, 4, 5, 0, 72, 0, 9, 1, 6, 13, 0, 
    
    -- channel=41
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 51, 0, 0, 0, 0, 
    0, 8, 0, 0, 0, 0, 0, 44, 37, 14, 48, 49, 5, 4, 1, 
    16, 15, 25, 32, 16, 7, 2, 0, 83, 89, 57, 130, 129, 54, 68, 
    109, 92, 94, 111, 114, 117, 101, 71, 23, 0, 13, 0, 0, 0, 73, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 18, 4, 0, 0, 0, 0, 0, 0, 0, 4, 0, 34, 55, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 21, 56, 20, 2, 0, 0, 
    13, 59, 35, 5, 11, 38, 29, 0, 0, 0, 0, 0, 0, 0, 40, 
    0, 0, 0, 12, 0, 0, 0, 23, 58, 3, 0, 9, 56, 70, 65, 
    13, 0, 0, 26, 62, 49, 6, 34, 18, 42, 71, 65, 43, 34, 28, 
    16, 12, 1, 14, 0, 1, 44, 21, 20, 26, 39, 38, 9, 20, 16, 
    40, 63, 70, 49, 57, 57, 25, 10, 42, 43, 13, 18, 22, 11, 3, 
    48, 52, 33, 23, 25, 38, 35, 19, 0, 0, 19, 12, 10, 0, 0, 
    8, 3, 0, 0, 0, 0, 6, 16, 36, 9, 8, 8, 6, 3, 13, 
    
    -- channel=42
    66, 86, 107, 111, 123, 130, 144, 135, 149, 151, 141, 156, 148, 152, 156, 
    77, 97, 124, 122, 136, 132, 137, 137, 149, 103, 118, 162, 149, 151, 159, 
    90, 102, 137, 135, 150, 134, 127, 116, 130, 44, 120, 139, 136, 145, 155, 
    87, 104, 130, 132, 141, 137, 123, 111, 35, 0, 19, 18, 76, 124, 132, 
    13, 27, 29, 54, 54, 61, 53, 31, 17, 25, 21, 69, 115, 84, 64, 
    33, 58, 41, 47, 68, 65, 52, 22, 33, 33, 88, 148, 103, 104, 43, 
    34, 24, 6, 40, 48, 41, 46, 46, 68, 75, 128, 125, 84, 105, 0, 
    45, 62, 78, 94, 86, 81, 75, 67, 61, 43, 66, 103, 101, 38, 90, 
    23, 9, 35, 53, 50, 37, 35, 46, 81, 72, 126, 110, 88, 83, 86, 
    5, 60, 64, 39, 34, 67, 78, 64, 53, 78, 90, 74, 45, 16, 21, 
    26, 37, 39, 23, 29, 39, 27, 0, 48, 58, 30, 7, 8, 3, 9, 
    36, 24, 2, 0, 15, 64, 17, 19, 28, 19, 8, 0, 0, 0, 0, 
    27, 8, 0, 0, 0, 0, 0, 18, 4, 0, 0, 10, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 17, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 4, 10, 5, 0, 21, 0, 0, 0, 0, 0, 0, 
    
    -- channel=43
    82, 26, 36, 62, 61, 66, 63, 83, 49, 65, 84, 63, 79, 69, 61, 
    83, 30, 34, 73, 58, 72, 63, 64, 56, 115, 17, 46, 84, 71, 57, 
    90, 38, 32, 75, 57, 69, 77, 55, 43, 171, 0, 45, 90, 66, 50, 
    94, 37, 49, 59, 75, 61, 84, 73, 89, 71, 0, 4, 0, 60, 56, 
    43, 33, 28, 9, 37, 35, 43, 76, 57, 43, 26, 0, 0, 53, 13, 
    0, 0, 45, 0, 0, 7, 17, 54, 29, 27, 0, 4, 89, 3, 94, 
    3, 28, 34, 0, 0, 39, 25, 32, 12, 14, 0, 39, 102, 40, 128, 
    19, 18, 8, 8, 26, 39, 48, 61, 54, 94, 13, 19, 50, 115, 0, 
    36, 52, 0, 28, 58, 64, 56, 48, 22, 69, 0, 31, 45, 56, 47, 
    38, 0, 25, 48, 35, 28, 40, 62, 48, 36, 37, 64, 72, 70, 26, 
    12, 35, 38, 64, 37, 26, 80, 62, 0, 27, 65, 63, 46, 33, 29, 
    0, 36, 71, 32, 6, 0, 85, 55, 18, 26, 40, 34, 21, 17, 21, 
    0, 49, 67, 41, 34, 25, 23, 16, 29, 25, 22, 4, 38, 4, 3, 
    15, 13, 11, 1, 10, 13, 9, 15, 0, 35, 13, 10, 9, 0, 1, 
    4, 0, 0, 0, 0, 0, 4, 19, 0, 62, 2, 6, 0, 0, 35, 
    
    -- channel=44
    165, 88, 125, 152, 159, 160, 166, 190, 151, 174, 183, 170, 182, 179, 165, 
    171, 98, 126, 166, 162, 167, 167, 172, 156, 218, 110, 156, 189, 183, 159, 
    177, 98, 122, 170, 161, 166, 181, 141, 133, 258, 31, 136, 193, 174, 150, 
    172, 94, 131, 147, 169, 149, 176, 159, 148, 145, 52, 67, 73, 151, 130, 
    101, 82, 95, 74, 110, 104, 112, 149, 108, 84, 63, 54, 38, 137, 76, 
    24, 35, 89, 38, 66, 63, 71, 104, 73, 79, 21, 80, 159, 93, 121, 
    42, 71, 74, 20, 64, 105, 90, 94, 79, 83, 50, 118, 190, 85, 155, 
    67, 75, 64, 60, 91, 109, 122, 128, 120, 157, 78, 101, 127, 176, 66, 
    86, 92, 53, 97, 124, 127, 124, 124, 93, 144, 59, 101, 118, 124, 107, 
    91, 41, 75, 104, 102, 100, 108, 121, 100, 111, 110, 135, 127, 122, 71, 
    64, 91, 98, 115, 80, 87, 149, 111, 17, 90, 118, 117, 90, 66, 57, 
    14, 90, 130, 78, 56, 29, 133, 87, 55, 76, 78, 66, 56, 39, 43, 
    24, 82, 100, 65, 63, 65, 64, 50, 54, 57, 54, 24, 59, 22, 20, 
    32, 33, 32, 21, 31, 35, 35, 46, 11, 59, 34, 28, 26, 13, 18, 
    19, 7, 11, 13, 17, 20, 24, 42, 0, 88, 18, 21, 12, 9, 49, 
    
    -- channel=45
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=46
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 26, 0, 0, 0, 0, 0, 
    7, 0, 15, 13, 8, 0, 0, 0, 58, 39, 26, 80, 30, 23, 30, 
    59, 50, 52, 60, 67, 62, 43, 25, 0, 0, 0, 0, 0, 14, 48, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 53, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 19, 0, 0, 0, 0, 
    0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 33, 47, 35, 
    0, 0, 0, 0, 14, 0, 0, 16, 0, 2, 34, 32, 16, 9, 21, 
    0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 9, 9, 0, 10, 12, 
    0, 21, 25, 16, 25, 23, 0, 0, 14, 15, 0, 1, 15, 1, 0, 
    32, 26, 10, 0, 4, 10, 6, 2, 0, 0, 5, 6, 1, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 10, 0, 10, 4, 4, 0, 0, 28, 
    
    -- channel=47
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 7, 0, 18, 21, 0, 0, 0, 
    5, 8, 21, 14, 0, 0, 0, 3, 13, 0, 0, 0, 32, 29, 22, 
    29, 27, 15, 32, 35, 38, 27, 17, 5, 2, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 0, 0, 0, 0, 0, 
    14, 16, 0, 0, 7, 10, 0, 0, 0, 0, 0, 0, 0, 2, 9, 
    0, 0, 2, 0, 0, 0, 0, 21, 20, 0, 0, 10, 23, 16, 9, 
    1, 0, 0, 17, 27, 5, 0, 0, 0, 18, 24, 6, 10, 2, 11, 
    0, 0, 0, 0, 0, 0, 24, 19, 0, 0, 10, 0, 0, 0, 0, 
    18, 32, 26, 25, 6, 0, 0, 3, 13, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=48
    35, 1, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 10, 3, 0, 
    29, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    26, 0, 0, 0, 0, 8, 0, 7, 0, 0, 0, 0, 0, 0, 0, 
    20, 2, 0, 2, 0, 0, 0, 8, 0, 0, 11, 5, 37, 0, 0, 
    8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 
    8, 0, 0, 7, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 0, 0, 0, 0, 12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 0, 0, 0, 0, 0, 11, 3, 0, 0, 0, 0, 0, 0, 0, 
    30, 0, 0, 0, 15, 0, 61, 136, 41, 0, 70, 31, 136, 31, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 
    0, 0, 0, 0, 0, 18, 3, 13, 1, 7, 0, 0, 22, 64, 0, 
    
    -- channel=49
    393, 439, 389, 366, 391, 411, 404, 400, 403, 407, 411, 406, 426, 456, 465, 
    394, 445, 436, 323, 315, 332, 324, 333, 339, 346, 349, 368, 452, 465, 471, 
    389, 432, 424, 310, 327, 315, 294, 323, 344, 346, 346, 354, 438, 468, 477, 
    386, 428, 400, 301, 331, 342, 329, 335, 345, 337, 342, 360, 385, 457, 466, 
    405, 426, 428, 387, 358, 355, 362, 376, 373, 366, 370, 421, 440, 457, 460, 
    438, 415, 382, 431, 427, 421, 433, 439, 427, 427, 432, 443, 455, 459, 465, 
    455, 409, 298, 253, 342, 440, 461, 467, 464, 453, 452, 451, 453, 455, 461, 
    471, 478, 451, 325, 176, 272, 406, 468, 462, 449, 450, 450, 453, 451, 454, 
    478, 490, 487, 468, 178, 134, 184, 257, 336, 397, 442, 457, 453, 450, 453, 
    478, 482, 485, 441, 153, 64, 100, 126, 146, 142, 180, 265, 348, 418, 451, 
    468, 475, 479, 437, 327, 210, 176, 275, 325, 228, 245, 214, 326, 403, 430, 
    342, 342, 327, 317, 312, 275, 267, 319, 329, 302, 327, 321, 341, 339, 344, 
    205, 212, 198, 185, 175, 165, 163, 183, 174, 165, 162, 163, 170, 164, 154, 
    102, 110, 101, 98, 90, 80, 80, 85, 85, 70, 68, 68, 68, 80, 155, 
    67, 73, 73, 74, 70, 88, 87, 95, 96, 88, 73, 70, 110, 175, 158, 
    
    -- channel=50
    103, 109, 68, 80, 95, 91, 83, 87, 81, 87, 88, 87, 96, 105, 108, 
    109, 120, 96, 60, 112, 121, 107, 121, 115, 116, 119, 118, 119, 117, 116, 
    107, 114, 114, 82, 64, 74, 62, 84, 74, 73, 77, 89, 123, 114, 120, 
    98, 112, 77, 62, 81, 84, 66, 82, 87, 81, 89, 83, 116, 116, 121, 
    93, 111, 101, 84, 89, 92, 89, 97, 97, 88, 92, 115, 105, 111, 115, 
    101, 107, 110, 101, 78, 79, 88, 91, 83, 81, 85, 105, 112, 110, 113, 
    109, 61, 20, 122, 158, 126, 117, 117, 111, 106, 113, 111, 114, 117, 122, 
    123, 116, 72, 0, 15, 148, 156, 123, 115, 109, 110, 108, 109, 107, 113, 
    126, 122, 114, 96, 0, 15, 76, 149, 154, 130, 124, 110, 111, 112, 114, 
    124, 120, 118, 110, 0, 1, 9, 3, 17, 60, 138, 158, 150, 127, 117, 
    129, 119, 120, 65, 0, 0, 0, 20, 0, 0, 0, 0, 53, 75, 114, 
    143, 141, 138, 141, 145, 105, 91, 122, 128, 99, 112, 98, 111, 127, 127, 
    31, 37, 28, 23, 20, 17, 24, 54, 54, 60, 62, 72, 78, 73, 73, 
    9, 27, 20, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=51
    32, 49, 48, 40, 39, 39, 35, 38, 37, 37, 36, 37, 39, 32, 33, 
    36, 49, 52, 38, 19, 26, 21, 25, 26, 25, 24, 36, 35, 40, 37, 
    37, 47, 54, 53, 28, 25, 30, 29, 35, 30, 32, 31, 31, 34, 39, 
    38, 51, 43, 26, 24, 26, 27, 24, 23, 22, 16, 20, 27, 37, 42, 
    36, 48, 56, 43, 43, 43, 47, 45, 42, 43, 37, 46, 43, 45, 45, 
    31, 39, 47, 55, 47, 50, 48, 48, 48, 45, 44, 40, 46, 44, 45, 
    28, 49, 34, 22, 42, 48, 47, 47, 46, 43, 43, 43, 43, 42, 44, 
    25, 41, 45, 31, 18, 27, 37, 40, 42, 43, 41, 43, 44, 45, 47, 
    20, 33, 35, 37, 36, 15, 9, 19, 30, 35, 47, 46, 43, 43, 47, 
    17, 31, 35, 25, 43, 20, 20, 18, 10, 16, 27, 24, 30, 39, 45, 
    22, 38, 35, 39, 54, 29, 33, 38, 24, 43, 29, 31, 26, 31, 37, 
    16, 31, 28, 27, 28, 40, 34, 34, 48, 56, 48, 56, 51, 61, 57, 
    25, 42, 38, 32, 25, 29, 33, 32, 35, 34, 34, 33, 34, 34, 32, 
    18, 24, 23, 20, 14, 18, 20, 17, 13, 13, 13, 13, 14, 13, 17, 
    13, 18, 17, 14, 15, 19, 16, 14, 13, 15, 11, 8, 11, 9, 0, 
    
    -- channel=52
    30, 13, 0, 19, 28, 16, 17, 21, 20, 20, 19, 20, 26, 32, 32, 
    21, 8, 5, 47, 66, 73, 70, 73, 73, 70, 70, 70, 34, 28, 28, 
    19, 5, 8, 64, 76, 79, 84, 91, 76, 74, 73, 69, 61, 27, 25, 
    15, 4, 19, 55, 57, 58, 53, 63, 52, 54, 65, 48, 57, 20, 20, 
    13, 6, 6, 15, 17, 15, 13, 23, 20, 20, 25, 34, 23, 18, 17, 
    22, 14, 16, 12, 12, 11, 18, 20, 16, 15, 20, 20, 16, 17, 17, 
    28, 0, 0, 43, 40, 23, 19, 18, 18, 18, 22, 19, 19, 20, 20, 
    32, 17, 16, 0, 24, 56, 47, 29, 22, 19, 22, 19, 18, 16, 14, 
    39, 29, 27, 29, 0, 32, 45, 55, 53, 39, 27, 18, 19, 17, 15, 
    43, 33, 28, 28, 0, 28, 33, 34, 32, 25, 41, 51, 51, 36, 23, 
    43, 28, 29, 10, 0, 0, 2, 35, 14, 6, 1, 1, 35, 31, 28, 
    56, 41, 40, 42, 43, 30, 38, 39, 22, 6, 24, 12, 17, 9, 10, 
    26, 18, 18, 23, 26, 25, 26, 32, 22, 26, 25, 27, 28, 25, 27, 
    24, 24, 20, 24, 24, 23, 22, 25, 25, 24, 25, 25, 25, 22, 16, 
    26, 24, 23, 26, 24, 24, 23, 27, 23, 22, 24, 30, 22, 13, 15, 
    
    -- channel=53
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 47, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 19, 47, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 31, 51, 45, 9, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 28, 28, 17, 28, 41, 53, 33, 8, 0, 0, 
    6, 0, 0, 0, 0, 0, 14, 22, 0, 0, 0, 6, 32, 6, 0, 
    15, 4, 6, 8, 9, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 1, 6, 3, 5, 14, 5, 12, 11, 15, 14, 10, 14, 
    20, 29, 27, 30, 31, 30, 30, 32, 31, 30, 33, 30, 29, 27, 38, 
    10, 24, 25, 30, 25, 26, 24, 28, 25, 27, 28, 34, 28, 52, 50, 
    
    -- channel=54
    133, 154, 134, 120, 124, 131, 126, 123, 124, 127, 128, 126, 127, 132, 137, 
    146, 171, 152, 76, 70, 80, 76, 80, 78, 80, 86, 90, 131, 142, 144, 
    146, 169, 158, 46, 46, 29, 25, 24, 38, 46, 46, 59, 123, 148, 149, 
    143, 165, 131, 27, 58, 72, 52, 60, 68, 66, 64, 71, 93, 151, 154, 
    144, 163, 153, 133, 125, 126, 129, 128, 128, 126, 124, 135, 133, 153, 154, 
    147, 156, 150, 145, 135, 131, 133, 133, 130, 134, 134, 144, 154, 150, 154, 
    147, 138, 111, 134, 142, 152, 153, 153, 150, 147, 149, 149, 153, 154, 154, 
    153, 160, 128, 58, 70, 133, 144, 150, 149, 144, 145, 146, 150, 149, 155, 
    154, 154, 150, 136, 43, 54, 92, 131, 132, 137, 145, 147, 150, 152, 155, 
    148, 147, 148, 147, 53, 39, 40, 35, 57, 95, 126, 136, 135, 139, 148, 
    147, 147, 149, 127, 52, 23, 45, 54, 52, 39, 39, 47, 87, 116, 141, 
    136, 142, 139, 139, 140, 119, 106, 128, 145, 121, 136, 123, 141, 150, 147, 
    69, 78, 74, 69, 66, 64, 66, 86, 89, 91, 93, 98, 102, 99, 98, 
    49, 63, 59, 52, 45, 44, 43, 42, 40, 33, 33, 32, 32, 32, 54, 
    17, 31, 31, 30, 26, 30, 27, 27, 29, 27, 25, 26, 33, 72, 91, 
    
    -- channel=55
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 35, 29, 34, 38, 42, 41, 32, 36, 41, 0, 0, 0, 
    0, 0, 0, 36, 12, 10, 33, 21, 12, 11, 10, 11, 4, 0, 0, 
    0, 0, 0, 12, 6, 10, 6, 7, 4, 11, 8, 1, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 31, 16, 15, 9, 3, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 35, 21, 20, 24, 20, 17, 6, 3, 0, 0, 0, 
    0, 0, 0, 5, 23, 18, 16, 14, 10, 28, 13, 20, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 2, 6, 8, 2, 0, 0, 1, 1, 1, 1, 1, 5, 
    38, 23, 24, 28, 32, 30, 26, 29, 28, 30, 30, 27, 27, 24, 16, 
    43, 25, 24, 26, 31, 30, 30, 33, 35, 34, 34, 32, 24, 10, 24, 
    
    -- channel=56
    48, 15, 0, 5, 27, 4, 0, 6, 0, 3, 1, 1, 18, 9, 5, 
    45, 29, 0, 0, 38, 43, 18, 45, 29, 33, 29, 51, 26, 9, 10, 
    46, 21, 3, 0, 0, 0, 0, 15, 0, 0, 0, 14, 44, 7, 12, 
    30, 22, 0, 0, 0, 0, 0, 7, 0, 0, 8, 0, 44, 11, 15, 
    3, 19, 1, 0, 10, 14, 14, 14, 8, 0, 14, 45, 1, 10, 10, 
    7, 0, 16, 18, 0, 0, 0, 0, 0, 0, 0, 11, 8, 5, 11, 
    21, 0, 0, 56, 109, 45, 12, 3, 0, 0, 7, 2, 8, 10, 16, 
    35, 0, 0, 0, 0, 125, 101, 21, 0, 0, 5, 1, 3, 1, 9, 
    35, 9, 0, 0, 0, 31, 83, 107, 89, 45, 40, 1, 0, 5, 10, 
    35, 10, 5, 0, 0, 22, 34, 18, 28, 38, 122, 102, 90, 52, 18, 
    43, 9, 6, 0, 0, 0, 0, 50, 0, 0, 0, 0, 68, 18, 20, 
    69, 44, 45, 50, 59, 3, 34, 78, 34, 23, 37, 22, 38, 41, 41, 
    6, 2, 0, 0, 0, 0, 6, 30, 8, 24, 25, 36, 36, 26, 37, 
    2, 27, 16, 21, 8, 13, 16, 17, 3, 0, 8, 5, 7, 9, 22, 
    0, 2, 2, 8, 0, 8, 0, 6, 0, 0, 0, 0, 19, 8, 0, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 38, 38, 33, 31, 35, 36, 37, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 8, 1, 0, 5, 3, 0, 0, 0, 0, 0, 
    0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 95, 125, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 116, 87, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 79, 152, 135, 63, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 24, 37, 24, 2, 25, 96, 173, 179, 133, 50, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    120, 124, 139, 149, 159, 127, 83, 91, 105, 68, 69, 51, 58, 79, 77, 
    5, 0, 0, 0, 0, 1, 5, 31, 49, 60, 68, 78, 84, 84, 92, 
    52, 55, 50, 41, 34, 34, 27, 25, 16, 13, 12, 9, 10, 3, 0, 
    7, 3, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 
    
    -- channel=58
    98, 104, 85, 98, 101, 104, 102, 105, 108, 107, 107, 106, 122, 136, 131, 
    88, 91, 92, 101, 99, 90, 88, 99, 100, 97, 97, 108, 113, 116, 123, 
    84, 85, 89, 121, 126, 142, 140, 152, 150, 151, 150, 155, 121, 118, 119, 
    85, 83, 87, 124, 106, 108, 115, 117, 104, 97, 105, 101, 128, 103, 109, 
    86, 85, 93, 88, 81, 79, 78, 93, 84, 82, 93, 111, 117, 110, 105, 
    98, 90, 72, 90, 115, 114, 121, 119, 114, 114, 120, 117, 103, 108, 111, 
    110, 71, 62, 46, 47, 89, 107, 109, 110, 107, 108, 105, 105, 105, 105, 
    117, 109, 117, 108, 66, 58, 83, 108, 109, 104, 109, 106, 107, 105, 103, 
    124, 123, 125, 118, 27, 49, 47, 39, 57, 79, 98, 110, 106, 103, 101, 
    126, 127, 123, 113, 0, 19, 38, 51, 46, 4, 3, 26, 58, 89, 104, 
    119, 123, 121, 85, 111, 93, 74, 135, 138, 96, 111, 92, 142, 131, 110, 
    65, 58, 49, 44, 40, 22, 57, 71, 39, 45, 60, 57, 62, 42, 49, 
    52, 52, 52, 53, 55, 45, 45, 42, 18, 14, 8, 7, 3, 0, 0, 
    7, 9, 4, 15, 20, 13, 16, 21, 24, 24, 26, 28, 29, 31, 69, 
    25, 31, 30, 36, 32, 40, 43, 51, 45, 46, 42, 41, 43, 82, 38, 
    
    -- channel=59
    1, 39, 74, 47, 30, 42, 49, 37, 43, 40, 42, 43, 27, 40, 54, 
    8, 37, 68, 116, 43, 78, 93, 72, 91, 83, 88, 70, 43, 58, 57, 
    9, 41, 65, 103, 65, 26, 61, 27, 45, 47, 41, 39, 51, 56, 56, 
    17, 40, 81, 39, 31, 37, 43, 29, 37, 57, 27, 38, 0, 53, 53, 
    38, 39, 51, 76, 44, 47, 43, 39, 51, 55, 38, 12, 56, 55, 58, 
    43, 63, 75, 49, 49, 47, 43, 52, 59, 52, 45, 46, 57, 56, 53, 
    33, 89, 72, 17, 29, 51, 54, 61, 64, 69, 59, 64, 60, 60, 57, 
    22, 63, 75, 112, 43, 0, 30, 61, 66, 67, 56, 61, 58, 59, 54, 
    24, 60, 67, 78, 193, 0, 0, 8, 51, 69, 50, 61, 62, 61, 59, 
    25, 58, 62, 85, 220, 5, 0, 9, 8, 21, 0, 38, 52, 59, 58, 
    19, 60, 61, 111, 49, 74, 0, 0, 26, 35, 0, 0, 0, 10, 33, 
    44, 84, 85, 82, 78, 104, 63, 36, 69, 69, 51, 61, 51, 53, 55, 
    29, 35, 38, 38, 34, 40, 33, 26, 58, 49, 54, 48, 53, 65, 56, 
    36, 21, 25, 15, 20, 13, 10, 9, 12, 13, 3, 5, 4, 0, 0, 
    33, 8, 5, 0, 8, 0, 5, 0, 7, 1, 7, 4, 0, 0, 51, 
    
    -- channel=60
    70, 127, 158, 125, 103, 135, 138, 124, 129, 127, 133, 132, 118, 133, 141, 
    74, 118, 158, 184, 110, 125, 143, 123, 139, 132, 137, 115, 122, 149, 148, 
    77, 119, 154, 156, 128, 89, 115, 79, 105, 113, 98, 95, 104, 149, 148, 
    84, 115, 180, 136, 119, 119, 132, 113, 126, 157, 124, 137, 79, 147, 142, 
    111, 116, 140, 156, 117, 119, 117, 115, 125, 133, 114, 95, 134, 141, 141, 
    122, 138, 138, 130, 128, 127, 123, 135, 139, 132, 127, 123, 143, 145, 139, 
    119, 173, 157, 71, 85, 126, 140, 149, 152, 154, 143, 148, 145, 147, 143, 
    112, 152, 176, 194, 73, 26, 95, 146, 154, 156, 144, 148, 144, 146, 138, 
    113, 151, 161, 175, 252, 35, 22, 62, 107, 132, 126, 149, 148, 147, 141, 
    114, 151, 157, 182, 271, 29, 28, 45, 42, 62, 32, 92, 106, 126, 136, 
    105, 153, 153, 207, 144, 132, 31, 0, 102, 91, 58, 61, 0, 85, 118, 
    93, 141, 141, 137, 130, 159, 100, 78, 129, 131, 105, 120, 103, 118, 121, 
    64, 81, 80, 77, 71, 70, 60, 51, 88, 74, 78, 72, 78, 90, 77, 
    61, 56, 62, 49, 55, 43, 41, 40, 48, 43, 33, 36, 32, 31, 0, 
    55, 37, 36, 29, 38, 24, 37, 28, 40, 35, 36, 34, 16, 14, 76, 
    
    -- channel=61
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=62
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 42, 52, 77, 77, 60, 71, 68, 59, 29, 0, 0, 0, 
    0, 0, 0, 33, 15, 0, 16, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 23, 10, 4, 7, 13, 22, 31, 19, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 64, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 17, 50, 16, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 12, 57, 82, 59, 21, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 67, 32, 15, 7, 29, 77, 101, 95, 53, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 71, 79, 83, 88, 63, 35, 41, 53, 23, 26, 9, 24, 37, 31, 
    0, 0, 0, 0, 0, 0, 0, 20, 36, 42, 49, 52, 58, 66, 67, 
    45, 48, 43, 34, 31, 28, 25, 21, 15, 13, 8, 7, 8, 0, 0, 
    12, 7, 4, 3, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    
    -- channel=63
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 10, 18, 11, 14, 17, 16, 19, 28, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 41, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 35, 35, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 38, 60, 32, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 0, 0, 4, 0, 0, 0, 32, 69, 63, 24, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    60, 71, 74, 77, 79, 70, 74, 62, 43, 51, 44, 44, 35, 29, 34, 
    0, 0, 3, 10, 13, 14, 19, 24, 25, 27, 28, 30, 32, 32, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=64
    12, 0, 47, 7, 0, 75, 0, 4, 1, 0, 0, 66, 0, 37, 16, 
    0, 0, 0, 10, 0, 37, 0, 44, 0, 13, 0, 100, 0, 71, 0, 
    0, 0, 0, 0, 0, 73, 43, 0, 2, 0, 63, 76, 0, 5, 14, 
    0, 114, 0, 0, 0, 78, 0, 0, 100, 0, 82, 58, 0, 0, 0, 
    0, 120, 0, 0, 65, 7, 0, 86, 11, 42, 4, 0, 0, 0, 0, 
    0, 107, 0, 0, 74, 6, 0, 47, 0, 0, 0, 63, 0, 0, 0, 
    0, 70, 13, 0, 0, 0, 0, 5, 0, 0, 0, 16, 0, 18, 0, 
    0, 45, 23, 0, 19, 0, 35, 9, 0, 14, 0, 14, 0, 1, 0, 
    10, 21, 0, 0, 3, 0, 3, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 39, 0, 0, 0, 19, 0, 0, 0, 0, 0, 2, 49, 
    0, 57, 0, 36, 12, 0, 86, 0, 0, 0, 0, 0, 0, 0, 24, 
    37, 76, 0, 22, 0, 29, 36, 1, 0, 0, 28, 0, 0, 3, 0, 
    0, 13, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 60, 9, 0, 0, 0, 0, 46, 4, 0, 0, 0, 76, 18, 
    0, 5, 64, 54, 0, 0, 0, 1, 0, 0, 0, 0, 0, 31, 131, 
    
    -- channel=65
    124, 47, 101, 113, 18, 51, 98, 102, 156, 162, 129, 184, 134, 87, 106, 
    181, 119, 135, 133, 4, 33, 69, 105, 155, 149, 129, 212, 199, 155, 173, 
    126, 117, 132, 107, 0, 73, 140, 121, 151, 76, 148, 249, 293, 223, 222, 
    82, 180, 147, 87, 41, 192, 168, 37, 128, 99, 212, 269, 319, 267, 183, 
    100, 271, 220, 88, 152, 235, 116, 107, 210, 223, 243, 251, 305, 281, 109, 
    76, 244, 305, 174, 219, 219, 158, 255, 249, 240, 215, 252, 286, 280, 94, 
    106, 212, 279, 295, 224, 220, 203, 231, 208, 219, 230, 266, 256, 283, 134, 
    140, 215, 253, 291, 288, 162, 244, 257, 263, 262, 243, 299, 262, 261, 85, 
    203, 247, 228, 250, 284, 252, 260, 280, 290, 294, 270, 275, 248, 190, 111, 
    232, 203, 140, 195, 220, 255, 286, 318, 315, 316, 269, 266, 191, 134, 202, 
    167, 187, 153, 216, 215, 204, 324, 356, 325, 282, 269, 258, 209, 204, 264, 
    267, 357, 250, 230, 224, 251, 320, 338, 323, 271, 299, 260, 210, 218, 265, 
    241, 356, 377, 301, 235, 259, 301, 222, 251, 302, 312, 252, 180, 155, 228, 
    131, 105, 316, 382, 326, 263, 258, 215, 232, 295, 296, 233, 98, 123, 250, 
    121, 49, 135, 343, 400, 369, 310, 291, 202, 229, 223, 205, 142, 193, 322, 
    
    -- channel=66
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 16, 22, 2, 0, 
    0, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 11, 19, 0, 
    0, 59, 18, 0, 0, 3, 0, 0, 0, 0, 0, 4, 0, 27, 0, 
    0, 16, 42, 6, 0, 12, 0, 10, 16, 24, 8, 12, 0, 13, 0, 
    0, 11, 12, 27, 7, 0, 33, 29, 4, 0, 18, 57, 0, 12, 0, 
    0, 0, 16, 19, 75, 0, 40, 34, 29, 47, 31, 39, 46, 12, 0, 
    9, 5, 0, 16, 4, 94, 29, 41, 52, 38, 31, 26, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 87, 56, 45, 49, 38, 26, 0, 0, 3, 
    0, 0, 0, 0, 0, 25, 56, 67, 57, 23, 38, 31, 0, 14, 0, 
    59, 104, 0, 0, 0, 35, 50, 46, 83, 40, 59, 12, 0, 2, 0, 
    0, 32, 92, 18, 0, 0, 3, 0, 15, 62, 44, 23, 0, 0, 0, 
    0, 0, 36, 85, 31, 0, 0, 0, 7, 56, 60, 7, 0, 0, 42, 
    
    -- channel=67
    0, 11, 0, 2, 10, 0, 0, 1, 0, 0, 0, 0, 0, 0, 5, 
    7, 1, 0, 3, 16, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 8, 22, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 7, 17, 0, 0, 8, 0, 18, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    10, 0, 0, 10, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    3, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 
    
    -- channel=68
    19, 12, 22, 5, 0, 31, 21, 27, 35, 29, 9, 41, 10, 34, 14, 
    23, 15, 17, 6, 0, 31, 16, 26, 21, 26, 15, 50, 11, 37, 17, 
    19, 13, 8, 13, 0, 28, 25, 22, 18, 5, 25, 57, 26, 20, 22, 
    1, 29, 20, 5, 14, 38, 19, 3, 38, 0, 53, 44, 33, 25, 8, 
    3, 48, 0, 29, 35, 32, 5, 26, 39, 41, 41, 47, 40, 23, 0, 
    5, 53, 24, 0, 36, 48, 50, 51, 30, 38, 35, 46, 37, 23, 0, 
    0, 42, 36, 19, 57, 74, 59, 67, 57, 67, 61, 58, 34, 29, 0, 
    6, 30, 20, 33, 46, 63, 69, 77, 74, 69, 70, 71, 37, 30, 0, 
    21, 32, 29, 30, 77, 25, 84, 72, 71, 69, 72, 71, 71, 46, 0, 
    25, 24, 3, 26, 21, 88, 61, 63, 76, 70, 61, 66, 36, 12, 35, 
    5, 26, 17, 35, 36, 8, 84, 74, 57, 69, 66, 65, 54, 36, 21, 
    24, 52, 22, 35, 11, 51, 68, 79, 69, 55, 73, 74, 61, 44, 13, 
    48, 73, 38, 35, 25, 45, 73, 76, 74, 63, 83, 63, 53, 42, 11, 
    8, 53, 67, 44, 38, 33, 46, 27, 61, 76, 62, 70, 33, 21, 18, 
    18, 10, 75, 78, 53, 32, 27, 35, 48, 76, 76, 45, 13, 27, 64, 
    
    -- channel=69
    38, 28, 58, 57, 33, 74, 51, 56, 74, 59, 42, 72, 21, 69, 40, 
    39, 36, 48, 54, 24, 74, 46, 68, 44, 63, 42, 84, 0, 61, 42, 
    54, 41, 41, 46, 18, 62, 64, 65, 53, 47, 62, 78, 22, 54, 54, 
    37, 71, 48, 28, 30, 90, 81, 33, 89, 5, 83, 84, 35, 45, 32, 
    38, 87, 10, 49, 55, 62, 25, 60, 66, 70, 79, 73, 44, 41, 10, 
    18, 94, 42, 4, 87, 52, 2, 44, 48, 57, 39, 68, 41, 46, 0, 
    12, 78, 63, 40, 35, 22, 5, 39, 27, 16, 6, 37, 19, 63, 0, 
    34, 62, 54, 49, 0, 16, 28, 18, 0, 11, 26, 5, 6, 39, 12, 
    38, 63, 48, 51, 62, 0, 25, 0, 15, 15, 5, 20, 18, 25, 4, 
    51, 42, 38, 68, 30, 61, 0, 5, 8, 2, 7, 10, 0, 32, 62, 
    28, 54, 36, 60, 75, 22, 53, 10, 0, 11, 9, 6, 9, 27, 60, 
    29, 48, 29, 75, 33, 69, 42, 14, 0, 0, 17, 10, 17, 33, 64, 
    79, 67, 29, 52, 52, 54, 46, 18, 23, 0, 12, 0, 10, 46, 79, 
    45, 102, 93, 43, 52, 64, 70, 15, 62, 22, 0, 9, 0, 76, 58, 
    40, 42, 129, 97, 39, 49, 64, 73, 51, 35, 26, 0, 13, 62, 111, 
    
    -- channel=70
    44, 16, 46, 66, 40, 32, 45, 42, 68, 63, 59, 58, 46, 46, 38, 
    62, 31, 60, 70, 25, 36, 45, 46, 54, 58, 56, 67, 43, 44, 63, 
    70, 50, 59, 63, 15, 25, 47, 64, 67, 54, 59, 72, 81, 77, 82, 
    47, 59, 60, 39, 10, 65, 78, 32, 64, 22, 67, 81, 104, 86, 86, 
    50, 102, 67, 44, 34, 73, 42, 24, 64, 61, 83, 75, 91, 98, 65, 
    34, 105, 104, 39, 74, 59, 11, 55, 61, 67, 53, 53, 86, 105, 44, 
    28, 85, 104, 92, 46, 20, 5, 43, 39, 29, 21, 45, 59, 97, 46, 
    56, 81, 89, 98, 37, 13, 35, 27, 13, 18, 35, 46, 45, 80, 49, 
    60, 85, 91, 93, 92, 19, 37, 31, 39, 46, 31, 47, 61, 56, 32, 
    86, 81, 64, 85, 68, 85, 39, 48, 48, 49, 37, 41, 29, 44, 70, 
    73, 60, 54, 79, 84, 53, 79, 68, 54, 55, 41, 35, 33, 55, 94, 
    58, 64, 45, 87, 82, 87, 75, 61, 58, 43, 46, 32, 22, 52, 109, 
    106, 111, 76, 67, 73, 87, 80, 49, 57, 44, 53, 29, 20, 46, 107, 
    60, 74, 107, 85, 70, 72, 80, 46, 58, 59, 41, 36, 16, 57, 84, 
    54, 15, 77, 105, 91, 79, 78, 88, 59, 57, 54, 30, 21, 61, 95, 
    
    -- channel=71
    28, 45, 27, 29, 37, 28, 38, 40, 40, 47, 45, 40, 55, 34, 43, 
    39, 49, 39, 27, 45, 27, 36, 37, 37, 38, 43, 34, 57, 32, 31, 
    29, 41, 39, 33, 48, 33, 43, 40, 37, 44, 31, 41, 43, 40, 36, 
    38, 23, 40, 39, 53, 35, 56, 65, 30, 52, 31, 52, 46, 40, 23, 
    44, 12, 37, 41, 38, 51, 61, 46, 42, 50, 53, 65, 54, 29, 36, 
    48, 12, 31, 53, 41, 68, 61, 35, 58, 69, 66, 57, 56, 31, 48, 
    48, 23, 36, 40, 65, 59, 68, 56, 60, 53, 51, 57, 60, 35, 54, 
    45, 29, 32, 30, 47, 63, 48, 59, 59, 62, 59, 41, 50, 38, 56, 
    41, 36, 42, 37, 36, 45, 48, 50, 50, 54, 62, 53, 45, 41, 47, 
    30, 43, 43, 26, 33, 37, 42, 39, 50, 44, 54, 52, 48, 33, 37, 
    41, 37, 52, 28, 40, 40, 34, 44, 40, 46, 48, 56, 57, 47, 20, 
    51, 45, 73, 53, 42, 34, 38, 51, 45, 48, 43, 53, 61, 50, 43, 
    32, 44, 70, 82, 65, 39, 38, 44, 42, 48, 43, 57, 52, 55, 43, 
    40, 44, 43, 73, 81, 73, 59, 58, 40, 43, 47, 57, 53, 31, 57, 
    44, 43, 38, 50, 68, 75, 73, 70, 66, 35, 34, 49, 56, 44, 41, 
    
    -- channel=72
    0, 0, 10, 5, 0, 75, 0, 35, 14, 35, 0, 109, 0, 69, 1, 
    0, 0, 0, 7, 0, 63, 13, 49, 0, 18, 0, 135, 0, 33, 0, 
    0, 30, 0, 0, 0, 43, 0, 0, 49, 0, 39, 121, 0, 0, 0, 
    0, 71, 0, 0, 0, 42, 0, 0, 76, 0, 37, 75, 0, 0, 0, 
    0, 115, 0, 0, 65, 5, 0, 48, 0, 13, 0, 72, 0, 0, 0, 
    0, 128, 1, 0, 37, 25, 0, 35, 0, 13, 0, 80, 0, 17, 0, 
    0, 67, 63, 0, 0, 11, 0, 5, 1, 16, 7, 16, 0, 24, 0, 
    0, 55, 31, 3, 0, 0, 46, 0, 0, 0, 0, 47, 0, 12, 0, 
    4, 14, 8, 18, 57, 0, 27, 2, 1, 13, 0, 17, 0, 0, 0, 
    0, 0, 0, 47, 21, 70, 7, 11, 0, 0, 0, 0, 0, 0, 38, 
    0, 55, 0, 36, 4, 0, 94, 0, 0, 0, 8, 0, 0, 0, 6, 
    0, 0, 0, 19, 0, 37, 51, 15, 0, 0, 9, 0, 0, 29, 0, 
    54, 114, 0, 0, 0, 44, 24, 0, 88, 0, 4, 0, 0, 44, 1, 
    0, 96, 152, 6, 0, 0, 0, 0, 47, 27, 11, 0, 0, 65, 34, 
    0, 0, 128, 136, 0, 0, 0, 0, 0, 30, 30, 0, 0, 0, 108, 
    
    -- channel=73
    0, 0, 0, 0, 0, 0, 0, 12, 16, 42, 2, 8, 0, 34, 0, 
    0, 0, 0, 0, 0, 28, 32, 0, 0, 0, 0, 2, 0, 0, 0, 
    43, 51, 3, 15, 5, 0, 0, 0, 38, 22, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 51, 0, 0, 0, 0, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 0, 0, 0, 
    12, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 0, 
    0, 0, 31, 0, 0, 0, 0, 0, 1, 1, 0, 0, 10, 0, 0, 
    3, 4, 0, 4, 0, 0, 0, 0, 0, 0, 0, 6, 0, 9, 25, 
    0, 0, 36, 33, 42, 0, 0, 0, 0, 0, 0, 0, 36, 59, 0, 
    0, 48, 22, 23, 25, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 6, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 3, 0, 0, 0, 7, 18, 15, 
    77, 113, 0, 0, 0, 10, 14, 69, 89, 0, 0, 0, 0, 63, 19, 
    0, 115, 123, 0, 0, 0, 0, 0, 0, 10, 0, 3, 53, 17, 0, 
    1, 0, 71, 97, 0, 0, 0, 0, 19, 51, 80, 40, 0, 0, 0, 
    
    -- channel=74
    52, 32, 63, 40, 0, 55, 51, 58, 76, 64, 38, 100, 37, 46, 52, 
    70, 72, 48, 47, 0, 40, 17, 70, 62, 78, 39, 119, 55, 104, 68, 
    43, 33, 40, 35, 0, 63, 87, 62, 46, 25, 55, 133, 97, 89, 84, 
    14, 94, 66, 27, 37, 116, 73, 0, 83, 26, 116, 140, 88, 98, 33, 
    38, 117, 58, 49, 96, 104, 31, 89, 101, 122, 111, 110, 106, 89, 0, 
    20, 101, 90, 61, 123, 104, 81, 133, 117, 107, 85, 149, 103, 78, 0, 
    43, 95, 98, 101, 109, 119, 109, 115, 94, 111, 114, 136, 90, 110, 20, 
    44, 83, 102, 97, 127, 100, 122, 134, 132, 140, 128, 125, 116, 87, 0, 
    82, 110, 73, 77, 125, 101, 140, 126, 141, 126, 121, 132, 86, 62, 25, 
    92, 58, 42, 75, 66, 103, 126, 142, 138, 133, 122, 118, 63, 51, 88, 
    30, 83, 58, 81, 105, 77, 148, 144, 126, 112, 112, 111, 93, 74, 109, 
    109, 186, 115, 104, 63, 107, 143, 139, 119, 110, 137, 126, 100, 95, 77, 
    88, 115, 145, 141, 92, 104, 131, 88, 87, 120, 136, 108, 90, 67, 80, 
    41, 62, 114, 146, 149, 119, 108, 75, 139, 126, 123, 107, 19, 75, 76, 
    36, 38, 104, 141, 149, 164, 142, 119, 89, 95, 89, 64, 69, 82, 183, 
    
    -- channel=75
    2, 20, 0, 0, 62, 0, 3, 0, 0, 0, 45, 0, 120, 0, 0, 
    13, 13, 16, 0, 71, 0, 1, 0, 12, 0, 46, 0, 110, 0, 23, 
    22, 16, 6, 19, 62, 0, 0, 10, 0, 50, 0, 0, 73, 2, 14, 
    39, 0, 21, 35, 0, 0, 23, 64, 0, 54, 0, 0, 61, 18, 90, 
    41, 0, 80, 22, 0, 4, 89, 0, 0, 0, 9, 0, 37, 19, 143, 
    76, 0, 20, 81, 0, 10, 47, 0, 29, 22, 41, 0, 57, 16, 149, 
    56, 0, 0, 40, 53, 22, 32, 11, 26, 20, 25, 7, 55, 0, 125, 
    41, 0, 0, 18, 35, 43, 0, 18, 44, 17, 16, 10, 69, 15, 125, 
    0, 0, 31, 20, 0, 71, 4, 38, 25, 25, 43, 24, 65, 55, 77, 
    8, 46, 40, 0, 25, 0, 35, 21, 33, 52, 36, 45, 83, 7, 0, 
    89, 0, 45, 0, 0, 32, 0, 47, 54, 53, 39, 43, 53, 13, 0, 
    0, 0, 68, 0, 49, 0, 0, 36, 46, 67, 16, 42, 58, 3, 23, 
    3, 0, 63, 47, 38, 0, 19, 75, 3, 45, 34, 66, 59, 0, 11, 
    48, 0, 0, 27, 58, 22, 3, 37, 0, 23, 36, 66, 113, 0, 0, 
    67, 8, 0, 0, 37, 45, 31, 12, 33, 13, 41, 53, 33, 0, 0, 
    
    -- channel=76
    51, 48, 4, 30, 95, 0, 43, 8, 43, 46, 102, 0, 187, 0, 36, 
    59, 55, 56, 37, 98, 0, 35, 0, 72, 27, 101, 0, 195, 0, 75, 
    74, 62, 51, 50, 83, 0, 15, 51, 29, 86, 30, 0, 168, 62, 90, 
    85, 0, 73, 74, 17, 0, 86, 89, 0, 99, 0, 12, 151, 88, 160, 
    79, 0, 159, 62, 0, 67, 138, 0, 53, 36, 80, 42, 116, 92, 204, 
    105, 0, 99, 145, 5, 70, 90, 35, 87, 82, 102, 0, 134, 86, 212, 
    102, 0, 42, 123, 112, 79, 89, 70, 90, 77, 79, 68, 122, 60, 187, 
    93, 20, 54, 104, 121, 78, 62, 91, 105, 84, 77, 76, 145, 77, 169, 
    54, 46, 81, 84, 51, 153, 58, 104, 97, 106, 119, 82, 134, 89, 133, 
    69, 95, 94, 43, 91, 40, 103, 98, 110, 126, 107, 116, 143, 62, 12, 
    143, 30, 97, 26, 38, 96, 22, 125, 135, 127, 106, 116, 113, 54, 64, 
    69, 71, 146, 31, 116, 33, 74, 122, 116, 140, 90, 114, 118, 50, 95, 
    64, 70, 171, 130, 112, 53, 90, 135, 58, 121, 104, 131, 126, 20, 85, 
    110, 0, 32, 134, 147, 98, 90, 114, 7, 95, 113, 130, 150, 0, 57, 
    121, 50, 0, 31, 146, 141, 126, 95, 104, 78, 95, 115, 94, 36, 0, 
    
    -- channel=77
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 
    
    -- channel=78
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 4, 0, 0, 5, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 11, 0, 0, 11, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 29, 
    0, 0, 0, 0, 8, 0, 0, 1, 0, 11, 2, 5, 39, 26, 0, 
    0, 1, 0, 0, 0, 17, 0, 0, 0, 3, 3, 8, 12, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 24, 18, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 9, 5, 0, 14, 20, 0, 0, 
    28, 2, 0, 0, 0, 0, 0, 73, 38, 0, 7, 16, 19, 0, 0, 
    0, 55, 0, 0, 0, 0, 0, 0, 0, 13, 2, 31, 64, 0, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 3, 31, 59, 15, 0, 0, 0, 
    
    -- channel=79
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 5, 16, 0, 
    0, 0, 0, 1, 0, 12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 20, 0, 0, 0, 0, 14, 35, 26, 0, 0, 0, 0, 0, 0, 
    0, 21, 20, 0, 0, 0, 0, 0, 0, 1, 0, 0, 3, 10, 0, 
    0, 0, 3, 22, 0, 0, 0, 0, 0, 29, 47, 0, 0, 0, 0, 
    
    -- channel=80
    0, 41, 0, 8, 0, 0, 0, 0, 0, 0, 2, 0, 13, 22, 0, 
    0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 20, 0, 12, 0, 0, 
    0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 1, 
    0, 19, 0, 0, 0, 0, 0, 23, 0, 16, 0, 0, 14, 0, 0, 
    90, 0, 40, 0, 0, 50, 0, 0, 0, 25, 0, 0, 19, 0, 11, 
    114, 21, 0, 0, 10, 7, 0, 0, 69, 25, 0, 0, 13, 16, 0, 
    0, 95, 0, 0, 38, 0, 0, 17, 0, 0, 0, 0, 8, 53, 0, 
    0, 74, 0, 0, 49, 0, 0, 0, 0, 0, 0, 0, 58, 73, 0, 
    0, 85, 0, 0, 59, 0, 0, 75, 0, 0, 0, 4, 40, 109, 0, 
    0, 31, 0, 0, 44, 0, 0, 25, 0, 0, 0, 5, 27, 85, 0, 
    0, 20, 0, 0, 0, 24, 22, 0, 0, 0, 0, 12, 39, 5, 7, 
    3, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 33, 35, 0, 48, 
    0, 14, 0, 0, 0, 26, 28, 0, 2, 0, 4, 39, 5, 24, 0, 
    4, 32, 0, 8, 0, 5, 0, 0, 0, 0, 12, 10, 0, 0, 16, 
    
    -- channel=81
    157, 172, 160, 163, 160, 142, 116, 119, 80, 50, 70, 62, 67, 97, 64, 
    220, 211, 169, 188, 187, 174, 141, 138, 91, 19, 65, 75, 109, 97, 79, 
    208, 222, 198, 204, 211, 199, 171, 154, 159, 106, 121, 82, 92, 95, 102, 
    197, 230, 208, 219, 220, 205, 185, 156, 172, 183, 154, 90, 74, 88, 108, 
    181, 220, 223, 221, 226, 210, 201, 210, 147, 169, 176, 100, 81, 94, 108, 
    149, 229, 251, 240, 213, 279, 256, 197, 152, 175, 149, 48, 67, 71, 100, 
    149, 251, 285, 251, 241, 295, 242, 209, 235, 237, 136, 31, 47, 73, 81, 
    112, 238, 270, 247, 320, 314, 259, 311, 311, 302, 168, 34, 60, 151, 65, 
    135, 252, 288, 188, 300, 281, 223, 208, 214, 174, 65, 0, 54, 210, 73, 
    143, 248, 315, 109, 192, 256, 171, 232, 127, 27, 15, 11, 58, 260, 144, 
    166, 216, 269, 73, 29, 52, 62, 133, 43, 0, 0, 28, 56, 232, 206, 
    159, 187, 225, 175, 92, 74, 94, 53, 0, 0, 0, 0, 46, 101, 209, 
    162, 195, 181, 230, 149, 131, 141, 90, 33, 6, 0, 0, 33, 33, 122, 
    151, 175, 168, 145, 134, 140, 177, 135, 112, 94, 82, 108, 91, 94, 102, 
    159, 185, 164, 169, 166, 182, 153, 141, 130, 111, 136, 163, 149, 123, 113, 
    
    -- channel=82
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 19, 3, 11, 10, 3, 0, 3, 0, 0, 0, 0, 1, 0, 0, 
    0, 21, 12, 18, 17, 10, 10, 0, 16, 5, 0, 0, 0, 0, 0, 
    15, 21, 13, 12, 16, 10, 7, 0, 0, 32, 12, 0, 0, 0, 0, 
    53, 3, 25, 17, 11, 29, 4, 53, 0, 19, 5, 0, 0, 0, 2, 
    42, 56, 34, 17, 13, 49, 23, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 73, 31, 35, 49, 27, 12, 55, 47, 31, 0, 0, 0, 0, 0, 
    0, 53, 35, 6, 74, 63, 26, 62, 60, 57, 0, 0, 0, 39, 0, 
    0, 72, 52, 0, 107, 56, 2, 20, 0, 0, 0, 0, 0, 63, 0, 
    8, 60, 52, 0, 0, 38, 21, 72, 0, 0, 0, 0, 0, 88, 0, 
    18, 28, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 35, 35, 
    15, 28, 17, 56, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 36, 
    17, 50, 13, 11, 0, 0, 34, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 21, 9, 12, 0, 16, 17, 20, 3, 1, 4, 11, 0, 0, 0, 
    
    -- channel=83
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 15, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 20, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 1, 7, 0, 1, 4, 6, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 13, 18, 14, 7, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 14, 14, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=84
    86, 104, 119, 118, 119, 120, 109, 104, 74, 70, 72, 62, 66, 81, 61, 
    102, 109, 116, 123, 126, 128, 128, 122, 93, 63, 74, 83, 89, 80, 77, 
    92, 106, 118, 126, 127, 131, 124, 137, 123, 72, 96, 89, 96, 90, 83, 
    85, 115, 118, 127, 130, 137, 134, 123, 126, 124, 112, 85, 82, 88, 88, 
    86, 104, 119, 125, 132, 132, 104, 100, 101, 126, 113, 73, 83, 88, 86, 
    88, 101, 114, 120, 120, 107, 73, 99, 81, 102, 89, 55, 76, 79, 87, 
    106, 109, 109, 98, 98, 104, 85, 56, 77, 84, 61, 40, 57, 76, 83, 
    85, 117, 97, 105, 100, 99, 110, 106, 90, 81, 53, 44, 60, 79, 67, 
    102, 116, 95, 85, 93, 98, 94, 114, 98, 92, 52, 36, 64, 96, 33, 
    97, 117, 84, 37, 115, 104, 80, 108, 91, 51, 43, 52, 74, 109, 25, 
    104, 115, 84, 35, 48, 62, 67, 119, 68, 48, 48, 59, 72, 115, 43, 
    109, 106, 86, 66, 85, 71, 93, 71, 26, 26, 25, 42, 67, 92, 81, 
    111, 114, 93, 106, 88, 99, 98, 77, 50, 36, 25, 32, 62, 57, 92, 
    102, 113, 101, 91, 68, 92, 116, 93, 83, 73, 73, 82, 74, 85, 79, 
    102, 111, 103, 110, 95, 114, 117, 110, 103, 99, 108, 112, 102, 92, 90, 
    
    -- channel=85
    0, 31, 4, 3, 2, 9, 0, 10, 0, 13, 9, 7, 14, 18, 0, 
    6, 7, 1, 9, 3, 3, 0, 0, 0, 10, 24, 9, 5, 0, 3, 
    2, 23, 9, 6, 3, 3, 0, 11, 0, 0, 15, 0, 9, 0, 0, 
    0, 28, 7, 7, 9, 0, 0, 0, 6, 0, 0, 0, 1, 12, 5, 
    4, 17, 10, 9, 9, 0, 0, 0, 3, 10, 0, 0, 19, 7, 5, 
    41, 3, 21, 6, 8, 3, 0, 19, 0, 10, 0, 0, 30, 12, 14, 
    80, 10, 6, 0, 4, 25, 0, 0, 18, 18, 0, 0, 28, 21, 14, 
    2, 41, 0, 5, 15, 0, 0, 3, 5, 0, 0, 0, 25, 13, 0, 
    0, 23, 0, 0, 37, 8, 0, 22, 11, 14, 0, 7, 47, 32, 0, 
    0, 31, 0, 0, 60, 19, 0, 0, 0, 0, 4, 12, 36, 36, 0, 
    0, 14, 7, 0, 47, 44, 7, 42, 0, 6, 29, 14, 26, 45, 0, 
    0, 0, 0, 0, 0, 0, 8, 0, 10, 26, 24, 50, 35, 38, 0, 
    0, 0, 10, 8, 0, 0, 0, 0, 0, 7, 19, 31, 43, 9, 53, 
    0, 1, 0, 4, 0, 7, 8, 0, 0, 0, 0, 8, 0, 16, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=86
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 16, 24, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 4, 0, 0, 28, 6, 0, 8, 13, 0, 0, 0, 0, 0, 
    0, 8, 3, 0, 18, 7, 0, 20, 37, 28, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 51, 18, 0, 13, 17, 20, 1, 0, 0, 14, 0, 
    0, 6, 34, 0, 44, 16, 0, 0, 0, 0, 0, 0, 0, 21, 5, 
    0, 0, 36, 0, 2, 27, 0, 7, 0, 0, 0, 0, 0, 26, 21, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 13, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=87
    100, 83, 91, 82, 93, 93, 97, 88, 77, 57, 53, 57, 59, 53, 58, 
    83, 87, 98, 92, 95, 98, 102, 97, 97, 66, 48, 58, 57, 60, 62, 
    79, 77, 93, 96, 94, 105, 103, 99, 103, 92, 72, 72, 57, 62, 61, 
    84, 75, 92, 94, 99, 105, 100, 96, 87, 96, 94, 83, 62, 60, 60, 
    71, 77, 88, 97, 99, 91, 72, 68, 78, 77, 83, 73, 56, 58, 58, 
    55, 83, 80, 88, 91, 79, 55, 50, 62, 56, 62, 65, 43, 58, 57, 
    35, 70, 74, 74, 81, 65, 85, 69, 46, 52, 62, 54, 41, 57, 53, 
    67, 48, 71, 74, 63, 76, 86, 65, 58, 59, 60, 49, 43, 52, 59, 
    74, 49, 64, 72, 42, 76, 71, 65, 62, 55, 57, 49, 41, 47, 57, 
    72, 55, 50, 62, 29, 49, 77, 57, 74, 58, 47, 43, 43, 45, 51, 
    71, 60, 52, 75, 38, 40, 47, 44, 61, 46, 34, 41, 47, 42, 54, 
    78, 61, 60, 77, 83, 71, 65, 54, 46, 37, 28, 22, 43, 49, 55, 
    73, 73, 66, 66, 75, 62, 62, 73, 63, 49, 47, 43, 36, 54, 38, 
    60, 62, 71, 68, 67, 65, 63, 75, 69, 66, 70, 66, 70, 64, 59, 
    74, 64, 74, 71, 72, 71, 72, 70, 71, 72, 68, 72, 75, 71, 69, 
    
    -- channel=88
    0, 3, 0, 1, 0, 0, 0, 10, 0, 8, 9, 0, 4, 26, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 13, 17, 0, 0, 
    0, 17, 0, 3, 0, 0, 0, 6, 0, 0, 6, 0, 8, 8, 2, 
    0, 14, 0, 12, 0, 0, 0, 0, 17, 0, 0, 0, 0, 19, 9, 
    18, 17, 0, 3, 0, 0, 0, 0, 0, 40, 6, 0, 27, 9, 12, 
    155, 0, 10, 0, 0, 34, 0, 3, 0, 33, 0, 0, 37, 10, 23, 
    122, 70, 0, 0, 14, 13, 0, 0, 0, 0, 0, 0, 24, 13, 11, 
    0, 126, 0, 6, 41, 0, 0, 12, 0, 0, 0, 0, 44, 22, 0, 
    0, 91, 0, 0, 55, 51, 0, 30, 32, 15, 0, 0, 84, 71, 0, 
    0, 104, 0, 0, 150, 49, 0, 35, 0, 0, 0, 0, 71, 109, 0, 
    0, 74, 0, 0, 45, 60, 36, 75, 0, 0, 18, 23, 34, 144, 0, 
    0, 14, 20, 0, 0, 0, 0, 0, 0, 6, 0, 43, 72, 73, 23, 
    11, 0, 2, 45, 0, 0, 12, 0, 0, 0, 0, 5, 42, 21, 53, 
    0, 58, 0, 29, 0, 7, 35, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 16, 0, 1, 0, 0, 0, 0, 0, 0, 10, 9, 0, 0, 12, 
    
    -- channel=89
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 16, 4, 1, 8, 9, 0, 
    49, 0, 0, 0, 9, 0, 0, 51, 30, 0, 5, 33, 12, 6, 1, 
    0, 34, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 8, 0, 13, 0, 0, 0, 0, 0, 0, 0, 5, 10, 0, 0, 
    0, 0, 0, 11, 25, 36, 0, 77, 67, 100, 112, 36, 3, 0, 0, 
    0, 1, 0, 0, 117, 30, 24, 0, 0, 37, 0, 0, 1, 0, 0, 
    0, 21, 23, 11, 0, 105, 78, 75, 87, 33, 46, 22, 0, 42, 0, 
    12, 0, 14, 0, 0, 0, 0, 0, 21, 21, 16, 36, 32, 47, 32, 
    0, 0, 0, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 23, 
    0, 25, 0, 7, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=90
    113, 169, 140, 148, 141, 140, 120, 119, 70, 65, 72, 69, 72, 95, 59, 
    152, 147, 147, 153, 158, 160, 150, 142, 96, 55, 72, 78, 98, 87, 77, 
    129, 148, 162, 162, 165, 167, 154, 159, 146, 101, 128, 99, 97, 87, 96, 
    112, 156, 154, 169, 167, 172, 156, 147, 152, 146, 134, 92, 75, 95, 95, 
    113, 151, 164, 165, 175, 165, 139, 151, 129, 144, 141, 75, 86, 88, 91, 
    112, 144, 172, 169, 156, 169, 138, 108, 90, 130, 108, 31, 77, 79, 92, 
    157, 149, 160, 145, 157, 168, 111, 103, 153, 147, 78, 31, 61, 84, 81, 
    93, 165, 144, 140, 177, 164, 175, 156, 145, 136, 90, 36, 62, 115, 74, 
    115, 168, 151, 122, 139, 136, 132, 111, 101, 80, 0, 2, 76, 134, 42, 
    104, 164, 140, 52, 98, 149, 81, 158, 108, 28, 42, 52, 80, 158, 48, 
    121, 144, 112, 7, 61, 28, 38, 98, 20, 24, 19, 37, 84, 148, 56, 
    108, 137, 109, 120, 94, 96, 120, 59, 4, 3, 0, 23, 57, 99, 82, 
    137, 125, 126, 123, 129, 107, 113, 91, 56, 40, 22, 33, 71, 50, 99, 
    113, 127, 110, 115, 73, 114, 136, 104, 97, 93, 91, 114, 100, 113, 69, 
    109, 150, 119, 138, 126, 139, 128, 109, 109, 100, 126, 132, 123, 106, 111, 
    
    -- channel=91
    79, 0, 32, 16, 33, 24, 39, 15, 58, 10, 8, 15, 0, 0, 45, 
    32, 49, 29, 25, 25, 25, 39, 25, 61, 19, 0, 11, 10, 31, 16, 
    65, 5, 23, 25, 24, 36, 41, 10, 40, 62, 0, 36, 11, 19, 17, 
    63, 15, 30, 18, 35, 39, 44, 37, 16, 37, 36, 54, 20, 0, 11, 
    39, 8, 27, 25, 25, 34, 29, 11, 41, 0, 26, 93, 0, 16, 14, 
    0, 41, 0, 29, 40, 0, 68, 38, 69, 0, 39, 75, 0, 10, 0, 
    0, 0, 48, 48, 7, 20, 79, 62, 0, 2, 82, 53, 0, 0, 6, 
    40, 0, 59, 35, 0, 60, 48, 25, 49, 55, 96, 59, 0, 0, 48, 
    42, 0, 40, 67, 1, 17, 84, 39, 45, 62, 119, 33, 0, 0, 112, 
    57, 0, 41, 156, 0, 14, 113, 0, 83, 44, 8, 13, 0, 0, 145, 
    57, 0, 52, 163, 0, 0, 21, 0, 89, 28, 1, 0, 0, 0, 135, 
    59, 13, 29, 52, 63, 16, 4, 55, 18, 0, 0, 0, 0, 0, 33, 
    22, 35, 23, 19, 64, 51, 6, 58, 41, 13, 8, 0, 0, 1, 0, 
    36, 0, 69, 19, 68, 3, 0, 66, 24, 36, 27, 2, 24, 0, 45, 
    27, 5, 48, 20, 38, 27, 30, 41, 37, 29, 12, 15, 36, 44, 3, 
    
    -- channel=92
    129, 39, 81, 72, 87, 72, 82, 47, 90, 31, 39, 46, 31, 21, 73, 
    98, 118, 82, 82, 84, 85, 88, 72, 100, 37, 18, 40, 42, 64, 46, 
    129, 83, 84, 89, 89, 99, 102, 61, 89, 96, 27, 60, 42, 52, 51, 
    119, 78, 95, 83, 99, 101, 102, 87, 70, 92, 78, 97, 54, 28, 48, 
    87, 79, 95, 87, 101, 95, 98, 85, 96, 56, 77, 138, 30, 48, 51, 
    0, 102, 80, 101, 105, 57, 135, 89, 122, 44, 90, 106, 14, 42, 36, 
    0, 62, 121, 121, 75, 90, 143, 123, 48, 63, 128, 77, 13, 32, 39, 
    70, 0, 132, 94, 74, 143, 111, 90, 117, 125, 158, 79, 5, 34, 75, 
    85, 3, 119, 114, 89, 88, 159, 89, 102, 107, 153, 50, 0, 13, 157, 
    101, 0, 119, 211, 0, 69, 172, 52, 114, 61, 34, 31, 0, 0, 208, 
    106, 25, 117, 209, 0, 23, 67, 18, 129, 41, 21, 27, 0, 0, 207, 
    99, 59, 84, 122, 78, 37, 22, 71, 34, 6, 8, 0, 0, 2, 94, 
    69, 83, 70, 77, 116, 83, 55, 89, 56, 24, 16, 0, 0, 25, 0, 
    86, 42, 117, 51, 120, 53, 42, 112, 58, 62, 52, 29, 51, 25, 71, 
    78, 54, 98, 63, 81, 77, 74, 85, 74, 68, 56, 60, 78, 86, 38, 
    
    -- channel=93
    27, 5, 27, 36, 34, 33, 30, 15, 3, 5, 8, 4, 4, 0, 3, 
    30, 34, 37, 32, 35, 40, 39, 36, 16, 1, 8, 8, 6, 7, 7, 
    18, 32, 37, 41, 39, 43, 43, 48, 32, 0, 0, 4, 12, 16, 8, 
    28, 22, 35, 39, 37, 48, 44, 41, 42, 35, 30, 17, 15, 14, 12, 
    23, 26, 36, 36, 46, 34, 38, 27, 29, 42, 35, 15, 14, 11, 12, 
    45, 21, 34, 32, 47, 13, 0, 6, 31, 19, 19, 14, 10, 12, 11, 
    0, 34, 16, 22, 27, 0, 19, 0, 0, 0, 3, 0, 4, 8, 8, 
    0, 14, 15, 17, 8, 16, 18, 0, 0, 0, 0, 0, 6, 0, 0, 
    12, 4, 11, 13, 4, 28, 22, 20, 15, 15, 17, 4, 4, 0, 0, 
    19, 4, 0, 0, 13, 13, 28, 5, 0, 7, 4, 0, 2, 0, 0, 
    15, 10, 0, 7, 0, 14, 35, 22, 37, 4, 0, 8, 0, 0, 0, 
    26, 8, 7, 12, 0, 0, 0, 0, 3, 0, 0, 0, 13, 9, 6, 
    28, 15, 7, 23, 24, 13, 22, 2, 0, 0, 0, 0, 0, 15, 0, 
    15, 29, 17, 15, 18, 13, 11, 19, 6, 0, 0, 0, 0, 0, 0, 
    18, 7, 24, 13, 12, 12, 19, 28, 16, 22, 20, 19, 16, 17, 10, 
    
    -- channel=94
    10, 0, 46, 42, 44, 52, 50, 41, 44, 41, 35, 31, 22, 29, 37, 
    29, 39, 38, 39, 40, 38, 51, 49, 41, 40, 38, 46, 37, 45, 35, 
    41, 20, 36, 43, 40, 46, 47, 56, 33, 0, 0, 38, 56, 51, 35, 
    35, 31, 41, 37, 48, 58, 63, 58, 56, 47, 45, 47, 50, 38, 44, 
    46, 23, 35, 42, 38, 46, 35, 10, 53, 61, 49, 57, 37, 49, 44, 
    19, 30, 12, 33, 56, 0, 7, 65, 58, 28, 54, 63, 35, 43, 43, 
    13, 33, 31, 30, 0, 21, 40, 0, 0, 0, 40, 38, 25, 28, 48, 
    46, 16, 34, 33, 0, 5, 22, 6, 12, 4, 19, 42, 23, 0, 41, 
    42, 11, 13, 52, 34, 39, 65, 92, 78, 107, 116, 52, 15, 2, 40, 
    62, 13, 11, 74, 49, 47, 72, 0, 59, 59, 13, 18, 26, 0, 15, 
    57, 46, 47, 62, 32, 93, 88, 100, 101, 57, 57, 35, 25, 24, 23, 
    68, 45, 30, 0, 23, 0, 12, 60, 45, 29, 27, 42, 32, 72, 29, 
    52, 51, 49, 44, 27, 57, 33, 24, 6, 0, 0, 0, 22, 40, 51, 
    67, 59, 64, 59, 55, 27, 45, 57, 23, 18, 7, 0, 1, 14, 40, 
    40, 36, 51, 34, 26, 42, 65, 67, 61, 56, 44, 40, 42, 45, 24, 
    
    -- channel=95
    0, 0, 0, 3, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 2, 0, 
    0, 0, 0, 0, 0, 0, 1, 2, 10, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 3, 3, 0, 0, 14, 8, 8, 11, 7, 0, 
    9, 0, 0, 0, 0, 0, 0, 37, 28, 5, 6, 0, 10, 4, 0, 
    3, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 
    0, 0, 0, 11, 17, 0, 17, 31, 29, 47, 29, 0, 0, 0, 0, 
    0, 0, 0, 6, 44, 39, 7, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 3, 4, 0, 0, 11, 27, 27, 38, 17, 17, 7, 0, 10, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 13, 5, 24, 0, 
    6, 0, 0, 9, 25, 21, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    6, 15, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 13, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=96
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 47, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 34, 0, 0, 40, 0, 
    0, 0, 0, 0, 4, 2, 16, 15, 10, 6, 0, 11, 11, 0, 0, 
    4, 0, 0, 0, 6, 17, 9, 11, 56, 44, 0, 3, 0, 0, 0, 
    1, 0, 0, 0, 14, 72, 82, 0, 0, 0, 75, 0, 9, 0, 0, 
    0, 0, 0, 8, 52, 0, 0, 0, 0, 115, 119, 0, 0, 2, 0, 
    0, 0, 26, 13, 0, 17, 0, 99, 181, 171, 0, 0, 0, 2, 121, 
    0, 17, 0, 0, 0, 0, 63, 153, 0, 0, 0, 0, 72, 117, 43, 
    11, 203, 0, 14, 0, 29, 114, 34, 0, 0, 0, 0, 39, 0, 0, 
    72, 0, 0, 0, 0, 92, 152, 6, 0, 0, 1, 94, 0, 0, 0, 
    20, 0, 45, 0, 37, 91, 130, 0, 0, 21, 0, 59, 26, 0, 0, 
    15, 16, 49, 0, 124, 83, 104, 0, 0, 53, 0, 0, 66, 0, 12, 
    16, 12, 0, 0, 0, 0, 0, 0, 0, 64, 0, 0, 0, 0, 9, 
    9, 0, 15, 20, 11, 19, 10, 3, 0, 37, 0, 0, 4, 7, 21, 
    
    -- channel=97
    100, 83, 94, 78, 65, 46, 53, 27, 26, 45, 12, 15, 0, 0, 0, 
    78, 69, 47, 21, 16, 8, 15, 4, 2, 0, 36, 0, 0, 7, 0, 
    37, 18, 2, 0, 0, 1, 4, 7, 10, 22, 84, 36, 10, 41, 6, 
    0, 0, 0, 0, 4, 14, 35, 48, 50, 55, 9, 1, 27, 14, 0, 
    0, 0, 0, 0, 17, 48, 88, 109, 172, 164, 64, 40, 34, 0, 0, 
    0, 0, 0, 0, 35, 147, 250, 260, 275, 277, 370, 47, 29, 43, 0, 
    2, 2, 0, 19, 87, 134, 135, 26, 22, 173, 495, 215, 0, 30, 0, 
    5, 6, 58, 92, 93, 88, 102, 164, 286, 431, 504, 261, 16, 1, 143, 
    1, 47, 54, 101, 59, 44, 160, 484, 506, 517, 450, 91, 120, 184, 331, 
    36, 284, 107, 64, 0, 0, 218, 462, 451, 358, 392, 343, 338, 340, 261, 
    72, 254, 150, 31, 0, 56, 265, 435, 317, 61, 70, 324, 346, 254, 53, 
    24, 61, 197, 8, 0, 147, 349, 447, 190, 36, 6, 113, 284, 99, 0, 
    0, 85, 210, 50, 170, 284, 403, 426, 157, 108, 73, 0, 183, 0, 0, 
    0, 53, 106, 23, 91, 137, 154, 153, 44, 99, 75, 0, 0, 0, 0, 
    24, 25, 41, 13, 0, 1, 0, 0, 0, 25, 17, 0, 0, 0, 0, 
    
    -- channel=98
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 26, 41, 91, 86, 10, 0, 9, 0, 0, 
    0, 0, 0, 0, 18, 49, 49, 15, 6, 53, 149, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 114, 30, 0, 0, 0, 
    0, 0, 0, 26, 0, 0, 36, 122, 130, 136, 87, 0, 0, 0, 55, 
    0, 45, 0, 1, 0, 0, 78, 133, 114, 126, 152, 0, 32, 59, 59, 
    48, 130, 0, 0, 0, 0, 76, 106, 77, 0, 52, 193, 81, 68, 0, 
    13, 0, 22, 0, 0, 30, 109, 98, 0, 0, 0, 72, 79, 0, 0, 
    0, 0, 38, 0, 0, 0, 97, 98, 0, 0, 0, 0, 94, 0, 0, 
    0, 7, 41, 4, 77, 121, 130, 129, 9, 25, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 
    
    -- channel=99
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 32, 19, 22, 0, 0, 
    0, 0, 0, 0, 0, 3, 16, 34, 22, 53, 12, 51, 22, 14, 5, 
    0, 0, 0, 0, 13, 18, 21, 46, 34, 4, 35, 26, 44, 29, 23, 
    0, 0, 0, 36, 20, 25, 56, 2, 20, 39, 20, 63, 30, 34, 17, 
    0, 0, 32, 34, 36, 25, 43, 25, 46, 19, 47, 54, 27, 32, 18, 
    0, 3, 51, 26, 38, 37, 38, 36, 10, 64, 16, 40, 41, 31, 34, 
    0, 40, 26, 35, 34, 20, 46, 38, 34, 30, 32, 24, 43, 31, 36, 
    7, 30, 28, 55, 42, 43, 22, 45, 46, 36, 34, 25, 12, 50, 16, 
    8, 17, 17, 40, 20, 27, 29, 33, 51, 23, 38, 30, 12, 37, 20, 
    9, 21, 41, 31, 34, 33, 30, 29, 26, 18, 25, 35, 21, 20, 20, 
    
    -- channel=100
    250, 249, 257, 253, 240, 222, 218, 200, 184, 164, 143, 130, 66, 63, 110, 
    237, 219, 219, 212, 199, 183, 181, 169, 160, 146, 135, 85, 33, 80, 125, 
    179, 171, 171, 169, 164, 156, 159, 155, 153, 151, 103, 35, 58, 115, 130, 
    142, 150, 153, 152, 157, 161, 158, 156, 152, 140, 43, 32, 102, 135, 133, 
    146, 155, 156, 155, 160, 158, 145, 140, 117, 75, 7, 50, 109, 126, 130, 
    155, 156, 155, 153, 147, 120, 98, 92, 94, 58, 11, 0, 61, 85, 116, 
    157, 156, 151, 142, 117, 75, 21, 2, 15, 32, 56, 0, 7, 52, 83, 
    155, 153, 134, 96, 51, 45, 19, 0, 22, 37, 27, 1, 0, 26, 35, 
    153, 136, 60, 28, 10, 17, 36, 62, 41, 26, 1, 0, 50, 27, 55, 
    148, 101, 0, 13, 0, 28, 36, 33, 12, 30, 51, 0, 29, 20, 22, 
    144, 80, 0, 0, 0, 8, 33, 16, 0, 0, 16, 49, 0, 8, 1, 
    108, 2, 6, 0, 8, 23, 29, 15, 0, 1, 4, 53, 7, 0, 10, 
    82, 22, 13, 0, 6, 0, 27, 2, 0, 21, 0, 11, 41, 0, 35, 
    72, 40, 26, 0, 28, 27, 23, 20, 0, 22, 0, 0, 29, 0, 25, 
    70, 24, 0, 0, 0, 0, 0, 2, 6, 44, 7, 0, 14, 15, 19, 
    
    -- channel=101
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 25, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 21, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 33, 3, 0, 
    0, 0, 0, 0, 0, 6, 13, 24, 26, 37, 51, 0, 24, 30, 8, 
    0, 0, 0, 0, 7, 15, 0, 0, 20, 35, 2, 0, 0, 13, 25, 
    0, 0, 0, 11, 13, 36, 32, 42, 2, 0, 0, 0, 1, 7, 22, 
    0, 0, 0, 32, 4, 42, 41, 26, 0, 13, 0, 0, 0, 5, 14, 
    0, 21, 0, 26, 10, 29, 66, 10, 12, 0, 68, 50, 0, 17, 0, 
    0, 1, 26, 6, 23, 55, 44, 0, 0, 21, 20, 75, 8, 0, 14, 
    0, 12, 35, 0, 32, 15, 47, 0, 0, 28, 5, 33, 62, 0, 39, 
    1, 12, 41, 14, 60, 51, 43, 37, 0, 43, 2, 12, 61, 16, 34, 
    0, 0, 20, 22, 27, 28, 31, 28, 31, 64, 13, 9, 34, 35, 37, 
    
    -- channel=102
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 61, 79, 84, 11, 3, 0, 0, 
    0, 0, 0, 0, 0, 25, 79, 64, 43, 58, 174, 38, 2, 16, 0, 
    0, 0, 0, 0, 14, 11, 25, 23, 37, 102, 166, 110, 3, 0, 13, 
    0, 0, 0, 45, 47, 41, 51, 141, 160, 167, 155, 24, 1, 18, 89, 
    0, 0, 24, 52, 15, 27, 77, 174, 161, 158, 138, 55, 84, 117, 108, 
    0, 107, 77, 46, 0, 26, 104, 161, 160, 68, 93, 157, 141, 129, 58, 
    0, 30, 101, 29, 11, 84, 132, 155, 93, 32, 24, 80, 123, 73, 0, 
    0, 41, 107, 27, 59, 94, 149, 157, 71, 48, 35, 26, 116, 28, 0, 
    0, 21, 90, 58, 109, 137, 141, 141, 67, 66, 54, 12, 51, 4, 0, 
    0, 0, 34, 24, 21, 24, 24, 18, 9, 49, 35, 0, 0, 0, 3, 
    
    -- channel=103
    179, 178, 174, 180, 172, 156, 147, 145, 123, 106, 113, 86, 30, 45, 85, 
    158, 151, 143, 137, 124, 116, 114, 113, 104, 106, 87, 66, 58, 50, 85, 
    108, 108, 105, 105, 105, 103, 103, 107, 106, 104, 37, 30, 58, 75, 88, 
    95, 98, 98, 99, 103, 103, 98, 102, 106, 92, 41, 42, 87, 92, 97, 
    92, 98, 98, 98, 98, 89, 77, 82, 74, 51, 33, 25, 52, 85, 87, 
    98, 97, 96, 96, 87, 59, 18, 6, 0, 4, 0, 44, 24, 46, 76, 
    98, 97, 95, 86, 44, 24, 16, 24, 22, 17, 0, 22, 29, 8, 42, 
    97, 95, 68, 38, 19, 26, 22, 22, 22, 0, 0, 9, 33, 30, 9, 
    94, 80, 31, 12, 13, 16, 25, 0, 0, 0, 0, 60, 24, 8, 0, 
    92, 13, 19, 4, 28, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    64, 0, 1, 5, 30, 8, 0, 0, 0, 29, 4, 0, 0, 0, 27, 
    59, 20, 0, 19, 17, 0, 0, 0, 12, 12, 19, 3, 0, 11, 36, 
    49, 9, 0, 19, 0, 0, 0, 0, 18, 4, 11, 15, 0, 30, 25, 
    49, 18, 0, 11, 0, 0, 0, 0, 17, 0, 14, 24, 13, 30, 21, 
    40, 22, 10, 8, 7, 6, 13, 16, 20, 9, 6, 28, 25, 24, 24, 
    
    -- channel=104
    0, 0, 12, 5, 0, 0, 10, 0, 14, 0, 0, 0, 0, 45, 0, 
    3, 0, 0, 0, 0, 0, 8, 0, 0, 0, 11, 0, 0, 54, 0, 
    13, 3, 6, 0, 5, 1, 1, 0, 0, 8, 1, 0, 0, 25, 0, 
    10, 7, 4, 0, 6, 2, 0, 0, 0, 0, 0, 63, 24, 0, 0, 
    9, 5, 4, 0, 13, 1, 13, 7, 1, 0, 0, 15, 0, 0, 0, 
    6, 1, 0, 0, 24, 23, 1, 0, 38, 11, 0, 0, 69, 0, 0, 
    3, 0, 0, 18, 21, 47, 6, 0, 26, 167, 93, 0, 0, 38, 8, 
    6, 0, 13, 0, 0, 27, 0, 0, 0, 57, 2, 0, 0, 27, 29, 
    1, 20, 0, 34, 0, 54, 120, 102, 22, 14, 0, 0, 16, 20, 23, 
    31, 63, 0, 38, 0, 62, 200, 49, 15, 0, 79, 0, 0, 0, 0, 
    96, 71, 0, 0, 0, 59, 169, 23, 0, 0, 89, 221, 0, 0, 0, 
    42, 14, 0, 0, 25, 84, 159, 0, 0, 18, 0, 164, 44, 0, 0, 
    30, 27, 34, 0, 66, 0, 84, 5, 0, 58, 0, 17, 116, 0, 34, 
    15, 31, 31, 12, 104, 100, 100, 87, 0, 92, 0, 0, 49, 0, 19, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 73, 0, 0, 1, 5, 19, 
    
    -- channel=105
    0, 0, 1, 18, 23, 23, 22, 19, 26, 49, 14, 4, 42, 37, 0, 
    17, 0, 14, 24, 25, 20, 14, 12, 6, 0, 0, 3, 4, 0, 0, 
    49, 50, 26, 16, 9, 0, 0, 0, 0, 0, 11, 21, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 20, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 89, 127, 0, 0, 67, 0, 0, 
    0, 0, 0, 0, 0, 93, 102, 112, 75, 18, 0, 0, 0, 56, 15, 
    0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 
    0, 0, 19, 60, 36, 55, 20, 0, 8, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 19, 35, 31, 4, 0, 85, 138, 0, 0, 0, 18, 
    31, 162, 14, 0, 20, 0, 0, 0, 28, 116, 97, 162, 34, 52, 113, 
    41, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 78, 31, 18, 3, 
    32, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 89, 47, 18, 
    0, 25, 71, 90, 144, 212, 232, 236, 140, 28, 29, 5, 71, 35, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 47, 24, 0, 0, 0, 
    
    -- channel=106
    249, 234, 248, 240, 221, 199, 199, 172, 159, 105, 109, 103, 33, 41, 90, 
    221, 210, 199, 179, 164, 149, 153, 137, 130, 118, 120, 72, 0, 83, 101, 
    149, 129, 134, 129, 129, 126, 131, 129, 129, 133, 96, 25, 61, 120, 106, 
    108, 119, 122, 122, 132, 133, 139, 148, 147, 138, 0, 21, 97, 105, 98, 
    117, 123, 123, 122, 133, 144, 138, 139, 156, 134, 26, 80, 105, 102, 101, 
    122, 123, 123, 119, 124, 140, 178, 168, 134, 54, 113, 41, 38, 90, 90, 
    125, 123, 116, 114, 125, 61, 0, 0, 0, 61, 156, 14, 24, 21, 63, 
    124, 121, 117, 118, 40, 59, 19, 64, 165, 230, 134, 12, 0, 17, 99, 
    120, 115, 56, 20, 0, 7, 68, 195, 144, 115, 83, 0, 61, 124, 131, 
    121, 194, 14, 17, 0, 12, 96, 113, 99, 75, 62, 103, 143, 95, 63, 
    140, 46, 0, 1, 0, 30, 129, 98, 39, 0, 1, 44, 47, 31, 0, 
    72, 6, 22, 0, 10, 59, 114, 111, 0, 7, 0, 58, 33, 0, 0, 
    50, 18, 32, 0, 75, 95, 140, 87, 0, 40, 21, 17, 27, 0, 14, 
    51, 21, 4, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 3, 
    58, 10, 0, 12, 2, 4, 3, 0, 0, 20, 0, 0, 0, 0, 8, 
    
    -- channel=107
    29, 39, 22, 31, 39, 30, 18, 36, 15, 31, 31, 13, 24, 0, 20, 
    19, 27, 34, 27, 23, 23, 14, 22, 15, 22, 0, 25, 44, 0, 15, 
    25, 36, 19, 23, 15, 17, 16, 15, 16, 10, 0, 54, 11, 0, 30, 
    11, 12, 15, 19, 12, 17, 8, 9, 11, 9, 76, 0, 18, 21, 25, 
    10, 15, 17, 21, 9, 5, 4, 8, 0, 1, 39, 0, 0, 14, 11, 
    15, 18, 19, 19, 0, 0, 0, 21, 44, 99, 25, 141, 0, 21, 9, 
    15, 21, 27, 4, 0, 27, 58, 59, 15, 0, 0, 230, 14, 0, 1, 
    18, 25, 0, 0, 23, 0, 42, 0, 0, 0, 48, 218, 107, 0, 0, 
    22, 0, 5, 0, 69, 0, 0, 0, 60, 73, 125, 192, 0, 0, 0, 
    0, 0, 159, 0, 70, 0, 0, 8, 49, 109, 63, 102, 0, 40, 72, 
    0, 39, 138, 27, 28, 0, 0, 34, 128, 135, 0, 0, 105, 83, 153, 
    0, 8, 3, 78, 0, 0, 0, 52, 237, 0, 14, 0, 17, 154, 12, 
    0, 0, 0, 67, 0, 0, 0, 49, 215, 0, 40, 0, 0, 143, 0, 
    0, 0, 22, 56, 0, 38, 52, 67, 144, 0, 55, 44, 0, 23, 0, 
    0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 39, 42, 0, 0, 0, 
    
    -- channel=108
    65, 79, 78, 81, 87, 73, 64, 74, 45, 60, 57, 39, 40, 17, 36, 
    74, 79, 77, 63, 59, 53, 46, 51, 42, 43, 18, 48, 46, 0, 36, 
    57, 68, 55, 48, 37, 38, 38, 39, 37, 31, 8, 79, 32, 10, 49, 
    34, 30, 32, 36, 32, 38, 41, 45, 43, 32, 78, 0, 42, 41, 46, 
    27, 31, 33, 38, 31, 36, 41, 53, 46, 84, 81, 7, 47, 44, 31, 
    30, 34, 37, 38, 19, 7, 27, 69, 78, 134, 107, 168, 0, 65, 33, 
    32, 38, 45, 23, 3, 39, 98, 91, 51, 0, 34, 324, 20, 15, 33, 
    35, 42, 10, 33, 60, 22, 68, 18, 0, 0, 138, 289, 125, 0, 0, 
    38, 15, 26, 34, 91, 0, 0, 17, 145, 174, 228, 253, 2, 0, 47, 
    9, 0, 190, 2, 83, 0, 0, 96, 140, 174, 127, 183, 59, 108, 137, 
    0, 52, 203, 50, 37, 0, 0, 118, 213, 163, 0, 0, 172, 148, 174, 
    0, 25, 64, 96, 0, 0, 0, 134, 306, 16, 37, 0, 83, 194, 32, 
    0, 7, 34, 96, 0, 36, 9, 139, 287, 0, 75, 0, 0, 165, 0, 
    0, 3, 39, 62, 0, 60, 79, 96, 181, 0, 88, 59, 0, 38, 0, 
    17, 23, 17, 25, 0, 0, 5, 7, 7, 0, 56, 51, 0, 0, 0, 
    
    -- channel=109
    100, 119, 140, 145, 138, 126, 123, 110, 89, 64, 59, 42, 2, 36, 39, 
    141, 121, 122, 118, 108, 95, 93, 84, 72, 63, 56, 16, 0, 15, 45, 
    92, 94, 95, 84, 75, 67, 69, 64, 59, 56, 0, 18, 6, 23, 37, 
    64, 62, 61, 62, 64, 62, 65, 60, 56, 39, 0, 4, 28, 46, 54, 
    55, 61, 62, 61, 64, 57, 51, 58, 48, 8, 0, 3, 53, 55, 49, 
    57, 61, 61, 61, 53, 29, 0, 0, 0, 0, 0, 0, 13, 40, 44, 
    61, 60, 56, 54, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 
    61, 59, 42, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    58, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=110
    127, 153, 161, 170, 166, 158, 151, 144, 138, 136, 106, 82, 75, 57, 78, 
    157, 137, 159, 162, 152, 140, 133, 125, 115, 102, 75, 64, 34, 37, 89, 
    147, 156, 142, 136, 123, 115, 114, 104, 98, 86, 43, 38, 20, 45, 89, 
    110, 112, 112, 111, 108, 109, 97, 84, 76, 71, 74, 39, 71, 106, 100, 
    105, 115, 119, 117, 109, 91, 83, 72, 10, 0, 0, 5, 73, 89, 95, 
    113, 116, 115, 114, 93, 8, 0, 0, 53, 52, 0, 23, 38, 57, 89, 
    115, 117, 116, 91, 44, 88, 84, 102, 65, 0, 0, 0, 12, 49, 71, 
    117, 114, 56, 27, 34, 2, 0, 0, 0, 0, 0, 56, 29, 1, 0, 
    119, 73, 56, 20, 40, 26, 0, 0, 0, 0, 8, 64, 0, 0, 0, 
    78, 0, 9, 4, 42, 11, 0, 0, 0, 59, 28, 0, 0, 0, 30, 
    61, 92, 17, 19, 26, 0, 0, 0, 49, 96, 75, 15, 14, 40, 115, 
    80, 8, 0, 22, 0, 0, 0, 0, 45, 0, 1, 25, 0, 58, 18, 
    57, 3, 0, 0, 0, 0, 0, 0, 18, 0, 0, 23, 23, 67, 34, 
    47, 25, 44, 58, 84, 127, 138, 145, 98, 6, 27, 29, 53, 32, 17, 
    37, 19, 0, 0, 0, 0, 0, 0, 4, 22, 44, 34, 6, 6, 0, 
    
    -- channel=111
    0, 8, 22, 25, 27, 29, 29, 24, 24, 5, 1, 3, 33, 26, 0, 
    28, 25, 32, 36, 35, 30, 27, 22, 18, 7, 0, 5, 0, 0, 0, 
    51, 39, 34, 30, 18, 12, 10, 4, 2, 0, 30, 29, 0, 0, 4, 
    12, 9, 9, 7, 7, 6, 3, 0, 0, 5, 1, 0, 0, 0, 5, 
    8, 10, 12, 11, 12, 21, 21, 0, 0, 0, 0, 5, 27, 15, 10, 
    7, 11, 12, 12, 5, 0, 21, 90, 119, 82, 0, 0, 28, 26, 11, 
    10, 10, 14, 6, 34, 39, 6, 1, 0, 0, 0, 0, 0, 28, 35, 
    12, 11, 6, 22, 5, 11, 0, 0, 0, 0, 0, 25, 6, 0, 0, 
    15, 0, 4, 12, 9, 0, 0, 4, 21, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 14, 0, 0, 64, 67, 0, 0, 0, 23, 
    32, 63, 7, 0, 0, 0, 0, 0, 28, 0, 5, 31, 17, 29, 19, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 21, 7, 5, 
    0, 4, 29, 41, 54, 66, 76, 77, 37, 3, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 4, 35, 0, 0, 0, 0, 
    
    -- channel=112
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 4, 16, 18, 18, 3, 
    0, 0, 0, 0, 0, 0, 0, 6, 13, 16, 0, 1, 0, 0, 0, 
    0, 4, 0, 0, 0, 17, 19, 9, 0, 0, 0, 0, 0, 0, 0, 
    50, 52, 0, 0, 6, 42, 16, 0, 2, 0, 1, 0, 3, 0, 1, 
    10, 0, 0, 0, 14, 60, 0, 0, 13, 0, 0, 9, 9, 0, 0, 
    0, 0, 0, 0, 18, 4, 0, 0, 17, 0, 0, 13, 0, 0, 0, 
    1, 9, 0, 0, 0, 53, 0, 13, 17, 0, 0, 0, 7, 0, 0, 
    15, 34, 43, 0, 9, 0, 24, 0, 8, 0, 0, 0, 13, 0, 0, 
    64, 29, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 42, 0, 18, 14, 14, 0, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 8, 33, 5, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 1, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 8, 12, 0, 0, 0, 1, 4, 0, 0, 0, 0, 
    
    -- channel=113
    148, 134, 149, 146, 151, 157, 127, 114, 96, 83, 62, 39, 21, 20, 12, 
    144, 131, 135, 104, 128, 134, 135, 112, 84, 87, 79, 78, 81, 88, 79, 
    128, 126, 87, 77, 92, 90, 101, 111, 125, 157, 152, 148, 127, 111, 81, 
    118, 130, 92, 43, 77, 94, 99, 115, 122, 149, 168, 144, 121, 103, 84, 
    215, 262, 222, 52, 72, 148, 172, 125, 121, 119, 140, 150, 149, 136, 127, 
    319, 328, 261, 59, 100, 172, 172, 138, 140, 124, 117, 139, 156, 164, 145, 
    298, 294, 285, 118, 92, 149, 151, 146, 168, 141, 118, 128, 142, 146, 110, 
    286, 305, 298, 252, 165, 137, 152, 152, 195, 170, 127, 111, 131, 118, 106, 
    329, 384, 425, 317, 335, 227, 211, 157, 187, 181, 148, 121, 133, 112, 70, 
    490, 532, 486, 386, 329, 267, 213, 163, 179, 188, 176, 133, 117, 64, 23, 
    570, 524, 275, 239, 188, 171, 149, 135, 172, 175, 161, 130, 101, 97, 38, 
    400, 328, 221, 201, 109, 85, 145, 82, 112, 146, 169, 157, 86, 114, 70, 
    200, 194, 188, 180, 146, 103, 133, 110, 116, 178, 214, 172, 107, 80, 108, 
    151, 155, 145, 104, 83, 106, 89, 102, 87, 115, 161, 148, 109, 60, 75, 
    106, 74, 59, 37, 50, 105, 90, 59, 39, 48, 63, 77, 56, 33, 33, 
    
    -- channel=114
    0, 0, 3, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    55, 51, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    35, 39, 37, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40, 48, 27, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    64, 96, 126, 36, 56, 2, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    136, 124, 16, 43, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    130, 101, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 25, 19, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=115
    12, 12, 13, 10, 0, 0, 0, 6, 10, 8, 12, 14, 15, 17, 19, 
    12, 11, 6, 11, 0, 0, 0, 0, 0, 7, 7, 9, 9, 10, 10, 
    10, 11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 6, 7, 
    9, 10, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 8, 2, 
    13, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 4, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 11, 14, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 8, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    4, 10, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 5, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 19, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 7, 11, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=116
    21, 20, 29, 28, 39, 40, 35, 28, 21, 23, 22, 18, 17, 20, 16, 
    20, 18, 28, 30, 44, 64, 53, 50, 35, 26, 27, 27, 31, 34, 32, 
    21, 21, 28, 30, 46, 58, 67, 71, 60, 45, 42, 46, 44, 40, 38, 
    22, 22, 11, 38, 45, 52, 60, 80, 81, 70, 57, 54, 42, 39, 46, 
    28, 36, 30, 25, 50, 60, 59, 64, 80, 79, 81, 67, 62, 60, 64, 
    45, 43, 17, 21, 36, 65, 57, 51, 67, 73, 77, 74, 80, 76, 67, 
    38, 35, 33, 0, 51, 62, 50, 64, 66, 59, 69, 79, 74, 72, 49, 
    36, 41, 45, 51, 20, 49, 53, 73, 67, 51, 63, 68, 65, 58, 47, 
    44, 44, 35, 41, 48, 41, 59, 67, 64, 49, 56, 62, 68, 62, 65, 
    50, 60, 66, 24, 74, 51, 79, 56, 59, 52, 58, 58, 61, 53, 64, 
    50, 45, 10, 42, 49, 65, 59, 58, 64, 62, 61, 53, 61, 64, 70, 
    42, 28, 9, 32, 28, 44, 56, 35, 49, 56, 55, 55, 67, 87, 61, 
    24, 30, 33, 41, 39, 45, 68, 42, 54, 61, 48, 59, 63, 84, 79, 
    34, 44, 53, 56, 59, 58, 54, 58, 55, 59, 53, 45, 64, 80, 86, 
    50, 55, 60, 66, 78, 76, 63, 71, 73, 66, 65, 64, 66, 82, 81, 
    
    -- channel=117
    31, 31, 32, 27, 48, 39, 34, 29, 29, 34, 31, 30, 31, 31, 27, 
    31, 30, 36, 37, 56, 71, 50, 48, 30, 32, 30, 27, 25, 23, 20, 
    34, 32, 38, 42, 67, 77, 86, 78, 38, 31, 27, 27, 22, 20, 20, 
    34, 33, 16, 61, 79, 85, 82, 83, 71, 55, 45, 33, 16, 19, 21, 
    25, 23, 20, 30, 80, 78, 67, 73, 82, 81, 81, 49, 28, 16, 18, 
    20, 19, 0, 27, 54, 88, 77, 72, 79, 82, 83, 76, 46, 14, 11, 
    19, 15, 9, 0, 70, 72, 63, 79, 73, 71, 78, 87, 51, 26, 11, 
    23, 20, 22, 0, 0, 61, 59, 76, 73, 68, 78, 84, 65, 40, 21, 
    22, 12, 0, 21, 11, 17, 38, 60, 79, 73, 77, 80, 79, 49, 20, 
    4, 1, 4, 0, 51, 10, 64, 49, 80, 78, 77, 78, 78, 35, 12, 
    0, 0, 0, 61, 67, 64, 73, 60, 78, 77, 71, 74, 66, 23, 12, 
    7, 11, 0, 22, 56, 83, 63, 44, 83, 78, 68, 66, 46, 36, 2, 
    23, 26, 26, 27, 15, 41, 63, 43, 76, 79, 64, 71, 35, 35, 18, 
    30, 33, 36, 30, 25, 26, 39, 56, 60, 76, 70, 70, 59, 27, 31, 
    31, 28, 27, 21, 25, 29, 33, 26, 25, 36, 55, 51, 33, 25, 17, 
    
    -- channel=118
    59, 54, 55, 55, 50, 38, 42, 44, 40, 37, 33, 28, 21, 17, 11, 
    58, 53, 53, 38, 33, 33, 23, 24, 29, 29, 19, 13, 10, 12, 12, 
    56, 53, 45, 24, 21, 9, 9, 3, 6, 31, 27, 27, 24, 26, 19, 
    46, 47, 25, 10, 11, 7, 0, 0, 0, 30, 37, 30, 24, 20, 5, 
    46, 54, 54, 0, 8, 22, 16, 0, 0, 0, 12, 13, 17, 1, 0, 
    82, 91, 73, 2, 7, 34, 38, 14, 4, 0, 0, 8, 11, 0, 0, 
    92, 88, 78, 10, 30, 33, 21, 15, 20, 8, 0, 3, 9, 16, 16, 
    83, 80, 79, 41, 3, 16, 11, 5, 28, 25, 3, 0, 16, 17, 10, 
    81, 85, 81, 58, 59, 37, 26, 3, 36, 35, 13, 4, 16, 11, 0, 
    101, 120, 134, 95, 91, 56, 43, 7, 32, 39, 25, 9, 12, 0, 0, 
    155, 151, 85, 96, 59, 49, 31, 13, 24, 30, 21, 8, 0, 0, 0, 
    150, 134, 63, 48, 29, 12, 23, 12, 27, 25, 24, 15, 0, 0, 0, 
    77, 71, 63, 47, 21, 7, 21, 12, 19, 32, 46, 31, 0, 0, 0, 
    46, 40, 36, 21, 4, 0, 0, 9, 0, 27, 47, 29, 2, 0, 0, 
    26, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=119
    25, 26, 25, 26, 40, 56, 49, 37, 30, 30, 33, 31, 32, 30, 33, 
    25, 26, 26, 42, 53, 70, 75, 72, 51, 35, 44, 42, 41, 36, 36, 
    27, 27, 31, 41, 68, 86, 95, 103, 83, 45, 41, 44, 40, 33, 38, 
    31, 30, 38, 54, 78, 89, 95, 101, 101, 79, 61, 62, 46, 41, 49, 
    33, 30, 27, 65, 75, 71, 78, 96, 107, 110, 102, 86, 64, 59, 60, 
    25, 26, 30, 61, 65, 70, 82, 92, 95, 105, 111, 98, 81, 61, 54, 
    22, 26, 31, 51, 49, 60, 86, 97, 87, 88, 102, 102, 80, 53, 42, 
    31, 32, 31, 49, 56, 60, 75, 91, 85, 85, 99, 103, 84, 68, 57, 
    32, 33, 35, 50, 43, 52, 56, 89, 86, 83, 95, 101, 91, 75, 62, 
    21, 13, 19, 33, 49, 55, 63, 94, 89, 86, 92, 102, 95, 79, 63, 
    12, 12, 53, 52, 64, 81, 82, 82, 86, 89, 90, 99, 95, 72, 65, 
    13, 24, 37, 38, 63, 82, 73, 65, 70, 86, 77, 85, 94, 70, 69, 
    34, 30, 36, 41, 52, 57, 63, 74, 72, 78, 67, 80, 90, 78, 66, 
    40, 43, 49, 59, 65, 58, 66, 76, 83, 75, 70, 83, 84, 83, 70, 
    46, 57, 66, 67, 65, 60, 67, 78, 77, 75, 75, 79, 80, 75, 68, 
    
    -- channel=120
    1, 0, 21, 2, 9, 1, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    1, 0, 13, 6, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 1, 0, 28, 0, 5, 12, 10, 8, 0, 0, 0, 0, 0, 0, 
    4, 7, 0, 1, 11, 5, 6, 11, 9, 22, 7, 0, 0, 0, 0, 
    1, 0, 0, 0, 12, 40, 0, 0, 0, 2, 18, 0, 3, 0, 0, 
    11, 6, 0, 0, 0, 46, 0, 0, 1, 0, 0, 25, 25, 0, 0, 
    14, 7, 0, 0, 22, 60, 0, 3, 6, 0, 0, 29, 3, 17, 0, 
    12, 8, 0, 0, 0, 19, 0, 13, 11, 0, 0, 1, 6, 9, 0, 
    18, 21, 0, 0, 0, 0, 1, 0, 16, 0, 0, 0, 17, 4, 0, 
    0, 2, 0, 0, 17, 0, 24, 0, 10, 0, 0, 0, 10, 0, 0, 
    3, 0, 0, 0, 24, 0, 19, 18, 11, 6, 0, 0, 1, 0, 0, 
    7, 4, 0, 0, 0, 23, 29, 0, 35, 25, 2, 0, 0, 33, 0, 
    5, 15, 6, 3, 0, 0, 31, 0, 12, 43, 0, 0, 0, 11, 7, 
    7, 8, 3, 4, 17, 0, 0, 1, 13, 44, 32, 0, 0, 1, 24, 
    2, 9, 9, 0, 27, 17, 0, 0, 0, 2, 28, 23, 0, 9, 4, 
    
    -- channel=121
    0, 1, 5, 11, 11, 1, 0, 4, 0, 1, 7, 6, 2, 0, 0, 
    1, 0, 4, 18, 2, 33, 12, 0, 5, 0, 0, 0, 0, 0, 0, 
    9, 6, 20, 26, 16, 10, 20, 9, 0, 0, 0, 0, 0, 5, 12, 
    0, 0, 0, 0, 14, 0, 0, 0, 16, 34, 5, 4, 0, 0, 0, 
    0, 0, 0, 0, 8, 1, 0, 0, 3, 8, 20, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 3, 0, 0, 4, 21, 5, 0, 0, 
    18, 14, 0, 0, 11, 57, 18, 2, 0, 0, 1, 16, 14, 29, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 15, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 11, 9, 32, 
    0, 0, 22, 1, 41, 0, 11, 0, 6, 0, 0, 0, 16, 8, 1, 
    0, 0, 58, 78, 64, 79, 44, 48, 13, 15, 16, 1, 0, 0, 0, 
    133, 127, 22, 0, 0, 32, 0, 0, 34, 17, 0, 0, 0, 10, 0, 
    48, 40, 18, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 1, 4, 
    5, 0, 19, 48, 38, 0, 0, 4, 17, 44, 65, 17, 12, 14, 18, 
    27, 48, 24, 0, 6, 4, 0, 5, 1, 0, 17, 29, 15, 7, 13, 
    
    -- channel=122
    50, 46, 56, 49, 69, 73, 55, 39, 38, 37, 24, 16, 13, 19, 16, 
    48, 44, 53, 46, 77, 89, 77, 69, 36, 41, 47, 54, 61, 64, 56, 
    43, 41, 36, 47, 69, 89, 97, 103, 88, 87, 85, 80, 68, 54, 41, 
    45, 50, 36, 64, 77, 95, 111, 128, 112, 81, 86, 72, 55, 56, 60, 
    102, 126, 99, 54, 89, 111, 128, 123, 124, 117, 110, 95, 85, 89, 95, 
    122, 113, 56, 58, 83, 128, 108, 105, 121, 131, 125, 111, 107, 102, 91, 
    92, 88, 84, 53, 80, 98, 97, 113, 118, 117, 117, 124, 104, 82, 52, 
    96, 110, 111, 95, 82, 117, 117, 132, 125, 111, 115, 116, 93, 73, 64, 
    125, 141, 158, 165, 137, 113, 115, 129, 116, 107, 117, 113, 107, 90, 56, 
    202, 208, 161, 96, 124, 85, 120, 111, 116, 114, 122, 113, 102, 61, 55, 
    169, 145, 44, 53, 84, 69, 91, 92, 118, 114, 107, 104, 99, 85, 72, 
    71, 33, 52, 79, 68, 82, 100, 70, 83, 102, 114, 114, 94, 100, 72, 
    45, 52, 55, 77, 74, 95, 98, 68, 98, 123, 116, 112, 97, 95, 85, 
    58, 76, 73, 52, 50, 72, 83, 86, 86, 91, 75, 93, 96, 82, 89, 
    58, 44, 53, 64, 81, 86, 84, 75, 76, 73, 78, 76, 70, 81, 70, 
    
    -- channel=123
    14, 17, 1, 24, 11, 14, 24, 20, 16, 11, 15, 16, 9, 0, 2, 
    14, 19, 4, 14, 12, 0, 25, 17, 19, 6, 2, 0, 0, 0, 9, 
    13, 15, 25, 5, 4, 0, 0, 0, 0, 4, 12, 14, 18, 24, 27, 
    8, 3, 30, 0, 0, 0, 0, 0, 0, 1, 13, 32, 18, 23, 17, 
    0, 0, 58, 49, 0, 0, 0, 8, 0, 0, 0, 11, 11, 21, 15, 
    18, 33, 105, 41, 0, 0, 7, 13, 0, 0, 0, 0, 0, 20, 26, 
    35, 41, 49, 95, 0, 0, 30, 0, 0, 2, 3, 0, 3, 8, 38, 
    21, 19, 39, 57, 89, 0, 9, 0, 0, 20, 7, 0, 0, 2, 16, 
    14, 7, 20, 39, 47, 61, 5, 19, 0, 12, 3, 1, 0, 8, 46, 
    2, 30, 89, 157, 30, 98, 0, 44, 0, 0, 4, 15, 0, 30, 12, 
    68, 100, 176, 40, 19, 44, 5, 10, 0, 2, 16, 8, 0, 10, 23, 
    124, 102, 77, 50, 38, 0, 0, 30, 0, 0, 0, 10, 18, 0, 46, 
    44, 37, 27, 19, 47, 17, 0, 25, 0, 0, 5, 13, 31, 0, 8, 
    13, 11, 30, 45, 25, 9, 2, 7, 4, 0, 5, 12, 12, 16, 0, 
    33, 36, 19, 13, 0, 0, 16, 25, 11, 3, 0, 7, 22, 2, 9, 
    
    -- channel=124
    57, 58, 42, 64, 60, 67, 66, 56, 50, 44, 40, 38, 28, 14, 21, 
    57, 62, 46, 47, 64, 42, 78, 58, 47, 42, 36, 32, 27, 26, 37, 
    52, 56, 59, 37, 57, 42, 42, 45, 35, 46, 58, 59, 54, 60, 60, 
    47, 44, 77, 16, 35, 34, 34, 40, 45, 51, 66, 79, 57, 59, 51, 
    40, 51, 128, 79, 22, 21, 56, 72, 52, 51, 46, 68, 53, 65, 56, 
    86, 105, 186, 74, 43, 1, 71, 84, 51, 57, 54, 39, 46, 70, 73, 
    104, 110, 122, 149, 18, 29, 93, 60, 48, 71, 68, 25, 60, 56, 78, 
    90, 91, 112, 120, 140, 0, 73, 44, 51, 91, 73, 46, 53, 44, 57, 
    87, 92, 125, 121, 142, 136, 82, 78, 49, 86, 74, 66, 33, 50, 74, 
    107, 133, 177, 264, 107, 186, 54, 111, 51, 69, 74, 80, 41, 71, 40, 
    182, 214, 241, 126, 91, 108, 62, 68, 58, 67, 79, 76, 47, 55, 47, 
    199, 180, 156, 106, 90, 33, 28, 68, 29, 42, 54, 79, 65, 24, 85, 
    104, 84, 81, 73, 95, 54, 29, 81, 29, 21, 76, 85, 90, 35, 51, 
    63, 57, 71, 78, 55, 55, 38, 52, 38, 24, 59, 75, 70, 50, 24, 
    65, 64, 52, 44, 14, 36, 57, 60, 37, 34, 20, 43, 59, 31, 34, 
    
    -- channel=125
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 17, 22, 19, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 18, 20, 28, 32, 17, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 9, 9, 9, 32, 34, 25, 14, 1, 0, 0, 0, 
    0, 0, 0, 7, 6, 0, 7, 28, 26, 40, 32, 17, 2, 3, 0, 
    0, 0, 0, 0, 0, 15, 19, 18, 8, 26, 32, 21, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 13, 23, 4, 14, 30, 24, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 20, 6, 13, 24, 23, 7, 0, 5, 
    0, 0, 0, 0, 0, 0, 4, 25, 5, 9, 17, 23, 10, 9, 11, 
    0, 0, 0, 4, 9, 18, 13, 32, 16, 10, 21, 26, 12, 5, 4, 
    0, 0, 0, 0, 11, 25, 0, 2, 23, 17, 11, 17, 16, 8, 11, 
    0, 0, 0, 0, 0, 0, 4, 4, 5, 4, 0, 15, 20, 12, 11, 
    0, 0, 0, 0, 7, 2, 4, 7, 11, 5, 7, 18, 20, 22, 12, 
    0, 4, 12, 13, 12, 3, 9, 20, 17, 11, 9, 14, 20, 23, 16, 
    
    -- channel=126
    0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 4, 7, 5, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 11, 0, 0, 0, 0, 0, 0, 0, 0, 3, 16, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 4, 6, 6, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 21, 
    0, 0, 0, 0, 4, 6, 0, 0, 0, 0, 0, 0, 2, 23, 37, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 60, 
    0, 0, 5, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 23, 36, 
    0, 0, 74, 36, 21, 29, 7, 9, 0, 0, 0, 0, 0, 0, 30, 
    77, 71, 5, 0, 3, 0, 0, 6, 0, 0, 0, 0, 6, 18, 26, 
    20, 18, 6, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 28, 19, 
    0, 0, 25, 56, 47, 9, 3, 5, 8, 14, 8, 0, 7, 36, 42, 
    38, 60, 44, 36, 34, 24, 22, 39, 37, 23, 26, 35, 37, 44, 50, 
    
    -- channel=127
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 6, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 27, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 8, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    54, 14, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=128
    0, 92, 52, 0, 0, 2, 0, 5, 0, 0, 93, 25, 0, 0, 0, 
    0, 47, 92, 0, 12, 0, 0, 7, 0, 0, 155, 0, 0, 0, 0, 
    0, 12, 137, 14, 48, 0, 0, 2, 0, 2, 74, 4, 0, 0, 0, 
    0, 102, 134, 0, 49, 0, 0, 0, 12, 61, 1, 50, 0, 0, 0, 
    0, 46, 0, 0, 77, 0, 0, 0, 11, 26, 22, 50, 0, 0, 4, 
    0, 0, 0, 0, 33, 0, 0, 0, 31, 36, 11, 62, 0, 0, 0, 
    0, 0, 0, 33, 0, 6, 0, 1, 0, 12, 14, 57, 0, 0, 0, 
    0, 0, 0, 99, 0, 0, 0, 0, 6, 0, 0, 0, 9, 0, 0, 
    0, 0, 0, 34, 0, 8, 0, 0, 15, 0, 11, 0, 30, 0, 29, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 0, 1, 12, 0, 0, 
    0, 0, 24, 0, 0, 0, 20, 0, 0, 0, 0, 16, 1, 0, 0, 
    0, 0, 43, 0, 0, 0, 17, 0, 0, 0, 43, 0, 11, 0, 0, 
    0, 0, 16, 0, 0, 0, 27, 0, 0, 0, 21, 0, 0, 0, 0, 
    0, 0, 13, 9, 0, 9, 0, 0, 0, 0, 12, 0, 0, 17, 6, 
    0, 0, 0, 29, 0, 0, 0, 0, 0, 21, 0, 2, 0, 11, 0, 
    
    -- channel=129
    0, 107, 301, 277, 271, 282, 288, 301, 282, 119, 235, 364, 348, 345, 334, 
    0, 37, 275, 275, 343, 287, 307, 346, 342, 183, 334, 419, 394, 379, 365, 
    0, 0, 248, 275, 402, 297, 217, 254, 255, 266, 399, 434, 440, 442, 428, 
    107, 141, 348, 283, 392, 375, 280, 219, 210, 302, 410, 470, 491, 448, 451, 
    347, 365, 403, 262, 357, 398, 354, 232, 221, 284, 405, 510, 510, 409, 406, 
    404, 400, 404, 302, 372, 376, 320, 228, 266, 297, 377, 516, 531, 436, 382, 
    410, 392, 322, 356, 338, 341, 310, 286, 326, 331, 370, 510, 534, 514, 425, 
    397, 380, 271, 400, 384, 369, 336, 284, 332, 321, 346, 369, 502, 502, 469, 
    386, 343, 350, 391, 431, 445, 382, 305, 282, 284, 333, 231, 312, 364, 443, 
    430, 376, 413, 400, 417, 423, 427, 393, 296, 316, 291, 275, 276, 298, 311, 
    456, 379, 426, 431, 432, 363, 384, 399, 383, 295, 254, 300, 320, 275, 249, 
    448, 385, 426, 456, 434, 353, 392, 388, 368, 248, 277, 294, 330, 280, 239, 
    430, 382, 410, 446, 366, 248, 379, 357, 314, 228, 270, 262, 268, 261, 252, 
    408, 350, 373, 454, 386, 314, 329, 289, 241, 195, 246, 239, 205, 235, 274, 
    348, 339, 312, 439, 408, 354, 248, 240, 183, 185, 222, 240, 218, 232, 255, 
    
    -- channel=130
    0, 51, 56, 28, 29, 39, 26, 33, 0, 0, 62, 51, 44, 41, 38, 
    0, 7, 83, 51, 42, 31, 58, 54, 55, 0, 79, 61, 56, 54, 52, 
    0, 0, 75, 43, 104, 10, 40, 81, 63, 30, 77, 88, 74, 72, 59, 
    0, 0, 46, 28, 124, 46, 0, 0, 24, 83, 85, 107, 95, 84, 98, 
    5, 33, 57, 0, 103, 92, 59, 8, 36, 71, 94, 111, 99, 41, 82, 
    58, 70, 62, 14, 85, 85, 50, 17, 29, 58, 84, 131, 97, 29, 41, 
    55, 61, 45, 59, 52, 71, 40, 55, 42, 62, 80, 124, 106, 69, 24, 
    50, 70, 9, 114, 60, 67, 57, 44, 71, 63, 66, 138, 132, 101, 79, 
    26, 57, 51, 96, 77, 63, 48, 20, 75, 33, 54, 0, 118, 97, 116, 
    40, 44, 84, 71, 96, 118, 100, 44, 0, 58, 43, 41, 24, 36, 73, 
    69, 42, 96, 75, 76, 45, 101, 99, 63, 42, 36, 46, 55, 33, 38, 
    77, 34, 105, 99, 89, 62, 71, 75, 66, 7, 48, 49, 65, 30, 12, 
    64, 43, 89, 97, 60, 71, 93, 75, 55, 18, 52, 40, 62, 45, 25, 
    55, 28, 71, 101, 46, 37, 59, 53, 35, 16, 39, 31, 14, 41, 40, 
    52, 27, 50, 115, 69, 59, 35, 42, 7, 20, 28, 31, 8, 31, 44, 
    
    -- channel=131
    25, 10, 0, 0, 0, 0, 0, 0, 0, 2, 16, 0, 0, 0, 0, 
    25, 15, 0, 2, 13, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 
    24, 18, 0, 0, 15, 18, 6, 0, 0, 22, 0, 0, 0, 0, 0, 
    4, 24, 0, 0, 10, 27, 18, 6, 11, 10, 0, 2, 3, 0, 0, 
    0, 0, 0, 1, 3, 18, 12, 13, 14, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 14, 13, 26, 12, 18, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 24, 12, 28, 8, 11, 10, 0, 0, 0, 0, 
    0, 0, 3, 0, 8, 9, 27, 9, 10, 6, 0, 0, 0, 0, 0, 
    0, 0, 12, 0, 18, 12, 20, 14, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 6, 21, 25, 4, 0, 0, 0, 2, 0, 0, 
    0, 0, 2, 3, 2, 3, 2, 9, 12, 0, 8, 0, 0, 3, 0, 
    0, 0, 0, 9, 2, 15, 0, 4, 0, 6, 0, 0, 0, 0, 2, 
    0, 0, 0, 5, 1, 28, 0, 0, 0, 1, 0, 2, 0, 5, 0, 
    0, 0, 0, 2, 12, 6, 0, 0, 0, 6, 0, 1, 2, 0, 0, 
    0, 0, 0, 4, 8, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    
    -- channel=132
    16, 79, 99, 84, 71, 91, 91, 90, 60, 30, 72, 94, 101, 102, 102, 
    17, 47, 104, 80, 45, 58, 75, 79, 76, 29, 87, 77, 84, 91, 94, 
    20, 27, 100, 76, 58, 18, 50, 72, 63, 45, 69, 64, 62, 68, 72, 
    15, 41, 86, 65, 69, 31, 32, 40, 49, 70, 56, 72, 63, 58, 68, 
    51, 66, 64, 41, 70, 48, 44, 31, 44, 57, 67, 78, 59, 51, 76, 
    63, 68, 63, 48, 68, 51, 38, 31, 40, 48, 55, 78, 58, 41, 64, 
    66, 65, 66, 62, 45, 39, 35, 46, 47, 45, 53, 81, 64, 52, 50, 
    62, 69, 51, 97, 51, 44, 35, 42, 53, 64, 54, 97, 80, 63, 54, 
    45, 62, 64, 89, 45, 45, 34, 29, 82, 50, 62, 41, 91, 65, 82, 
    52, 59, 68, 53, 60, 57, 44, 38, 32, 62, 68, 72, 62, 68, 75, 
    57, 45, 63, 57, 55, 44, 64, 56, 48, 65, 60, 74, 66, 57, 65, 
    61, 43, 72, 56, 56, 56, 69, 62, 58, 48, 74, 64, 66, 57, 54, 
    57, 59, 73, 52, 42, 65, 75, 68, 61, 51, 71, 59, 69, 61, 57, 
    56, 55, 71, 54, 50, 64, 77, 66, 61, 57, 67, 57, 53, 68, 63, 
    56, 54, 67, 59, 46, 58, 59, 70, 53, 58, 63, 62, 54, 66, 66, 
    
    -- channel=133
    26, 75, 30, 0, 16, 13, 8, 8, 0, 0, 39, 21, 3, 6, 3, 
    26, 57, 60, 0, 0, 15, 11, 11, 5, 0, 59, 9, 4, 6, 1, 
    24, 38, 76, 5, 6, 0, 16, 35, 8, 0, 48, 20, 4, 3, 0, 
    5, 28, 66, 1, 18, 0, 0, 0, 15, 33, 17, 17, 0, 2, 13, 
    0, 24, 25, 0, 35, 0, 0, 0, 13, 20, 27, 27, 5, 6, 42, 
    10, 20, 19, 0, 16, 1, 0, 0, 13, 17, 26, 37, 13, 5, 38, 
    20, 17, 14, 2, 8, 6, 0, 0, 4, 11, 24, 39, 14, 3, 10, 
    21, 15, 0, 24, 0, 1, 0, 12, 4, 18, 17, 48, 18, 16, 11, 
    11, 21, 0, 21, 0, 0, 0, 0, 40, 0, 14, 0, 68, 27, 42, 
    12, 13, 9, 0, 19, 12, 0, 0, 0, 12, 10, 8, 4, 15, 40, 
    16, 8, 17, 5, 0, 0, 23, 4, 0, 10, 1, 15, 7, 0, 14, 
    24, 4, 31, 0, 0, 0, 11, 0, 4, 0, 27, 7, 9, 0, 0, 
    24, 24, 30, 3, 0, 0, 15, 5, 0, 0, 25, 5, 21, 3, 6, 
    21, 30, 36, 13, 0, 0, 11, 7, 5, 4, 24, 10, 5, 24, 10, 
    23, 31, 34, 24, 0, 7, 0, 9, 2, 22, 17, 16, 3, 22, 16, 
    
    -- channel=134
    8, 26, 31, 19, 31, 16, 13, 19, 17, 10, 40, 45, 20, 19, 16, 
    8, 17, 52, 29, 70, 54, 49, 51, 59, 10, 63, 70, 52, 42, 32, 
    5, 11, 50, 32, 103, 69, 55, 68, 59, 37, 100, 101, 86, 80, 69, 
    0, 5, 67, 50, 109, 83, 42, 40, 46, 72, 107, 107, 109, 111, 105, 
    51, 60, 89, 37, 99, 106, 84, 49, 55, 70, 101, 120, 119, 90, 97, 
    84, 90, 91, 45, 89, 100, 83, 48, 66, 73, 97, 131, 127, 90, 81, 
    84, 80, 66, 64, 86, 91, 82, 58, 83, 87, 96, 129, 129, 112, 80, 
    86, 78, 30, 78, 89, 96, 84, 76, 77, 77, 91, 105, 120, 129, 104, 
    83, 75, 50, 83, 99, 99, 91, 73, 63, 47, 71, 25, 95, 102, 105, 
    92, 74, 93, 85, 114, 126, 110, 84, 49, 59, 61, 39, 30, 52, 73, 
    105, 89, 105, 97, 94, 88, 102, 103, 85, 65, 38, 50, 60, 47, 45, 
    108, 88, 109, 110, 105, 65, 80, 83, 84, 37, 46, 57, 67, 47, 35, 
    102, 88, 100, 116, 95, 40, 82, 76, 65, 34, 53, 48, 65, 48, 41, 
    94, 76, 86, 119, 79, 31, 66, 55, 43, 26, 47, 42, 35, 42, 47, 
    83, 72, 73, 126, 96, 82, 44, 38, 27, 26, 39, 43, 29, 40, 50, 
    
    -- channel=135
    20, 23, 51, 63, 40, 60, 65, 60, 55, 48, 36, 49, 70, 72, 76, 
    21, 20, 34, 62, 18, 36, 40, 48, 51, 59, 20, 46, 58, 62, 65, 
    24, 20, 22, 58, 10, 27, 33, 31, 37, 40, 18, 41, 42, 38, 44, 
    52, 48, 19, 54, 11, 24, 34, 34, 30, 24, 20, 32, 28, 32, 42, 
    58, 40, 43, 64, 17, 18, 26, 34, 23, 22, 25, 32, 38, 60, 54, 
    52, 47, 47, 62, 23, 19, 27, 39, 17, 20, 22, 29, 38, 60, 65, 
    58, 58, 64, 42, 34, 28, 23, 26, 18, 19, 27, 29, 43, 47, 60, 
    58, 53, 58, 22, 30, 18, 25, 19, 29, 43, 29, 41, 39, 42, 53, 
    58, 53, 41, 23, 28, 19, 24, 26, 39, 52, 35, 59, 44, 50, 49, 
    56, 53, 29, 32, 31, 22, 20, 28, 38, 38, 43, 49, 50, 44, 45, 
    49, 50, 32, 35, 35, 40, 26, 30, 33, 40, 50, 39, 35, 47, 43, 
    49, 53, 33, 25, 27, 47, 30, 39, 36, 55, 41, 42, 33, 45, 48, 
    51, 61, 47, 27, 30, 56, 28, 46, 46, 51, 39, 45, 36, 44, 44, 
    55, 65, 57, 25, 35, 38, 39, 50, 50, 54, 40, 45, 47, 41, 42, 
    57, 60, 61, 17, 34, 36, 50, 46, 49, 45, 44, 42, 48, 40, 42, 
    
    -- channel=136
    0, 176, 48, 0, 0, 19, 0, 4, 0, 0, 134, 8, 0, 0, 0, 
    3, 108, 107, 29, 0, 0, 25, 19, 0, 0, 144, 0, 0, 0, 0, 
    2, 40, 155, 23, 50, 0, 9, 56, 12, 20, 55, 31, 0, 0, 0, 
    0, 31, 71, 0, 90, 0, 0, 0, 11, 98, 9, 63, 0, 0, 36, 
    0, 27, 0, 0, 89, 12, 0, 0, 22, 72, 44, 58, 0, 0, 43, 
    0, 9, 0, 0, 43, 5, 0, 0, 0, 50, 44, 82, 0, 0, 0, 
    0, 5, 0, 21, 0, 22, 0, 37, 0, 30, 35, 75, 6, 0, 0, 
    0, 18, 0, 100, 0, 1, 0, 0, 37, 16, 1, 94, 77, 0, 12, 
    0, 21, 0, 45, 0, 0, 0, 0, 74, 0, 0, 0, 113, 27, 96, 
    0, 0, 8, 0, 23, 20, 9, 0, 0, 25, 0, 10, 9, 0, 57, 
    0, 0, 45, 0, 0, 0, 55, 22, 0, 0, 14, 15, 9, 0, 0, 
    0, 0, 70, 3, 0, 0, 17, 0, 0, 0, 50, 1, 17, 0, 0, 
    0, 0, 58, 3, 0, 37, 36, 4, 0, 0, 41, 2, 11, 12, 0, 
    0, 0, 65, 21, 0, 0, 0, 3, 0, 0, 26, 5, 0, 44, 8, 
    0, 0, 44, 57, 0, 0, 0, 13, 0, 37, 14, 8, 0, 17, 19, 
    
    -- channel=137
    0, 38, 0, 0, 0, 2, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    1, 28, 30, 21, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 16, 0, 0, 0, 28, 64, 69, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 1, 29, 0, 0, 0, 0, 1, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 3, 2, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 1, 0, 0, 0, 0, 15, 0, 7, 111, 56, 4, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 19, 1, 0, 0, 81, 83, 47, 
    0, 0, 0, 0, 4, 33, 8, 0, 0, 0, 7, 0, 0, 0, 39, 
    0, 0, 0, 0, 0, 0, 13, 12, 0, 0, 15, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 12, 0, 0, 45, 3, 14, 17, 7, 6, 9, 29, 25, 0, 
    0, 0, 29, 0, 0, 0, 4, 20, 20, 23, 0, 0, 0, 6, 0, 
    33, 0, 32, 14, 0, 0, 30, 25, 14, 2, 7, 0, 0, 0, 15, 
    
    -- channel=138
    0, 108, 161, 131, 137, 152, 156, 158, 129, 70, 124, 183, 181, 181, 175, 
    0, 62, 146, 117, 124, 136, 137, 156, 140, 53, 189, 177, 175, 178, 174, 
    4, 22, 141, 137, 129, 86, 81, 100, 81, 95, 176, 156, 165, 176, 177, 
    81, 104, 211, 123, 121, 107, 119, 90, 87, 138, 134, 178, 177, 150, 155, 
    139, 185, 157, 93, 134, 120, 112, 68, 83, 115, 145, 194, 173, 137, 163, 
    152, 156, 147, 120, 141, 120, 87, 67, 102, 120, 138, 188, 179, 152, 161, 
    159, 151, 124, 131, 110, 105, 95, 106, 112, 114, 136, 192, 181, 176, 172, 
    152, 147, 106, 163, 135, 119, 90, 116, 101, 129, 118, 142, 162, 163, 164, 
    137, 132, 130, 172, 133, 153, 131, 83, 136, 107, 125, 107, 129, 104, 170, 
    153, 157, 152, 137, 139, 123, 117, 122, 135, 135, 109, 117, 134, 133, 133, 
    161, 136, 143, 156, 155, 114, 129, 127, 117, 115, 97, 139, 132, 103, 112, 
    161, 126, 159, 149, 145, 117, 155, 140, 130, 84, 137, 117, 126, 115, 96, 
    156, 138, 155, 138, 102, 95, 140, 130, 105, 88, 120, 104, 102, 93, 106, 
    148, 135, 150, 144, 122, 160, 127, 110, 93, 81, 111, 101, 83, 110, 117, 
    121, 130, 136, 136, 130, 128, 92, 100, 73, 97, 99, 105, 95, 117, 103, 
    
    -- channel=139
    0, 0, 0, 45, 20, 15, 32, 16, 57, 73, 0, 13, 37, 37, 45, 
    0, 0, 0, 26, 28, 35, 25, 27, 55, 134, 0, 41, 46, 41, 48, 
    0, 0, 0, 7, 3, 120, 37, 4, 54, 24, 0, 27, 47, 38, 47, 
    38, 0, 0, 74, 0, 87, 62, 53, 7, 0, 42, 0, 65, 91, 39, 
    73, 0, 39, 111, 0, 47, 79, 102, 10, 0, 10, 1, 67, 110, 13, 
    56, 38, 60, 75, 4, 56, 92, 60, 9, 0, 12, 0, 66, 104, 37, 
    55, 46, 89, 26, 44, 18, 72, 19, 54, 18, 9, 0, 59, 79, 70, 
    66, 43, 115, 0, 69, 54, 66, 45, 34, 31, 57, 18, 34, 84, 53, 
    91, 27, 53, 0, 60, 49, 60, 101, 0, 66, 38, 65, 0, 61, 0, 
    74, 38, 35, 59, 37, 54, 67, 78, 60, 4, 74, 29, 16, 40, 11, 
    58, 78, 16, 48, 49, 99, 10, 47, 86, 81, 35, 10, 30, 64, 34, 
    52, 94, 0, 56, 72, 96, 24, 52, 67, 105, 0, 43, 28, 59, 56, 
    59, 72, 7, 55, 109, 43, 18, 60, 81, 71, 2, 43, 38, 44, 40, 
    69, 69, 0, 35, 94, 30, 62, 53, 61, 46, 8, 31, 53, 0, 24, 
    66, 51, 10, 14, 73, 70, 85, 39, 66, 0, 22, 22, 40, 8, 28, 
    
    -- channel=140
    4, 0, 82, 109, 102, 95, 111, 95, 136, 115, 0, 103, 125, 122, 129, 
    1, 0, 32, 77, 108, 107, 100, 104, 133, 190, 0, 143, 145, 138, 141, 
    4, 0, 0, 68, 83, 198, 93, 73, 122, 89, 49, 127, 151, 144, 150, 
    80, 0, 0, 138, 60, 179, 132, 110, 64, 10, 135, 95, 166, 188, 136, 
    163, 64, 134, 180, 27, 134, 164, 160, 68, 38, 98, 105, 184, 213, 104, 
    152, 124, 157, 153, 74, 132, 169, 119, 77, 49, 92, 97, 185, 222, 133, 
    153, 134, 165, 115, 119, 101, 154, 75, 124, 86, 90, 97, 173, 201, 169, 
    164, 128, 195, 33, 152, 128, 145, 110, 109, 90, 132, 87, 133, 197, 161, 
    194, 109, 147, 57, 155, 142, 142, 186, 33, 130, 126, 128, 26, 153, 88, 
    183, 121, 125, 146, 123, 145, 158, 163, 140, 87, 141, 102, 81, 113, 76, 
    165, 169, 109, 141, 145, 180, 92, 130, 180, 150, 101, 80, 103, 135, 99, 
    155, 195, 75, 154, 167, 171, 106, 133, 151, 173, 47, 109, 106, 130, 117, 
    162, 171, 87, 152, 205, 93, 107, 138, 157, 134, 67, 106, 100, 109, 105, 
    166, 164, 74, 135, 193, 106, 132, 125, 128, 95, 69, 93, 110, 52, 95, 
    152, 147, 74, 106, 167, 157, 150, 98, 122, 48, 77, 85, 98, 66, 87, 
    
    -- channel=141
    0, 0, 15, 0, 14, 20, 15, 7, 0, 0, 0, 0, 9, 10, 12, 
    0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 10, 
    0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=142
    13, 13, 5, 10, 12, 6, 5, 0, 0, 17, 0, 0, 0, 0, 5, 
    12, 24, 17, 4, 0, 0, 3, 0, 2, 12, 0, 0, 0, 0, 3, 
    13, 22, 0, 0, 0, 3, 38, 46, 52, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 20, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 29, 0, 0, 0, 0, 3, 0, 0, 13, 50, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 11, 0, 9, 40, 41, 0, 
    0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 30, 6, 0, 0, 32, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 29, 9, 0, 0, 15, 14, 
    0, 0, 0, 0, 0, 8, 0, 0, 2, 24, 0, 8, 0, 6, 7, 
    0, 0, 0, 0, 28, 50, 3, 15, 28, 25, 4, 13, 33, 20, 5, 
    0, 0, 0, 0, 0, 0, 25, 27, 34, 26, 5, 10, 20, 7, 0, 
    6, 0, 0, 0, 0, 6, 42, 29, 37, 4, 13, 4, 1, 1, 17, 
    
    -- channel=143
    0, 16, 2, 0, 3, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 17, 10, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 17, 23, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 4, 41, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 2, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 6, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=144
    0, 0, 0, 0, 0, 3, 9, 41, 23, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 16, 
    0, 0, 0, 0, 48, 32, 15, 0, 3, 18, 64, 11, 0, 0, 16, 
    0, 0, 0, 0, 106, 0, 0, 0, 0, 0, 0, 46, 0, 0, 0, 
    0, 0, 0, 0, 61, 0, 0, 0, 0, 0, 0, 62, 10, 0, 29, 
    6, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 80, 0, 0, 
    4, 0, 0, 0, 17, 0, 0, 0, 8, 0, 0, 18, 12, 0, 7, 
    0, 0, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 15, 109, 
    0, 0, 69, 0, 47, 0, 0, 0, 90, 79, 3, 65, 103, 0, 64, 
    0, 0, 14, 0, 1, 0, 0, 29, 0, 0, 0, 0, 0, 0, 113, 
    0, 0, 12, 0, 0, 3, 49, 0, 47, 0, 2, 71, 0, 59, 49, 
    0, 0, 34, 40, 0, 0, 1, 0, 82, 0, 3, 8, 0, 0, 102, 
    0, 0, 32, 5, 0, 0, 0, 6, 18, 188, 0, 0, 0, 30, 123, 
    5, 0, 0, 0, 0, 0, 5, 21, 33, 26, 0, 0, 0, 61, 87, 
    0, 0, 0, 0, 0, 0, 0, 11, 11, 13, 8, 0, 0, 48, 150, 
    
    -- channel=145
    495, 489, 480, 368, 370, 382, 414, 460, 514, 513, 489, 503, 468, 455, 412, 
    547, 547, 514, 289, 284, 302, 299, 327, 382, 428, 446, 497, 502, 441, 467, 
    553, 552, 499, 227, 245, 288, 280, 272, 265, 284, 414, 513, 465, 385, 426, 
    551, 537, 468, 248, 322, 404, 346, 329, 331, 341, 363, 463, 475, 411, 354, 
    548, 529, 370, 202, 291, 300, 284, 298, 324, 331, 360, 445, 526, 499, 455, 
    514, 488, 343, 169, 186, 240, 227, 220, 227, 257, 282, 352, 518, 554, 554, 
    448, 371, 300, 218, 214, 235, 221, 184, 209, 243, 196, 258, 387, 449, 551, 
    389, 208, 293, 262, 178, 165, 143, 100, 74, 82, 68, 76, 180, 269, 518, 
    387, 184, 289, 117, 186, 203, 229, 200, 216, 249, 252, 213, 269, 273, 456, 
    418, 151, 203, 49, 129, 108, 128, 197, 271, 251, 244, 242, 276, 167, 355, 
    428, 168, 141, 86, 34, 85, 179, 95, 193, 179, 170, 251, 143, 214, 325, 
    406, 110, 149, 195, 53, 20, 88, 35, 141, 209, 244, 265, 68, 132, 267, 
    375, 247, 196, 243, 109, 13, 0, 10, 54, 328, 373, 246, 27, 78, 276, 
    373, 343, 232, 212, 145, 42, 8, 32, 88, 233, 283, 204, 0, 91, 278, 
    343, 319, 259, 136, 124, 68, 47, 60, 79, 120, 177, 165, 14, 86, 311, 
    
    -- channel=146
    87, 83, 91, 58, 70, 68, 58, 60, 94, 103, 95, 109, 56, 68, 37, 
    118, 117, 108, 41, 95, 117, 122, 141, 157, 132, 98, 119, 112, 69, 96, 
    131, 133, 104, 0, 74, 66, 56, 40, 64, 88, 124, 115, 96, 55, 105, 
    130, 125, 108, 9, 130, 122, 80, 111, 96, 94, 86, 152, 89, 45, 53, 
    133, 118, 94, 38, 116, 120, 99, 109, 116, 114, 93, 137, 121, 64, 45, 
    149, 115, 48, 5, 95, 82, 81, 94, 95, 107, 126, 125, 167, 131, 132, 
    130, 90, 89, 17, 40, 84, 72, 54, 78, 85, 44, 97, 159, 170, 146, 
    100, 41, 93, 26, 72, 36, 46, 39, 56, 50, 42, 66, 102, 117, 192, 
    71, 0, 89, 23, 64, 66, 43, 0, 0, 0, 0, 0, 24, 69, 180, 
    82, 0, 80, 0, 62, 17, 56, 108, 81, 108, 96, 96, 112, 43, 162, 
    104, 0, 9, 0, 0, 28, 22, 0, 83, 31, 40, 54, 29, 48, 124, 
    109, 0, 51, 7, 0, 0, 81, 0, 93, 51, 48, 102, 0, 72, 132, 
    112, 0, 8, 60, 0, 0, 0, 0, 1, 93, 43, 0, 0, 4, 115, 
    107, 96, 37, 48, 26, 0, 0, 0, 7, 110, 119, 21, 0, 27, 117, 
    104, 83, 42, 18, 23, 0, 0, 0, 0, 32, 76, 31, 0, 17, 122, 
    
    -- channel=147
    13, 9, 11, 14, 21, 25, 19, 9, 1, 6, 0, 8, 13, 0, 5, 
    18, 17, 13, 39, 42, 52, 58, 47, 33, 13, 5, 3, 4, 0, 0, 
    20, 20, 25, 59, 88, 88, 96, 92, 85, 60, 29, 3, 0, 0, 0, 
    20, 16, 35, 63, 72, 75, 78, 102, 100, 97, 38, 18, 19, 0, 0, 
    20, 19, 36, 91, 73, 84, 101, 98, 92, 95, 84, 39, 18, 21, 20, 
    21, 18, 61, 67, 76, 94, 93, 90, 90, 85, 76, 56, 25, 20, 20, 
    21, 29, 35, 80, 78, 92, 97, 93, 89, 73, 68, 51, 32, 39, 24, 
    15, 35, 43, 24, 83, 84, 79, 66, 58, 66, 58, 49, 67, 71, 32, 
    28, 50, 11, 61, 61, 53, 72, 72, 53, 56, 49, 46, 45, 57, 37, 
    33, 45, 25, 59, 49, 63, 56, 70, 59, 69, 69, 67, 56, 77, 54, 
    34, 62, 34, 50, 47, 59, 70, 43, 64, 59, 64, 62, 59, 66, 53, 
    51, 58, 46, 50, 49, 34, 36, 64, 28, 55, 45, 23, 72, 35, 69, 
    67, 83, 43, 42, 63, 40, 34, 38, 49, 32, 34, 31, 46, 53, 57, 
    60, 63, 65, 42, 57, 50, 35, 38, 38, 28, 64, 45, 51, 43, 69, 
    73, 75, 64, 59, 50, 50, 41, 43, 46, 49, 51, 56, 45, 42, 66, 
    
    -- channel=148
    41, 42, 40, 38, 43, 46, 45, 47, 55, 50, 51, 53, 34, 55, 36, 
    45, 45, 44, 11, 16, 11, 17, 25, 35, 43, 50, 56, 54, 46, 62, 
    44, 45, 36, 0, 0, 0, 0, 0, 0, 0, 39, 60, 50, 40, 72, 
    43, 39, 33, 0, 23, 17, 0, 0, 0, 0, 10, 54, 45, 46, 56, 
    47, 41, 16, 0, 4, 0, 0, 0, 0, 0, 0, 47, 50, 28, 39, 
    56, 40, 4, 0, 10, 0, 0, 0, 0, 0, 0, 16, 51, 44, 45, 
    58, 34, 38, 0, 0, 0, 0, 0, 0, 0, 0, 18, 44, 46, 46, 
    56, 23, 51, 19, 0, 0, 0, 0, 5, 1, 0, 16, 17, 2, 57, 
    46, 7, 60, 11, 8, 29, 9, 0, 5, 19, 0, 3, 25, 18, 69, 
    33, 0, 45, 0, 24, 0, 3, 17, 4, 0, 0, 0, 5, 0, 45, 
    38, 0, 26, 0, 4, 15, 1, 0, 15, 0, 0, 0, 5, 0, 47, 
    21, 0, 28, 9, 0, 10, 32, 0, 60, 18, 18, 44, 0, 29, 32, 
    12, 0, 13, 16, 0, 0, 13, 13, 19, 54, 33, 0, 3, 16, 38, 
    14, 8, 0, 13, 2, 0, 12, 17, 20, 45, 12, 0, 0, 26, 30, 
    2, 0, 0, 4, 5, 0, 8, 8, 11, 14, 20, 2, 0, 20, 30, 
    
    -- channel=149
    0, 0, 0, 0, 0, 0, 0, 5, 15, 3, 6, 3, 0, 22, 0, 
    0, 0, 0, 0, 0, 0, 5, 10, 14, 20, 13, 17, 2, 10, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 26, 8, 4, 7, 45, 
    0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 25, 28, 0, 0, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 
    0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 6, 22, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 39, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 7, 0, 10, 16, 6, 2, 32, 
    0, 0, 34, 0, 3, 0, 0, 0, 0, 0, 0, 0, 2, 0, 38, 
    0, 0, 22, 0, 20, 0, 16, 9, 0, 1, 0, 0, 0, 0, 38, 
    0, 0, 19, 0, 8, 7, 0, 0, 8, 0, 0, 0, 0, 0, 26, 
    0, 0, 4, 0, 0, 20, 46, 0, 62, 0, 0, 30, 0, 35, 24, 
    0, 0, 4, 0, 0, 5, 18, 19, 19, 30, 0, 0, 0, 7, 31, 
    0, 0, 0, 0, 0, 0, 16, 20, 12, 47, 0, 0, 0, 23, 15, 
    0, 0, 0, 0, 1, 0, 9, 11, 11, 11, 12, 0, 0, 19, 25, 
    
    -- channel=150
    121, 119, 124, 94, 92, 92, 93, 102, 130, 131, 127, 129, 105, 109, 94, 
    143, 143, 141, 89, 122, 132, 130, 145, 153, 137, 122, 134, 130, 110, 113, 
    152, 153, 136, 70, 118, 131, 120, 120, 132, 139, 120, 134, 122, 97, 111, 
    151, 151, 131, 90, 144, 139, 142, 166, 152, 144, 148, 140, 114, 91, 84, 
    149, 148, 123, 96, 147, 156, 143, 158, 162, 156, 152, 141, 133, 112, 85, 
    141, 142, 85, 90, 123, 129, 134, 139, 141, 149, 155, 151, 162, 152, 152, 
    127, 108, 95, 66, 92, 128, 127, 109, 114, 126, 97, 115, 154, 148, 156, 
    98, 61, 72, 75, 109, 102, 100, 92, 89, 85, 85, 90, 114, 130, 170, 
    86, 32, 92, 57, 94, 83, 81, 52, 38, 43, 41, 31, 78, 105, 153, 
    106, 48, 86, 19, 85, 72, 92, 97, 126, 131, 130, 126, 132, 91, 130, 
    116, 35, 63, 43, 41, 58, 65, 68, 98, 93, 95, 98, 79, 88, 111, 
    130, 49, 61, 67, 28, 38, 90, 41, 82, 76, 88, 120, 36, 101, 100, 
    135, 56, 62, 107, 46, 22, 21, 28, 38, 93, 92, 79, 31, 42, 104, 
    133, 130, 96, 95, 74, 30, 17, 27, 40, 124, 128, 102, 13, 53, 112, 
    138, 125, 105, 72, 72, 40, 29, 37, 48, 69, 96, 83, 17, 52, 120, 
    
    -- channel=151
    24, 23, 18, 33, 21, 11, 17, 14, 14, 23, 29, 27, 32, 34, 46, 
    12, 13, 13, 21, 0, 0, 0, 0, 0, 2, 37, 20, 28, 43, 44, 
    11, 11, 15, 20, 0, 0, 0, 0, 0, 0, 0, 18, 26, 43, 43, 
    11, 9, 18, 4, 0, 0, 0, 0, 0, 0, 0, 9, 29, 37, 41, 
    12, 11, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 21, 25, 
    9, 10, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 10, 
    6, 19, 16, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 29, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 28, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 26, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 31, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 
    0, 17, 0, 0, 4, 2, 0, 11, 0, 0, 0, 0, 16, 0, 0, 
    0, 0, 0, 0, 0, 9, 9, 6, 6, 0, 0, 0, 12, 0, 0, 
    0, 0, 0, 0, 0, 5, 13, 7, 0, 0, 0, 0, 18, 0, 0, 
    0, 0, 0, 0, 0, 2, 6, 1, 0, 0, 0, 0, 14, 0, 0, 
    
    -- channel=152
    0, 0, 0, 0, 3, 0, 0, 3, 18, 0, 0, 14, 0, 0, 0, 
    0, 0, 0, 0, 28, 60, 65, 61, 77, 68, 21, 34, 6, 0, 34, 
    2, 4, 0, 0, 42, 0, 0, 0, 0, 48, 119, 17, 0, 0, 77, 
    2, 0, 0, 0, 106, 37, 0, 13, 1, 5, 24, 100, 0, 0, 13, 
    11, 0, 0, 0, 77, 53, 0, 25, 29, 33, 0, 97, 34, 0, 0, 
    52, 0, 0, 0, 84, 32, 0, 24, 28, 44, 42, 85, 107, 0, 4, 
    41, 0, 8, 0, 3, 14, 0, 0, 31, 14, 3, 91, 116, 92, 41, 
    0, 0, 87, 0, 2, 0, 4, 0, 31, 41, 9, 53, 114, 92, 155, 
    0, 0, 78, 0, 50, 20, 1, 0, 0, 0, 0, 0, 11, 0, 171, 
    0, 0, 64, 0, 61, 0, 60, 111, 3, 55, 20, 38, 42, 0, 204, 
    0, 0, 0, 0, 0, 52, 38, 0, 104, 0, 3, 47, 0, 29, 148, 
    0, 0, 71, 0, 0, 27, 100, 0, 145, 12, 4, 41, 0, 57, 206, 
    11, 0, 0, 0, 0, 0, 7, 23, 47, 133, 0, 0, 0, 50, 181, 
    17, 0, 0, 0, 0, 0, 0, 18, 46, 112, 74, 0, 0, 80, 159, 
    0, 0, 0, 0, 5, 0, 0, 6, 21, 35, 61, 0, 0, 63, 174, 
    
    -- channel=153
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 38, 72, 81, 108, 135, 122, 84, 35, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 29, 0, 0, 14, 41, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 50, 0, 0, 6, 
    0, 0, 55, 39, 7, 32, 44, 6, 7, 14, 0, 0, 0, 0, 0, 
    20, 2, 0, 0, 62, 11, 0, 33, 41, 21, 52, 41, 4, 0, 0, 
    7, 36, 39, 0, 0, 0, 0, 0, 0, 17, 28, 58, 105, 105, 8, 
    7, 61, 14, 0, 34, 0, 0, 12, 76, 77, 45, 91, 103, 52, 33, 
    0, 0, 0, 100, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 48, 
    0, 0, 64, 0, 52, 23, 56, 69, 56, 63, 74, 70, 60, 50, 38, 
    0, 0, 0, 0, 7, 35, 0, 0, 44, 0, 0, 0, 0, 0, 12, 
    5, 17, 40, 0, 0, 19, 107, 65, 58, 48, 0, 34, 59, 80, 58, 
    3, 0, 0, 0, 0, 0, 7, 8, 7, 0, 0, 0, 8, 8, 0, 
    0, 8, 0, 4, 0, 0, 0, 0, 0, 81, 83, 2, 7, 8, 21, 
    12, 0, 0, 19, 7, 0, 0, 0, 0, 9, 39, 17, 0, 5, 0, 
    
    -- channel=154
    159, 166, 146, 113, 114, 132, 150, 185, 189, 164, 160, 157, 151, 178, 136, 
    166, 168, 149, 53, 44, 42, 49, 44, 69, 110, 129, 162, 154, 143, 162, 
    158, 159, 127, 11, 11, 38, 34, 31, 26, 57, 139, 165, 150, 118, 159, 
    158, 148, 121, 0, 71, 80, 34, 9, 24, 45, 103, 137, 137, 150, 139, 
    157, 144, 69, 0, 34, 30, 0, 8, 25, 26, 36, 155, 170, 145, 179, 
    146, 125, 68, 0, 0, 0, 0, 0, 0, 1, 10, 65, 157, 158, 159, 
    136, 73, 69, 5, 41, 19, 0, 0, 17, 20, 17, 55, 89, 103, 152, 
    114, 25, 95, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 151, 
    127, 41, 118, 0, 16, 51, 37, 32, 106, 130, 92, 107, 121, 67, 144, 
    110, 9, 43, 0, 7, 0, 0, 36, 10, 17, 0, 3, 24, 0, 114, 
    114, 3, 49, 0, 0, 0, 36, 13, 1, 5, 0, 40, 7, 33, 121, 
    91, 0, 20, 54, 7, 3, 0, 0, 72, 25, 53, 77, 0, 0, 79, 
    61, 31, 93, 34, 0, 3, 0, 0, 16, 137, 126, 44, 0, 11, 107, 
    83, 46, 17, 24, 10, 0, 8, 19, 39, 49, 27, 0, 0, 33, 78, 
    43, 42, 29, 3, 5, 0, 15, 15, 16, 17, 21, 0, 1, 20, 98, 
    
    -- channel=155
    59, 48, 66, 93, 46, 37, 39, 21, 32, 66, 67, 54, 80, 39, 74, 
    69, 65, 91, 154, 48, 28, 36, 53, 42, 45, 58, 31, 66, 92, 27, 
    72, 69, 110, 189, 0, 14, 24, 39, 20, 0, 0, 39, 78, 94, 0, 
    72, 83, 85, 204, 0, 48, 111, 58, 58, 38, 23, 0, 78, 80, 47, 
    68, 89, 131, 156, 0, 28, 91, 44, 40, 47, 66, 0, 40, 97, 29, 
    40, 109, 121, 151, 0, 33, 46, 50, 53, 27, 46, 16, 0, 74, 70, 
    34, 125, 69, 111, 11, 36, 75, 46, 16, 50, 60, 0, 0, 37, 50, 
    83, 132, 0, 110, 64, 57, 23, 46, 45, 42, 33, 28, 0, 0, 0, 
    75, 139, 0, 144, 0, 26, 57, 75, 0, 0, 63, 0, 0, 42, 0, 
    95, 167, 2, 80, 0, 44, 0, 0, 77, 17, 59, 39, 34, 87, 0, 
    68, 195, 5, 46, 22, 0, 0, 67, 0, 51, 25, 0, 71, 0, 0, 
    73, 202, 0, 9, 77, 0, 0, 102, 0, 63, 32, 11, 144, 3, 0, 
    63, 126, 0, 40, 72, 39, 1, 0, 0, 0, 65, 135, 70, 0, 0, 
    37, 88, 97, 55, 34, 77, 0, 0, 0, 0, 17, 138, 51, 0, 0, 
    67, 62, 81, 73, 25, 47, 4, 0, 0, 0, 0, 87, 48, 0, 0, 
    
    -- channel=156
    165, 153, 175, 174, 129, 114, 117, 107, 126, 172, 170, 159, 185, 136, 164, 
    178, 175, 200, 207, 106, 92, 91, 116, 122, 136, 155, 137, 169, 197, 129, 
    183, 180, 212, 243, 38, 66, 75, 95, 73, 57, 66, 144, 181, 190, 88, 
    183, 194, 178, 261, 0, 101, 149, 110, 112, 87, 90, 102, 179, 180, 115, 
    176, 200, 193, 201, 25, 69, 139, 84, 89, 91, 137, 58, 141, 213, 138, 
    140, 211, 187, 176, 8, 70, 87, 78, 83, 70, 90, 77, 86, 184, 180, 
    120, 205, 129, 153, 32, 61, 110, 68, 46, 79, 86, 32, 67, 124, 162, 
    158, 175, 47, 160, 84, 86, 51, 76, 50, 46, 53, 34, 7, 45, 55, 
    160, 175, 26, 162, 24, 54, 80, 106, 33, 13, 115, 43, 0, 79, 6, 
    183, 208, 50, 103, 3, 74, 21, 10, 120, 73, 114, 92, 98, 120, 0, 
    156, 241, 36, 71, 33, 7, 15, 91, 6, 92, 68, 39, 95, 50, 0, 
    152, 243, 20, 55, 96, 5, 0, 129, 0, 100, 76, 58, 164, 24, 0, 
    130, 199, 25, 94, 110, 57, 8, 0, 0, 0, 119, 198, 76, 0, 0, 
    107, 151, 150, 105, 66, 103, 6, 0, 0, 0, 79, 209, 68, 0, 0, 
    126, 123, 142, 101, 54, 72, 21, 16, 13, 19, 28, 134, 58, 0, 0, 
    
    -- channel=157
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=158
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 43, 40, 38, 56, 73, 54, 24, 0, 0, 0, 0, 0, 
    0, 0, 0, 17, 0, 0, 0, 0, 0, 6, 0, 0, 0, 9, 0, 
    0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 3, 
    0, 0, 44, 36, 0, 16, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 31, 27, 0, 6, 22, 27, 9, 21, 15, 0, 0, 0, 
    3, 43, 40, 0, 0, 0, 7, 2, 0, 9, 28, 24, 47, 29, 0, 
    26, 85, 0, 13, 30, 23, 16, 40, 69, 60, 51, 72, 49, 27, 0, 
    0, 17, 3, 91, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 49, 37, 26, 26, 31, 44, 19, 52, 37, 55, 44, 29, 51, 0, 
    0, 19, 3, 10, 29, 14, 0, 34, 7, 8, 5, 0, 30, 0, 0, 
    3, 78, 0, 0, 11, 31, 75, 60, 18, 24, 0, 30, 71, 60, 0, 
    0, 0, 0, 2, 0, 9, 17, 13, 1, 0, 0, 0, 40, 0, 0, 
    0, 13, 11, 12, 8, 17, 0, 0, 0, 48, 33, 44, 26, 0, 0, 
    5, 0, 0, 33, 13, 12, 0, 0, 2, 11, 29, 25, 18, 0, 0, 
    
    -- channel=159
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 20, 40, 40, 48, 56, 58, 37, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 22, 25, 1, 5, 0, 0, 8, 6, 0, 0, 0, 
    0, 0, 19, 16, 6, 19, 18, 6, 11, 14, 0, 10, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 14, 7, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 19, 11, 27, 47, 27, 31, 38, 37, 1, 
    7, 7, 1, 5, 9, 0, 0, 0, 21, 6, 14, 40, 13, 13, 3, 
    0, 4, 11, 6, 5, 27, 17, 0, 0, 0, 0, 0, 0, 10, 17, 
    0, 1, 21, 3, 7, 2, 0, 35, 9, 2, 12, 3, 20, 3, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    10, 12, 0, 0, 0, 8, 32, 10, 42, 35, 0, 41, 32, 5, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 3, 0, 4, 
    2, 2, 0, 1, 1, 0, 0, 0, 14, 13, 9, 0, 0, 0, 3, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    
    
    others => 0);
end gold_package;
