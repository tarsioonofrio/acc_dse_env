library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 0, 291, 0, 0, 0, 459, 98, 382, 258, 0, 0, 0, 0, 29, 177, 0, 403, 0, 0, 183, 0, 3, 39, 489, 0, 17, 0, 374, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 313, 0, 249, 160, 168, 239, 0, 0, 0, 0, 0, 0, 0, 282, 90, 181, 287, 269, 67, 0, 80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 312, 0, 0, 355, 0, 281, 6, 207, 0, 178, 187, 458, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 130, 0, 117, 0, 0, 0, 0, 370, 303, 152, 237, 0, 136, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 78, 0, 203, 257, 0, 172, 0, 66, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 5, 0, 0, 0, 435, 54, 586, 206, 250, 199, 197, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 254, 330, 203, 279, 124, 11, 0, 0, 0, 157, 0, 54, 177, 79, 0, 0, 0, 0, 85, 31, 0, 0, 0, 0, 0, 319, 309, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 555, 494, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 350, 0, 0, 0, 0, 0, 0, 0, 155, 0, 0, 0, 0, 0, 0, 0, 0, 0, 304, 549, 0, 0, 80, 124, 23, 145, 0, 0, 0, 0, 68, 227, 0, 0, 0, 0, 0, 0, 589, 188, 347, 235, 0, 52, 80, 0, 0, 82, 97, 365, 471, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 171, 55, 0, 260, 2, 0, 140, 0, 59, 0, 0, 0, 0, 0, 287, 106, 159, 0, 0, 0, 347, 128, 196, 368, 249, 0, 0, 62, 168, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 111, 0, 0, 50, 0, 0, 0, 128, 85, 0, 0, 0, 0, 0, 0, 0, 11, 0, 162, 160, 0, 0, 0, 0, 0, 67, 0, 125, 105, 0, 68, 0, 0, 0, 134, 0, 258, 0, 0, 0, 0, 0, 244, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 167, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 112, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 89, 0, 25, 186, 0, 0, 0, 258, 477, 72, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 148, 101, 0, 0, 28, 20, 0, 0, 150, 0, 0, 0, 0, 0, 55, 103, 109, 172, 511, 273, 314, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 79, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 206, 211, 137, 335, 0, 0, 0, 0, 0, 0, 0, 0, 9, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 86, 131, 0, 236, 138, 259, 118, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 271, 263, 242, 448, 0, 0, 76, 0, 67, 0, 0, 0, 201, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 329, 0, 54, 0, 251, 255, 0, 0, 0, 0, 0, 0, 0, 0, 494, 0, 0, 0, 0, 0, 0, 0, 156, 210, 172, 141, 249, 93, 200, 0, 182, 109, 223, 0, 148, 235, 55, 0, 20, 94, 158, 258, 0, 0, 0, 0, 0, 0, 0, 0, 0, 81, 17, 16, 0, 0, 74, 0, 0, 0, 0, 0, 0, 22, 0, 200, 59, 269, 135, 26, 0, 0, 0, 0, 102, 456, 270, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 380, 35, 198, 156, 331, 132, 0, 0, 0, 0, 60, 217, 395, 295, 151, 0, 49, 27, 0, 0, 0, 0, 0, 0, 0, 11, 0, 30, 0, 148, 261, 43, 118, 16, 0, 0, 0, 0, 0, 155, 146, 67, 517, 0, 0, 316, 345, 154, 406, 44, 0, 411, 59, 319, 0, 65, 0, 0, 173, 0, 0, 44, 0, 0, 215, 0, 0, 0, 46, 0, 55, 110, 0, 0, 0, 42, 0, 0, 0, 181, 0, 321, 0, 214, 0, 0, 0, 0, 0, 51, 0, 0, 203, 82, 332, 0, 0, 0, 0, 254, 410, 483, 429, 436, 126, 0, 0, 0, 313, 312, 149, 326, 0, 0, 0, 0, 0, 0, 223, 0, 206, 98, 32, 0, 0, 0, 137, 127, 349, 589, 98, 0, 402, 0, 0, 0, 151, 27, 164, 178, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 503, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 94, 57, 0, 246, 0, 0, 0, 116, 115, 0, 0, 0, 0, 0, 0, 159, 0, 0, 0, 0, 130, 65, 55, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 278, 88, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 369, 310, 0, 0, 0, 97, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 111, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 92, 91, 451, 324, 191, 304, 0, 0, 0, 0, 0, 0, 0, 43, 0, 0, 0, 31, 0, 10, 0, 80, 68, 0, 0, 0, 0, 0, 276, 265, 0, 223, 122, 262, 148, 0, 262, 5, 0, 0, 129, 27, 132, 423, 60, 0, 6, 0, 0, 96, 0, 196, 484, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end ifmap_package;
