library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 4, 3, 0, 0, 0, 0, 0, 0, 0, 
    24, 13, 9, 0, 49, 33, 2, 0, 0, 0, 0, 9, 0, 2, 0, 
    0, 0, 13, 0, 0, 0, 11, 3, 1, 0, 7, 0, 0, 0, 2, 
    5, 0, 0, 0, 0, 0, 2, 5, 4, 0, 0, 0, 0, 0, 5, 
    4, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 9, 0, 3, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 68, 37, 11, 0, 11, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    4, 2, 0, 0, 0, 0, 0, 1, 0, 8, 15, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 23, 0, 0, 0, 14, 11, 0, 
    19, 27, 0, 0, 0, 42, 13, 17, 0, 0, 0, 0, 0, 19, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 11, 2, 2, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 12, 
    5, 0, 0, 13, 59, 18, 0, 0, 0, 0, 0, 7, 2, 0, 0, 
    0, 0, 25, 0, 16, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 11, 23, 3, 3, 0, 1, 6, 8, 1, 
    0, 0, 0, 0, 0, 41, 9, 0, 0, 0, 40, 28, 15, 0, 0, 
    2, 0, 0, 0, 5, 0, 0, 0, 0, 34, 19, 9, 0, 0, 1, 
    2, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 2, 2, 
    55, 17, 0, 0, 43, 53, 35, 33, 14, 0, 0, 0, 0, 0, 0, 
    0, 42, 5, 2, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 44, 29, 5, 0, 0, 0, 0, 0, 0, 8, 0, 0, 18, 
    0, 0, 1, 44, 11, 18, 16, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 26, 4, 7, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 17, 0, 0, 24, 3, 19, 0, 0, 0, 12, 0, 0, 0, 0, 
    0, 26, 0, 0, 3, 7, 27, 0, 0, 7, 4, 0, 0, 0, 0, 
    0, 18, 0, 0, 0, 29, 12, 0, 0, 7, 3, 0, 0, 0, 0, 
    15, 21, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 18, 7, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 
    22, 16, 8, 8, 22, 0, 14, 19, 0, 0, 0, 0, 0, 0, 0, 
    2, 11, 4, 42, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    3, 0, 1, 1, 3, 2, 0, 0, 3, 5, 6, 5, 4, 7, 8, 
    4, 1, 0, 0, 1, 0, 7, 1, 5, 13, 21, 24, 18, 9, 7, 
    4, 2, 1, 0, 1, 0, 3, 22, 25, 9, 7, 11, 22, 25, 5, 
    20, 25, 5, 1, 2, 10, 6, 19, 18, 7, 0, 12, 15, 29, 15, 
    8, 8, 6, 5, 0, 6, 0, 12, 17, 20, 4, 16, 16, 23, 33, 
    9, 0, 0, 4, 0, 0, 0, 11, 19, 7, 0, 10, 14, 18, 30, 
    11, 0, 5, 0, 0, 0, 0, 0, 10, 0, 0, 16, 21, 15, 18, 
    1, 0, 26, 6, 15, 0, 0, 0, 6, 0, 0, 14, 16, 7, 9, 
    0, 0, 11, 0, 13, 3, 7, 9, 14, 15, 3, 10, 19, 10, 7, 
    0, 0, 0, 9, 4, 16, 8, 0, 20, 0, 12, 28, 22, 7, 5, 
    0, 0, 0, 0, 0, 17, 0, 0, 3, 26, 35, 31, 29, 21, 24, 
    6, 0, 0, 0, 0, 8, 18, 18, 22, 25, 25, 24, 23, 24, 22, 
    30, 14, 0, 0, 2, 22, 23, 25, 27, 28, 27, 25, 20, 20, 21, 
    25, 29, 11, 0, 15, 23, 25, 26, 24, 23, 24, 21, 24, 23, 15, 
    23, 24, 26, 12, 27, 23, 18, 21, 22, 23, 25, 26, 21, 17, 27, 
    
    -- channel=7
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 1, 0, 1, 35, 0, 0, 0, 6, 0, 0, 3, 5, 0, 
    0, 15, 0, 0, 1, 16, 0, 0, 0, 45, 0, 0, 0, 3, 19, 
    0, 65, 0, 3, 0, 1, 0, 0, 0, 44, 0, 0, 0, 0, 44, 
    0, 55, 0, 20, 18, 0, 0, 0, 0, 47, 0, 0, 2, 0, 10, 
    0, 22, 0, 0, 57, 0, 0, 0, 0, 126, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 63, 31, 0, 0, 0, 115, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 23, 64, 0, 0, 0, 74, 0, 0, 11, 2, 0, 
    0, 1, 0, 30, 0, 0, 0, 1, 13, 0, 13, 0, 9, 19, 12, 
    0, 0, 0, 47, 0, 0, 7, 2, 0, 0, 0, 0, 36, 35, 0, 
    61, 0, 0, 109, 0, 0, 35, 0, 0, 0, 0, 9, 8, 6, 0, 
    46, 13, 0, 98, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 37, 24, 7, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 3, 
    0, 0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 24, 0, 0, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=9
    25, 26, 24, 26, 26, 23, 27, 31, 28, 22, 17, 16, 19, 25, 27, 
    25, 29, 27, 28, 24, 0, 25, 20, 23, 0, 0, 1, 5, 12, 22, 
    16, 10, 26, 29, 28, 25, 15, 13, 0, 0, 0, 0, 4, 5, 10, 
    16, 0, 24, 24, 19, 5, 0, 0, 0, 0, 0, 1, 1, 5, 2, 
    0, 0, 21, 0, 0, 0, 0, 0, 2, 0, 0, 3, 0, 4, 5, 
    0, 0, 16, 23, 0, 0, 0, 1, 7, 0, 0, 1, 0, 0, 0, 
    0, 0, 2, 31, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 9, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 13, 0, 9, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 1, 0, 2, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=12
    3, 0, 0, 0, 0, 0, 0, 0, 0, 7, 13, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 22, 0, 0, 0, 12, 4, 0, 
    23, 17, 0, 0, 0, 46, 11, 13, 0, 0, 0, 0, 0, 18, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 14, 1, 5, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 16, 
    7, 0, 0, 27, 49, 12, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 17, 0, 15, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 21, 25, 0, 6, 0, 4, 2, 11, 0, 
    0, 0, 0, 0, 0, 41, 4, 0, 0, 0, 35, 31, 15, 0, 0, 
    0, 0, 0, 0, 3, 2, 0, 0, 7, 32, 23, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 
    54, 6, 0, 0, 60, 48, 34, 31, 10, 0, 0, 0, 0, 0, 0, 
    0, 43, 0, 13, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 41, 31, 1, 0, 0, 0, 0, 0, 0, 8, 0, 0, 29, 
    0, 0, 7, 41, 14, 17, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 6, 0, 0, 
    19, 9, 0, 0, 0, 35, 4, 4, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 11, 0, 3, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 14, 
    7, 0, 0, 29, 37, 5, 0, 0, 0, 0, 2, 2, 0, 0, 0, 
    0, 4, 7, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 21, 20, 0, 5, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 27, 25, 11, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 9, 25, 19, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 
    51, 3, 0, 0, 62, 40, 30, 26, 7, 0, 0, 0, 0, 0, 0, 
    1, 42, 0, 21, 30, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 41, 30, 1, 0, 0, 0, 0, 0, 3, 10, 0, 0, 36, 
    0, 0, 13, 32, 15, 17, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    31, 34, 33, 32, 31, 33, 34, 34, 32, 29, 27, 28, 29, 30, 28, 
    29, 36, 34, 33, 31, 26, 33, 34, 29, 15, 11, 16, 21, 23, 27, 
    30, 23, 33, 34, 33, 31, 23, 19, 15, 7, 10, 6, 9, 15, 22, 
    14, 8, 30, 33, 31, 20, 17, 12, 6, 11, 12, 15, 8, 10, 17, 
    5, 7, 27, 25, 18, 24, 20, 14, 10, 7, 13, 14, 8, 6, 16, 
    11, 5, 27, 38, 20, 26, 16, 13, 8, 7, 16, 12, 8, 6, 9, 
    11, 9, 21, 32, 18, 16, 15, 12, 11, 5, 12, 10, 6, 6, 9, 
    14, 5, 12, 16, 17, 17, 15, 13, 10, 13, 10, 11, 8, 11, 14, 
    10, 7, 11, 6, 19, 15, 13, 10, 6, 16, 19, 12, 9, 12, 25, 
    7, 6, 6, 3, 15, 16, 8, 8, 14, 17, 9, 7, 7, 20, 26, 
    0, 10, 7, 1, 0, 9, 9, 8, 6, 2, 0, 0, 0, 0, 0, 
    0, 0, 4, 6, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    24, 23, 24, 27, 28, 21, 27, 29, 29, 24, 19, 15, 19, 26, 27, 
    27, 25, 23, 29, 21, 22, 40, 26, 21, 4, 21, 20, 10, 13, 24, 
    27, 0, 27, 29, 26, 2, 34, 16, 7, 0, 15, 9, 28, 6, 9, 
    51, 0, 31, 23, 34, 5, 21, 18, 12, 0, 30, 10, 19, 23, 0, 
    38, 1, 45, 0, 16, 20, 28, 26, 17, 0, 16, 36, 7, 25, 3, 
    27, 0, 48, 27, 0, 8, 33, 23, 38, 0, 35, 31, 0, 14, 22, 
    25, 27, 20, 42, 0, 0, 11, 26, 32, 0, 37, 28, 6, 0, 23, 
    25, 14, 29, 30, 0, 0, 32, 8, 21, 0, 25, 29, 0, 4, 17, 
    24, 0, 52, 0, 30, 0, 18, 17, 0, 30, 0, 23, 0, 2, 20, 
    3, 0, 49, 0, 25, 8, 0, 20, 19, 5, 22, 2, 0, 8, 28, 
    0, 4, 43, 0, 59, 26, 0, 0, 28, 19, 2, 0, 0, 0, 11, 
    0, 0, 11, 0, 48, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 15, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 22, 6, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=20
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 0, 0, 29, 20, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 7, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 5, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 2, 38, 19, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 56, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 20, 
    0, 0, 0, 23, 0, 0, 0, 0, 0, 85, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 139, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 70, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 1, 0, 0, 0, 0, 0, 12, 0, 0, 
    0, 0, 0, 100, 0, 0, 0, 0, 0, 0, 0, 11, 1, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 22, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 99, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 
    
    -- channel=23
    4, 7, 11, 12, 10, 10, 8, 8, 10, 0, 0, 0, 8, 10, 9, 
    12, 14, 12, 10, 15, 51, 17, 2, 0, 14, 29, 8, 0, 0, 11, 
    0, 0, 9, 10, 6, 0, 0, 0, 14, 27, 16, 23, 15, 0, 7, 
    28, 28, 11, 13, 11, 19, 35, 19, 11, 0, 12, 0, 2, 1, 0, 
    46, 50, 16, 32, 89, 50, 15, 14, 0, 18, 34, 23, 19, 23, 0, 
    4, 14, 17, 0, 0, 0, 36, 27, 23, 36, 7, 0, 7, 20, 28, 
    25, 3, 0, 11, 0, 29, 9, 24, 17, 15, 7, 15, 10, 24, 20, 
    23, 32, 23, 28, 19, 11, 0, 0, 7, 0, 4, 3, 5, 0, 10, 
    24, 18, 10, 20, 11, 0, 2, 17, 23, 0, 0, 0, 0, 15, 22, 
    6, 11, 20, 19, 13, 2, 24, 51, 2, 0, 0, 1, 23, 20, 6, 
    8, 14, 8, 58, 103, 66, 18, 0, 9, 15, 30, 41, 19, 0, 0, 
    0, 0, 36, 38, 0, 0, 0, 0, 0, 5, 8, 6, 14, 10, 10, 
    9, 0, 14, 0, 0, 12, 8, 7, 9, 14, 19, 22, 8, 6, 30, 
    9, 8, 0, 0, 3, 12, 17, 9, 9, 12, 4, 0, 6, 20, 0, 
    10, 9, 0, 0, 0, 0, 0, 11, 22, 24, 11, 11, 40, 27, 13, 
    
    -- channel=24
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=28
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 18, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 21, 0, 0, 
    59, 0, 0, 0, 0, 0, 21, 0, 0, 0, 17, 0, 9, 2, 0, 
    31, 6, 0, 0, 44, 0, 9, 9, 6, 0, 8, 14, 7, 30, 0, 
    0, 0, 0, 0, 0, 0, 38, 12, 54, 0, 0, 0, 0, 11, 13, 
    0, 31, 0, 24, 0, 0, 0, 4, 36, 0, 7, 10, 0, 0, 4, 
    0, 33, 0, 27, 0, 0, 0, 0, 6, 0, 0, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 18, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 43, 0, 0, 0, 0, 49, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 33, 0, 85, 10, 0, 0, 7, 22, 13, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 4, 0, 2, 
    9, 0, 0, 0, 0, 2, 3, 2, 5, 4, 6, 4, 0, 0, 5, 
    13, 0, 0, 46, 0, 0, 13, 1, 0, 0, 0, 0, 5, 0, 0, 
    15, 4, 0, 0, 0, 0, 0, 0, 3, 13, 7, 0, 0, 25, 30, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=30
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 20, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 46, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 29, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 49, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=32
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=33
    58, 59, 60, 61, 60, 58, 62, 65, 61, 51, 43, 44, 49, 52, 52, 
    60, 63, 63, 63, 63, 63, 57, 53, 38, 29, 23, 20, 25, 43, 51, 
    37, 46, 63, 63, 64, 48, 33, 20, 22, 27, 21, 18, 17, 22, 43, 
    20, 34, 58, 64, 52, 43, 36, 22, 16, 28, 21, 20, 11, 11, 34, 
    23, 38, 52, 64, 58, 44, 25, 16, 9, 27, 31, 22, 18, 14, 18, 
    16, 27, 50, 45, 27, 33, 32, 25, 12, 40, 25, 13, 18, 16, 15, 
    20, 18, 36, 46, 35, 41, 35, 26, 16, 34, 20, 15, 15, 21, 21, 
    24, 20, 26, 37, 44, 44, 17, 18, 19, 35, 24, 13, 17, 21, 32, 
    23, 22, 11, 27, 30, 18, 22, 21, 27, 26, 24, 5, 11, 32, 52, 
    25, 25, 12, 20, 22, 19, 27, 31, 18, 21, 6, 7, 23, 47, 50, 
    22, 26, 10, 39, 36, 30, 26, 14, 8, 3, 2, 5, 0, 3, 4, 
    0, 12, 26, 47, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 21, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=34
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=35
    3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 4, 23, 0, 0, 2, 0, 14, 0, 
    0, 0, 0, 0, 0, 16, 0, 22, 0, 7, 0, 0, 0, 1, 0, 
    18, 0, 18, 63, 0, 46, 0, 0, 0, 52, 0, 6, 0, 0, 29, 
    92, 0, 29, 38, 0, 57, 0, 0, 0, 12, 7, 19, 0, 0, 14, 
    119, 0, 22, 0, 0, 9, 0, 11, 0, 0, 1, 3, 2, 0, 2, 
    87, 0, 67, 0, 24, 0, 15, 0, 0, 0, 0, 0, 0, 0, 14, 
    33, 0, 50, 0, 46, 11, 0, 0, 11, 0, 0, 2, 2, 0, 0, 
    0, 0, 0, 0, 0, 71, 35, 0, 36, 0, 0, 3, 0, 0, 0, 
    0, 5, 0, 10, 0, 21, 1, 0, 9, 2, 2, 6, 4, 0, 3, 
    0, 0, 24, 0, 0, 25, 0, 0, 1, 2, 0, 0, 0, 0, 0, 
    3, 0, 74, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 
    0, 0, 55, 0, 16, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 1, 0, 0, 4, 0, 0, 0, 7, 5, 0, 0, 
    
    -- channel=36
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=37
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=38
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=39
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 35, 4, 0, 0, 0, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 7, 3, 0, 0, 
    8, 17, 0, 0, 0, 3, 18, 6, 0, 0, 0, 0, 0, 0, 0, 
    23, 35, 2, 14, 66, 43, 0, 1, 0, 5, 13, 9, 4, 9, 0, 
    0, 0, 1, 0, 0, 0, 15, 8, 9, 26, 0, 0, 0, 6, 16, 
    7, 0, 0, 0, 0, 12, 0, 10, 0, 6, 0, 0, 0, 7, 7, 
    7, 7, 8, 8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 4, 0, 0, 1, 5, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 4, 0, 0, 8, 29, 0, 0, 0, 0, 10, 12, 0, 
    0, 0, 0, 38, 80, 47, 12, 0, 0, 3, 12, 28, 6, 0, 0, 
    0, 0, 12, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 6, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 0, 0, 21, 11, 0, 
    
    -- channel=40
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=41
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=42
    63, 65, 65, 65, 64, 63, 70, 72, 63, 54, 51, 54, 57, 60, 56, 
    64, 70, 68, 67, 64, 54, 65, 60, 49, 27, 21, 27, 37, 50, 56, 
    47, 58, 67, 68, 66, 58, 40, 29, 20, 18, 17, 18, 21, 32, 51, 
    24, 32, 66, 66, 56, 40, 30, 19, 15, 24, 24, 22, 14, 17, 44, 
    14, 30, 62, 50, 42, 40, 31, 19, 16, 17, 25, 23, 17, 17, 29, 
    9, 23, 61, 42, 27, 35, 29, 25, 17, 14, 26, 19, 18, 15, 18, 
    9, 20, 49, 55, 34, 24, 31, 24, 21, 18, 21, 15, 14, 12, 22, 
    11, 18, 26, 43, 32, 29, 28, 23, 22, 27, 20, 16, 14, 24, 39, 
    9, 13, 9, 22, 25, 27, 24, 15, 23, 35, 20, 20, 17, 34, 53, 
    12, 12, 11, 11, 22, 23, 21, 21, 20, 26, 20, 12, 23, 50, 55, 
    8, 16, 14, 6, 13, 11, 12, 16, 13, 7, 0, 0, 0, 0, 0, 
    0, 4, 17, 19, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=43
    47, 49, 50, 50, 51, 45, 53, 61, 56, 40, 28, 30, 34, 40, 43, 
    50, 54, 54, 53, 51, 30, 39, 41, 29, 0, 0, 0, 5, 26, 37, 
    25, 36, 54, 57, 57, 45, 20, 6, 0, 0, 0, 0, 0, 0, 23, 
    0, 0, 43, 55, 40, 20, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 26, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 38, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 32, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=44
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 3, 4, 
    0, 0, 0, 1, 0, 0, 25, 3, 0, 0, 17, 12, 0, 0, 1, 
    11, 0, 0, 0, 0, 0, 30, 4, 0, 0, 14, 8, 29, 0, 0, 
    69, 0, 2, 0, 16, 0, 12, 21, 8, 0, 40, 0, 22, 24, 0, 
    63, 0, 37, 0, 8, 23, 35, 38, 16, 0, 9, 50, 0, 32, 0, 
    52, 0, 51, 12, 0, 4, 40, 25, 52, 0, 50, 48, 0, 16, 28, 
    57, 20, 3, 35, 0, 0, 0, 37, 42, 0, 55, 39, 0, 0, 26, 
    51, 13, 36, 22, 0, 0, 54, 0, 25, 0, 31, 39, 0, 0, 9, 
    45, 0, 94, 0, 39, 0, 12, 10, 0, 20, 0, 34, 0, 0, 0, 
    0, 0, 83, 0, 31, 11, 0, 15, 22, 0, 28, 0, 0, 0, 6, 
    0, 0, 68, 0, 100, 39, 0, 0, 50, 30, 1, 0, 0, 0, 7, 
    0, 0, 16, 0, 68, 36, 0, 0, 6, 0, 0, 0, 0, 0, 5, 
    21, 0, 0, 1, 78, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 31, 23, 0, 14, 0, 0, 0, 0, 0, 2, 0, 6, 
    29, 0, 0, 0, 6, 0, 0, 0, 0, 2, 10, 0, 0, 16, 39, 
    
    -- channel=45
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=46
    51, 51, 50, 51, 51, 47, 55, 60, 53, 47, 46, 46, 44, 47, 47, 
    50, 53, 51, 54, 49, 12, 50, 49, 51, 11, 0, 10, 25, 40, 45, 
    43, 51, 54, 55, 52, 47, 39, 27, 6, 0, 0, 0, 3, 21, 34, 
    13, 0, 51, 51, 42, 26, 0, 4, 0, 0, 8, 6, 7, 8, 21, 
    0, 0, 49, 27, 0, 0, 9, 5, 6, 0, 0, 7, 0, 3, 15, 
    2, 0, 50, 34, 0, 17, 0, 3, 1, 0, 8, 18, 0, 0, 0, 
    0, 0, 38, 51, 0, 0, 0, 4, 8, 0, 10, 1, 0, 0, 3, 
    0, 0, 6, 25, 5, 0, 25, 10, 12, 0, 3, 5, 0, 4, 26, 
    0, 0, 1, 0, 9, 18, 9, 0, 0, 16, 4, 30, 3, 7, 24, 
    0, 0, 0, 0, 4, 12, 0, 0, 0, 23, 27, 6, 0, 18, 44, 
    0, 0, 1, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=47
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    8, 0, 0, 0, 28, 14, 8, 0, 0, 0, 3, 0, 0, 0, 0, 
    4, 8, 4, 0, 0, 8, 18, 0, 0, 0, 15, 0, 0, 0, 0, 
    8, 13, 0, 0, 0, 0, 16, 6, 0, 0, 10, 0, 0, 0, 0, 
    15, 20, 0, 0, 0, 4, 16, 0, 0, 0, 1, 0, 0, 0, 0, 
    24, 17, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 14, 14, 0, 1, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    3, 15, 12, 0, 44, 8, 2, 14, 3, 0, 0, 0, 0, 0, 0, 
    0, 5, 14, 20, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 30, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=48
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 14, 0, 0, 25, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 33, 16, 29, 0, 0, 0, 0, 12, 24, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 
    
    -- channel=49
    0, 0, 3, 4, 5, 3, 3, 2, 3, 0, 0, 0, 0, 6, 4, 
    5, 6, 5, 5, 3, 26, 22, 1, 0, 0, 22, 13, 0, 0, 4, 
    0, 0, 4, 3, 3, 0, 0, 0, 4, 6, 10, 4, 19, 0, 0, 
    32, 17, 8, 3, 10, 0, 24, 16, 6, 0, 5, 0, 0, 5, 0, 
    24, 38, 21, 0, 52, 59, 13, 11, 0, 0, 18, 27, 6, 15, 4, 
    9, 0, 16, 8, 0, 0, 17, 16, 25, 0, 13, 0, 0, 8, 24, 
    16, 9, 0, 6, 0, 3, 0, 14, 8, 0, 1, 12, 4, 4, 17, 
    20, 2, 30, 15, 7, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    14, 0, 24, 0, 27, 0, 0, 9, 0, 20, 0, 0, 0, 0, 16, 
    0, 0, 12, 1, 5, 8, 0, 30, 21, 0, 0, 0, 7, 13, 2, 
    0, 1, 5, 2, 73, 61, 13, 0, 0, 14, 14, 27, 13, 0, 0, 
    0, 0, 5, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 6, 9, 3, 0, 7, 18, 2, 
    
    -- channel=50
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 4, 0, 0, 0, 13, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    26, 9, 0, 0, 0, 0, 14, 5, 0, 0, 0, 0, 0, 3, 0, 
    14, 26, 3, 0, 35, 30, 0, 5, 0, 0, 7, 17, 1, 13, 0, 
    0, 0, 1, 0, 0, 0, 9, 7, 24, 0, 0, 0, 0, 1, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 6, 0, 0, 11, 
    1, 0, 14, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 0, 10, 0, 0, 4, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 7, 0, 0, 0, 0, 21, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 66, 48, 0, 0, 0, 4, 13, 22, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 0, 0, 4, 13, 3, 
    
    -- channel=51
    27, 26, 27, 27, 27, 22, 29, 34, 30, 24, 21, 21, 21, 24, 27, 
    27, 27, 28, 28, 26, 0, 18, 21, 28, 0, 0, 0, 5, 19, 22, 
    18, 30, 28, 31, 30, 23, 16, 9, 0, 0, 0, 0, 0, 4, 14, 
    0, 0, 22, 27, 16, 7, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 13, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 8, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=52
    0, 2, 7, 6, 4, 5, 4, 2, 4, 0, 0, 0, 3, 1, 1, 
    6, 7, 7, 5, 9, 48, 7, 3, 0, 3, 11, 0, 0, 0, 4, 
    0, 0, 4, 4, 2, 0, 0, 0, 2, 16, 2, 5, 0, 0, 0, 
    0, 18, 1, 7, 8, 6, 22, 8, 0, 0, 0, 0, 0, 0, 0, 
    17, 35, 3, 24, 80, 41, 0, 3, 0, 7, 11, 6, 4, 3, 0, 
    0, 4, 5, 0, 0, 0, 22, 4, 1, 44, 0, 0, 0, 3, 9, 
    6, 0, 0, 2, 0, 30, 0, 12, 0, 15, 0, 0, 0, 8, 4, 
    15, 6, 2, 8, 6, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 4, 0, 8, 11, 0, 0, 4, 7, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 1, 9, 29, 0, 0, 0, 0, 11, 15, 0, 
    1, 2, 0, 55, 79, 51, 30, 0, 0, 0, 7, 27, 3, 0, 0, 
    0, 0, 14, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 17, 1, 0, 
    
    -- channel=53
    41, 44, 43, 43, 41, 40, 46, 52, 43, 30, 26, 29, 33, 37, 36, 
    41, 48, 46, 45, 43, 20, 31, 32, 26, 0, 0, 0, 8, 26, 31, 
    18, 36, 45, 48, 46, 39, 17, 6, 0, 0, 0, 0, 0, 3, 25, 
    0, 0, 38, 44, 26, 16, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    0, 0, 25, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 25, 31, 10, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 31, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 8, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=54
    17, 15, 17, 19, 20, 13, 18, 22, 23, 15, 10, 9, 12, 17, 19, 
    21, 16, 17, 19, 16, 12, 24, 15, 8, 0, 3, 3, 0, 8, 17, 
    10, 2, 20, 21, 19, 0, 18, 5, 1, 0, 0, 0, 4, 0, 4, 
    16, 0, 18, 19, 20, 6, 0, 2, 0, 0, 3, 0, 1, 6, 0, 
    9, 0, 25, 0, 0, 0, 0, 4, 0, 0, 0, 8, 0, 7, 0, 
    0, 0, 26, 9, 0, 0, 0, 0, 9, 0, 0, 8, 0, 0, 7, 
    3, 0, 5, 24, 0, 0, 0, 3, 2, 0, 2, 4, 0, 0, 2, 
    0, 0, 7, 11, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 7, 
    0, 0, 14, 0, 9, 0, 0, 0, 0, 4, 0, 4, 0, 0, 8, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 16, 
    0, 0, 0, 0, 15, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=55
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=56
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 0, 4, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 23, 12, 0, 0, 0, 0, 0, 0, 
    19, 2, 0, 0, 71, 27, 8, 7, 2, 0, 0, 2, 0, 3, 6, 
    14, 7, 0, 31, 41, 0, 2, 0, 0, 0, 0, 0, 11, 10, 0, 
    18, 4, 0, 56, 7, 0, 0, 0, 0, 1, 9, 13, 10, 2, 38, 
    21, 8, 6, 20, 7, 3, 9, 0, 0, 0, 8, 0, 0, 18, 21, 
    
    -- channel=58
    48, 49, 51, 50, 50, 46, 53, 57, 50, 35, 28, 33, 39, 43, 42, 
    51, 52, 53, 51, 51, 48, 45, 38, 23, 17, 6, 9, 18, 32, 40, 
    22, 37, 52, 54, 53, 36, 26, 15, 7, 6, 0, 4, 0, 11, 34, 
    3, 24, 48, 52, 41, 31, 14, 2, 0, 4, 8, 2, 0, 0, 24, 
    0, 11, 42, 42, 23, 17, 10, 4, 0, 13, 11, 3, 3, 0, 8, 
    0, 7, 41, 27, 12, 16, 15, 9, 0, 10, 4, 2, 1, 0, 1, 
    0, 0, 28, 36, 15, 19, 6, 10, 0, 5, 4, 1, 2, 2, 4, 
    0, 3, 7, 24, 16, 4, 4, 4, 7, 15, 7, 2, 0, 3, 27, 
    0, 0, 0, 8, 10, 8, 12, 4, 10, 17, 3, 0, 2, 23, 37, 
    3, 0, 0, 1, 0, 5, 14, 5, 1, 2, 0, 0, 2, 29, 35, 
    0, 1, 0, 10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=59
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 5, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 3, 0, 4, 0, 0, 15, 15, 0, 0, 0, 0, 1, 4, 0, 
    30, 15, 0, 21, 20, 0, 5, 3, 1, 6, 9, 10, 10, 11, 10, 
    14, 20, 3, 24, 0, 5, 7, 5, 5, 7, 10, 12, 16, 15, 13, 
    15, 11, 21, 25, 4, 8, 5, 6, 8, 10, 14, 16, 13, 17, 26, 
    15, 13, 10, 15, 7, 10, 13, 8, 8, 9, 10, 10, 13, 20, 10, 
    
    -- channel=60
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 4, 0, 0, 23, 7, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 7, 0, 0, 0, 0, 7, 0, 0, 0, 1, 0, 0, 0, 0, 
    3, 3, 0, 0, 0, 7, 12, 2, 0, 0, 0, 0, 0, 0, 0, 
    9, 10, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 9, 2, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    12, 7, 4, 0, 0, 0, 7, 21, 5, 0, 0, 0, 0, 0, 0, 
    24, 20, 1, 2, 37, 22, 12, 11, 5, 0, 1, 3, 3, 3, 5, 
    5, 17, 8, 25, 21, 2, 2, 1, 0, 0, 0, 1, 8, 9, 3, 
    9, 5, 19, 35, 4, 1, 0, 0, 2, 3, 7, 11, 7, 6, 23, 
    10, 8, 8, 13, 2, 6, 9, 3, 0, 0, 4, 2, 0, 7, 6, 
    
    -- channel=61
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 13, 0, 0, 0, 0, 13, 10, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 11, 15, 15, 15, 14, 15, 
    24, 6, 0, 0, 0, 10, 14, 10, 10, 14, 16, 20, 22, 19, 17, 
    22, 20, 6, 0, 0, 10, 11, 13, 14, 17, 19, 19, 17, 26, 30, 
    23, 22, 16, 0, 7, 11, 13, 11, 15, 14, 18, 12, 16, 27, 21, 
    
    -- channel=62
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 14, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 13, 1, 3, 5, 13, 10, 10, 
    48, 11, 0, 0, 26, 46, 37, 38, 37, 35, 38, 40, 38, 38, 41, 
    49, 40, 0, 0, 44, 34, 37, 35, 35, 36, 37, 36, 44, 47, 34, 
    56, 45, 30, 34, 34, 33, 32, 35, 39, 40, 47, 53, 50, 44, 67, 
    54, 51, 44, 47, 43, 47, 49, 38, 31, 31, 42, 42, 26, 39, 54, 
    
    -- channel=63
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 12, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 21, 0, 0, 0, 3, 0, 0, 
    21, 17, 0, 0, 0, 34, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 7, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 14, 34, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 12, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 23, 17, 0, 2, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 21, 23, 6, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 1, 34, 21, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 26, 6, 0, 0, 0, 0, 0, 0, 
    48, 6, 0, 0, 46, 23, 13, 11, 0, 0, 0, 0, 0, 0, 0, 
    0, 34, 0, 10, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 39, 27, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 25, 
    0, 0, 0, 23, 3, 9, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=64
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=65
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=66
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 4, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 31, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=67
    3, 8, 6, 3, 2, 7, 5, 5, 3, 0, 0, 10, 7, 0, 0, 
    6, 10, 8, 2, 9, 26, 0, 1, 0, 18, 0, 0, 8, 14, 2, 
    0, 33, 6, 5, 7, 30, 0, 0, 0, 37, 0, 0, 0, 3, 25, 
    0, 43, 0, 11, 0, 15, 0, 0, 0, 42, 0, 0, 0, 0, 46, 
    0, 19, 0, 33, 0, 0, 0, 0, 0, 51, 0, 0, 2, 0, 3, 
    0, 15, 0, 0, 77, 0, 0, 0, 0, 98, 0, 0, 10, 0, 0, 
    0, 0, 0, 0, 61, 30, 0, 0, 0, 89, 0, 0, 1, 9, 0, 
    0, 0, 0, 0, 19, 46, 0, 0, 0, 58, 0, 0, 14, 0, 0, 
    0, 1, 0, 32, 0, 9, 0, 0, 14, 0, 19, 0, 16, 22, 5, 
    0, 0, 0, 41, 0, 0, 20, 0, 0, 0, 0, 1, 25, 25, 0, 
    58, 0, 0, 86, 0, 0, 12, 0, 0, 0, 0, 0, 0, 3, 0, 
    38, 26, 0, 60, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 28, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 10, 0, 3, 0, 0, 0, 0, 0, 0, 12, 0, 0, 
    
    -- channel=68
    74, 76, 77, 77, 76, 72, 80, 84, 77, 64, 56, 60, 64, 68, 67, 
    76, 79, 79, 79, 77, 70, 69, 68, 52, 34, 20, 24, 37, 57, 65, 
    53, 64, 80, 81, 80, 62, 50, 30, 25, 18, 16, 15, 14, 30, 57, 
    19, 35, 74, 79, 67, 49, 33, 19, 15, 22, 25, 22, 16, 17, 42, 
    12, 24, 64, 61, 42, 30, 26, 21, 14, 22, 24, 20, 17, 14, 23, 
    9, 23, 65, 57, 38, 38, 33, 22, 13, 24, 24, 19, 17, 13, 14, 
    12, 13, 53, 63, 33, 38, 29, 25, 17, 17, 21, 16, 14, 16, 21, 
    16, 12, 19, 44, 34, 32, 22, 23, 26, 29, 26, 16, 15, 23, 43, 
    12, 10, 11, 24, 33, 24, 28, 21, 23, 28, 31, 18, 18, 38, 59, 
    21, 13, 11, 6, 20, 21, 23, 18, 17, 30, 14, 9, 19, 51, 61, 
    12, 16, 10, 17, 13, 7, 7, 8, 6, 0, 0, 0, 0, 0, 0, 
    0, 4, 14, 19, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=69
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=70
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=71
    1, 1, 2, 0, 0, 4, 0, 0, 0, 0, 0, 4, 1, 0, 0, 
    1, 4, 5, 0, 7, 11, 0, 0, 0, 12, 0, 0, 8, 10, 0, 
    0, 25, 1, 0, 4, 20, 0, 0, 6, 40, 0, 0, 0, 13, 14, 
    0, 52, 0, 7, 0, 15, 0, 0, 0, 56, 0, 0, 0, 0, 47, 
    0, 31, 0, 52, 0, 0, 0, 0, 0, 64, 0, 0, 0, 0, 19, 
    0, 12, 0, 0, 55, 0, 0, 0, 0, 116, 0, 0, 12, 0, 0, 
    0, 0, 0, 0, 58, 31, 0, 0, 0, 100, 0, 0, 4, 11, 0, 
    0, 0, 0, 0, 38, 55, 0, 0, 0, 63, 0, 0, 19, 2, 0, 
    0, 6, 0, 25, 0, 10, 0, 0, 22, 0, 15, 0, 15, 17, 8, 
    0, 4, 0, 48, 0, 0, 25, 0, 0, 0, 0, 0, 30, 26, 0, 
    48, 0, 0, 104, 0, 0, 33, 0, 0, 0, 5, 9, 14, 15, 0, 
    56, 26, 0, 77, 0, 0, 4, 2, 0, 2, 3, 6, 4, 4, 0, 
    0, 48, 53, 0, 0, 0, 0, 0, 0, 3, 7, 6, 1, 4, 9, 
    0, 3, 86, 0, 0, 5, 0, 0, 4, 4, 2, 3, 0, 18, 0, 
    0, 2, 5, 3, 0, 11, 4, 0, 6, 0, 0, 4, 28, 0, 0, 
    
    -- channel=72
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 1, 0, 0, 2, 40, 0, 0, 0, 6, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 17, 0, 7, 0, 0, 0, 
    1, 24, 0, 1, 0, 7, 17, 3, 0, 0, 0, 0, 0, 0, 0, 
    17, 31, 0, 20, 62, 21, 0, 0, 0, 16, 12, 2, 7, 8, 0, 
    0, 0, 0, 0, 0, 0, 14, 6, 4, 41, 0, 0, 0, 5, 15, 
    0, 0, 0, 0, 0, 20, 0, 3, 0, 9, 0, 0, 0, 13, 4, 
    0, 6, 0, 7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 4, 12, 0, 0, 0, 0, 7, 8, 
    0, 0, 0, 6, 0, 0, 13, 27, 0, 0, 0, 0, 16, 11, 0, 
    0, 0, 0, 55, 66, 38, 1, 0, 0, 0, 19, 30, 4, 0, 0, 
    0, 0, 10, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 2, 6, 7, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 0, 0, 27, 3, 0, 
    
    -- channel=73
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 8, 30, 14, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 40, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 16, 0, 28, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 65, 17, 6, 0, 4, 19, 0, 0, 0, 
    0, 0, 33, 0, 0, 31, 0, 0, 0, 0, 0, 88, 0, 0, 0, 
    0, 0, 34, 0, 0, 0, 0, 0, 0, 25, 76, 0, 0, 0, 0, 
    0, 0, 48, 0, 0, 0, 0, 5, 30, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 157, 120, 38, 35, 11, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 149, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 106, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 
    3, 0, 0, 54, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    
    -- channel=74
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 0, 2, 4, 
    0, 0, 0, 1, 0, 0, 17, 3, 13, 0, 8, 6, 0, 0, 1, 
    13, 0, 0, 0, 0, 0, 26, 13, 0, 0, 11, 6, 25, 0, 0, 
    68, 0, 1, 0, 10, 0, 9, 10, 1, 0, 32, 0, 21, 13, 0, 
    56, 0, 24, 0, 4, 0, 33, 24, 15, 0, 9, 35, 0, 26, 0, 
    28, 0, 31, 0, 0, 0, 31, 24, 44, 0, 36, 40, 0, 13, 11, 
    22, 25, 2, 39, 0, 0, 15, 22, 49, 0, 50, 27, 0, 0, 14, 
    13, 27, 11, 25, 0, 0, 48, 4, 25, 0, 25, 34, 0, 0, 5, 
    22, 0, 54, 0, 3, 0, 17, 5, 0, 18, 0, 38, 0, 0, 0, 
    0, 0, 70, 0, 33, 0, 0, 20, 0, 4, 36, 2, 0, 0, 6, 
    0, 0, 65, 0, 60, 14, 0, 12, 44, 23, 0, 0, 0, 0, 8, 
    0, 0, 16, 0, 79, 37, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 9, 80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 62, 17, 0, 5, 0, 0, 0, 0, 0, 0, 0, 8, 
    18, 0, 0, 10, 5, 0, 0, 0, 0, 0, 4, 0, 0, 8, 34, 
    
    -- channel=75
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 7, 10, 8, 8, 
    13, 0, 0, 0, 0, 5, 3, 4, 5, 9, 13, 13, 7, 9, 17, 
    16, 13, 0, 0, 0, 6, 7, 4, 7, 9, 10, 9, 14, 19, 2, 
    14, 17, 6, 0, 0, 2, 2, 6, 8, 11, 8, 12, 18, 12, 15, 
    
    -- channel=76
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=77
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=78
    15, 14, 13, 14, 16, 11, 17, 22, 20, 18, 16, 12, 10, 13, 15, 
    15, 15, 14, 17, 11, 0, 21, 20, 24, 0, 0, 0, 1, 6, 11, 
    21, 8, 17, 18, 17, 8, 20, 8, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 15, 15, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=79
    23, 24, 26, 26, 26, 23, 27, 28, 26, 17, 11, 13, 18, 21, 22, 
    26, 27, 27, 27, 27, 33, 21, 19, 4, 3, 0, 0, 1, 13, 21, 
    10, 13, 27, 27, 27, 8, 2, 0, 0, 1, 0, 0, 0, 0, 15, 
    0, 14, 24, 27, 22, 10, 9, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 10, 17, 17, 22, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 8, 0, 0, 2, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 0, 5, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 4, 3, 0, 0, 0, 3, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 6, 22, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 17, 15, 
    0, 0, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=80
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=81
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=82
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=83
    19, 19, 21, 22, 22, 19, 23, 25, 23, 15, 8, 9, 13, 19, 19, 
    23, 24, 23, 23, 21, 24, 23, 18, 3, 0, 0, 0, 0, 7, 18, 
    11, 2, 23, 24, 23, 3, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    5, 8, 21, 23, 21, 2, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 18, 4, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 8, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=84
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=85
    2, 0, 0, 0, 0, 0, 0, 0, 0, 5, 14, 13, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 21, 0, 0, 0, 19, 15, 0, 
    14, 36, 0, 0, 0, 31, 12, 17, 0, 0, 0, 0, 0, 22, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 6, 0, 0, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 0, 0, 0, 0, 16, 
    0, 0, 0, 5, 56, 16, 0, 0, 0, 0, 0, 2, 2, 0, 0, 
    0, 0, 30, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 5, 20, 0, 2, 0, 0, 5, 7, 0, 
    0, 0, 0, 0, 0, 40, 6, 0, 0, 0, 29, 23, 18, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 28, 17, 9, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 13, 10, 
    55, 25, 0, 0, 24, 50, 34, 33, 13, 2, 0, 0, 0, 0, 0, 
    0, 44, 19, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 50, 22, 2, 0, 0, 0, 0, 0, 0, 6, 0, 0, 15, 
    0, 0, 5, 39, 9, 16, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=86
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 8, 13, 16, 14, 0, 0, 
    14, 0, 0, 0, 0, 0, 1, 11, 13, 1, 9, 7, 14, 15, 0, 
    21, 8, 0, 0, 2, 3, 8, 13, 14, 6, 7, 13, 13, 19, 4, 
    12, 7, 0, 0, 0, 0, 7, 11, 19, 0, 4, 12, 11, 16, 21, 
    15, 10, 0, 0, 0, 0, 0, 8, 16, 0, 9, 14, 13, 12, 13, 
    12, 16, 8, 0, 0, 0, 6, 3, 11, 0, 6, 12, 12, 8, 1, 
    13, 11, 17, 8, 0, 1, 5, 6, 9, 0, 0, 12, 12, 4, 0, 
    5, 8, 20, 13, 11, 7, 7, 13, 8, 0, 14, 19, 16, 0, 0, 
    5, 6, 18, 5, 24, 18, 9, 11, 22, 21, 27, 31, 26, 12, 10, 
    18, 13, 16, 0, 3, 23, 25, 26, 32, 32, 36, 37, 40, 38, 39, 
    44, 20, 9, 0, 25, 37, 38, 37, 37, 38, 41, 41, 39, 39, 43, 
    47, 43, 12, 14, 29, 37, 39, 38, 39, 40, 41, 40, 43, 42, 40, 
    47, 47, 37, 27, 32, 33, 35, 38, 39, 40, 41, 42, 41, 44, 50, 
    
    -- channel=87
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 17, 14, 5, 3, 
    13, 0, 0, 0, 0, 1, 4, 6, 17, 20, 25, 24, 27, 25, 26, 
    35, 12, 0, 0, 0, 21, 22, 21, 22, 26, 29, 29, 28, 28, 32, 
    37, 32, 9, 0, 13, 21, 22, 22, 24, 26, 28, 30, 31, 36, 31, 
    34, 34, 27, 8, 19, 23, 23, 23, 23, 24, 26, 28, 29, 29, 35, 
    
    -- channel=88
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 77, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=89
    17, 13, 17, 19, 20, 13, 18, 20, 21, 16, 10, 8, 12, 18, 21, 
    20, 15, 16, 19, 16, 12, 28, 14, 8, 2, 14, 12, 4, 6, 18, 
    14, 0, 18, 19, 19, 0, 15, 9, 8, 0, 7, 7, 18, 4, 3, 
    33, 0, 19, 16, 21, 7, 14, 17, 9, 0, 13, 3, 10, 16, 0, 
    24, 0, 29, 0, 8, 18, 10, 16, 9, 0, 7, 24, 6, 19, 7, 
    15, 0, 28, 15, 0, 0, 8, 15, 25, 0, 14, 16, 0, 12, 19, 
    17, 0, 3, 26, 0, 0, 0, 13, 18, 0, 13, 17, 5, 1, 17, 
    10, 0, 22, 18, 0, 0, 11, 0, 8, 0, 5, 15, 0, 0, 12, 
    4, 0, 29, 0, 22, 0, 4, 8, 0, 16, 0, 10, 0, 0, 14, 
    0, 0, 21, 0, 9, 10, 0, 8, 14, 0, 10, 3, 0, 5, 17, 
    0, 0, 16, 0, 33, 23, 0, 0, 11, 16, 8, 6, 0, 0, 3, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    
    -- channel=90
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=91
    9, 11, 10, 11, 10, 10, 12, 13, 11, 10, 10, 7, 10, 14, 12, 
    10, 13, 10, 12, 7, 0, 23, 12, 16, 0, 9, 10, 4, 5, 9, 
    12, 0, 10, 13, 8, 0, 21, 13, 3, 0, 9, 7, 18, 2, 1, 
    36, 0, 13, 8, 12, 0, 8, 11, 4, 0, 19, 7, 13, 15, 0, 
    34, 0, 25, 0, 5, 13, 23, 17, 10, 0, 10, 26, 1, 18, 0, 
    22, 0, 31, 4, 0, 16, 21, 19, 23, 0, 22, 26, 0, 10, 16, 
    24, 11, 16, 26, 0, 0, 7, 15, 27, 0, 29, 18, 0, 0, 14, 
    18, 12, 21, 16, 0, 0, 23, 6, 17, 0, 16, 21, 0, 0, 12, 
    15, 0, 34, 0, 8, 4, 15, 2, 0, 14, 0, 22, 0, 0, 6, 
    0, 0, 36, 0, 23, 3, 0, 9, 8, 5, 20, 7, 0, 0, 14, 
    0, 0, 33, 0, 34, 14, 0, 2, 26, 13, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 33, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    
    -- channel=92
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 21, 2, 0, 0, 0, 0, 0, 0, 
    1, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 13, 6, 0, 17, 4, 0, 1, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 20, 19, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=93
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 
    0, 0, 0, 0, 0, 33, 0, 13, 0, 0, 0, 0, 0, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 0, 20, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 40, 0, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 0, 0, 0, 0, 19, 34, 32, 0, 0, 0, 0, 0, 0, 0, 
    0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 33, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=94
    50, 52, 53, 53, 53, 49, 55, 59, 54, 42, 35, 38, 42, 44, 45, 
    52, 55, 55, 55, 54, 53, 47, 45, 31, 19, 8, 9, 18, 35, 43, 
    31, 42, 55, 56, 55, 42, 28, 13, 8, 9, 2, 4, 2, 10, 36, 
    7, 20, 50, 56, 46, 33, 20, 5, 2, 7, 11, 4, 2, 0, 24, 
    2, 13, 42, 45, 35, 19, 12, 5, 0, 8, 12, 5, 5, 2, 5, 
    0, 8, 40, 31, 15, 16, 18, 10, 2, 12, 8, 3, 3, 2, 1, 
    0, 1, 26, 43, 19, 21, 15, 12, 4, 9, 5, 1, 0, 3, 5, 
    0, 5, 3, 29, 19, 17, 8, 6, 8, 16, 9, 1, 0, 6, 23, 
    0, 0, 0, 10, 12, 6, 10, 7, 9, 16, 7, 2, 1, 20, 38, 
    6, 0, 0, 0, 1, 6, 12, 10, 0, 11, 1, 0, 4, 33, 40, 
    2, 3, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=95
    0, 2, 0, 4, 4, 0, 0, 3, 7, 6, 4, 0, 1, 4, 8, 
    2, 0, 0, 5, 0, 0, 19, 8, 13, 0, 12, 5, 0, 0, 4, 
    15, 0, 0, 5, 0, 0, 31, 13, 0, 0, 9, 6, 21, 0, 0, 
    62, 0, 1, 0, 17, 0, 11, 13, 2, 0, 31, 0, 20, 13, 0, 
    56, 0, 22, 0, 10, 2, 29, 26, 11, 0, 9, 34, 0, 25, 0, 
    31, 0, 31, 0, 0, 5, 33, 23, 39, 0, 33, 39, 0, 13, 13, 
    31, 14, 1, 39, 0, 0, 7, 23, 42, 0, 45, 27, 0, 0, 13, 
    24, 19, 14, 21, 0, 0, 39, 0, 23, 0, 27, 31, 0, 0, 5, 
    27, 0, 57, 0, 12, 0, 16, 8, 0, 11, 0, 32, 0, 0, 0, 
    1, 0, 65, 0, 28, 0, 0, 16, 0, 2, 29, 1, 0, 0, 10, 
    0, 0, 57, 0, 67, 18, 0, 3, 41, 22, 0, 0, 0, 0, 6, 
    0, 0, 15, 0, 62, 33, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 74, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 42, 18, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 24, 
    
    -- channel=96
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=97
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=98
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 28, 23, 0, 0, 0, 0, 15, 21, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 3, 1, 
    10, 0, 0, 0, 0, 0, 0, 0, 2, 8, 11, 13, 0, 0, 15, 
    6, 5, 0, 0, 0, 1, 7, 2, 0, 3, 0, 0, 0, 13, 0, 
    7, 6, 0, 0, 0, 0, 0, 0, 8, 14, 7, 5, 22, 19, 9, 
    
    -- channel=99
    43, 42, 44, 45, 45, 40, 46, 50, 45, 35, 28, 31, 35, 38, 39, 
    46, 45, 46, 46, 45, 43, 38, 36, 22, 16, 8, 10, 16, 32, 38, 
    25, 34, 47, 47, 48, 29, 21, 9, 11, 10, 3, 3, 4, 15, 32, 
    3, 28, 44, 46, 38, 26, 17, 7, 6, 10, 6, 7, 3, 6, 24, 
    0, 16, 35, 34, 20, 12, 3, 5, 3, 14, 8, 5, 7, 4, 13, 
    0, 7, 33, 32, 6, 6, 10, 6, 3, 22, 2, 0, 6, 3, 5, 
    0, 0, 23, 32, 16, 20, 6, 7, 0, 14, 0, 3, 5, 8, 9, 
    0, 0, 5, 23, 20, 13, 0, 3, 7, 18, 6, 1, 5, 9, 21, 
    0, 0, 0, 9, 17, 2, 8, 10, 10, 14, 11, 0, 7, 20, 35, 
    1, 0, 0, 0, 0, 6, 8, 7, 5, 7, 0, 0, 10, 33, 34, 
    3, 0, 0, 13, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=100
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 21, 24, 5, 5, 7, 1, 2, 2, 0, 1, 4, 
    13, 0, 0, 0, 30, 0, 2, 1, 2, 0, 0, 0, 5, 7, 0, 
    16, 7, 0, 17, 7, 0, 1, 0, 1, 1, 6, 9, 10, 0, 22, 
    15, 7, 7, 11, 9, 5, 8, 3, 0, 0, 5, 3, 0, 1, 21, 
    
    -- channel=101
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=102
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=103
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=104
    24, 22, 24, 26, 29, 19, 26, 35, 34, 24, 14, 12, 13, 18, 25, 
    29, 26, 27, 29, 27, 0, 18, 22, 14, 0, 0, 0, 0, 11, 21, 
    13, 19, 29, 31, 32, 10, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 23, 30, 21, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=105
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 14, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 53, 24, 11, 8, 0, 0, 0, 0, 6, 1, 0, 0, 
    1, 4, 2, 41, 0, 0, 0, 0, 0, 0, 2, 5, 12, 12, 8, 
    11, 1, 21, 0, 0, 3, 1, 0, 1, 7, 15, 19, 11, 11, 29, 
    12, 12, 16, 0, 0, 8, 5, 3, 5, 10, 9, 9, 10, 28, 0, 
    8, 15, 5, 0, 0, 0, 0, 3, 13, 16, 8, 12, 38, 25, 5, 
    
    -- channel=106
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 7, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 3, 0, 
    3, 8, 0, 0, 0, 7, 0, 0, 0, 5, 0, 0, 3, 0, 0, 
    9, 17, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 15, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 9, 0, 35, 4, 4, 20, 13, 2, 1, 16, 24, 26, 14, 6, 
    48, 29, 5, 26, 3, 22, 31, 32, 33, 35, 42, 45, 49, 49, 48, 
    54, 45, 28, 15, 13, 41, 40, 39, 41, 45, 51, 53, 51, 52, 59, 
    58, 52, 48, 22, 30, 44, 41, 41, 44, 48, 53, 55, 55, 66, 56, 
    56, 58, 48, 36, 36, 45, 45, 43, 45, 49, 48, 51, 60, 59, 50, 
    
    -- channel=107
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=108
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    
    -- channel=109
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=110
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 55, 11, 0, 0, 0, 0, 0, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 5, 2, 3, 
    13, 0, 0, 0, 0, 1, 0, 0, 0, 4, 9, 12, 4, 2, 18, 
    15, 6, 0, 0, 0, 0, 7, 0, 0, 4, 2, 0, 7, 13, 0, 
    16, 10, 0, 0, 0, 0, 0, 2, 9, 12, 5, 3, 17, 24, 20, 
    
    -- channel=111
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=112
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=113
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 4, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 6, 9, 15, 15, 12, 8, 3, 
    11, 5, 0, 0, 0, 0, 2, 9, 16, 7, 11, 11, 17, 20, 5, 
    15, 15, 0, 0, 0, 1, 7, 15, 17, 11, 4, 12, 13, 23, 11, 
    10, 12, 1, 0, 0, 0, 0, 10, 16, 8, 3, 12, 14, 19, 20, 
    9, 6, 0, 0, 0, 0, 0, 7, 15, 10, 2, 10, 15, 15, 19, 
    5, 5, 8, 0, 0, 0, 2, 3, 13, 6, 3, 12, 14, 14, 16, 
    3, 0, 15, 8, 6, 6, 0, 5, 10, 0, 1, 11, 15, 12, 4, 
    0, 1, 11, 9, 10, 1, 5, 10, 14, 1, 13, 11, 14, 6, 2, 
    0, 0, 8, 5, 17, 10, 2, 5, 14, 13, 15, 22, 22, 6, 3, 
    6, 0, 5, 1, 0, 21, 15, 8, 19, 18, 28, 30, 30, 29, 30, 
    29, 8, 6, 0, 3, 18, 19, 20, 28, 31, 32, 30, 29, 30, 31, 
    37, 27, 6, 0, 12, 27, 28, 28, 30, 32, 32, 32, 32, 31, 30, 
    36, 34, 24, 8, 26, 27, 28, 30, 29, 30, 31, 33, 32, 35, 35, 
    33, 33, 30, 25, 32, 32, 31, 29, 27, 26, 31, 30, 27, 29, 36, 
    
    -- channel=114
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 7, 0, 0, 0, 0, 0, 0, 2, 0, 3, 0, 0, 0, 0, 
    7, 17, 0, 0, 0, 0, 1, 0, 1, 0, 3, 0, 0, 0, 0, 
    12, 16, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 18, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 15, 18, 8, 3, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    16, 11, 15, 8, 26, 14, 18, 19, 15, 7, 14, 23, 25, 15, 13, 
    34, 22, 10, 14, 29, 28, 29, 29, 33, 34, 40, 42, 46, 47, 47, 
    55, 32, 12, 26, 28, 39, 39, 37, 38, 42, 46, 49, 49, 49, 53, 
    59, 50, 26, 37, 33, 39, 41, 39, 41, 45, 50, 52, 52, 59, 59, 
    59, 55, 46, 32, 36, 39, 40, 40, 42, 46, 48, 46, 50, 62, 56, 
    
    -- channel=115
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 0, 0, 11, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 8, 0, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 27, 0, 0, 0, 0, 0, 
    5, 11, 0, 0, 0, 10, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    12, 19, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 14, 0, 21, 0, 0, 1, 7, 0, 0, 0, 0, 0, 0, 0, 
    24, 11, 0, 53, 30, 17, 24, 2, 0, 0, 8, 21, 19, 4, 0, 
    24, 22, 9, 46, 0, 0, 5, 6, 11, 17, 24, 28, 34, 33, 30, 
    35, 23, 30, 11, 0, 25, 23, 22, 22, 28, 36, 40, 34, 35, 49, 
    37, 35, 34, 0, 10, 29, 26, 24, 27, 32, 34, 33, 35, 51, 29, 
    35, 39, 29, 5, 11, 20, 21, 26, 34, 37, 30, 34, 55, 48, 29, 
    
    -- channel=116
    46, 48, 47, 47, 46, 44, 51, 54, 47, 38, 33, 35, 36, 39, 37, 
    45, 48, 49, 50, 46, 35, 42, 43, 31, 6, 0, 2, 17, 29, 35, 
    37, 40, 50, 51, 52, 50, 31, 8, 0, 0, 0, 0, 0, 8, 28, 
    0, 4, 45, 47, 42, 18, 5, 0, 0, 4, 10, 5, 0, 0, 15, 
    0, 0, 40, 23, 8, 10, 13, 2, 0, 0, 1, 0, 0, 0, 4, 
    3, 12, 43, 47, 33, 27, 14, 0, 0, 0, 19, 5, 0, 0, 0, 
    0, 10, 32, 36, 15, 16, 20, 9, 0, 0, 11, 0, 0, 0, 0, 
    6, 0, 0, 16, 5, 19, 27, 15, 6, 16, 13, 1, 0, 8, 18, 
    6, 3, 4, 1, 16, 17, 9, 0, 0, 15, 14, 9, 0, 10, 30, 
    16, 8, 0, 0, 2, 8, 0, 0, 7, 18, 3, 0, 0, 23, 36, 
    1, 10, 3, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 10, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=117
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=118
    0, 0, 2, 3, 4, 1, 0, 0, 5, 0, 0, 0, 0, 2, 4, 
    5, 4, 2, 1, 4, 42, 11, 0, 0, 11, 27, 12, 0, 0, 2, 
    0, 0, 2, 3, 1, 0, 0, 0, 12, 17, 5, 9, 10, 0, 0, 
    26, 25, 3, 5, 9, 12, 27, 9, 4, 0, 3, 0, 0, 1, 0, 
    26, 32, 6, 12, 54, 32, 6, 10, 0, 11, 24, 16, 12, 15, 0, 
    0, 0, 2, 0, 0, 0, 25, 18, 22, 21, 0, 0, 0, 11, 22, 
    13, 0, 0, 6, 0, 19, 0, 12, 6, 2, 0, 13, 9, 16, 10, 
    13, 15, 15, 17, 6, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    12, 2, 10, 3, 13, 0, 0, 19, 6, 10, 0, 0, 0, 5, 13, 
    0, 0, 12, 15, 0, 0, 12, 37, 1, 0, 0, 0, 6, 8, 0, 
    0, 2, 2, 37, 77, 47, 0, 0, 0, 14, 28, 31, 13, 0, 2, 
    0, 0, 8, 20, 0, 0, 0, 0, 0, 1, 2, 2, 9, 6, 5, 
    6, 0, 0, 0, 0, 5, 2, 3, 6, 10, 13, 15, 0, 0, 20, 
    3, 4, 0, 0, 0, 6, 13, 5, 2, 5, 1, 0, 2, 14, 0, 
    4, 3, 0, 0, 0, 0, 0, 0, 13, 19, 7, 6, 28, 20, 5, 
    
    -- channel=119
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=120
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=121
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 32, 10, 0, 0, 0, 30, 14, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 13, 0, 0, 0, 10, 10, 32, 0, 0, 
    78, 0, 0, 0, 17, 0, 31, 8, 7, 0, 34, 0, 16, 12, 0, 
    56, 11, 14, 0, 61, 12, 31, 27, 12, 0, 20, 36, 10, 37, 0, 
    0, 0, 19, 0, 0, 0, 56, 26, 65, 0, 24, 22, 0, 18, 26, 
    0, 42, 0, 36, 0, 0, 8, 27, 47, 0, 33, 28, 0, 0, 18, 
    0, 41, 3, 39, 0, 0, 18, 0, 17, 0, 17, 26, 0, 0, 0, 
    19, 0, 43, 0, 4, 0, 5, 23, 0, 20, 0, 9, 0, 0, 0, 
    0, 0, 71, 0, 17, 0, 0, 54, 0, 0, 16, 0, 0, 0, 0, 
    0, 0, 58, 0, 122, 38, 0, 0, 33, 33, 16, 17, 2, 0, 11, 
    0, 0, 9, 0, 28, 0, 0, 0, 0, 0, 0, 0, 2, 0, 4, 
    16, 0, 0, 13, 25, 4, 4, 2, 3, 2, 3, 3, 0, 0, 5, 
    17, 2, 0, 51, 9, 0, 17, 2, 0, 0, 0, 0, 3, 0, 0, 
    22, 1, 0, 0, 0, 0, 0, 0, 2, 13, 9, 0, 0, 28, 36, 
    
    -- channel=122
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 9, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 5, 4, 22, 0, 0, 
    62, 0, 0, 0, 5, 0, 12, 0, 0, 0, 29, 0, 16, 9, 0, 
    49, 0, 17, 0, 21, 0, 25, 18, 9, 0, 9, 28, 0, 27, 0, 
    0, 0, 25, 0, 0, 0, 39, 20, 47, 0, 22, 27, 0, 10, 12, 
    0, 30, 0, 34, 0, 0, 9, 18, 44, 0, 38, 20, 0, 0, 12, 
    0, 32, 0, 29, 0, 0, 25, 0, 20, 0, 18, 25, 0, 0, 2, 
    9, 0, 38, 0, 0, 0, 10, 7, 0, 12, 0, 21, 0, 0, 0, 
    0, 0, 65, 0, 21, 0, 0, 31, 0, 0, 23, 0, 0, 0, 0, 
    0, 0, 57, 0, 80, 12, 0, 0, 34, 19, 0, 0, 0, 0, 0, 
    0, 0, 11, 0, 49, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 3, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 59, 7, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 32, 
    
    -- channel=123
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 2, 7, 13, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 18, 2, 0, 0, 0, 0, 0, 0, 
    2, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 12, 8, 0, 0, 0, 7, 
    0, 0, 0, 15, 0, 0, 0, 0, 7, 1, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 11, 3, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 7, 0, 13, 0, 0, 0, 
    0, 0, 0, 0, 4, 2, 17, 13, 0, 30, 5, 0, 7, 7, 0, 
    0, 0, 0, 21, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 24, 22, 0, 0, 0, 0, 1, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 7, 1, 0, 0, 0, 0, 5, 2, 4, 4, 1, 0, 
    
    -- channel=124
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 18, 7, 0, 0, 
    18, 0, 0, 0, 0, 15, 0, 0, 0, 0, 2, 0, 4, 20, 0, 
    0, 6, 0, 0, 0, 0, 0, 2, 0, 7, 0, 13, 0, 8, 0, 
    0, 12, 1, 0, 0, 33, 0, 0, 3, 0, 0, 5, 0, 0, 52, 
    16, 0, 0, 68, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 5, 0, 0, 4, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 0, 30, 0, 12, 0, 0, 0, 0, 23, 0, 0, 0, 4, 0, 
    0, 0, 12, 0, 41, 0, 0, 0, 0, 34, 14, 0, 0, 0, 1, 
    0, 0, 0, 0, 2, 16, 0, 0, 65, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 33, 17, 0, 0, 0, 0, 0, 15, 0, 0, 
    37, 0, 0, 20, 29, 0, 8, 1, 0, 0, 0, 0, 0, 2, 0, 
    13, 42, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 2, 68, 0, 0, 0, 0, 4, 0, 0, 3, 0, 0, 0, 24, 
    0, 0, 20, 0, 5, 2, 0, 0, 0, 0, 7, 0, 0, 12, 0, 
    
    -- channel=125
    6, 5, 10, 5, 5, 9, 6, 5, 5, 0, 0, 7, 7, 1, 0, 
    9, 10, 11, 3, 14, 34, 0, 1, 0, 19, 0, 0, 9, 12, 3, 
    0, 23, 8, 4, 10, 0, 0, 0, 13, 45, 0, 0, 0, 10, 18, 
    0, 69, 3, 14, 0, 23, 0, 0, 0, 47, 0, 0, 0, 0, 44, 
    0, 38, 0, 61, 16, 3, 0, 0, 0, 73, 0, 0, 4, 0, 20, 
    0, 9, 0, 1, 35, 0, 0, 0, 0, 134, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 46, 46, 0, 0, 0, 102, 0, 0, 6, 16, 0, 
    0, 0, 0, 0, 35, 48, 0, 0, 0, 60, 0, 0, 16, 0, 0, 
    0, 0, 0, 25, 0, 0, 0, 0, 24, 0, 5, 0, 12, 18, 16, 
    0, 0, 0, 46, 0, 2, 32, 0, 0, 0, 0, 0, 32, 32, 0, 
    43, 0, 0, 123, 0, 0, 34, 0, 0, 0, 11, 20, 14, 11, 0, 
    28, 17, 0, 80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 30, 59, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 9, 
    0, 0, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 4, 0, 0, 0, 31, 0, 0, 
    
    -- channel=126
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=127
    38, 39, 40, 39, 39, 35, 45, 49, 40, 28, 24, 29, 31, 35, 32, 
    40, 44, 42, 41, 38, 17, 33, 34, 23, 0, 0, 0, 11, 26, 31, 
    22, 36, 44, 44, 43, 29, 12, 1, 0, 0, 0, 0, 0, 5, 24, 
    0, 3, 40, 41, 30, 9, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 27, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 24, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=128
    0, 1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 2, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=129
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=130
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 43, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=131
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=132
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=133
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=134
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=135
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 16, 1, 5, 0, 9, 7, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 25, 7, 0, 0, 9, 1, 25, 0, 0, 
    68, 0, 0, 0, 9, 0, 7, 8, 0, 0, 30, 0, 18, 17, 0, 
    52, 0, 23, 0, 0, 0, 29, 23, 13, 0, 6, 35, 0, 26, 0, 
    24, 0, 32, 0, 0, 0, 31, 20, 46, 0, 33, 37, 0, 9, 13, 
    20, 27, 3, 33, 0, 0, 7, 18, 46, 0, 47, 27, 0, 0, 15, 
    14, 19, 15, 21, 0, 0, 38, 0, 21, 0, 23, 33, 0, 0, 1, 
    20, 0, 59, 0, 6, 0, 14, 5, 0, 14, 0, 32, 0, 0, 0, 
    0, 0, 71, 0, 33, 0, 0, 17, 1, 0, 30, 0, 0, 0, 4, 
    0, 0, 63, 0, 66, 18, 0, 1, 43, 19, 0, 0, 0, 0, 6, 
    0, 0, 10, 0, 75, 33, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 5, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 53, 13, 0, 4, 0, 0, 0, 0, 0, 0, 0, 6, 
    17, 0, 0, 0, 2, 0, 0, 0, 0, 0, 3, 0, 0, 7, 35, 
    
    -- channel=136
    22, 23, 23, 24, 23, 23, 23, 24, 24, 20, 15, 14, 16, 17, 15, 
    21, 22, 24, 25, 25, 34, 28, 21, 14, 13, 15, 7, 5, 11, 16, 
    16, 11, 24, 24, 25, 28, 23, 7, 6, 19, 29, 20, 11, 1, 10, 
    17, 3, 23, 25, 24, 20, 27, 17, 11, 19, 31, 17, 11, 0, 0, 
    42, 30, 31, 33, 54, 44, 37, 19, 6, 12, 37, 23, 11, 4, 0, 
    51, 44, 36, 29, 41, 51, 47, 27, 9, 21, 51, 24, 13, 13, 3, 
    53, 43, 24, 20, 18, 44, 54, 39, 20, 26, 46, 21, 11, 18, 16, 
    60, 49, 30, 22, 24, 51, 48, 29, 21, 27, 42, 21, 12, 19, 17, 
    66, 57, 42, 28, 31, 25, 27, 22, 19, 22, 22, 10, 1, 12, 22, 
    62, 59, 44, 27, 35, 19, 27, 40, 25, 22, 7, 0, 1, 18, 24, 
    45, 58, 43, 47, 72, 43, 42, 48, 30, 8, 2, 7, 12, 17, 19, 
    25, 48, 53, 70, 75, 30, 16, 16, 15, 12, 12, 14, 18, 20, 20, 
    19, 21, 49, 75, 42, 15, 14, 12, 12, 13, 16, 20, 21, 22, 26, 
    21, 14, 31, 54, 25, 17, 17, 13, 13, 16, 18, 19, 18, 23, 24, 
    23, 15, 16, 16, 12, 11, 15, 16, 18, 21, 19, 16, 27, 35, 18, 
    
    -- channel=137
    29, 28, 30, 30, 30, 27, 31, 34, 31, 22, 17, 21, 25, 26, 28, 
    32, 32, 32, 30, 32, 33, 19, 21, 14, 14, 5, 4, 10, 23, 27, 
    10, 30, 32, 32, 33, 22, 8, 5, 6, 15, 0, 1, 0, 9, 27, 
    0, 28, 29, 32, 23, 22, 10, 1, 5, 12, 0, 1, 0, 0, 25, 
    0, 14, 17, 27, 13, 2, 0, 0, 0, 18, 1, 0, 7, 2, 9, 
    0, 0, 11, 15, 4, 0, 0, 0, 0, 29, 0, 0, 6, 2, 2, 
    0, 0, 6, 20, 21, 11, 0, 0, 0, 25, 0, 0, 4, 7, 2, 
    0, 0, 0, 15, 18, 8, 0, 0, 0, 21, 0, 0, 4, 5, 14, 
    0, 0, 0, 8, 0, 0, 0, 5, 8, 10, 1, 0, 8, 18, 24, 
    0, 0, 0, 7, 0, 0, 8, 4, 0, 0, 0, 2, 13, 27, 20, 
    5, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=138
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=139
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=140
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 3, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 1, 0, 0, 
    13, 0, 0, 0, 0, 0, 5, 0, 4, 0, 0, 2, 0, 2, 0, 
    12, 8, 0, 0, 0, 0, 2, 0, 7, 0, 10, 7, 0, 0, 0, 
    4, 24, 0, 0, 0, 0, 11, 0, 13, 0, 15, 3, 0, 0, 0, 
    6, 19, 0, 0, 0, 0, 15, 4, 1, 0, 3, 7, 0, 0, 0, 
    15, 15, 17, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 
    7, 10, 27, 0, 16, 0, 0, 5, 0, 0, 11, 0, 0, 0, 0, 
    7, 7, 27, 0, 15, 7, 4, 26, 26, 8, 6, 8, 16, 15, 15, 
    36, 17, 13, 0, 51, 37, 30, 29, 31, 25, 29, 30, 32, 33, 34, 
    44, 27, 0, 25, 43, 28, 31, 28, 27, 27, 30, 32, 38, 36, 33, 
    48, 38, 10, 52, 26, 27, 30, 30, 29, 31, 36, 40, 39, 34, 55, 
    48, 41, 35, 42, 30, 29, 32, 29, 26, 30, 37, 32, 23, 45, 52, 
    
    -- channel=141
    15, 13, 15, 17, 18, 13, 16, 18, 18, 12, 6, 6, 11, 15, 17, 
    18, 16, 16, 17, 16, 23, 17, 10, 3, 6, 12, 8, 2, 8, 16, 
    6, 2, 17, 17, 18, 5, 5, 2, 6, 8, 8, 5, 13, 4, 10, 
    18, 15, 18, 16, 16, 9, 17, 9, 9, 0, 7, 4, 6, 8, 4, 
    10, 20, 16, 5, 20, 11, 5, 6, 6, 0, 11, 12, 10, 13, 4, 
    0, 3, 12, 9, 0, 0, 11, 11, 17, 4, 3, 0, 5, 9, 11, 
    0, 10, 0, 17, 3, 4, 4, 7, 11, 5, 3, 8, 7, 9, 12, 
    0, 5, 5, 17, 11, 0, 0, 0, 5, 6, 4, 7, 3, 5, 9, 
    0, 0, 4, 3, 10, 0, 4, 13, 4, 15, 1, 0, 2, 9, 17, 
    0, 0, 7, 3, 2, 0, 0, 20, 5, 0, 0, 2, 9, 16, 12, 
    0, 0, 5, 2, 25, 17, 0, 0, 0, 6, 9, 10, 3, 0, 0, 
    0, 0, 1, 11, 0, 0, 0, 0, 0, 0, 2, 0, 2, 3, 2, 
    5, 0, 0, 5, 0, 0, 1, 2, 4, 5, 4, 4, 1, 0, 2, 
    1, 0, 0, 0, 0, 1, 4, 2, 0, 1, 1, 0, 0, 2, 0, 
    3, 0, 0, 0, 2, 0, 0, 0, 4, 5, 5, 2, 6, 9, 4, 
    
    -- channel=142
    8, 9, 10, 7, 6, 11, 9, 7, 5, 5, 10, 13, 12, 10, 7, 
    7, 10, 10, 6, 9, 4, 6, 8, 11, 14, 7, 12, 17, 12, 6, 
    5, 16, 8, 7, 7, 7, 5, 13, 18, 19, 5, 9, 2, 16, 12, 
    0, 20, 6, 8, 3, 14, 3, 9, 7, 25, 1, 12, 7, 8, 23, 
    0, 7, 2, 24, 0, 18, 6, 8, 7, 35, 6, 4, 10, 2, 23, 
    11, 6, 4, 19, 24, 25, 0, 5, 0, 38, 1, 5, 13, 6, 11, 
    16, 0, 14, 0, 21, 20, 0, 5, 0, 29, 0, 5, 13, 12, 6, 
    16, 0, 11, 0, 17, 15, 1, 11, 4, 21, 2, 3, 16, 12, 10, 
    7, 11, 1, 12, 11, 21, 8, 3, 14, 5, 12, 6, 19, 13, 9, 
    6, 10, 0, 22, 3, 23, 23, 0, 13, 10, 4, 15, 17, 13, 6, 
    12, 12, 0, 34, 0, 2, 17, 6, 1, 8, 11, 12, 11, 6, 3, 
    17, 17, 6, 16, 0, 7, 15, 15, 8, 8, 6, 8, 7, 6, 5, 
    0, 20, 31, 0, 0, 9, 8, 9, 6, 6, 6, 6, 5, 7, 6, 
    0, 7, 39, 0, 1, 9, 5, 8, 10, 9, 6, 5, 4, 7, 0, 
    0, 7, 11, 1, 3, 9, 7, 7, 9, 6, 3, 7, 10, 0, 0, 
    
    -- channel=143
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=144
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 3, 5, 
    0, 0, 0, 2, 0, 0, 14, 1, 8, 0, 4, 4, 0, 0, 2, 
    8, 0, 0, 2, 0, 0, 23, 10, 0, 0, 8, 6, 19, 0, 0, 
    56, 0, 1, 0, 7, 0, 5, 7, 1, 0, 31, 0, 18, 10, 0, 
    45, 0, 23, 0, 0, 0, 30, 22, 14, 0, 5, 30, 0, 22, 0, 
    25, 0, 32, 0, 0, 0, 28, 20, 39, 0, 34, 37, 0, 11, 10, 
    22, 18, 0, 36, 0, 0, 5, 22, 40, 0, 43, 23, 0, 0, 13, 
    12, 21, 7, 20, 0, 0, 51, 4, 23, 0, 22, 30, 0, 0, 9, 
    20, 0, 51, 0, 6, 0, 13, 2, 0, 20, 0, 38, 0, 0, 0, 
    0, 0, 61, 0, 21, 0, 0, 12, 1, 0, 34, 0, 0, 0, 3, 
    0, 0, 58, 0, 51, 3, 0, 6, 36, 21, 0, 0, 0, 0, 0, 
    0, 0, 11, 0, 63, 31, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 1, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 52, 12, 0, 2, 0, 0, 0, 0, 0, 0, 0, 3, 
    14, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 3, 25, 
    
    -- channel=145
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 25, 6, 0, 0, 3, 19, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 7, 9, 0, 0, 5, 0, 0, 
    17, 29, 0, 0, 0, 2, 15, 0, 0, 0, 0, 0, 0, 2, 0, 
    7, 28, 1, 0, 20, 18, 0, 3, 0, 11, 20, 9, 6, 6, 0, 
    0, 0, 0, 0, 0, 0, 11, 13, 16, 15, 0, 0, 0, 1, 17, 
    7, 0, 0, 0, 0, 9, 0, 0, 0, 1, 0, 11, 10, 11, 6, 
    6, 5, 17, 6, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    1, 0, 4, 0, 9, 0, 5, 15, 1, 17, 0, 0, 0, 5, 8, 
    0, 0, 1, 19, 0, 0, 6, 23, 8, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 30, 40, 30, 0, 0, 0, 6, 24, 17, 7, 0, 0, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 6, 8, 3, 
    6, 0, 0, 0, 0, 2, 0, 2, 4, 7, 10, 11, 0, 0, 14, 
    1, 5, 0, 0, 0, 4, 10, 5, 0, 2, 0, 0, 1, 11, 0, 
    0, 2, 3, 0, 0, 0, 0, 0, 6, 16, 7, 7, 22, 16, 1, 
    
    -- channel=146
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 9, 7, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 7, 7, 1, 3, 7, 1, 0, 
    10, 0, 0, 0, 0, 0, 0, 2, 7, 8, 0, 0, 4, 1, 0, 
    25, 15, 0, 0, 14, 1, 0, 0, 0, 13, 8, 6, 7, 6, 1, 
    21, 17, 0, 0, 0, 2, 5, 4, 1, 18, 10, 7, 9, 9, 0, 
    24, 19, 2, 0, 0, 9, 11, 9, 0, 0, 8, 6, 11, 3, 0, 
    29, 31, 20, 10, 0, 7, 0, 5, 2, 0, 3, 6, 6, 0, 0, 
    25, 27, 19, 24, 8, 5, 8, 5, 6, 4, 8, 10, 0, 0, 0, 
    36, 24, 19, 27, 15, 15, 33, 34, 25, 21, 30, 37, 44, 44, 42, 
    69, 48, 19, 24, 42, 58, 56, 56, 56, 57, 61, 65, 67, 66, 67, 
    76, 63, 42, 33, 51, 58, 57, 56, 57, 61, 67, 69, 69, 73, 75, 
    81, 72, 64, 50, 54, 59, 58, 57, 61, 65, 73, 76, 76, 83, 81, 
    77, 76, 69, 58, 58, 63, 63, 59, 59, 64, 66, 68, 71, 76, 72, 
    
    -- channel=147
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=148
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=149
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 10, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 10, 0, 0, 0, 0, 1, 0, 0, 6, 2, 0, 0, 0, 0, 
    8, 12, 0, 0, 0, 1, 8, 2, 0, 0, 0, 0, 0, 0, 0, 
    14, 19, 2, 1, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 18, 6, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 13, 8, 10, 3, 0, 11, 20, 6, 0, 0, 1, 9, 9, 4, 
    38, 31, 10, 16, 27, 28, 26, 25, 21, 19, 23, 27, 30, 31, 30, 
    35, 34, 24, 22, 24, 24, 23, 23, 22, 23, 28, 29, 32, 34, 35, 
    38, 32, 33, 34, 19, 25, 23, 22, 25, 28, 33, 36, 36, 36, 44, 
    38, 36, 33, 31, 22, 27, 28, 26, 25, 28, 29, 31, 32, 38, 35, 
    
    -- channel=150
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 2, 0, 0, 2, 38, 6, 0, 0, 13, 24, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 15, 0, 6, 3, 0, 0, 
    12, 28, 1, 3, 5, 15, 21, 4, 0, 0, 0, 0, 0, 0, 0, 
    23, 31, 2, 23, 63, 30, 0, 1, 0, 15, 17, 7, 6, 8, 0, 
    0, 0, 1, 0, 0, 0, 16, 9, 7, 29, 0, 0, 0, 6, 17, 
    7, 0, 0, 0, 0, 20, 0, 8, 0, 6, 0, 3, 2, 11, 2, 
    9, 11, 13, 19, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 2, 0, 10, 4, 0, 0, 7, 12, 0, 0, 0, 0, 2, 7, 
    0, 0, 0, 13, 0, 0, 16, 28, 0, 0, 0, 0, 12, 8, 0, 
    0, 0, 0, 42, 68, 41, 2, 0, 0, 10, 24, 31, 14, 7, 9, 
    0, 0, 11, 18, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 2, 5, 7, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 8, 0, 0, 22, 4, 0, 
    
    -- channel=151
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 26, 0, 0, 0, 14, 0, 0, 0, 27, 0, 0, 0, 10, 0, 
    0, 36, 0, 0, 0, 0, 0, 0, 0, 66, 0, 0, 0, 0, 51, 
    0, 0, 0, 33, 0, 0, 0, 0, 0, 68, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 73, 0, 0, 0, 0, 122, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 60, 6, 0, 0, 0, 105, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 24, 44, 0, 0, 0, 63, 0, 0, 15, 0, 0, 
    0, 0, 0, 10, 0, 16, 0, 0, 9, 0, 16, 0, 21, 5, 0, 
    0, 0, 0, 36, 0, 0, 11, 0, 0, 0, 0, 0, 21, 1, 0, 
    44, 0, 0, 94, 0, 0, 17, 0, 0, 0, 0, 0, 0, 7, 0, 
    89, 30, 0, 48, 0, 0, 16, 14, 0, 3, 5, 9, 4, 3, 0, 
    0, 75, 58, 0, 0, 0, 0, 0, 0, 3, 7, 3, 2, 9, 5, 
    0, 4, 120, 0, 0, 5, 0, 0, 6, 5, 6, 12, 0, 21, 0, 
    0, 6, 9, 22, 0, 28, 18, 0, 2, 0, 0, 9, 25, 0, 0, 
    
    -- channel=152
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=153
    9, 9, 12, 11, 12, 8, 13, 15, 12, 3, 0, 4, 7, 9, 11, 
    16, 14, 13, 11, 12, 26, 0, 6, 0, 0, 0, 0, 0, 8, 11, 
    0, 9, 14, 13, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 30, 11, 15, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 4, 0, 4, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 16, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=154
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=155
    4, 2, 0, 0, 0, 0, 0, 1, 0, 7, 15, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 26, 0, 0, 0, 16, 10, 0, 
    17, 29, 0, 0, 1, 49, 20, 25, 0, 0, 0, 0, 0, 17, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 9, 6, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 12, 
    5, 0, 0, 16, 59, 17, 0, 0, 0, 0, 0, 11, 1, 0, 0, 
    0, 0, 22, 0, 18, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 22, 27, 4, 2, 4, 4, 3, 6, 3, 
    0, 0, 0, 0, 0, 51, 12, 0, 0, 4, 29, 36, 19, 0, 0, 
    4, 0, 0, 0, 0, 1, 0, 0, 0, 28, 28, 10, 0, 0, 1, 
    0, 0, 1, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 6, 5, 
    51, 18, 0, 0, 50, 62, 42, 40, 15, 1, 0, 0, 0, 0, 0, 
    0, 39, 3, 0, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 33, 39, 5, 0, 0, 0, 0, 0, 0, 7, 0, 0, 19, 
    0, 0, 4, 51, 14, 16, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=156
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 2, 0, 3, 38, 0, 0, 0, 10, 0, 0, 0, 3, 0, 
    0, 10, 0, 0, 2, 2, 0, 0, 3, 45, 0, 0, 0, 0, 14, 
    0, 64, 0, 4, 0, 6, 0, 0, 0, 41, 0, 0, 0, 0, 37, 
    0, 47, 0, 32, 19, 0, 0, 0, 0, 57, 0, 0, 2, 0, 9, 
    0, 14, 0, 0, 46, 0, 0, 0, 0, 132, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 53, 41, 0, 0, 0, 108, 0, 0, 1, 13, 0, 
    0, 0, 0, 0, 26, 56, 0, 0, 0, 67, 0, 0, 12, 0, 0, 
    0, 0, 0, 27, 0, 0, 0, 2, 14, 0, 9, 0, 8, 17, 14, 
    0, 0, 0, 45, 0, 0, 14, 0, 0, 0, 0, 0, 32, 31, 0, 
    53, 0, 0, 118, 0, 0, 35, 0, 0, 0, 5, 16, 10, 3, 0, 
    30, 12, 0, 92, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 28, 36, 0, 0, 0, 0, 0, 0, 0, 3, 4, 0, 0, 7, 
    0, 0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 4, 0, 0, 0, 30, 0, 0, 
    
    -- channel=157
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 4, 20, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 13, 2, 0, 
    27, 0, 0, 0, 4, 0, 0, 18, 0, 0, 0, 0, 0, 18, 0, 
    0, 0, 21, 0, 0, 49, 0, 11, 0, 0, 0, 29, 0, 0, 35, 
    46, 0, 12, 66, 0, 0, 0, 0, 14, 0, 16, 2, 0, 0, 19, 
    42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 9, 
    36, 0, 52, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    2, 0, 66, 0, 65, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 37, 0, 0, 59, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 46, 0, 0, 0, 12, 1, 3, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=158
    36, 35, 37, 37, 37, 33, 39, 42, 36, 26, 19, 22, 26, 32, 31, 
    38, 38, 40, 38, 37, 31, 30, 25, 11, 4, 0, 4, 12, 23, 29, 
    15, 27, 39, 39, 42, 24, 6, 1, 4, 4, 0, 0, 0, 13, 24, 
    0, 29, 37, 38, 25, 14, 5, 0, 0, 9, 0, 0, 0, 1, 25, 
    0, 15, 27, 28, 2, 5, 0, 0, 0, 12, 0, 0, 0, 0, 15, 
    0, 0, 21, 24, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 
    0, 0, 16, 15, 16, 8, 0, 0, 0, 15, 0, 0, 0, 0, 2, 
    0, 0, 1, 7, 17, 5, 0, 0, 0, 19, 0, 0, 0, 2, 14, 
    0, 0, 0, 0, 4, 0, 0, 0, 5, 6, 2, 0, 3, 18, 34, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 9, 28, 23, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=159
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=160
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=161
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=162
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=163
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=164
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=165
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 1, 0, 0, 0, 
    1, 20, 0, 0, 0, 0, 13, 1, 0, 0, 0, 0, 0, 0, 0, 
    6, 26, 0, 1, 51, 20, 0, 0, 0, 0, 3, 3, 2, 7, 0, 
    0, 0, 0, 0, 0, 0, 7, 0, 7, 24, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 4, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 11, 
    0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 7, 5, 0, 
    0, 0, 0, 32, 62, 38, 0, 0, 0, 0, 11, 23, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 
    
    -- channel=166
    11, 12, 7, 7, 7, 5, 11, 13, 7, 16, 25, 20, 10, 8, 8, 
    3, 5, 6, 10, 3, 0, 4, 17, 41, 0, 0, 0, 7, 12, 8, 
    33, 32, 8, 9, 7, 37, 25, 9, 0, 0, 0, 0, 0, 5, 7, 
    0, 0, 6, 3, 7, 0, 0, 0, 0, 0, 8, 4, 7, 0, 0, 
    0, 0, 11, 0, 0, 0, 3, 0, 9, 0, 0, 0, 0, 0, 0, 
    2, 0, 15, 12, 20, 13, 0, 0, 0, 0, 13, 18, 0, 0, 0, 
    0, 2, 18, 22, 0, 0, 11, 0, 8, 0, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 47, 21, 10, 0, 8, 2, 0, 5, 5, 
    0, 0, 2, 0, 0, 26, 0, 0, 0, 0, 6, 44, 0, 0, 0, 
    0, 0, 7, 0, 3, 1, 0, 0, 0, 37, 44, 1, 0, 0, 13, 
    0, 0, 14, 0, 0, 0, 0, 33, 26, 0, 0, 0, 0, 0, 0, 
    8, 1, 0, 0, 66, 36, 2, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=167
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=168
    20, 22, 23, 23, 23, 21, 24, 28, 25, 15, 9, 11, 16, 20, 22, 
    24, 26, 26, 24, 24, 15, 18, 15, 10, 0, 0, 0, 0, 9, 18, 
    2, 11, 23, 26, 25, 6, 1, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 18, 25, 14, 8, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 12, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=169
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=170
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 1, 0, 0, 1, 36, 0, 0, 0, 11, 12, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 20, 0, 0, 0, 0, 0, 
    0, 47, 0, 2, 0, 11, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 22, 0, 21, 17, 7, 0, 0, 0, 39, 5, 0, 5, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 30, 0, 0, 0, 26, 0, 0, 7, 13, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 7, 0, 0, 7, 8, 0, 0, 0, 0, 11, 10, 
    0, 0, 0, 19, 0, 0, 17, 1, 0, 0, 0, 0, 9, 7, 0, 
    0, 0, 0, 72, 12, 14, 0, 0, 0, 0, 23, 21, 4, 0, 0, 
    0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17, 0, 0, 0, 0, 0, 0, 1, 3, 4, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 0, 0, 24, 0, 0, 
    
    -- channel=171
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=172
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=173
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=174
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 4, 
    36, 5, 0, 0, 0, 21, 23, 22, 18, 19, 21, 23, 22, 24, 22, 
    31, 33, 4, 0, 10, 17, 19, 19, 19, 21, 23, 22, 25, 28, 22, 
    31, 29, 35, 0, 13, 20, 16, 19, 21, 22, 29, 31, 30, 28, 38, 
    28, 30, 31, 23, 24, 27, 26, 20, 17, 17, 23, 26, 19, 20, 27, 
    
    -- channel=175
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 7, 5, 0, 0, 0, 0, 22, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 
    0, 0, 3, 5, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 38, 
    7, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 0, 15, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=176
    5, 3, 2, 0, 2, 0, 5, 11, 5, 1, 3, 5, 0, 3, 7, 
    5, 3, 3, 2, 0, 0, 0, 0, 5, 0, 0, 0, 0, 7, 3, 
    0, 23, 5, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=177
    15, 17, 15, 14, 14, 13, 17, 20, 15, 10, 9, 10, 8, 7, 9, 
    13, 15, 16, 16, 16, 0, 0, 11, 13, 0, 0, 0, 0, 8, 6, 
    6, 25, 17, 18, 19, 31, 6, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 9, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 17, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 4, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=178
    70, 74, 74, 73, 72, 70, 77, 82, 73, 59, 51, 55, 59, 63, 61, 
    72, 77, 77, 76, 73, 72, 65, 66, 47, 25, 11, 17, 31, 50, 59, 
    51, 59, 77, 78, 78, 64, 43, 19, 13, 16, 8, 6, 6, 21, 51, 
    5, 32, 70, 76, 66, 40, 26, 9, 6, 19, 20, 16, 5, 5, 37, 
    0, 23, 60, 54, 39, 33, 22, 12, 6, 18, 18, 11, 8, 1, 19, 
    0, 22, 60, 65, 41, 36, 31, 13, 3, 28, 22, 8, 8, 2, 2, 
    1, 18, 44, 57, 36, 40, 28, 20, 4, 26, 12, 6, 6, 7, 11, 
    11, 7, 11, 34, 28, 36, 21, 21, 13, 36, 21, 6, 6, 18, 33, 
    10, 11, 3, 20, 29, 20, 18, 15, 12, 30, 22, 8, 10, 30, 57, 
    20, 14, 1, 7, 7, 18, 17, 13, 14, 23, 5, 0, 10, 52, 58, 
    14, 17, 1, 19, 8, 0, 12, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 2, 36, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=179
    0, 2, 0, 0, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 1, 0, 2, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 3, 51, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 9, 3, 20, 0, 0, 10, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 34, 5, 1, 0, 10, 0, 0, 0, 0, 0, 
    0, 12, 0, 0, 0, 10, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    17, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 12, 0, 6, 0, 0, 5, 19, 0, 0, 0, 0, 0, 0, 0, 
    13, 20, 0, 35, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 19, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=180
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=181
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 7, 6, 1, 2, 
    9, 0, 0, 0, 0, 0, 1, 4, 6, 9, 10, 5, 0, 3, 0, 
    10, 14, 0, 0, 0, 0, 0, 5, 6, 6, 9, 9, 11, 12, 0, 
    3, 15, 9, 0, 6, 13, 4, 0, 0, 0, 4, 11, 1, 0, 7, 
    
    -- channel=182
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 8, 5, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 5, 0, 0, 3, 3, 0, 
    2, 6, 0, 0, 0, 0, 0, 0, 7, 2, 0, 0, 3, 3, 0, 
    12, 14, 0, 0, 3, 0, 0, 0, 3, 11, 1, 0, 6, 5, 2, 
    6, 19, 0, 0, 0, 0, 0, 0, 0, 18, 1, 2, 7, 6, 0, 
    9, 12, 0, 0, 0, 5, 4, 4, 0, 3, 0, 2, 8, 4, 0, 
    16, 22, 12, 6, 0, 0, 0, 1, 1, 0, 0, 1, 6, 0, 0, 
    13, 19, 12, 20, 2, 0, 0, 2, 7, 0, 5, 7, 6, 0, 0, 
    26, 13, 12, 19, 9, 12, 28, 24, 18, 15, 26, 34, 41, 34, 27, 
    65, 35, 11, 22, 27, 39, 47, 46, 48, 51, 58, 61, 63, 64, 63, 
    76, 60, 27, 25, 31, 54, 55, 54, 55, 59, 65, 67, 68, 68, 71, 
    78, 70, 57, 39, 44, 57, 56, 55, 57, 62, 70, 72, 72, 78, 82, 
    75, 74, 68, 53, 55, 60, 60, 56, 57, 62, 65, 66, 67, 76, 72, 
    
    -- channel=183
    6, 4, 6, 6, 7, 3, 6, 7, 6, 7, 6, 4, 4, 6, 7, 
    7, 3, 6, 7, 5, 0, 6, 4, 6, 0, 0, 0, 0, 4, 8, 
    8, 6, 6, 6, 7, 1, 0, 0, 0, 0, 0, 0, 8, 4, 4, 
    7, 3, 6, 4, 4, 0, 0, 4, 5, 0, 0, 0, 0, 6, 3, 
    0, 4, 8, 0, 0, 0, 0, 0, 4, 0, 0, 2, 1, 7, 5, 
    0, 0, 3, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 3, 4, 
    0, 0, 0, 4, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 6, 6, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 2, 2, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    
    -- channel=184
    35, 36, 34, 33, 32, 30, 39, 41, 33, 30, 33, 34, 30, 31, 29, 
    32, 35, 35, 35, 31, 0, 25, 33, 39, 0, 0, 0, 18, 30, 27, 
    31, 47, 35, 37, 35, 42, 25, 13, 0, 0, 0, 0, 0, 17, 26, 
    0, 0, 32, 32, 21, 6, 0, 0, 0, 2, 0, 3, 0, 1, 24, 
    0, 0, 24, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 27, 24, 22, 13, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 33, 27, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 8, 9, 3, 0, 0, 0, 0, 2, 17, 
    0, 0, 0, 0, 0, 21, 1, 0, 0, 0, 11, 22, 6, 5, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 17, 1, 0, 8, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=185
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 29, 0, 0, 26, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 13, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 55, 42, 39, 3, 0, 0, 0, 19, 34, 16, 0, 0, 
    0, 0, 0, 31, 0, 0, 0, 0, 0, 5, 13, 14, 23, 21, 17, 
    23, 0, 0, 0, 0, 13, 11, 10, 13, 22, 29, 34, 17, 14, 41, 
    20, 23, 0, 0, 0, 17, 18, 15, 14, 20, 17, 11, 16, 42, 0, 
    18, 25, 11, 0, 0, 0, 0, 10, 27, 31, 20, 22, 54, 39, 16, 
    
    -- channel=186
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 38, 0, 0, 0, 0, 0, 0, 12, 20, 16, 0, 0, 
    13, 0, 0, 8, 0, 0, 2, 2, 7, 15, 20, 23, 27, 26, 21, 
    27, 19, 5, 0, 0, 18, 16, 17, 19, 26, 31, 32, 22, 23, 36, 
    25, 30, 32, 0, 0, 21, 18, 19, 22, 26, 28, 25, 26, 46, 14, 
    20, 34, 27, 0, 10, 22, 15, 16, 25, 27, 22, 28, 45, 27, 14, 
    
    -- channel=187
    0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 3, 39, 0, 0, 0, 24, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 7, 
    0, 54, 0, 6, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 34, 0, 0, 0, 0, 0, 52, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 14, 0, 
    0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 59, 0, 0, 0, 0, 0, 0, 15, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=188
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=189
    2, 2, 5, 1, 2, 5, 3, 3, 5, 3, 7, 11, 9, 3, 2, 
    5, 5, 6, 0, 7, 0, 0, 4, 9, 13, 0, 0, 7, 13, 2, 
    0, 26, 4, 2, 3, 0, 0, 2, 11, 3, 0, 0, 0, 7, 9, 
    0, 18, 0, 8, 0, 18, 0, 0, 0, 10, 0, 0, 0, 0, 24, 
    0, 0, 0, 41, 0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 4, 5, 0, 0, 0, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 7, 14, 0, 0, 0, 0, 7, 9, 3, 0, 
    0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=190
    11, 9, 15, 13, 13, 12, 12, 15, 15, 0, 0, 0, 7, 11, 13, 
    16, 16, 15, 11, 16, 20, 3, 0, 0, 5, 0, 0, 0, 5, 9, 
    0, 1, 15, 15, 16, 0, 0, 0, 10, 0, 0, 0, 0, 0, 6, 
    0, 31, 8, 17, 3, 12, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 27, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 7, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 0, 
    0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=191
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 7, 0, 0, 13, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 24, 24, 23, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=192
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 28, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 42, 22, 23, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=193
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 7, 16, 25, 27, 29, 31, 30, 
    54, 7, 0, 0, 0, 16, 19, 20, 25, 32, 36, 36, 32, 32, 34, 
    56, 43, 0, 0, 0, 20, 20, 24, 25, 30, 40, 42, 44, 49, 46, 
    49, 49, 34, 3, 25, 31, 26, 21, 20, 24, 36, 40, 31, 36, 52, 
    
    -- channel=194
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=195
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 24, 0, 0, 0, 2, 0, 0, 0, 1, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 1, 10, 
    0, 55, 0, 1, 0, 1, 0, 0, 0, 31, 0, 0, 0, 0, 33, 
    0, 40, 0, 25, 12, 0, 0, 0, 0, 45, 0, 0, 0, 0, 10, 
    0, 4, 0, 0, 22, 0, 0, 0, 0, 107, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 37, 26, 0, 0, 0, 85, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 19, 40, 0, 0, 0, 48, 0, 0, 5, 0, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 10, 0, 0, 0, 2, 11, 10, 
    0, 0, 0, 32, 0, 0, 7, 0, 0, 0, 0, 0, 28, 26, 0, 
    33, 0, 0, 92, 0, 0, 23, 0, 0, 0, 1, 10, 4, 0, 0, 
    17, 0, 0, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 17, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 
    
    -- channel=196
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 0, 39, 21, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 12, 1, 3, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 7, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 50, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=197
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 18, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 10, 9, 8, 5, 5, 
    7, 0, 0, 0, 0, 7, 8, 10, 11, 14, 14, 9, 2, 5, 5, 
    6, 14, 0, 0, 0, 7, 6, 10, 13, 11, 8, 5, 9, 10, 0, 
    2, 14, 9, 0, 6, 11, 6, 9, 9, 4, 5, 14, 10, 0, 7, 
    
    -- channel=198
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=199
    6, 5, 0, 0, 1, 1, 3, 6, 2, 9, 15, 10, 0, 1, 2, 
    0, 0, 0, 2, 0, 0, 0, 5, 27, 0, 0, 0, 13, 7, 0, 
    21, 21, 1, 3, 5, 48, 20, 21, 0, 0, 0, 0, 0, 15, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 9, 0, 11, 5, 2, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 11, 
    8, 0, 0, 24, 46, 15, 0, 0, 0, 0, 1, 11, 0, 0, 0, 
    0, 0, 21, 1, 12, 0, 1, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 23, 25, 2, 0, 5, 7, 0, 6, 3, 
    0, 0, 0, 0, 0, 45, 11, 0, 0, 8, 28, 34, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 26, 4, 0, 0, 5, 
    0, 0, 5, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 
    39, 4, 0, 0, 62, 53, 33, 31, 7, 0, 0, 0, 0, 0, 0, 
    0, 29, 0, 7, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 21, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 41, 9, 9, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=200
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=201
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=202
    36, 39, 41, 39, 40, 37, 42, 45, 42, 29, 22, 28, 32, 34, 34, 
    43, 43, 44, 40, 42, 46, 29, 32, 17, 15, 2, 3, 13, 27, 32, 
    17, 33, 41, 43, 43, 26, 10, 2, 4, 12, 0, 0, 0, 9, 31, 
    0, 35, 36, 44, 33, 24, 8, 0, 0, 10, 0, 0, 0, 0, 30, 
    0, 15, 21, 40, 16, 7, 0, 0, 0, 22, 0, 0, 1, 0, 12, 
    0, 0, 14, 23, 7, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 
    0, 0, 10, 20, 24, 17, 0, 0, 0, 27, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 19, 9, 0, 0, 0, 22, 0, 0, 0, 0, 12, 
    0, 0, 0, 8, 0, 0, 0, 0, 6, 5, 0, 0, 1, 17, 32, 
    0, 0, 0, 4, 0, 0, 8, 0, 0, 0, 0, 0, 13, 35, 28, 
    0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=203
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 1, 3, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 8, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 0, 
    8, 9, 0, 0, 0, 0, 6, 0, 8, 0, 5, 0, 0, 1, 0, 
    6, 24, 0, 0, 0, 0, 4, 0, 4, 5, 4, 3, 1, 2, 0, 
    13, 18, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 
    21, 20, 15, 2, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    12, 16, 19, 13, 4, 0, 0, 15, 3, 0, 0, 0, 0, 0, 0, 
    18, 14, 16, 11, 33, 21, 21, 16, 13, 9, 17, 25, 28, 15, 13, 
    30, 18, 10, 22, 29, 20, 27, 26, 30, 31, 37, 40, 43, 44, 44, 
    53, 30, 7, 31, 17, 37, 38, 35, 36, 39, 44, 47, 46, 45, 50, 
    54, 48, 24, 31, 27, 37, 40, 38, 38, 43, 47, 47, 48, 54, 55, 
    54, 52, 46, 27, 32, 35, 35, 36, 40, 45, 46, 43, 48, 61, 52, 
    
    -- channel=204
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=205
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=206
    1, 0, 5, 0, 0, 4, 1, 0, 0, 0, 0, 2, 1, 0, 0, 
    3, 4, 7, 0, 9, 20, 0, 0, 0, 14, 0, 0, 5, 8, 0, 
    0, 18, 3, 0, 7, 2, 0, 0, 11, 43, 0, 0, 0, 9, 12, 
    0, 62, 0, 8, 0, 17, 0, 0, 0, 52, 0, 0, 0, 0, 42, 
    0, 34, 0, 57, 3, 2, 0, 0, 0, 72, 0, 0, 0, 0, 20, 
    0, 6, 0, 10, 41, 0, 0, 0, 0, 134, 0, 0, 8, 0, 0, 
    0, 0, 0, 0, 50, 44, 0, 0, 0, 105, 0, 0, 4, 14, 0, 
    0, 0, 0, 0, 41, 53, 0, 0, 0, 63, 0, 0, 17, 0, 0, 
    0, 1, 0, 22, 0, 0, 0, 0, 20, 0, 11, 0, 12, 14, 12, 
    0, 0, 0, 47, 0, 0, 27, 0, 0, 0, 0, 0, 30, 27, 0, 
    44, 0, 0, 119, 0, 0, 38, 0, 0, 0, 7, 17, 13, 8, 0, 
    37, 18, 0, 85, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 
    0, 37, 58, 0, 0, 0, 0, 0, 0, 2, 5, 5, 0, 0, 9, 
    0, 0, 87, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 20, 0, 
    0, 0, 3, 0, 0, 6, 0, 0, 6, 0, 0, 1, 32, 0, 0, 
    
    -- channel=207
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 3, 0, 
    0, 22, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 2, 6, 
    0, 39, 0, 0, 0, 7, 0, 0, 0, 32, 0, 0, 0, 0, 36, 
    0, 0, 0, 36, 0, 0, 0, 0, 0, 59, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 31, 0, 0, 0, 0, 95, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 29, 15, 0, 0, 0, 66, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 10, 0, 0, 0, 32, 0, 0, 4, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 5, 0, 0, 0, 9, 6, 0, 
    0, 0, 0, 21, 0, 0, 14, 0, 0, 0, 0, 0, 14, 4, 0, 
    17, 0, 0, 72, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 4, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    
    -- channel=208
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 5, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    13, 13, 0, 0, 11, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 
    14, 13, 0, 0, 0, 5, 2, 0, 0, 25, 0, 0, 2, 5, 0, 
    18, 15, 0, 0, 0, 14, 0, 0, 0, 8, 0, 0, 4, 0, 0, 
    24, 28, 7, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 26, 6, 24, 0, 0, 4, 5, 3, 0, 0, 0, 0, 0, 0, 
    31, 21, 6, 41, 15, 15, 27, 20, 6, 4, 17, 25, 30, 20, 14, 
    53, 35, 14, 38, 21, 28, 36, 36, 35, 36, 42, 46, 50, 51, 50, 
    55, 50, 36, 29, 21, 41, 40, 39, 40, 45, 51, 54, 52, 54, 60, 
    59, 53, 56, 25, 32, 45, 42, 42, 44, 49, 54, 56, 55, 67, 58, 
    56, 58, 51, 37, 37, 45, 44, 42, 46, 50, 50, 52, 61, 63, 50, 
    
    -- channel=209
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 1, 40, 3, 0, 0, 0, 16, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 16, 4, 9, 4, 0, 0, 
    11, 22, 0, 0, 0, 1, 23, 10, 1, 0, 0, 0, 0, 0, 0, 
    23, 41, 2, 12, 72, 40, 0, 4, 0, 7, 16, 12, 9, 13, 0, 
    0, 0, 1, 0, 0, 0, 19, 11, 13, 35, 0, 0, 0, 8, 21, 
    6, 0, 0, 0, 0, 17, 0, 9, 0, 7, 0, 2, 0, 12, 12, 
    8, 7, 8, 9, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 2, 6, 0, 0, 6, 8, 0, 0, 0, 0, 3, 14, 
    0, 0, 0, 3, 0, 0, 6, 34, 0, 0, 0, 0, 15, 13, 0, 
    0, 0, 0, 49, 85, 58, 12, 0, 0, 1, 20, 36, 10, 0, 0, 
    0, 0, 12, 27, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 5, 8, 12, 0, 0, 18, 
    0, 0, 0, 0, 0, 1, 6, 0, 0, 2, 0, 0, 0, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 13, 13, 0, 0, 29, 15, 0, 
    
    -- channel=210
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 15, 1, 0, 0, 11, 8, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 22, 6, 0, 0, 10, 5, 25, 0, 0, 
    68, 0, 0, 0, 13, 0, 12, 7, 1, 0, 33, 0, 17, 13, 0, 
    48, 0, 22, 0, 11, 0, 32, 25, 15, 0, 9, 34, 0, 27, 0, 
    17, 0, 30, 0, 0, 0, 37, 22, 51, 0, 34, 34, 0, 11, 14, 
    14, 32, 0, 36, 0, 0, 7, 22, 46, 0, 43, 27, 0, 0, 16, 
    10, 26, 9, 24, 0, 0, 43, 0, 20, 0, 22, 33, 0, 0, 3, 
    21, 0, 55, 0, 7, 0, 11, 10, 0, 20, 0, 31, 0, 0, 0, 
    0, 0, 70, 0, 25, 0, 0, 23, 3, 0, 28, 0, 0, 0, 2, 
    0, 0, 62, 0, 72, 16, 0, 0, 36, 22, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 65, 23, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 12, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 56, 10, 0, 5, 0, 0, 0, 0, 0, 0, 0, 3, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 12, 30, 
    
    -- channel=211
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=212
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 16, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 28, 0, 0, 0, 6, 7, 0, 
    20, 29, 0, 0, 0, 34, 2, 2, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 7, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 9, 
    1, 0, 0, 10, 38, 13, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 13, 0, 13, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 22, 18, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 21, 26, 8, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 36, 25, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 28, 8, 0, 0, 0, 0, 0, 0, 
    48, 12, 0, 0, 41, 29, 14, 13, 0, 0, 0, 0, 0, 0, 0, 
    0, 31, 0, 1, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 36, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 26, 3, 8, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=213
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 7, 14, 13, 6, 8, 8, 10, 5, 8, 9, 
    17, 16, 0, 0, 0, 3, 7, 6, 8, 8, 7, 6, 11, 10, 0, 
    17, 14, 7, 0, 0, 4, 3, 9, 7, 8, 14, 17, 13, 11, 28, 
    15, 15, 16, 17, 16, 16, 11, 2, 0, 1, 12, 9, 0, 7, 16, 
    
    -- channel=214
    0, 0, 2, 3, 3, 0, 2, 3, 4, 0, 0, 0, 0, 2, 4, 
    5, 4, 3, 2, 3, 11, 1, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=215
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=216
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 16, 0, 0, 0, 0, 0, 
    0, 15, 0, 0, 0, 0, 33, 38, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 9, 0, 24, 0, 0, 
    36, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 1, 0, 
    7, 0, 4, 0, 0, 17, 0, 2, 0, 0, 0, 33, 0, 4, 0, 
    29, 0, 18, 3, 0, 0, 0, 5, 4, 0, 26, 4, 0, 0, 0, 
    0, 14, 0, 8, 0, 0, 12, 2, 23, 0, 18, 14, 0, 0, 27, 
    0, 0, 0, 0, 0, 33, 33, 0, 0, 0, 0, 42, 1, 6, 0, 
    3, 0, 17, 0, 0, 0, 26, 0, 0, 0, 31, 20, 0, 0, 0, 
    0, 0, 29, 0, 0, 0, 0, 0, 6, 24, 0, 0, 0, 0, 3, 
    0, 4, 15, 0, 0, 85, 26, 29, 19, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 0, 108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 25, 24, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 0, 0, 41, 5, 0, 0, 0, 0, 0, 0, 5, 0, 0, 17, 
    
    -- channel=217
    0, 2, 5, 6, 5, 3, 3, 3, 4, 0, 0, 0, 1, 3, 4, 
    6, 6, 5, 6, 6, 44, 10, 0, 0, 0, 12, 0, 0, 0, 3, 
    0, 0, 3, 6, 2, 0, 0, 0, 0, 2, 3, 6, 8, 0, 0, 
    21, 0, 0, 4, 8, 0, 21, 8, 2, 0, 12, 0, 0, 0, 0, 
    32, 24, 11, 0, 68, 40, 8, 9, 0, 0, 11, 18, 2, 14, 0, 
    0, 0, 14, 0, 0, 0, 32, 10, 20, 0, 8, 0, 0, 7, 15, 
    7, 3, 0, 14, 0, 10, 0, 19, 7, 0, 1, 4, 0, 2, 10, 
    14, 10, 3, 12, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    17, 0, 16, 0, 11, 0, 0, 6, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 21, 0, 0, 0, 0, 33, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 5, 4, 102, 43, 6, 0, 4, 2, 0, 18, 0, 0, 0, 
    0, 0, 10, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 0, 
    
    -- channel=218
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=219
    7, 3, 8, 3, 4, 7, 5, 4, 2, 0, 0, 8, 6, 1, 0, 
    7, 7, 9, 1, 11, 14, 0, 0, 0, 13, 0, 0, 9, 13, 0, 
    0, 29, 7, 3, 10, 5, 0, 0, 11, 38, 0, 0, 0, 14, 15, 
    0, 57, 2, 11, 0, 19, 0, 0, 0, 53, 0, 0, 0, 0, 45, 
    0, 26, 0, 57, 0, 1, 0, 0, 0, 74, 0, 0, 0, 0, 24, 
    0, 9, 0, 11, 42, 2, 0, 0, 0, 120, 0, 0, 10, 0, 0, 
    0, 0, 1, 0, 46, 41, 0, 0, 0, 93, 0, 0, 7, 13, 0, 
    0, 0, 0, 0, 39, 44, 0, 0, 0, 59, 0, 0, 19, 4, 0, 
    0, 4, 0, 23, 0, 9, 0, 0, 24, 0, 8, 0, 17, 19, 13, 
    0, 5, 0, 45, 0, 11, 33, 0, 0, 0, 0, 0, 29, 27, 0, 
    39, 3, 0, 106, 0, 0, 35, 0, 0, 0, 5, 13, 13, 9, 0, 
    41, 28, 0, 71, 0, 0, 0, 0, 0, 0, 2, 4, 3, 2, 0, 
    0, 42, 68, 0, 0, 0, 0, 0, 0, 3, 6, 6, 0, 3, 10, 
    0, 3, 88, 0, 0, 5, 0, 0, 3, 3, 1, 0, 0, 17, 0, 
    0, 1, 8, 0, 0, 10, 3, 0, 7, 0, 0, 5, 29, 0, 0, 
    
    -- channel=220
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 0, 0, 0, 0, 41, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=221
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 17, 0, 8, 0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 108, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 3, 0, 
    0, 0, 0, 76, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=222
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=223
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=224
    52, 52, 52, 52, 53, 48, 56, 60, 52, 42, 37, 40, 42, 45, 45, 
    53, 53, 54, 54, 52, 38, 42, 42, 35, 17, 3, 11, 27, 40, 43, 
    34, 51, 55, 56, 57, 55, 33, 20, 7, 8, 1, 3, 5, 23, 41, 
    0, 27, 51, 53, 42, 28, 8, 2, 6, 18, 10, 12, 7, 9, 37, 
    0, 8, 41, 34, 0, 2, 6, 3, 8, 16, 4, 0, 5, 1, 21, 
    0, 13, 39, 41, 34, 17, 7, 4, 0, 13, 5, 5, 8, 1, 0, 
    0, 7, 37, 35, 30, 16, 10, 6, 0, 16, 4, 1, 7, 3, 6, 
    0, 0, 4, 20, 19, 12, 10, 18, 10, 28, 12, 5, 7, 14, 31, 
    0, 0, 0, 12, 10, 25, 16, 7, 11, 25, 18, 13, 16, 29, 39, 
    6, 2, 0, 4, 0, 8, 10, 0, 6, 16, 10, 1, 8, 35, 40, 
    5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=225
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 27, 9, 0, 0, 0, 17, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 9, 0, 0, 
    24, 10, 0, 0, 3, 0, 16, 9, 1, 0, 3, 0, 0, 0, 0, 
    26, 19, 9, 0, 41, 38, 2, 8, 0, 0, 11, 18, 2, 12, 0, 
    4, 0, 9, 0, 0, 0, 16, 10, 20, 0, 2, 0, 0, 6, 20, 
    19, 0, 0, 2, 0, 3, 0, 13, 1, 0, 0, 10, 0, 3, 10, 
    18, 0, 17, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 23, 0, 19, 0, 0, 6, 0, 6, 0, 0, 0, 0, 5, 
    0, 0, 13, 0, 0, 0, 0, 22, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 79, 44, 0, 0, 0, 11, 14, 22, 4, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 3, 8, 0, 0, 10, 12, 2, 
    
    -- channel=226
    34, 34, 33, 33, 33, 30, 37, 39, 33, 29, 27, 27, 27, 32, 32, 
    31, 35, 34, 36, 31, 6, 33, 30, 33, 2, 0, 7, 15, 22, 29, 
    27, 28, 34, 36, 35, 34, 24, 17, 2, 0, 0, 0, 8, 13, 21, 
    14, 0, 32, 31, 26, 10, 1, 3, 1, 0, 7, 7, 6, 8, 13, 
    0, 0, 32, 7, 0, 2, 9, 5, 8, 0, 0, 8, 0, 5, 12, 
    0, 0, 30, 29, 0, 8, 0, 5, 7, 0, 6, 11, 0, 1, 2, 
    0, 0, 19, 36, 3, 0, 0, 0, 10, 0, 6, 1, 0, 0, 4, 
    0, 0, 0, 14, 3, 0, 17, 8, 8, 0, 3, 6, 0, 5, 18, 
    0, 0, 0, 0, 4, 14, 6, 0, 0, 19, 2, 21, 5, 7, 21, 
    0, 0, 0, 0, 1, 5, 0, 0, 1, 12, 19, 4, 0, 10, 25, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=227
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 5, 25, 1, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 12, 17, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 43, 43, 22, 21, 21, 17, 17, 18, 13, 14, 18, 
    28, 14, 0, 0, 51, 13, 18, 15, 16, 13, 13, 9, 22, 24, 4, 
    35, 21, 0, 48, 23, 11, 13, 15, 17, 16, 24, 30, 28, 10, 52, 
    34, 26, 20, 39, 29, 26, 31, 19, 7, 6, 21, 18, 0, 15, 41, 
    
    -- channel=228
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=229
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 1, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    13, 4, 0, 0, 0, 0, 0, 0, 2, 0, 8, 4, 0, 0, 0, 
    6, 17, 0, 0, 0, 0, 7, 0, 7, 0, 8, 1, 0, 0, 0, 
    7, 11, 0, 0, 0, 0, 13, 2, 0, 0, 0, 3, 0, 0, 0, 
    15, 15, 16, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    6, 9, 21, 0, 14, 0, 0, 0, 1, 3, 9, 1, 0, 0, 0, 
    8, 7, 19, 0, 10, 13, 16, 30, 27, 10, 12, 17, 26, 25, 24, 
    46, 22, 10, 0, 47, 38, 32, 33, 36, 34, 39, 39, 40, 41, 44, 
    54, 38, 2, 26, 43, 35, 38, 35, 35, 36, 40, 43, 48, 47, 44, 
    58, 48, 28, 50, 33, 35, 37, 37, 37, 41, 46, 50, 48, 50, 64, 
    56, 50, 43, 44, 37, 39, 42, 37, 34, 38, 44, 40, 34, 54, 57, 
    
    -- channel=230
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=231
    0, 0, 3, 3, 4, 2, 0, 2, 4, 0, 0, 0, 3, 2, 4, 
    9, 6, 2, 1, 6, 47, 3, 0, 0, 17, 24, 5, 0, 0, 4, 
    0, 0, 3, 4, 0, 0, 0, 0, 9, 18, 0, 11, 3, 0, 4, 
    14, 31, 2, 6, 5, 19, 21, 2, 3, 0, 5, 0, 1, 0, 0, 
    27, 27, 1, 15, 55, 18, 0, 6, 0, 21, 19, 7, 11, 14, 0, 
    0, 1, 4, 0, 0, 0, 25, 12, 16, 24, 0, 0, 0, 10, 21, 
    7, 0, 0, 3, 0, 22, 0, 13, 1, 1, 0, 8, 8, 17, 6, 
    5, 18, 5, 22, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 6, 
    4, 0, 0, 13, 0, 0, 3, 12, 13, 0, 0, 0, 0, 13, 7, 
    0, 0, 7, 17, 0, 0, 22, 32, 0, 0, 0, 0, 12, 9, 0, 
    2, 0, 0, 42, 76, 25, 0, 0, 0, 14, 25, 27, 4, 0, 0, 
    0, 0, 11, 9, 0, 0, 0, 0, 0, 0, 0, 0, 7, 1, 1, 
    0, 0, 9, 0, 0, 3, 0, 0, 3, 7, 10, 9, 0, 0, 20, 
    0, 0, 0, 0, 0, 2, 9, 0, 0, 1, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 14, 0, 5, 28, 7, 1, 
    
    -- channel=232
    0, 0, 1, 0, 1, 0, 1, 4, 1, 0, 0, 0, 0, 1, 4, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 3, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=233
    18, 23, 24, 26, 24, 22, 25, 29, 26, 10, 0, 2, 12, 15, 15, 
    25, 28, 27, 27, 28, 48, 23, 13, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 25, 28, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 21, 28, 19, 8, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 12, 18, 27, 57, 16, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 21, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 17, 0, 14, 7, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 12, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 10, 13, 
    0, 0, 0, 15, 52, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=234
    0, 1, 0, 0, 0, 0, 0, 0, 0, 6, 7, 0, 0, 1, 4, 
    0, 0, 0, 2, 0, 0, 13, 7, 22, 0, 3, 7, 0, 0, 0, 
    27, 0, 0, 0, 0, 15, 33, 17, 0, 0, 14, 4, 27, 0, 0, 
    63, 0, 0, 0, 12, 0, 4, 7, 4, 0, 35, 9, 24, 17, 0, 
    41, 0, 21, 0, 0, 0, 35, 23, 24, 0, 4, 31, 0, 23, 0, 
    27, 0, 25, 4, 0, 3, 29, 20, 44, 0, 42, 42, 0, 11, 4, 
    11, 44, 5, 37, 0, 0, 25, 18, 49, 0, 52, 25, 0, 0, 12, 
    7, 26, 7, 16, 0, 0, 61, 20, 25, 0, 32, 38, 0, 0, 5, 
    22, 0, 54, 0, 2, 9, 20, 9, 0, 28, 2, 50, 0, 0, 0, 
    8, 0, 70, 0, 32, 0, 0, 13, 6, 16, 47, 2, 0, 0, 7, 
    0, 0, 70, 0, 36, 0, 0, 25, 45, 21, 0, 0, 0, 0, 13, 
    0, 0, 8, 0, 113, 54, 16, 15, 15, 1, 0, 0, 0, 0, 4, 
    14, 0, 0, 36, 89, 0, 6, 2, 2, 0, 0, 0, 2, 0, 0, 
    19, 0, 0, 90, 20, 0, 7, 2, 0, 0, 1, 4, 6, 0, 31, 
    25, 0, 1, 31, 16, 0, 2, 0, 0, 0, 10, 0, 0, 14, 38, 
    
    -- channel=235
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=236
    25, 25, 21, 23, 25, 19, 24, 31, 26, 29, 33, 26, 22, 23, 26, 
    20, 19, 22, 27, 20, 0, 28, 22, 56, 0, 0, 0, 10, 18, 21, 
    28, 35, 21, 27, 21, 49, 45, 36, 0, 0, 0, 9, 16, 9, 9, 
    35, 0, 20, 20, 15, 13, 0, 6, 2, 0, 25, 10, 23, 7, 0, 
    38, 0, 35, 1, 0, 0, 22, 8, 15, 0, 0, 15, 0, 13, 0, 
    32, 0, 37, 7, 0, 30, 0, 15, 12, 0, 28, 45, 0, 12, 0, 
    21, 0, 28, 40, 0, 0, 14, 14, 33, 0, 44, 9, 0, 0, 1, 
    0, 8, 11, 17, 0, 0, 69, 28, 24, 0, 26, 23, 0, 2, 28, 
    1, 0, 23, 0, 0, 47, 21, 0, 0, 29, 0, 65, 1, 0, 0, 
    1, 0, 33, 0, 11, 9, 0, 0, 0, 29, 65, 16, 0, 0, 29, 
    0, 0, 45, 0, 0, 0, 0, 28, 41, 22, 0, 0, 0, 0, 3, 
    0, 0, 15, 0, 78, 53, 7, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 95, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 58, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 29, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    
    -- channel=237
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 
    0, 0, 0, 0, 11, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 7, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    76, 0, 0, 0, 0, 0, 8, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 103, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 2, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=238
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 7, 0, 0, 4, 
    71, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 13, 0, 0, 8, 
    88, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 0, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 50, 0, 18, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 38, 0, 0, 16, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 0, 0, 10, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    
    -- channel=239
    11, 5, 7, 9, 10, 6, 8, 9, 11, 12, 10, 8, 8, 10, 12, 
    11, 6, 7, 8, 8, 0, 12, 6, 9, 11, 14, 16, 14, 12, 11, 
    8, 10, 9, 9, 10, 4, 11, 19, 16, 4, 6, 9, 15, 18, 7, 
    16, 14, 12, 9, 8, 12, 6, 12, 13, 5, 5, 10, 13, 18, 12, 
    11, 4, 13, 8, 0, 0, 1, 8, 12, 11, 6, 12, 11, 15, 19, 
    12, 0, 10, 7, 0, 0, 0, 10, 13, 0, 2, 12, 10, 13, 16, 
    11, 0, 12, 8, 0, 0, 0, 5, 10, 0, 7, 13, 14, 11, 13, 
    3, 0, 18, 12, 11, 0, 0, 5, 9, 0, 4, 14, 10, 7, 11, 
    0, 0, 12, 1, 12, 9, 11, 9, 11, 17, 7, 12, 12, 8, 8, 
    0, 0, 6, 5, 7, 10, 7, 1, 12, 3, 13, 17, 10, 8, 12, 
    0, 0, 8, 0, 0, 9, 0, 0, 7, 19, 21, 15, 16, 19, 22, 
    9, 0, 3, 0, 1, 17, 16, 16, 17, 18, 17, 16, 15, 16, 16, 
    22, 11, 2, 0, 15, 14, 14, 16, 18, 18, 18, 16, 14, 15, 14, 
    20, 18, 5, 0, 16, 15, 17, 16, 14, 14, 17, 16, 19, 15, 14, 
    17, 15, 17, 17, 22, 17, 15, 14, 13, 14, 17, 18, 13, 13, 21, 
    
    -- channel=240
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=241
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=242
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 9, 11, 0, 0, 0, 0, 0, 16, 0, 0, 
    45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 12, 11, 0, 
    10, 0, 0, 0, 0, 0, 10, 5, 19, 0, 0, 11, 0, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 16, 21, 0, 0, 0, 
    0, 28, 0, 21, 0, 0, 9, 0, 36, 0, 23, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 38, 6, 10, 0, 8, 19, 0, 0, 0, 
    0, 0, 21, 0, 0, 0, 0, 0, 0, 7, 0, 41, 0, 0, 0, 
    0, 0, 42, 0, 13, 0, 0, 0, 0, 13, 42, 0, 0, 0, 0, 
    0, 0, 42, 0, 0, 0, 0, 13, 30, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 89, 32, 4, 2, 4, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 16, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 80, 9, 0, 0, 0, 0, 0, 0, 1, 0, 0, 33, 
    16, 0, 0, 30, 13, 0, 3, 0, 0, 0, 3, 0, 0, 4, 30, 
    
    -- channel=243
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=244
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=245
    39, 39, 39, 38, 39, 37, 42, 43, 40, 38, 40, 38, 35, 37, 35, 
    37, 38, 40, 40, 36, 7, 43, 42, 47, 12, 5, 18, 29, 31, 33, 
    42, 38, 39, 40, 40, 38, 35, 28, 13, 0, 3, 4, 13, 26, 25, 
    12, 3, 36, 38, 36, 20, 3, 14, 8, 8, 12, 17, 11, 16, 21, 
    0, 0, 39, 24, 0, 21, 17, 14, 14, 1, 0, 15, 3, 7, 30, 
    20, 0, 38, 49, 4, 29, 0, 8, 5, 0, 20, 21, 5, 6, 9, 
    15, 0, 32, 34, 11, 0, 4, 10, 9, 0, 14, 9, 5, 0, 9, 
    11, 0, 22, 14, 12, 0, 31, 19, 9, 0, 10, 11, 5, 13, 21, 
    1, 0, 17, 0, 22, 28, 11, 0, 1, 25, 9, 31, 13, 6, 23, 
    0, 0, 2, 0, 9, 30, 4, 0, 20, 25, 28, 12, 1, 18, 36, 
    0, 0, 6, 0, 0, 0, 0, 8, 14, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 22, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=246
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=247
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=248
    34, 33, 32, 30, 29, 30, 35, 36, 29, 28, 30, 34, 28, 27, 26, 
    31, 32, 34, 31, 32, 5, 9, 25, 29, 12, 0, 0, 26, 37, 27, 
    23, 58, 33, 32, 36, 52, 8, 11, 8, 14, 0, 0, 0, 32, 37, 
    0, 31, 30, 32, 14, 17, 0, 0, 2, 45, 0, 11, 0, 5, 56, 
    0, 0, 6, 34, 0, 0, 0, 0, 4, 34, 0, 0, 1, 0, 31, 
    0, 4, 0, 24, 58, 1, 0, 0, 0, 51, 0, 0, 14, 0, 0, 
    0, 0, 26, 5, 49, 6, 0, 0, 0, 48, 0, 0, 3, 2, 0, 
    0, 0, 0, 0, 25, 32, 0, 12, 0, 43, 0, 0, 17, 17, 16, 
    0, 0, 0, 14, 0, 29, 0, 0, 13, 0, 32, 3, 27, 26, 24, 
    0, 0, 0, 9, 0, 2, 5, 0, 0, 24, 2, 12, 23, 30, 20, 
    17, 0, 0, 20, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 9, 0, 10, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 29, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=249
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=250
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=251
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 13, 4, 0, 
    8, 12, 0, 0, 0, 25, 8, 17, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 3, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 13, 
    0, 0, 0, 18, 39, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 29, 4, 0, 0, 0, 24, 13, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 4, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 0, 0, 0, 11, 36, 30, 27, 5, 0, 0, 0, 0, 0, 0, 
    0, 25, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 24, 4, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=252
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=253
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=254
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 2, 8, 0, 0, 
    11, 0, 0, 0, 0, 0, 14, 9, 3, 0, 0, 0, 0, 0, 0, 
    19, 26, 0, 0, 62, 38, 0, 0, 0, 0, 0, 11, 0, 12, 0, 
    0, 0, 0, 0, 0, 0, 11, 0, 12, 6, 0, 0, 0, 6, 14, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 2, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 3, 0, 0, 0, 0, 22, 0, 0, 0, 0, 9, 6, 0, 
    0, 0, 0, 2, 81, 48, 29, 0, 10, 3, 4, 32, 11, 0, 0, 
    0, 0, 2, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 8, 4, 0, 0, 9, 10, 0, 
    
    -- channel=255
    28, 32, 31, 31, 30, 30, 32, 36, 31, 22, 18, 20, 23, 27, 27, 
    30, 36, 33, 32, 31, 25, 23, 25, 17, 4, 0, 0, 8, 18, 24, 
    15, 22, 32, 34, 32, 27, 7, 6, 0, 0, 0, 0, 0, 4, 20, 
    0, 9, 27, 33, 23, 14, 1, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 15, 21, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 9, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 23, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 8, 0, 0, 0, 0, 3, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 7, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end gold_package;
