library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package inmem_package is
  type mem is array(0 to 4000000) of integer;

  constant input_mem : mem := (
    -- bias
    -397, 1301, -3042, 3806, -4800, -4379, -4224, -2063, 1200, 1395, 4454, 5171, -2890, -3671, -3224, -1145, -3536, -6192, -658, 222, 5085, 937, 919, 3182, -3213, 2796, -3730, 2439, 6655, -5784, -5038, -674, 2868, 4796, -894, 3888, -2801, 3200, -2791, -4402, 999, -2773, 931, -655, -4903, 2194, -3935, -102, 5819, 5494, -2015, 431, 1055, -3539, -1444, 5310, -846, -3780, -2406, -2883, -2554, 525, -513, 1192,

    -- weights
    -- filter=0 channel=0
    -11, 13, -5, -3, -3, 0, -2, -11, 8,
    -- filter=0 channel=1
    -7, 0, 7, -3, -7, 2, -1, 12, -11,
    -- filter=0 channel=2
    -6, -10, -10, 0, -8, -20, -10, 6, -12,
    -- filter=0 channel=3
    11, -7, -6, 0, -3, 0, -7, -4, -7,
    -- filter=0 channel=4
    8, 17, 0, 1, -2, 10, 5, -9, 7,
    -- filter=0 channel=5
    11, 5, 10, -16, -12, 10, 4, -15, -1,
    -- filter=0 channel=6
    -11, -2, -12, -4, -7, -8, -7, 0, -15,
    -- filter=0 channel=7
    -7, -6, 7, 8, -3, -13, 3, -11, 13,
    -- filter=0 channel=8
    20, 8, -11, -8, -10, -8, 14, 15, -2,
    -- filter=0 channel=9
    3, -3, -9, 5, 6, 4, 2, -17, 4,
    -- filter=0 channel=10
    -9, 2, -4, -7, 0, -12, -9, -7, 8,
    -- filter=0 channel=11
    -2, 0, 14, -7, 11, 2, 12, 6, -8,
    -- filter=0 channel=12
    0, -7, -10, 4, 14, 7, -7, -10, 13,
    -- filter=0 channel=13
    -5, -4, 5, -14, 3, -2, 12, -8, 0,
    -- filter=0 channel=14
    0, -6, 4, 0, 15, -3, 4, 8, 6,
    -- filter=0 channel=15
    12, -11, 0, 0, -13, 8, 7, -6, -10,
    -- filter=0 channel=16
    -5, 3, 9, 2, 4, 12, 9, -9, 4,
    -- filter=0 channel=17
    -3, 7, -4, -12, 4, -12, -3, 12, 5,
    -- filter=0 channel=18
    7, 9, -10, 9, 12, 8, 12, -12, -5,
    -- filter=0 channel=19
    -12, -5, -8, -7, -2, -6, -5, 1, 10,
    -- filter=0 channel=20
    -1, -1, -8, -16, -4, -9, -1, 2, -13,
    -- filter=0 channel=21
    -1, -9, -1, -3, 11, -12, -3, 6, 7,
    -- filter=0 channel=22
    14, 0, -9, 3, -13, 10, 0, -5, 13,
    -- filter=0 channel=23
    19, 15, -3, 19, 11, 11, 9, -5, -3,
    -- filter=0 channel=24
    -7, 7, -10, -7, -13, -6, 6, -2, 0,
    -- filter=0 channel=25
    2, 6, -4, -11, 0, -12, 7, -8, -14,
    -- filter=0 channel=26
    0, 9, -7, -13, -7, -15, -15, -3, 11,
    -- filter=0 channel=27
    12, 0, -14, 4, -6, -5, -11, 8, 13,
    -- filter=0 channel=28
    13, -5, -9, -8, -11, -10, 0, 10, 11,
    -- filter=0 channel=29
    2, 0, 0, 5, 0, 7, -14, 13, 12,
    -- filter=0 channel=30
    -10, -8, 12, -2, 3, 8, 8, -2, -14,
    -- filter=0 channel=31
    -10, 7, 2, 6, -8, 9, -11, -8, 12,
    -- filter=1 channel=0
    -5, 9, 9, 13, 10, 14, -8, 14, 4,
    -- filter=1 channel=1
    9, -10, -8, -2, 3, -7, 13, -13, -4,
    -- filter=1 channel=2
    0, 1, -4, -2, -12, -12, 10, 1, 2,
    -- filter=1 channel=3
    -3, 0, -9, -1, -8, -12, -3, -10, 10,
    -- filter=1 channel=4
    0, -5, -5, 4, -2, -13, -13, -14, -3,
    -- filter=1 channel=5
    10, -7, -6, -14, 0, -11, 3, 11, -11,
    -- filter=1 channel=6
    1, -12, 6, 14, -12, 5, -11, 0, 9,
    -- filter=1 channel=7
    -7, -2, -2, 2, 8, -2, 5, -10, 13,
    -- filter=1 channel=8
    8, 13, -4, 13, -4, 1, -1, 7, 2,
    -- filter=1 channel=9
    0, -6, 14, 10, -5, -6, -13, -1, 2,
    -- filter=1 channel=10
    6, 0, 2, 2, -4, -2, 7, 5, 13,
    -- filter=1 channel=11
    -1, -14, -2, 0, 8, 10, -12, -3, 1,
    -- filter=1 channel=12
    0, 8, -4, 0, 6, -13, 13, -4, 3,
    -- filter=1 channel=13
    8, -14, -5, 6, -14, 13, 0, -5, -1,
    -- filter=1 channel=14
    -11, -9, 5, -4, -14, -9, 0, -10, 10,
    -- filter=1 channel=15
    -3, -14, 4, 10, 2, -9, 14, -3, -10,
    -- filter=1 channel=16
    -4, 10, 0, -1, 6, -12, -14, -2, 4,
    -- filter=1 channel=17
    -3, -9, 2, -14, -11, 4, 11, 10, -10,
    -- filter=1 channel=18
    11, -7, 1, 11, 13, 4, 10, 11, 5,
    -- filter=1 channel=19
    -12, 12, 8, 12, -4, 0, -1, -6, -10,
    -- filter=1 channel=20
    -11, 2, -5, -5, 3, -2, 8, -11, 14,
    -- filter=1 channel=21
    2, 10, -12, -10, 3, -9, 5, 1, -12,
    -- filter=1 channel=22
    -1, -3, -10, 10, 5, -5, 11, -13, -13,
    -- filter=1 channel=23
    12, -6, 2, -13, 2, -3, -14, -4, -8,
    -- filter=1 channel=24
    8, -4, -8, -5, -9, -8, -1, 2, 12,
    -- filter=1 channel=25
    -5, -7, 7, 6, 1, -7, 11, -4, -9,
    -- filter=1 channel=26
    -11, -8, -10, -11, -7, -10, 8, 13, 0,
    -- filter=1 channel=27
    13, -7, 4, 5, 14, 9, 2, -13, -9,
    -- filter=1 channel=28
    -13, 12, 15, -13, 8, 14, -7, -9, 10,
    -- filter=1 channel=29
    14, 12, 8, 4, 12, -5, 7, 7, 7,
    -- filter=1 channel=30
    8, -7, 9, 10, 6, 0, -11, -6, 10,
    -- filter=1 channel=31
    8, 14, -14, 14, -9, 12, 12, 3, 0,
    -- filter=2 channel=0
    -3, 3, 8, 5, -12, -7, 13, 9, 2,
    -- filter=2 channel=1
    13, -10, 6, -10, 7, -3, 9, -5, -7,
    -- filter=2 channel=2
    5, -2, -10, 5, -13, -14, -12, -1, 10,
    -- filter=2 channel=3
    -10, -7, -5, 6, 10, -8, -5, 11, -5,
    -- filter=2 channel=4
    3, 2, -4, 3, -4, -9, 7, -13, -11,
    -- filter=2 channel=5
    -11, 2, 6, 0, 13, 5, -4, 2, -13,
    -- filter=2 channel=6
    16, 4, -4, 3, -5, 8, 10, 10, 11,
    -- filter=2 channel=7
    2, 1, -7, -2, -11, -3, 7, 8, 3,
    -- filter=2 channel=8
    13, 2, -2, -6, 11, 9, -4, 0, 10,
    -- filter=2 channel=9
    -2, -14, 12, -11, 0, -7, -6, -15, 3,
    -- filter=2 channel=10
    -2, -5, -13, 4, 10, 4, -2, -12, -5,
    -- filter=2 channel=11
    0, 13, -1, 5, -8, -5, 5, -2, 11,
    -- filter=2 channel=12
    16, 0, 11, -14, -6, -7, 7, 11, 0,
    -- filter=2 channel=13
    16, -11, 0, 3, 14, 9, 8, 1, 1,
    -- filter=2 channel=14
    14, -4, 8, 7, 10, -2, 9, -7, -12,
    -- filter=2 channel=15
    -14, 5, 9, 11, -11, 5, 10, -1, -2,
    -- filter=2 channel=16
    -3, -1, -11, 0, 2, -1, 2, -3, -14,
    -- filter=2 channel=17
    4, 13, 13, 14, -14, -2, -3, -8, -14,
    -- filter=2 channel=18
    -10, -13, -10, 9, -13, 0, 14, 9, 13,
    -- filter=2 channel=19
    14, -6, 0, 13, -6, -4, -8, -3, -14,
    -- filter=2 channel=20
    14, -7, 7, -8, 11, -13, 13, -1, 11,
    -- filter=2 channel=21
    -2, -1, -3, -2, 1, -3, -10, -5, 10,
    -- filter=2 channel=22
    -4, -12, -4, -13, -14, 6, -6, -10, 7,
    -- filter=2 channel=23
    -9, 5, -14, 7, -16, -10, 4, -2, 9,
    -- filter=2 channel=24
    -6, 2, 11, 14, 0, 0, 5, -5, 5,
    -- filter=2 channel=25
    13, -6, -6, -3, 10, 11, 0, -1, -12,
    -- filter=2 channel=26
    0, 1, 13, 5, 8, -6, 10, 2, -1,
    -- filter=2 channel=27
    11, 4, -6, 0, -1, -10, 8, -10, 5,
    -- filter=2 channel=28
    3, -14, -10, -4, 13, -14, 11, -10, 14,
    -- filter=2 channel=29
    -12, -1, 7, -4, 4, -12, -9, 9, -2,
    -- filter=2 channel=30
    7, 14, 0, 8, 13, -6, 7, -10, -11,
    -- filter=2 channel=31
    -12, 6, 2, 5, 9, 10, 13, 4, 8,
    -- filter=3 channel=0
    11, -5, 13, 13, -5, -3, -9, -1, -1,
    -- filter=3 channel=1
    -3, 1, -6, -8, -1, -8, -11, 8, 8,
    -- filter=3 channel=2
    -36, -18, 21, -38, -3, 16, -6, 5, 9,
    -- filter=3 channel=3
    -10, -12, 14, 2, 7, 2, 14, -4, -6,
    -- filter=3 channel=4
    -15, 0, 13, -21, 11, 21, 7, -5, 18,
    -- filter=3 channel=5
    13, 17, 20, 5, 16, 19, -12, -8, -10,
    -- filter=3 channel=6
    -15, 8, 20, -17, -9, 0, -5, -9, 13,
    -- filter=3 channel=7
    -22, -6, 19, -22, -16, 0, -17, 1, -7,
    -- filter=3 channel=8
    4, 11, 8, -3, -7, 20, 13, 13, 9,
    -- filter=3 channel=9
    -15, -3, 19, -23, -13, 2, 0, -7, 13,
    -- filter=3 channel=10
    -3, 1, -11, -11, 3, -12, -4, 0, -11,
    -- filter=3 channel=11
    -12, -2, 10, -13, 10, 0, 1, -12, 3,
    -- filter=3 channel=12
    -5, -11, 14, 4, 15, -3, -3, -8, 0,
    -- filter=3 channel=13
    -16, -9, -7, 0, 9, 1, -4, 4, -10,
    -- filter=3 channel=14
    -22, 7, 17, -6, 15, 9, -8, 8, 6,
    -- filter=3 channel=15
    14, 12, -12, -13, -14, 0, -2, 1, -4,
    -- filter=3 channel=16
    4, -5, 22, -10, -7, 20, 16, 2, 9,
    -- filter=3 channel=17
    5, -14, 8, -8, 0, 23, -13, -10, 2,
    -- filter=3 channel=18
    2, 1, 9, 0, 16, 1, 10, -3, -8,
    -- filter=3 channel=19
    0, 21, 21, 15, 20, 17, 17, 1, 20,
    -- filter=3 channel=20
    4, 6, 18, 0, 0, 12, -7, -6, -4,
    -- filter=3 channel=21
    -17, -6, 9, -16, -7, 12, -11, -10, -10,
    -- filter=3 channel=22
    -15, 0, 3, -11, -2, 0, 2, -9, 15,
    -- filter=3 channel=23
    -27, -1, 33, -15, -2, 15, -11, 14, 3,
    -- filter=3 channel=24
    -28, 4, 22, -1, -3, -5, 7, 2, 7,
    -- filter=3 channel=25
    -9, 7, 3, -7, 5, 9, -12, 10, -13,
    -- filter=3 channel=26
    -2, -20, 9, 6, 5, -8, 10, 0, 0,
    -- filter=3 channel=27
    -9, -14, 12, 9, 9, -6, -10, 4, 11,
    -- filter=3 channel=28
    -13, 7, 1, 10, 9, -10, -5, 14, 19,
    -- filter=3 channel=29
    -8, 9, -8, 4, 11, -4, 5, 0, -7,
    -- filter=3 channel=30
    5, 6, 7, -7, 3, -1, 3, -9, -15,
    -- filter=3 channel=31
    8, -11, 14, -14, 12, -9, 0, 10, 11,
    -- filter=4 channel=0
    -5, 3, -6, 3, -14, -3, 0, -1, 3,
    -- filter=4 channel=1
    0, -4, -13, -1, 3, 5, -11, -14, -12,
    -- filter=4 channel=2
    18, 9, -4, 4, 17, -13, -3, 15, 3,
    -- filter=4 channel=3
    -15, -13, -9, 9, -16, 1, -10, -16, 5,
    -- filter=4 channel=4
    -8, -11, 13, 1, 7, 18, 3, 4, -1,
    -- filter=4 channel=5
    -15, 5, -10, 9, -5, -9, -2, -11, 4,
    -- filter=4 channel=6
    -5, -3, -11, 4, 4, -8, -2, 8, 6,
    -- filter=4 channel=7
    12, -3, -6, -5, -12, -15, -6, 6, 5,
    -- filter=4 channel=8
    1, -5, 6, -7, 11, 7, 14, 19, 13,
    -- filter=4 channel=9
    17, 7, -7, 3, 10, 5, 13, -13, -12,
    -- filter=4 channel=10
    5, 7, -3, 0, 0, 9, -4, -4, 3,
    -- filter=4 channel=11
    -1, 6, 11, 5, 7, -4, -14, -2, -14,
    -- filter=4 channel=12
    -3, 4, 0, 1, -10, 15, 1, 1, -6,
    -- filter=4 channel=13
    13, 0, 0, -14, 3, 8, -6, -2, -8,
    -- filter=4 channel=14
    -14, 14, 9, -20, 13, 15, -1, -1, 3,
    -- filter=4 channel=15
    11, 7, -8, 14, -13, -14, -1, 2, 0,
    -- filter=4 channel=16
    -13, -8, -8, -8, 0, 7, -12, 0, 1,
    -- filter=4 channel=17
    5, -4, 9, -12, -12, -12, -18, -15, -8,
    -- filter=4 channel=18
    0, -1, -6, 8, 9, -6, 5, 3, 11,
    -- filter=4 channel=19
    -3, -21, -10, -25, -7, 10, -19, -3, -2,
    -- filter=4 channel=20
    -1, 10, 2, 12, -6, -2, -15, -6, 7,
    -- filter=4 channel=21
    13, 9, -11, -2, 0, -9, -12, 9, 2,
    -- filter=4 channel=22
    0, 3, -12, -13, -8, 8, -12, 0, 1,
    -- filter=4 channel=23
    12, 5, 3, -12, 17, 22, -7, 10, 16,
    -- filter=4 channel=24
    5, -6, -10, -13, 0, 7, 3, -1, 5,
    -- filter=4 channel=25
    2, 12, 6, 4, -12, 2, -6, -5, -5,
    -- filter=4 channel=26
    10, 1, -11, -17, -12, -17, -12, -15, -14,
    -- filter=4 channel=27
    0, -4, 0, 12, 2, -9, -15, -4, 1,
    -- filter=4 channel=28
    3, 1, 9, -14, 12, 4, -12, 4, -3,
    -- filter=4 channel=29
    -10, 2, 5, 0, -7, -12, 3, -6, -4,
    -- filter=4 channel=30
    4, 7, 1, 11, -11, 4, -11, 7, 1,
    -- filter=4 channel=31
    0, 0, 11, -2, -1, -1, 2, 8, 14,
    -- filter=5 channel=0
    -1, -5, 0, 10, 5, 8, 3, 12, -11,
    -- filter=5 channel=1
    -3, -2, -13, 2, -2, -7, -14, -8, 0,
    -- filter=5 channel=2
    -14, -9, -11, 4, -15, -4, 3, 3, -12,
    -- filter=5 channel=3
    0, 2, 2, -3, 10, 2, 0, -9, -14,
    -- filter=5 channel=4
    -8, 2, -14, -3, -9, -10, 4, 9, 10,
    -- filter=5 channel=5
    -3, 9, 7, 13, -5, 1, 1, 2, -12,
    -- filter=5 channel=6
    10, 8, -4, -2, 11, 0, 0, 1, 0,
    -- filter=5 channel=7
    -3, 9, 3, -12, 12, -4, 7, -15, -11,
    -- filter=5 channel=8
    5, -12, -8, 13, 5, -2, -13, 14, 12,
    -- filter=5 channel=9
    11, 4, -7, -4, 8, -5, 9, 6, 13,
    -- filter=5 channel=10
    13, -10, 4, -11, 0, 13, 6, 3, -12,
    -- filter=5 channel=11
    8, -11, 11, 5, 8, -12, 0, -4, -7,
    -- filter=5 channel=12
    -11, 13, 6, -6, 12, -4, 9, 2, 0,
    -- filter=5 channel=13
    -6, -4, 9, 8, 2, 10, -7, -8, 14,
    -- filter=5 channel=14
    -14, 1, -14, 4, 7, -5, -3, 11, -7,
    -- filter=5 channel=15
    3, 0, -2, 0, 0, 13, 2, -11, -6,
    -- filter=5 channel=16
    10, -10, -5, -6, -13, 3, -9, 1, -10,
    -- filter=5 channel=17
    -3, -1, 14, 11, -14, -3, 7, -9, -14,
    -- filter=5 channel=18
    6, -6, -10, -6, -8, 11, 5, 0, 7,
    -- filter=5 channel=19
    -3, -10, 13, 8, 3, -9, -7, 0, -14,
    -- filter=5 channel=20
    -11, -12, -2, -7, 3, -1, -2, -15, 8,
    -- filter=5 channel=21
    -7, -8, -8, 6, -3, 9, -13, -5, -7,
    -- filter=5 channel=22
    -12, 0, -7, -9, -6, 7, 3, -12, -7,
    -- filter=5 channel=23
    -8, 5, -4, 16, 8, 15, -5, -13, 4,
    -- filter=5 channel=24
    7, -13, -8, 4, 8, -7, 13, 3, -9,
    -- filter=5 channel=25
    2, 1, 0, 8, 2, -8, 0, 11, 14,
    -- filter=5 channel=26
    9, -3, 12, -14, -15, 13, -4, -9, -10,
    -- filter=5 channel=27
    9, -7, -13, 5, 0, 2, 0, 6, 8,
    -- filter=5 channel=28
    9, -14, 12, 13, 11, 13, -7, 0, -14,
    -- filter=5 channel=29
    -11, -14, -5, 0, 6, -12, -9, -7, 1,
    -- filter=5 channel=30
    -11, -11, 2, 14, 8, 0, 10, -7, -5,
    -- filter=5 channel=31
    -3, 5, 0, 3, 13, 14, -3, 14, 10,
    -- filter=6 channel=0
    2, -13, -4, 12, 13, -4, 13, -15, 5,
    -- filter=6 channel=1
    7, 3, 9, -2, 0, -12, -9, 5, -14,
    -- filter=6 channel=2
    -26, -1, -3, 0, -4, -10, 33, 37, 35,
    -- filter=6 channel=3
    -7, 3, 6, -4, -2, -7, 10, 5, -8,
    -- filter=6 channel=4
    -22, 0, 8, -22, -26, -24, 8, -18, -9,
    -- filter=6 channel=5
    6, -5, -10, 0, 11, 3, -11, 8, 9,
    -- filter=6 channel=6
    -9, -13, -5, 5, 3, 1, 21, 11, 7,
    -- filter=6 channel=7
    -23, -10, -7, 13, -9, 12, 0, 20, 31,
    -- filter=6 channel=8
    1, -5, -6, -3, -15, -6, -4, -5, -11,
    -- filter=6 channel=9
    -22, 0, 5, 1, 2, -16, 13, 3, 12,
    -- filter=6 channel=10
    11, -5, 14, 8, 6, 7, 16, -3, 19,
    -- filter=6 channel=11
    -10, 4, 3, 2, -15, -6, -4, 0, 14,
    -- filter=6 channel=12
    11, -19, -5, -16, -15, 1, 17, -8, -5,
    -- filter=6 channel=13
    -10, 1, 3, 12, 4, 14, 3, 12, 12,
    -- filter=6 channel=14
    -5, -9, -11, 0, -20, -12, 4, 0, -7,
    -- filter=6 channel=15
    -10, -10, -7, 11, -5, -3, -7, -9, 6,
    -- filter=6 channel=16
    10, 0, -8, 16, 3, 7, 4, 5, 0,
    -- filter=6 channel=17
    3, -7, 4, 17, -5, 0, 29, 20, 20,
    -- filter=6 channel=18
    3, -7, -11, 13, -2, 7, 6, 10, -8,
    -- filter=6 channel=19
    9, 2, 6, 14, 3, -18, -9, 5, 4,
    -- filter=6 channel=20
    -17, 11, 2, 11, -7, 4, 18, 12, 19,
    -- filter=6 channel=21
    -3, 10, 5, -8, -2, 20, 24, 1, 15,
    -- filter=6 channel=22
    10, -17, 6, 11, 5, 5, 11, -16, -11,
    -- filter=6 channel=23
    -1, -9, -3, -15, -28, -11, -6, 0, -10,
    -- filter=6 channel=24
    -10, -7, 3, -9, -7, 4, 18, 20, 24,
    -- filter=6 channel=25
    9, 5, 6, 11, 4, 13, -12, 10, 0,
    -- filter=6 channel=26
    -18, 6, -1, -7, 13, -5, 7, 3, 16,
    -- filter=6 channel=27
    10, -2, 11, 5, -6, 11, 0, 12, 14,
    -- filter=6 channel=28
    16, 2, -6, 5, 9, 13, -7, -5, 4,
    -- filter=6 channel=29
    8, 6, -14, 12, 3, -12, 11, 0, -7,
    -- filter=6 channel=30
    9, 0, -9, -5, -1, 10, -4, 15, 1,
    -- filter=6 channel=31
    -6, 0, -9, 10, -11, -13, -12, -4, 9,
    -- filter=7 channel=0
    2, 5, 8, 10, 1, -6, -10, -2, -13,
    -- filter=7 channel=1
    -10, -13, 7, 8, 7, 14, -8, -3, -13,
    -- filter=7 channel=2
    -14, 25, 23, 9, -4, -2, -9, -8, -23,
    -- filter=7 channel=3
    9, 2, -12, -14, 5, -9, 10, -9, 13,
    -- filter=7 channel=4
    12, 17, 0, 8, 9, 13, -14, -13, 4,
    -- filter=7 channel=5
    14, 16, 4, -11, -9, -6, 3, 3, 10,
    -- filter=7 channel=6
    11, -1, -4, -5, -7, -8, -6, 9, 2,
    -- filter=7 channel=7
    -1, 13, 1, 0, -10, 4, 12, -17, 0,
    -- filter=7 channel=8
    -6, -10, 15, 6, 16, 3, 0, -3, 3,
    -- filter=7 channel=9
    -9, 1, 19, 2, 0, -12, -4, -9, -13,
    -- filter=7 channel=10
    -13, 4, -9, 10, 9, 8, -11, 0, 3,
    -- filter=7 channel=11
    2, 3, -1, 6, 4, 14, 10, -5, -2,
    -- filter=7 channel=12
    -11, 10, -11, -1, -6, -5, -12, 7, -5,
    -- filter=7 channel=13
    -9, -10, -9, 14, 2, -11, 1, -14, -15,
    -- filter=7 channel=14
    -7, 13, -7, 14, -6, 0, -9, -11, 3,
    -- filter=7 channel=15
    0, -7, -14, -7, 1, -5, -10, 1, 2,
    -- filter=7 channel=16
    9, -10, 0, 3, 9, 12, -10, -16, -17,
    -- filter=7 channel=17
    4, -5, -1, 9, -2, 10, 14, 3, 0,
    -- filter=7 channel=18
    13, 4, -10, -4, 0, 10, -14, -13, -1,
    -- filter=7 channel=19
    -10, 3, -9, -7, -10, -3, -7, -11, -6,
    -- filter=7 channel=20
    5, 10, 9, -4, -2, 13, -13, -6, 7,
    -- filter=7 channel=21
    -16, 9, 7, -1, 11, -13, 8, -8, -16,
    -- filter=7 channel=22
    -8, -7, 15, -12, -7, 7, -2, 15, -12,
    -- filter=7 channel=23
    -5, -4, -6, 8, 14, 15, -17, 0, -1,
    -- filter=7 channel=24
    8, 13, -4, 10, -2, 12, 11, -5, -14,
    -- filter=7 channel=25
    13, -9, 3, 6, -4, -5, -4, 13, 9,
    -- filter=7 channel=26
    0, -9, 9, 11, 2, 5, -4, -3, -4,
    -- filter=7 channel=27
    0, 13, 7, -13, -1, -13, -1, 10, -4,
    -- filter=7 channel=28
    -6, -6, 4, 10, 7, 5, -4, 10, 13,
    -- filter=7 channel=29
    13, 7, 9, -6, 1, 9, 0, -2, 2,
    -- filter=7 channel=30
    6, 3, -8, -8, 13, -2, 7, 8, -2,
    -- filter=7 channel=31
    -4, 5, 11, 7, -9, 12, -3, 8, -7,
    -- filter=8 channel=0
    0, 12, 15, -14, 8, -2, -7, -8, -1,
    -- filter=8 channel=1
    -3, 4, 5, 15, 3, -12, 8, 3, 10,
    -- filter=8 channel=2
    -13, -7, -19, -12, 0, -23, 6, -17, -7,
    -- filter=8 channel=3
    -4, 6, -5, 11, 11, 0, -7, -2, 10,
    -- filter=8 channel=4
    20, -1, 10, 6, 8, 6, 10, -3, 0,
    -- filter=8 channel=5
    -5, -7, -16, 4, -14, -10, -1, -13, -14,
    -- filter=8 channel=6
    -6, -12, 9, -6, -10, 11, -9, 13, 8,
    -- filter=8 channel=7
    3, 8, -10, 1, -19, 3, -3, -11, -15,
    -- filter=8 channel=8
    1, 14, -5, 9, 1, -8, 14, -6, 8,
    -- filter=8 channel=9
    0, 0, -10, 9, -17, -19, -17, -1, -2,
    -- filter=8 channel=10
    -15, -5, -11, 1, -11, -6, -6, -13, -9,
    -- filter=8 channel=11
    -10, 0, -13, -8, 9, 8, 4, 2, 8,
    -- filter=8 channel=12
    14, 18, 11, 5, 2, -1, -10, -9, 6,
    -- filter=8 channel=13
    8, -10, 4, -16, -1, -12, 9, -18, 0,
    -- filter=8 channel=14
    21, 8, 16, 7, 15, 5, 13, -7, 19,
    -- filter=8 channel=15
    11, -2, -9, -11, 14, 13, 0, -5, -8,
    -- filter=8 channel=16
    -4, 6, -13, 3, 3, 8, 11, -10, 3,
    -- filter=8 channel=17
    14, 19, 10, -10, -4, 0, -6, -13, 12,
    -- filter=8 channel=18
    13, 12, 1, -7, 8, -4, -13, 15, 12,
    -- filter=8 channel=19
    -8, 17, -7, 4, 18, -2, 9, 14, -4,
    -- filter=8 channel=20
    10, 11, 3, -6, -11, -2, 0, 1, -3,
    -- filter=8 channel=21
    -8, 9, -10, -8, -10, 5, 11, 3, -1,
    -- filter=8 channel=22
    -5, 2, 2, 4, 0, 11, 11, -2, -3,
    -- filter=8 channel=23
    16, 21, -4, -3, -4, 10, 13, 11, 1,
    -- filter=8 channel=24
    -6, -13, -6, -3, -4, -23, -10, 5, -15,
    -- filter=8 channel=25
    8, 5, 1, -5, 12, -12, 12, -10, -8,
    -- filter=8 channel=26
    -3, -13, -4, 5, 3, -18, 7, -4, 2,
    -- filter=8 channel=27
    -2, 0, -6, 14, -7, -6, -9, 5, 14,
    -- filter=8 channel=28
    5, -8, -1, -8, 13, -7, -10, -7, 7,
    -- filter=8 channel=29
    -2, 5, -1, -3, 4, 7, 1, 4, 6,
    -- filter=8 channel=30
    10, 13, 5, 8, -11, 14, -10, 9, -14,
    -- filter=8 channel=31
    5, -7, -13, 9, -2, 13, -4, -8, -6,
    -- filter=9 channel=0
    6, -10, -13, -5, 11, 14, -1, 3, 9,
    -- filter=9 channel=1
    6, -8, 8, -11, 2, -5, 0, -8, 10,
    -- filter=9 channel=2
    -19, -46, -37, -4, -17, 6, 23, 38, 33,
    -- filter=9 channel=3
    -13, -9, -8, -1, -3, 11, 3, 0, -14,
    -- filter=9 channel=4
    6, -10, -9, -6, -7, -17, 1, 3, 10,
    -- filter=9 channel=5
    -13, -3, -6, -4, 0, -4, -6, -5, -11,
    -- filter=9 channel=6
    14, 4, -20, -15, 13, 12, 3, -7, 3,
    -- filter=9 channel=7
    -14, -19, -20, -10, -15, 6, -5, 4, 30,
    -- filter=9 channel=8
    1, 1, 2, 1, -19, -2, 4, 0, -1,
    -- filter=9 channel=9
    5, -15, -29, -4, -7, 13, 4, 27, 24,
    -- filter=9 channel=10
    4, -4, -5, -13, -14, 8, 1, -1, 17,
    -- filter=9 channel=11
    8, 13, -12, -9, 1, -2, -2, -9, 11,
    -- filter=9 channel=12
    4, -17, -5, 15, 3, 3, -2, -1, 23,
    -- filter=9 channel=13
    3, 0, -11, -2, 0, 17, 5, 8, 25,
    -- filter=9 channel=14
    0, -18, -5, 14, 0, -3, 5, 4, 22,
    -- filter=9 channel=15
    9, 2, 7, -7, -3, 10, 5, -14, 8,
    -- filter=9 channel=16
    0, -6, -9, -13, 16, 0, 8, 22, 0,
    -- filter=9 channel=17
    9, -7, -17, 8, -11, 0, 12, 22, 1,
    -- filter=9 channel=18
    12, 8, -13, 4, -2, 15, -4, 13, -8,
    -- filter=9 channel=19
    3, 15, -3, -10, -9, 15, 2, -14, 9,
    -- filter=9 channel=20
    -3, -16, -15, 0, 7, -6, 3, 7, 13,
    -- filter=9 channel=21
    -19, -7, 4, 0, 4, -3, 7, 11, 22,
    -- filter=9 channel=22
    6, -8, 3, -9, -6, 8, 0, 5, 9,
    -- filter=9 channel=23
    -13, -1, -11, -6, -15, -19, 3, 15, 19,
    -- filter=9 channel=24
    4, -15, -16, -16, -12, 20, 21, 23, 26,
    -- filter=9 channel=25
    6, -1, 0, -11, -10, 1, 5, -10, 12,
    -- filter=9 channel=26
    -11, 2, -19, -18, 3, -9, 15, 19, 27,
    -- filter=9 channel=27
    -1, -6, -8, 14, 12, -1, 8, 9, -4,
    -- filter=9 channel=28
    -11, 0, -2, -10, 8, -13, 1, 14, 14,
    -- filter=9 channel=29
    -3, -13, 0, 13, 11, 8, 6, 5, -4,
    -- filter=9 channel=30
    -7, -11, -4, 10, 12, -11, 12, -4, 13,
    -- filter=9 channel=31
    12, 4, 7, -13, -12, 0, -2, -13, 7,
    -- filter=10 channel=0
    6, -5, -2, 9, -12, 0, 5, 5, -13,
    -- filter=10 channel=1
    7, 4, 10, 1, 2, -4, 4, 0, -10,
    -- filter=10 channel=2
    -2, 4, 8, 15, 12, 2, 12, 0, 20,
    -- filter=10 channel=3
    -7, -5, 6, -2, -20, 0, -9, -19, 7,
    -- filter=10 channel=4
    4, 6, 31, 15, 19, 14, -14, 8, 33,
    -- filter=10 channel=5
    -21, 4, -20, -7, -6, -7, -8, 7, 2,
    -- filter=10 channel=6
    -15, -25, 0, -18, -7, 4, -24, 5, 14,
    -- filter=10 channel=7
    1, -1, -17, -20, 7, -7, -17, -7, -5,
    -- filter=10 channel=8
    -2, 21, 29, -4, 4, 17, -10, 6, 31,
    -- filter=10 channel=9
    10, 2, -4, 11, 10, -11, -3, 12, -3,
    -- filter=10 channel=10
    -9, -14, -24, -17, -18, -2, -7, -3, -6,
    -- filter=10 channel=11
    0, -15, -4, -11, -8, 5, -12, -6, 10,
    -- filter=10 channel=12
    -1, 6, -1, -3, -7, 17, -6, -3, 16,
    -- filter=10 channel=13
    -13, 6, -14, 8, 1, -5, -14, 0, 4,
    -- filter=10 channel=14
    -13, 21, 25, 10, 10, 5, -6, 7, 26,
    -- filter=10 channel=15
    13, 2, 6, 6, 0, 2, -14, -9, 8,
    -- filter=10 channel=16
    -19, -2, 16, -8, -18, 12, 4, -3, -2,
    -- filter=10 channel=17
    -30, -8, 4, -14, -21, 4, -31, -3, 1,
    -- filter=10 channel=18
    -7, -1, -6, -10, -12, -13, 7, -3, 5,
    -- filter=10 channel=19
    -31, -9, -19, -20, -32, -1, -18, -26, -12,
    -- filter=10 channel=20
    -15, -18, -11, -2, -19, -19, -6, -15, 4,
    -- filter=10 channel=21
    -3, -2, -22, 4, -17, -9, -14, 2, -18,
    -- filter=10 channel=22
    -4, 6, 8, -10, 10, 4, 2, 6, 10,
    -- filter=10 channel=23
    16, 17, 36, 14, 27, 27, 4, 37, 22,
    -- filter=10 channel=24
    -4, -11, -20, 6, -18, -2, 3, 10, -7,
    -- filter=10 channel=25
    -11, -1, 4, 4, -12, -9, -3, 7, -2,
    -- filter=10 channel=26
    -8, -10, -20, -19, -11, -10, -3, -18, -16,
    -- filter=10 channel=27
    11, 3, -14, -16, -5, 9, -5, 0, 3,
    -- filter=10 channel=28
    -20, 3, 0, -1, -11, -13, -4, -13, 6,
    -- filter=10 channel=29
    -9, -8, -7, 3, 9, 7, 8, 10, -9,
    -- filter=10 channel=30
    -23, -19, -6, -9, 0, 5, -4, -21, -17,
    -- filter=10 channel=31
    6, -9, -1, -14, 4, -6, 11, -10, 8,
    -- filter=11 channel=0
    4, -7, 5, 14, 6, 5, 6, 6, -12,
    -- filter=11 channel=1
    11, -6, 4, 0, -7, -7, 7, 11, -4,
    -- filter=11 channel=2
    17, -20, -14, 12, 0, -33, 26, -2, -35,
    -- filter=11 channel=3
    13, 0, 11, 2, -6, 5, 16, -1, 13,
    -- filter=11 channel=4
    0, -13, -5, 3, -7, 9, 25, -8, -12,
    -- filter=11 channel=5
    4, -4, 12, 1, 8, 4, -6, -6, -13,
    -- filter=11 channel=6
    4, 0, 11, 14, -1, 9, 19, 3, 0,
    -- filter=11 channel=7
    0, -11, 0, 20, -4, -3, 23, 2, -21,
    -- filter=11 channel=8
    5, 5, 3, -1, -11, -18, 12, 0, 7,
    -- filter=11 channel=9
    4, -20, 7, 0, -11, 0, 12, -17, -24,
    -- filter=11 channel=10
    17, 5, -7, 3, -12, 2, -1, 0, -9,
    -- filter=11 channel=11
    6, -8, 3, 6, -2, 9, 11, -4, -6,
    -- filter=11 channel=12
    6, 11, -5, 20, -11, -5, 7, 16, -12,
    -- filter=11 channel=13
    13, 9, -14, 5, 2, -12, 7, -1, 3,
    -- filter=11 channel=14
    -3, -10, 9, 20, -6, 3, 14, 3, -4,
    -- filter=11 channel=15
    10, -1, 0, 0, -9, 10, -3, 7, -11,
    -- filter=11 channel=16
    -4, -5, -3, 11, 1, -8, -3, -9, 6,
    -- filter=11 channel=17
    1, -5, 6, 32, 13, 10, 29, 15, 15,
    -- filter=11 channel=18
    -9, 6, -9, 4, -13, -4, 9, 3, -11,
    -- filter=11 channel=19
    0, 4, 21, 24, 10, 4, 29, 2, 16,
    -- filter=11 channel=20
    -9, 2, 0, -6, 13, -17, 13, 3, -8,
    -- filter=11 channel=21
    14, -8, -19, 10, 0, -12, -9, -17, 6,
    -- filter=11 channel=22
    -8, -5, -9, 6, 3, -3, -8, 9, -14,
    -- filter=11 channel=23
    -16, -17, -11, -3, -16, -20, 15, -1, -1,
    -- filter=11 channel=24
    14, -4, -6, -1, -12, -26, 8, -11, 3,
    -- filter=11 channel=25
    -9, 3, 8, -8, -6, -5, 11, -13, -7,
    -- filter=11 channel=26
    -6, -8, -7, 19, -7, -10, 19, 14, -4,
    -- filter=11 channel=27
    -1, 8, -9, -9, -4, 12, 14, 12, 13,
    -- filter=11 channel=28
    0, -6, -2, 4, 14, -4, -8, 17, -3,
    -- filter=11 channel=29
    -4, -4, -8, -3, 7, 6, 7, -1, -13,
    -- filter=11 channel=30
    11, -6, -6, 2, 10, 8, -5, 13, 4,
    -- filter=11 channel=31
    -12, -10, -11, -7, 9, -14, 9, 11, -12,
    -- filter=12 channel=0
    0, 11, 3, 10, 14, 6, -10, 4, -5,
    -- filter=12 channel=1
    -7, 10, 6, 5, -10, 1, 10, -6, -5,
    -- filter=12 channel=2
    -1, 7, -1, -8, -2, 6, -10, 7, -6,
    -- filter=12 channel=3
    3, -6, -11, -4, -3, 14, -3, 1, -3,
    -- filter=12 channel=4
    -2, 14, 8, -5, 7, 8, 2, -13, -13,
    -- filter=12 channel=5
    9, 0, -11, 0, -1, 8, -11, 1, 4,
    -- filter=12 channel=6
    10, -4, 13, 6, 0, 5, -5, 12, 1,
    -- filter=12 channel=7
    -2, 0, -2, -14, -6, 11, 2, -9, -5,
    -- filter=12 channel=8
    -11, -14, 7, -1, 3, 11, 12, -14, 0,
    -- filter=12 channel=9
    2, -8, 4, 3, -7, 4, -15, -5, 11,
    -- filter=12 channel=10
    -9, -1, 0, 0, 1, 7, 8, 3, 10,
    -- filter=12 channel=11
    9, -4, -11, 4, 10, -5, -12, 2, -7,
    -- filter=12 channel=12
    13, 9, -1, 8, 2, -11, -8, -8, 0,
    -- filter=12 channel=13
    3, 2, 0, 0, -17, -14, -5, -4, -8,
    -- filter=12 channel=14
    -7, -10, -3, 1, -6, 11, 5, 8, 5,
    -- filter=12 channel=15
    -9, -11, 14, -6, 9, 12, 11, 1, -14,
    -- filter=12 channel=16
    -10, -5, 2, 5, 2, 9, 5, -9, -1,
    -- filter=12 channel=17
    -3, 8, -13, 8, 7, -11, -15, -1, -14,
    -- filter=12 channel=18
    0, -3, 8, 11, -6, 9, -1, -5, 1,
    -- filter=12 channel=19
    -2, 3, -4, 3, 7, -6, 3, 12, -7,
    -- filter=12 channel=20
    -7, 0, -11, 1, -7, 10, -8, 9, -8,
    -- filter=12 channel=21
    -9, -2, 3, 1, -17, -6, 12, 14, 7,
    -- filter=12 channel=22
    12, 9, 8, 5, 8, -14, 11, 4, -13,
    -- filter=12 channel=23
    16, 1, -15, 16, -10, 6, -9, -12, -10,
    -- filter=12 channel=24
    11, 15, -10, 9, -6, -5, 1, 1, 10,
    -- filter=12 channel=25
    -1, 2, 6, -11, 5, 0, 6, 5, 12,
    -- filter=12 channel=26
    9, 11, 14, -16, -11, 0, 9, 0, -5,
    -- filter=12 channel=27
    -8, -1, -8, 10, 11, 0, -2, 0, -1,
    -- filter=12 channel=28
    6, -3, -9, -9, -2, -5, -1, 1, -6,
    -- filter=12 channel=29
    13, 6, -8, 11, -8, -14, 9, 10, 10,
    -- filter=12 channel=30
    4, -9, -11, -1, -14, -11, -11, -5, 5,
    -- filter=12 channel=31
    -3, 12, -14, 0, 9, 1, -2, -1, -8,
    -- filter=13 channel=0
    3, -5, -2, -9, 11, -4, 0, 11, 0,
    -- filter=13 channel=1
    3, 0, -13, -2, -3, 7, 0, -10, 0,
    -- filter=13 channel=2
    8, -12, -14, 2, -12, 12, -10, -13, -12,
    -- filter=13 channel=3
    14, 12, -10, 0, 2, 12, 12, -7, -4,
    -- filter=13 channel=4
    -8, -5, -1, 1, -11, 8, -3, -2, -7,
    -- filter=13 channel=5
    -8, -7, 2, -7, 9, -1, -13, -12, -14,
    -- filter=13 channel=6
    5, -6, 14, -7, 3, 14, -7, 8, -2,
    -- filter=13 channel=7
    -8, -9, 5, 1, -12, 3, 0, 8, -12,
    -- filter=13 channel=8
    9, 8, 4, 14, -13, 4, -7, 13, -3,
    -- filter=13 channel=9
    11, -9, 2, 0, -3, 2, 6, 0, 0,
    -- filter=13 channel=10
    4, 4, 4, 6, -10, -4, 8, 1, 1,
    -- filter=13 channel=11
    -12, 1, -6, -7, 9, -8, -2, -1, -5,
    -- filter=13 channel=12
    -4, 6, 14, 14, 8, 2, -14, -13, 2,
    -- filter=13 channel=13
    9, 12, 12, 9, 0, 11, 5, 6, -3,
    -- filter=13 channel=14
    4, -14, -14, -6, 4, 11, -2, -9, 6,
    -- filter=13 channel=15
    12, 0, 8, 4, 0, -1, -5, -14, 14,
    -- filter=13 channel=16
    -10, -11, -9, 0, 14, 5, 0, 6, -3,
    -- filter=13 channel=17
    -7, -1, 3, -10, -7, -1, 11, 6, 2,
    -- filter=13 channel=18
    0, 10, -9, -3, 4, -4, -12, 8, -14,
    -- filter=13 channel=19
    6, 13, 9, -2, -14, -11, 0, 11, -7,
    -- filter=13 channel=20
    11, 7, 3, 0, 11, 13, 12, -5, -11,
    -- filter=13 channel=21
    7, 10, 14, -11, -9, -13, -11, -13, 4,
    -- filter=13 channel=22
    -10, 0, -1, -6, -3, 0, 6, 5, 3,
    -- filter=13 channel=23
    9, -9, -13, -11, -5, 11, -11, -3, 11,
    -- filter=13 channel=24
    -2, -5, -3, -14, 14, 2, -13, 3, -3,
    -- filter=13 channel=25
    -9, 13, 9, -5, -8, 15, 3, 11, -8,
    -- filter=13 channel=26
    0, 1, -9, 0, -2, -2, -11, 12, -11,
    -- filter=13 channel=27
    -4, 8, -14, -11, -12, 1, 5, -13, 0,
    -- filter=13 channel=28
    -9, 6, -13, -10, 11, -4, 0, -1, 12,
    -- filter=13 channel=29
    -14, -9, 2, 0, -11, 0, -2, 14, 4,
    -- filter=13 channel=30
    9, 11, -2, 0, 13, -10, -8, 13, 0,
    -- filter=13 channel=31
    5, 13, -2, -4, -12, 0, 13, -8, 3,
    -- filter=14 channel=0
    3, -11, -11, 9, -13, -9, -1, -3, 10,
    -- filter=14 channel=1
    13, 5, -10, 6, 14, -12, 1, 6, 13,
    -- filter=14 channel=2
    38, 35, 26, -10, 0, -15, 7, -4, -19,
    -- filter=14 channel=3
    -14, -9, -13, -6, -10, -16, -3, 7, 9,
    -- filter=14 channel=4
    11, 20, 14, 14, 11, 8, 4, -4, 5,
    -- filter=14 channel=5
    -6, 8, -12, -1, -15, 6, -2, 10, -7,
    -- filter=14 channel=6
    7, -14, 0, -23, -20, -3, -11, -19, -6,
    -- filter=14 channel=7
    13, 1, 18, -19, -16, -7, -8, -13, 0,
    -- filter=14 channel=8
    11, 10, 9, -2, -4, 8, -6, 9, 5,
    -- filter=14 channel=9
    6, 2, 3, 7, -14, -13, 1, -1, -17,
    -- filter=14 channel=10
    -2, 0, -1, 4, -5, -10, 1, 12, -1,
    -- filter=14 channel=11
    9, 7, -6, -2, -4, -11, 12, 2, 13,
    -- filter=14 channel=12
    19, 18, 4, -13, -6, -9, -14, 1, 3,
    -- filter=14 channel=13
    7, 6, 0, -5, -6, -3, -3, -7, -14,
    -- filter=14 channel=14
    -9, -8, 0, -16, -6, -10, -7, 2, -15,
    -- filter=14 channel=15
    3, -3, -5, -6, -6, -9, -2, -8, 12,
    -- filter=14 channel=16
    4, -13, 10, -5, -21, 0, 1, -3, 7,
    -- filter=14 channel=17
    7, -10, -6, -7, -32, -19, -13, -16, 2,
    -- filter=14 channel=18
    -7, 2, 4, -10, -1, -19, 2, -9, 3,
    -- filter=14 channel=19
    -22, -33, -24, -17, -2, -8, -3, -19, -19,
    -- filter=14 channel=20
    11, 9, -2, -13, -11, 4, -2, -13, -4,
    -- filter=14 channel=21
    -5, 3, -5, -6, -15, 3, 10, 1, -5,
    -- filter=14 channel=22
    2, -4, -11, 6, -9, -6, -14, -6, 12,
    -- filter=14 channel=23
    40, 22, 35, 0, 19, 8, -2, 10, 0,
    -- filter=14 channel=24
    23, 19, 20, -22, -7, 5, 10, -4, 8,
    -- filter=14 channel=25
    4, -11, 9, 10, 8, 8, -4, -8, -10,
    -- filter=14 channel=26
    6, -9, 6, -14, -8, -10, -10, -15, -2,
    -- filter=14 channel=27
    -14, -6, -14, 11, -5, 5, 4, 3, -13,
    -- filter=14 channel=28
    2, -14, -2, -12, -6, 4, -13, 4, -8,
    -- filter=14 channel=29
    -1, 2, -5, -6, 8, 8, 3, 7, -11,
    -- filter=14 channel=30
    -16, -12, 0, 4, -2, 7, -15, 6, 5,
    -- filter=14 channel=31
    -7, 0, 0, 4, 10, 5, 11, -4, -6,
    -- filter=15 channel=0
    -12, -3, -14, 13, -1, 1, -3, -4, 10,
    -- filter=15 channel=1
    -1, 10, -11, -2, -1, 7, -10, 9, -6,
    -- filter=15 channel=2
    -3, 4, 5, -17, 4, -2, 14, 3, 9,
    -- filter=15 channel=3
    -5, -5, 3, -2, 14, -12, 7, -8, 0,
    -- filter=15 channel=4
    -11, -9, -14, -28, -13, 2, -15, 3, -13,
    -- filter=15 channel=5
    8, -2, -6, -3, 7, 1, -2, 14, -12,
    -- filter=15 channel=6
    0, 0, 16, 3, -9, 11, -5, -9, 7,
    -- filter=15 channel=7
    20, 24, 24, 12, 8, 21, 17, 12, 4,
    -- filter=15 channel=8
    2, -21, -6, -22, -8, 10, -6, 3, 2,
    -- filter=15 channel=9
    10, 8, 11, 3, -9, 2, 11, 11, 8,
    -- filter=15 channel=10
    3, 4, 7, 10, 2, 19, -5, -6, 7,
    -- filter=15 channel=11
    9, 0, 0, 0, 12, 1, -5, 13, -13,
    -- filter=15 channel=12
    -12, -18, -17, -1, -15, -3, -14, -8, -6,
    -- filter=15 channel=13
    12, -3, 18, -9, 16, 10, 1, 3, 2,
    -- filter=15 channel=14
    -5, -18, 3, -22, -1, -13, -6, -18, 9,
    -- filter=15 channel=15
    -12, 10, 11, -13, 8, 13, -2, 12, -6,
    -- filter=15 channel=16
    6, -2, -9, 9, -11, -3, 5, 14, -9,
    -- filter=15 channel=17
    6, -3, -1, 19, 5, 12, 13, -5, -10,
    -- filter=15 channel=18
    2, -9, 12, 9, 0, 5, -1, -14, 14,
    -- filter=15 channel=19
    11, -12, -8, -17, -12, 0, -16, -1, -8,
    -- filter=15 channel=20
    -2, 19, 7, -6, 3, -1, 12, 2, 15,
    -- filter=15 channel=21
    18, 12, 9, 2, -4, 0, 14, -6, 2,
    -- filter=15 channel=22
    2, 3, -7, -11, 6, 6, 5, -4, -4,
    -- filter=15 channel=23
    -29, -11, -18, -14, -21, 2, -6, -26, -14,
    -- filter=15 channel=24
    10, 20, 0, 16, -10, 6, 10, -10, -4,
    -- filter=15 channel=25
    -14, 4, 3, 7, -5, 11, 12, 7, 2,
    -- filter=15 channel=26
    21, 14, -1, 13, 15, 6, 13, -5, 3,
    -- filter=15 channel=27
    3, 13, -14, 5, 5, -11, -5, -8, -6,
    -- filter=15 channel=28
    -14, 1, 13, -4, 0, 0, -13, 0, -12,
    -- filter=15 channel=29
    12, 0, -4, 8, 3, 14, 8, -2, 11,
    -- filter=15 channel=30
    17, -1, 13, -6, 11, -3, 6, -12, 14,
    -- filter=15 channel=31
    -1, 5, -3, -12, 11, 13, -12, 4, 14,
    -- filter=16 channel=0
    12, 4, -4, 1, 0, 8, 9, 12, -14,
    -- filter=16 channel=1
    -2, -9, -7, 10, 10, 7, -9, 8, -2,
    -- filter=16 channel=2
    -6, 2, -7, 12, 9, 3, -14, 6, 2,
    -- filter=16 channel=3
    7, -6, 8, 3, -5, -1, 9, -4, -6,
    -- filter=16 channel=4
    14, -11, 8, -14, 14, -14, -4, -5, -14,
    -- filter=16 channel=5
    0, -1, 7, -13, -8, -9, 0, 8, 9,
    -- filter=16 channel=6
    -4, -9, 10, 3, -3, -12, -4, -6, 4,
    -- filter=16 channel=7
    -4, 2, -7, 1, -5, -16, 9, 13, 11,
    -- filter=16 channel=8
    13, 4, -4, 10, 6, -12, 0, -2, -2,
    -- filter=16 channel=9
    -3, -8, 8, 1, -8, -16, 8, 0, 2,
    -- filter=16 channel=10
    -7, 6, -12, -13, 8, 7, -12, 8, 4,
    -- filter=16 channel=11
    4, 6, 2, -2, 4, 4, 1, 9, -1,
    -- filter=16 channel=12
    -4, 7, 9, -7, 4, -6, -2, 0, -5,
    -- filter=16 channel=13
    9, 8, -6, 7, -11, 10, 9, 4, -13,
    -- filter=16 channel=14
    14, 5, 11, -8, 6, -12, -5, -12, -15,
    -- filter=16 channel=15
    -2, -12, -1, -10, -9, 3, -2, 3, -10,
    -- filter=16 channel=16
    -5, -1, -2, -7, 1, 12, -11, -1, 0,
    -- filter=16 channel=17
    8, -5, -10, -3, -10, 1, 2, 2, -4,
    -- filter=16 channel=18
    3, 9, -6, 9, -3, 5, 2, -2, -6,
    -- filter=16 channel=19
    -13, -5, -2, 8, -5, -10, 5, -8, 5,
    -- filter=16 channel=20
    -5, -2, 0, 4, 0, 12, -5, -13, 0,
    -- filter=16 channel=21
    6, 0, 13, -15, -1, -1, -7, 2, 12,
    -- filter=16 channel=22
    -13, -13, -13, 3, 11, -3, 13, -7, 0,
    -- filter=16 channel=23
    -14, -13, 0, -11, 0, 9, -4, 9, 4,
    -- filter=16 channel=24
    -14, 12, 0, 11, 12, 2, 5, 15, -7,
    -- filter=16 channel=25
    5, -4, -13, -2, -7, 14, 11, -12, -1,
    -- filter=16 channel=26
    -1, -6, -10, -14, 14, -15, 5, 7, -8,
    -- filter=16 channel=27
    2, -13, -1, 3, -11, 6, 3, 2, -9,
    -- filter=16 channel=28
    -7, 8, 4, 5, 2, 6, 0, 2, 2,
    -- filter=16 channel=29
    12, -4, 14, 4, -13, -8, 12, 1, -3,
    -- filter=16 channel=30
    -5, 7, 2, 0, 4, -13, -12, 10, 3,
    -- filter=16 channel=31
    3, 1, 3, 7, 1, -1, -9, 5, -1,
    -- filter=17 channel=0
    2, -11, -9, 0, 6, -1, 11, 9, 0,
    -- filter=17 channel=1
    -4, 3, -14, 0, -10, -8, 0, -11, 4,
    -- filter=17 channel=2
    0, 29, 29, -28, -7, -25, 14, 1, 9,
    -- filter=17 channel=3
    3, -5, -14, 11, 1, 8, 6, -2, 2,
    -- filter=17 channel=4
    4, 14, 17, -16, 12, 8, -16, -1, 16,
    -- filter=17 channel=5
    16, -9, 14, -9, -10, 3, -14, -13, -2,
    -- filter=17 channel=6
    9, -3, -12, 7, 6, 11, -10, 9, -4,
    -- filter=17 channel=7
    4, 11, -8, -17, -19, -23, 15, -2, -15,
    -- filter=17 channel=8
    -5, -3, 24, -8, -10, -1, -7, -11, -9,
    -- filter=17 channel=9
    7, 0, 9, -9, -20, 7, 11, 4, -12,
    -- filter=17 channel=10
    12, 1, 2, -14, -1, 9, 1, 4, 8,
    -- filter=17 channel=11
    1, 7, 15, -2, 0, -15, 8, -3, -3,
    -- filter=17 channel=12
    7, 2, -1, -22, -4, -9, 11, 1, 5,
    -- filter=17 channel=13
    -3, -9, 3, -14, -19, -9, 0, -11, -2,
    -- filter=17 channel=14
    3, 10, 22, -26, 4, 13, -7, -8, 16,
    -- filter=17 channel=15
    -13, 11, 9, 5, -12, -7, 3, 6, 11,
    -- filter=17 channel=16
    -4, 0, 3, -13, -3, 5, 10, -3, 0,
    -- filter=17 channel=17
    0, 0, -4, -10, -27, -12, 10, -11, -12,
    -- filter=17 channel=18
    -15, 5, 0, -15, -1, 9, 3, -8, -9,
    -- filter=17 channel=19
    0, -10, 0, 7, -10, 7, 2, -3, -5,
    -- filter=17 channel=20
    -8, 10, -11, -14, -16, -10, 11, 0, 2,
    -- filter=17 channel=21
    4, -10, 13, -5, 0, 0, 10, -8, 6,
    -- filter=17 channel=22
    15, 15, 11, -4, -13, 12, -6, 2, 13,
    -- filter=17 channel=23
    5, 32, 32, 2, 2, 19, -4, -8, 0,
    -- filter=17 channel=24
    9, 16, 11, 7, -24, -14, 2, -15, 6,
    -- filter=17 channel=25
    -5, 5, 6, 10, -14, 2, -1, -13, 10,
    -- filter=17 channel=26
    16, -3, -5, 5, 3, -4, 1, 10, -11,
    -- filter=17 channel=27
    -2, 4, -1, 2, 8, 5, -11, -9, 7,
    -- filter=17 channel=28
    -11, -3, -7, 10, 3, -6, 5, -2, 7,
    -- filter=17 channel=29
    13, -11, -5, 5, -1, -8, 4, 0, -5,
    -- filter=17 channel=30
    -1, 3, -8, 8, -9, -14, -9, -14, 8,
    -- filter=17 channel=31
    11, -14, -4, -6, 1, -12, 6, 10, -11,
    -- filter=18 channel=0
    -4, 0, 13, 2, -5, 7, 4, 0, 3,
    -- filter=18 channel=1
    -8, 1, -8, -12, -3, 14, -10, 8, -12,
    -- filter=18 channel=2
    -19, -7, -4, 8, 8, 9, 17, 10, -2,
    -- filter=18 channel=3
    15, -11, 4, -5, 14, 10, 6, 6, 2,
    -- filter=18 channel=4
    -19, 1, -10, -11, -7, 1, 12, 3, -8,
    -- filter=18 channel=5
    3, -3, 5, 11, 9, 2, -8, 7, -3,
    -- filter=18 channel=6
    -3, 9, 0, 14, 9, 3, -3, 0, -2,
    -- filter=18 channel=7
    8, 11, 18, 2, 1, 3, 12, 14, 25,
    -- filter=18 channel=8
    -6, -12, 1, -12, -8, -16, 0, 2, -3,
    -- filter=18 channel=9
    -7, -10, 2, 0, 0, -11, -1, -6, 9,
    -- filter=18 channel=10
    -8, -1, -6, 13, -8, 15, 0, -2, -1,
    -- filter=18 channel=11
    6, 13, -12, 9, 9, 0, 9, 7, 3,
    -- filter=18 channel=12
    0, 3, 0, 11, 3, 14, 0, -3, -4,
    -- filter=18 channel=13
    9, 2, 14, -6, 13, 17, 12, 15, 0,
    -- filter=18 channel=14
    0, -2, 0, -1, -5, -4, 12, -13, 10,
    -- filter=18 channel=15
    0, -9, 5, -6, 5, -6, -14, 8, 0,
    -- filter=18 channel=16
    -9, -10, -10, -8, -5, -7, 0, 4, -15,
    -- filter=18 channel=17
    13, -9, 0, 1, 3, 20, 0, 7, 3,
    -- filter=18 channel=18
    0, -5, 9, 10, -8, 1, 9, -3, 11,
    -- filter=18 channel=19
    3, 6, -3, 19, -2, -17, -5, -10, -15,
    -- filter=18 channel=20
    7, -1, 6, -2, 2, -2, 8, 4, 2,
    -- filter=18 channel=21
    14, 4, 2, 15, 9, 6, 17, -1, 15,
    -- filter=18 channel=22
    -2, -16, -1, 4, 12, -11, -11, 9, -3,
    -- filter=18 channel=23
    -30, -4, 3, -26, -10, -18, 4, 9, -4,
    -- filter=18 channel=24
    9, -2, 1, 7, 12, -4, 8, 17, 10,
    -- filter=18 channel=25
    -8, -3, 0, 3, 8, 7, 13, 15, 0,
    -- filter=18 channel=26
    -8, 10, 5, 10, -2, 21, -3, 1, 19,
    -- filter=18 channel=27
    -7, 7, -4, 2, 3, 3, 8, 10, 7,
    -- filter=18 channel=28
    15, 11, -4, 11, 5, 16, 0, -3, -8,
    -- filter=18 channel=29
    -12, -6, 10, 11, -2, 10, -10, 2, 14,
    -- filter=18 channel=30
    10, 4, -3, 13, 7, 11, -13, -4, 10,
    -- filter=18 channel=31
    -2, 11, 5, 12, 12, 9, -6, 9, 10,
    -- filter=19 channel=0
    1, 6, 7, -4, 0, 0, 12, 6, 0,
    -- filter=19 channel=1
    4, 11, -6, -12, 4, 7, 1, 2, 14,
    -- filter=19 channel=2
    -39, 7, 45, -31, -6, 14, -16, -4, 6,
    -- filter=19 channel=3
    -6, -6, 9, -12, -3, 6, 4, 10, 0,
    -- filter=19 channel=4
    3, 12, 29, -8, 4, 27, -10, -19, 14,
    -- filter=19 channel=5
    6, 21, 2, 0, 10, 19, -10, 0, 7,
    -- filter=19 channel=6
    -14, -8, 17, 14, -13, 13, 10, 3, 3,
    -- filter=19 channel=7
    -12, -13, 21, -4, -20, -6, 4, -8, -4,
    -- filter=19 channel=8
    -19, -6, 11, -12, -17, 16, 6, 5, 6,
    -- filter=19 channel=9
    -10, 7, 22, -8, 1, 16, -6, -8, -8,
    -- filter=19 channel=10
    0, 0, 14, 9, -8, 14, -2, 5, 0,
    -- filter=19 channel=11
    -12, 3, 12, -12, -6, -13, -12, 5, -9,
    -- filter=19 channel=12
    -10, -2, 23, -19, -3, -1, -19, -12, -6,
    -- filter=19 channel=13
    -20, -13, 5, -15, 1, 14, 12, -5, -1,
    -- filter=19 channel=14
    -8, 1, 19, -28, 7, 5, -1, -14, -4,
    -- filter=19 channel=15
    4, -2, -2, 6, -14, -13, 6, 0, -5,
    -- filter=19 channel=16
    -3, 13, 3, 10, -12, 9, 0, -13, -4,
    -- filter=19 channel=17
    -6, 3, 18, -17, -5, 19, -3, 3, 3,
    -- filter=19 channel=18
    12, 1, 0, 5, -4, -12, 2, -14, 9,
    -- filter=19 channel=19
    8, 4, 9, -9, 12, 21, 0, -8, 7,
    -- filter=19 channel=20
    -12, -5, 2, -1, -8, 4, 12, 5, 6,
    -- filter=19 channel=21
    -4, -2, 15, 6, -5, 4, -12, 6, 1,
    -- filter=19 channel=22
    10, 0, -8, -8, -1, 4, -5, 0, 11,
    -- filter=19 channel=23
    -31, 18, 39, -36, 6, 20, -11, -6, -1,
    -- filter=19 channel=24
    -1, -6, 5, -12, -18, 9, 15, -2, 4,
    -- filter=19 channel=25
    6, -13, 0, -9, 5, -5, 0, 8, -5,
    -- filter=19 channel=26
    -16, -12, 7, 5, 0, 0, 17, 3, -4,
    -- filter=19 channel=27
    -10, -2, 0, 5, -7, 12, -12, -4, 11,
    -- filter=19 channel=28
    1, 9, 10, -12, -1, -11, -7, -8, -10,
    -- filter=19 channel=29
    -11, 5, 2, 14, 4, 10, -12, 10, -1,
    -- filter=19 channel=30
    0, -11, 7, 1, -5, -10, 7, -6, 12,
    -- filter=19 channel=31
    -8, -8, -4, -10, 12, 0, -5, 2, -9,
    -- filter=20 channel=0
    8, 0, 0, -10, 5, -4, -5, 8, -8,
    -- filter=20 channel=1
    -12, 0, -3, 12, 1, -3, -2, -12, -11,
    -- filter=20 channel=2
    -21, -7, -2, -12, 0, 5, -6, -32, 1,
    -- filter=20 channel=3
    -12, 4, 2, -7, -6, 11, -9, -11, -6,
    -- filter=20 channel=4
    -5, 16, 23, 6, -3, 17, 6, 12, 15,
    -- filter=20 channel=5
    5, -2, 0, -9, -14, 12, -14, -13, -1,
    -- filter=20 channel=6
    -4, -15, -12, 1, 7, 6, 8, 1, -1,
    -- filter=20 channel=7
    -4, -10, 11, -10, -22, -13, -7, -8, -1,
    -- filter=20 channel=8
    6, -6, 15, 7, 15, 16, -9, 13, -8,
    -- filter=20 channel=9
    -5, -4, -6, -18, -19, 6, 0, -15, -8,
    -- filter=20 channel=10
    -17, -7, 7, -7, -6, -1, 12, 11, -1,
    -- filter=20 channel=11
    0, 3, 15, 0, -11, 13, -10, 7, -11,
    -- filter=20 channel=12
    -2, 0, -4, 8, 13, 19, -12, 1, 15,
    -- filter=20 channel=13
    1, 1, 3, 4, -9, -15, 13, -2, -15,
    -- filter=20 channel=14
    -2, 12, 9, 9, 21, 5, -4, 16, -6,
    -- filter=20 channel=15
    -12, -14, -7, 0, 5, 13, 2, -13, 4,
    -- filter=20 channel=16
    -13, -10, 12, -13, 12, -1, -14, -6, 7,
    -- filter=20 channel=17
    6, 0, 21, -5, -18, 5, 5, 2, -10,
    -- filter=20 channel=18
    10, -5, 15, -9, -9, 10, 10, 15, -7,
    -- filter=20 channel=19
    6, 2, 10, 18, 6, 20, 3, 1, 23,
    -- filter=20 channel=20
    10, 12, -7, 10, -5, 3, -3, -2, 0,
    -- filter=20 channel=21
    -12, -1, -18, 6, 2, -12, 1, -5, -16,
    -- filter=20 channel=22
    8, -11, 12, 14, 13, -7, -4, -3, 0,
    -- filter=20 channel=23
    -2, 15, 30, -16, 3, 17, 5, 0, 17,
    -- filter=20 channel=24
    -19, -3, 9, -9, -6, -11, 3, -17, -9,
    -- filter=20 channel=25
    -14, 11, 14, -6, 7, 0, 13, 4, 8,
    -- filter=20 channel=26
    -7, 4, -6, -1, 2, 2, -8, 2, -3,
    -- filter=20 channel=27
    4, 1, 3, -6, -7, 0, 0, 8, 9,
    -- filter=20 channel=28
    5, 2, 3, -14, -5, 0, 11, -11, -8,
    -- filter=20 channel=29
    -11, 3, 5, -4, 13, 1, 10, -1, 0,
    -- filter=20 channel=30
    -6, -7, -9, -13, 9, 4, 3, -2, -2,
    -- filter=20 channel=31
    5, 14, -6, 14, -3, 9, 12, -1, 12,
    -- filter=21 channel=0
    -3, 10, -10, 8, 0, 4, 1, 14, -4,
    -- filter=21 channel=1
    9, -5, 2, 5, 10, -12, -9, 15, 1,
    -- filter=21 channel=2
    0, 2, 13, -25, 16, 25, -6, -3, 5,
    -- filter=21 channel=3
    -7, 16, -5, -2, -11, 15, 7, 13, 10,
    -- filter=21 channel=4
    0, -13, -11, -1, 2, 0, 6, 4, 0,
    -- filter=21 channel=5
    -1, 5, -3, -9, -2, 9, -15, -6, 9,
    -- filter=21 channel=6
    0, -4, -5, -10, 11, 15, -12, -11, 9,
    -- filter=21 channel=7
    -7, 2, -4, 2, -6, 10, -17, 9, 3,
    -- filter=21 channel=8
    1, -19, -15, 2, 4, 8, -8, -1, 12,
    -- filter=21 channel=9
    6, -9, 10, -14, -7, 13, -13, 10, 0,
    -- filter=21 channel=10
    3, 12, 0, 3, -7, 10, 5, 9, 14,
    -- filter=21 channel=11
    15, 14, -8, -11, 3, 14, 8, -8, 12,
    -- filter=21 channel=12
    0, -11, 5, -16, 1, 9, 0, -7, 18,
    -- filter=21 channel=13
    3, -7, -11, 0, 9, -4, -3, -6, 13,
    -- filter=21 channel=14
    4, -12, -13, -12, 9, 0, -7, -12, -8,
    -- filter=21 channel=15
    -10, -5, -2, 5, 5, 4, 7, -6, 10,
    -- filter=21 channel=16
    2, 0, -5, 5, -3, 1, -16, 8, -9,
    -- filter=21 channel=17
    7, 4, 14, 10, 15, 18, -8, 12, 24,
    -- filter=21 channel=18
    9, 7, -3, 14, 0, 2, -8, 0, 6,
    -- filter=21 channel=19
    15, -1, -8, -1, 3, 3, 11, 21, 14,
    -- filter=21 channel=20
    -12, 14, 9, -3, 16, -9, -5, -3, 14,
    -- filter=21 channel=21
    11, 3, 18, -12, -4, 7, 10, 12, 0,
    -- filter=21 channel=22
    5, -15, -13, -4, -9, 4, 14, -8, 8,
    -- filter=21 channel=23
    -6, -26, -18, -3, -13, -7, -7, 5, -1,
    -- filter=21 channel=24
    -5, -3, 16, 0, 11, 14, -16, -8, 13,
    -- filter=21 channel=25
    0, 12, -4, 5, -11, -10, 0, -13, -11,
    -- filter=21 channel=26
    14, -11, -5, -6, -1, -3, -8, 14, 12,
    -- filter=21 channel=27
    9, -1, 8, 14, 13, -14, 4, 6, 11,
    -- filter=21 channel=28
    -11, 0, -4, -11, 15, 17, 9, 1, -2,
    -- filter=21 channel=29
    -5, -13, 13, 1, -3, 2, 1, -8, -7,
    -- filter=21 channel=30
    10, 13, 10, -7, -5, -10, -3, 0, 15,
    -- filter=21 channel=31
    6, -11, -6, 15, -6, -2, -10, -2, 12,
    -- filter=22 channel=0
    -2, -9, -12, 4, -11, 0, -3, -4, -6,
    -- filter=22 channel=1
    11, 12, -1, 15, 0, 4, -11, 9, 7,
    -- filter=22 channel=2
    -23, 9, 22, -16, 16, 12, -3, -3, 15,
    -- filter=22 channel=3
    11, -2, -10, 16, 14, 4, 15, -2, -5,
    -- filter=22 channel=4
    -11, -12, -5, 8, -28, -8, 2, -3, -3,
    -- filter=22 channel=5
    4, 2, 14, 1, -1, 13, 6, 10, 5,
    -- filter=22 channel=6
    9, 14, 19, -8, -4, 21, -7, 15, -4,
    -- filter=22 channel=7
    -10, 8, 25, -12, -5, 17, -1, 0, 23,
    -- filter=22 channel=8
    0, -18, -4, 0, 0, -4, -11, 8, -17,
    -- filter=22 channel=9
    -4, 7, 9, -8, 10, 17, 2, 4, -5,
    -- filter=22 channel=10
    3, 6, 6, 0, 10, 0, 11, 15, 3,
    -- filter=22 channel=11
    6, -2, 7, 13, 14, -6, 6, 9, 15,
    -- filter=22 channel=12
    -14, -12, 9, -13, -6, -9, -4, -15, -7,
    -- filter=22 channel=13
    11, 9, 18, -1, -6, -3, -1, 0, 10,
    -- filter=22 channel=14
    -6, -17, -14, 2, -17, -6, -5, -18, -2,
    -- filter=22 channel=15
    -2, -8, -11, 1, 0, 8, 9, 12, 5,
    -- filter=22 channel=16
    0, 5, 16, -6, 16, 14, 4, -3, 5,
    -- filter=22 channel=17
    3, -10, 6, 16, 11, 5, 6, 17, 3,
    -- filter=22 channel=18
    14, -9, -1, -4, -3, -7, 1, 11, -3,
    -- filter=22 channel=19
    20, -2, 15, -7, 9, -3, -5, 9, 2,
    -- filter=22 channel=20
    -10, -3, 7, 0, 9, -6, 8, 15, -6,
    -- filter=22 channel=21
    -13, -5, 7, 7, 14, 17, 1, 8, 24,
    -- filter=22 channel=22
    0, 1, -3, 10, -2, 4, -3, -5, 6,
    -- filter=22 channel=23
    4, -2, 3, 1, -23, -18, -8, 1, -16,
    -- filter=22 channel=24
    -11, 11, 9, -1, 12, 8, -12, 1, 13,
    -- filter=22 channel=25
    0, 3, -11, 2, -7, 1, -6, -10, -3,
    -- filter=22 channel=26
    14, -7, 13, -11, 11, 18, 7, 9, 21,
    -- filter=22 channel=27
    14, -14, 10, 12, -7, -5, 7, -10, 12,
    -- filter=22 channel=28
    14, -10, -7, 0, 8, -9, 5, -14, -9,
    -- filter=22 channel=29
    -10, -1, 11, -6, -9, -3, -1, -2, 1,
    -- filter=22 channel=30
    -3, 17, -7, 1, 13, 0, -9, 5, 14,
    -- filter=22 channel=31
    5, 4, 2, -6, -4, -1, 6, 7, -10,
    -- filter=23 channel=0
    13, 5, 5, 0, 10, -4, 5, 7, -13,
    -- filter=23 channel=1
    -5, -9, 4, -4, 8, -4, -12, -9, -8,
    -- filter=23 channel=2
    -11, 18, -18, -2, 9, -19, -18, 11, -12,
    -- filter=23 channel=3
    0, 4, 2, 6, 0, -4, 16, 5, -9,
    -- filter=23 channel=4
    7, 6, -8, 2, -2, 6, -5, -13, 1,
    -- filter=23 channel=5
    16, 19, -5, -7, 2, -11, 17, 14, 7,
    -- filter=23 channel=6
    -4, -7, 7, 0, 22, 1, 1, 8, -5,
    -- filter=23 channel=7
    -3, 4, 7, -4, 17, 8, 2, -1, 6,
    -- filter=23 channel=8
    5, -11, -3, -18, 4, 2, 7, 11, 4,
    -- filter=23 channel=9
    -16, -5, -17, -9, 13, -10, -13, 8, -2,
    -- filter=23 channel=10
    2, -8, 0, 0, 3, -2, 0, 13, -3,
    -- filter=23 channel=11
    -1, -4, 11, 1, -11, -12, -6, 3, 15,
    -- filter=23 channel=12
    7, 13, 15, 7, 6, 1, -12, -12, 13,
    -- filter=23 channel=13
    5, 18, 6, -13, 0, 5, -2, 0, 2,
    -- filter=23 channel=14
    11, 18, 0, 1, 3, -4, 3, -11, -1,
    -- filter=23 channel=15
    -12, 2, -6, 13, 6, 13, 5, -9, -12,
    -- filter=23 channel=16
    -5, 13, 14, 18, 13, -8, -7, 10, 6,
    -- filter=23 channel=17
    4, 21, 8, -9, 16, -1, 5, 15, 14,
    -- filter=23 channel=18
    -6, 3, 1, -2, -10, 9, -4, 3, 1,
    -- filter=23 channel=19
    14, -5, 9, 28, 12, 6, -1, -4, 5,
    -- filter=23 channel=20
    14, -3, -1, 16, 14, -3, 16, 10, 8,
    -- filter=23 channel=21
    -17, -10, 4, 3, -1, -16, -12, 0, -8,
    -- filter=23 channel=22
    5, -12, -5, 12, 3, -9, 5, 0, -7,
    -- filter=23 channel=23
    0, -2, 0, -14, -18, -22, -19, -12, -16,
    -- filter=23 channel=24
    8, 7, -5, 0, 15, -11, 2, 17, -11,
    -- filter=23 channel=25
    -2, 6, -2, 2, -5, -7, -13, 3, -9,
    -- filter=23 channel=26
    12, 8, 2, 6, 20, 12, 5, 10, 8,
    -- filter=23 channel=27
    0, -3, -11, -3, 1, -4, 0, 0, 4,
    -- filter=23 channel=28
    -3, -1, -5, -12, 8, 7, -2, 7, 9,
    -- filter=23 channel=29
    -13, 0, 13, 11, -14, 9, 13, 7, -12,
    -- filter=23 channel=30
    11, 3, 14, 14, 10, 8, 7, 11, 17,
    -- filter=23 channel=31
    -11, 6, 10, -5, -11, 11, 9, 9, -7,
    -- filter=24 channel=0
    -14, 7, -11, 5, 2, -14, -11, -7, 5,
    -- filter=24 channel=1
    2, -10, 9, 0, 14, 2, -9, -12, 9,
    -- filter=24 channel=2
    9, -10, 11, -14, -11, -14, 3, -14, -7,
    -- filter=24 channel=3
    8, 2, -12, 0, 0, 8, -1, 10, 11,
    -- filter=24 channel=4
    16, -5, 19, 9, -3, 0, 18, -14, -13,
    -- filter=24 channel=5
    -4, 13, 10, 1, -12, 9, -14, 13, -2,
    -- filter=24 channel=6
    9, 9, 10, -12, -3, 1, 6, -6, -8,
    -- filter=24 channel=7
    -15, -5, 0, -1, -15, -3, -10, 0, 0,
    -- filter=24 channel=8
    -9, 15, 1, 14, -8, -6, -8, 1, -4,
    -- filter=24 channel=9
    -2, 5, 3, -9, 12, -12, 9, -14, 3,
    -- filter=24 channel=10
    9, -13, 14, 8, 12, 0, 14, -1, 2,
    -- filter=24 channel=11
    -4, 9, 0, -1, -11, -2, 0, -4, -1,
    -- filter=24 channel=12
    -10, 1, -11, 10, -12, 3, -9, -4, 11,
    -- filter=24 channel=13
    -13, 0, 2, -9, -8, -2, -3, 15, -10,
    -- filter=24 channel=14
    -2, 18, 8, 7, 2, -9, 17, 6, -13,
    -- filter=24 channel=15
    3, -4, -12, 12, 14, 14, 3, 1, -14,
    -- filter=24 channel=16
    -4, 4, 14, -13, -1, 6, 0, 2, 10,
    -- filter=24 channel=17
    -14, -8, -3, 2, -9, 0, -7, 16, 15,
    -- filter=24 channel=18
    10, -11, 0, 10, -5, -12, -9, -9, -3,
    -- filter=24 channel=19
    14, -7, -13, 11, 9, -6, 0, -8, 8,
    -- filter=24 channel=20
    8, 0, 1, 1, 12, -14, 0, 6, 2,
    -- filter=24 channel=21
    -3, 11, 0, 8, -3, 0, 6, 6, 2,
    -- filter=24 channel=22
    -6, -13, 4, 3, 8, -2, -3, 10, -14,
    -- filter=24 channel=23
    11, 19, 4, -3, 14, 12, 16, -13, -16,
    -- filter=24 channel=24
    11, -5, 2, 5, -4, -16, -3, 8, -1,
    -- filter=24 channel=25
    7, -2, 8, 6, -4, -9, -3, -8, 10,
    -- filter=24 channel=26
    12, 8, 8, -12, -9, 4, 2, -3, 14,
    -- filter=24 channel=27
    -4, -14, -7, -3, -12, 4, -7, -14, 8,
    -- filter=24 channel=28
    6, -5, 5, 1, 14, 0, 13, -10, -2,
    -- filter=24 channel=29
    0, -3, 5, -1, 8, 0, 14, 14, -9,
    -- filter=24 channel=30
    -3, -3, 12, 1, -7, 12, -9, 3, -2,
    -- filter=24 channel=31
    5, -10, -9, 2, -7, -3, 5, -12, -5,
    -- filter=25 channel=0
    9, -11, 2, 15, -13, 2, -11, -7, -14,
    -- filter=25 channel=1
    11, -13, 6, 0, -11, -6, 7, 11, 9,
    -- filter=25 channel=2
    -1, 4, 14, 4, 1, 1, 21, 2, -4,
    -- filter=25 channel=3
    2, -13, -6, -11, -8, 4, 0, 7, 7,
    -- filter=25 channel=4
    10, -1, -3, 10, 3, 1, -3, 9, -3,
    -- filter=25 channel=5
    14, 1, -5, -2, 7, 13, -4, -9, -14,
    -- filter=25 channel=6
    0, -3, 8, -5, 10, 0, -5, 15, -8,
    -- filter=25 channel=7
    -10, -15, -13, 6, -5, -8, -10, -5, 0,
    -- filter=25 channel=8
    -2, 0, -13, -1, 2, 1, 14, 4, -10,
    -- filter=25 channel=9
    -14, 6, 5, -8, -11, -14, -3, 6, -16,
    -- filter=25 channel=10
    -13, -10, 12, -14, 0, -5, 12, 0, 5,
    -- filter=25 channel=11
    -3, -13, 11, -4, 6, 3, -3, -10, -2,
    -- filter=25 channel=12
    1, 7, 14, -11, -10, -1, -1, 6, -7,
    -- filter=25 channel=13
    -10, -8, 6, -6, 0, 4, -3, 8, 12,
    -- filter=25 channel=14
    -12, -9, 10, 14, -1, 10, -3, -8, -9,
    -- filter=25 channel=15
    -5, -12, -11, 13, 3, -8, 12, -9, -12,
    -- filter=25 channel=16
    5, 9, -6, -5, -5, 3, 4, 8, -8,
    -- filter=25 channel=17
    -12, 5, -4, -11, -14, 5, -7, 12, -6,
    -- filter=25 channel=18
    -12, -14, -8, 2, 1, 8, 14, 9, 6,
    -- filter=25 channel=19
    5, -2, 3, -8, 16, -4, -1, -2, -2,
    -- filter=25 channel=20
    0, 2, -7, -11, -12, -4, -5, -3, 9,
    -- filter=25 channel=21
    0, 9, -1, 2, -4, -10, 5, 7, -14,
    -- filter=25 channel=22
    -8, -4, 14, 0, -13, 5, 0, 16, 9,
    -- filter=25 channel=23
    -3, -6, -5, 6, -6, 3, 12, 13, 5,
    -- filter=25 channel=24
    -5, -7, 14, 7, -9, 4, 11, 13, 1,
    -- filter=25 channel=25
    -7, 0, -10, -11, 6, 8, 10, -14, -1,
    -- filter=25 channel=26
    6, -4, 7, -4, -6, -7, 12, -12, 8,
    -- filter=25 channel=27
    12, 2, 5, -13, -9, 12, 4, 9, -13,
    -- filter=25 channel=28
    0, -14, 3, -11, 0, -1, -13, -8, -11,
    -- filter=25 channel=29
    -4, -2, 2, -5, -3, -11, -5, 2, 6,
    -- filter=25 channel=30
    1, -7, -14, 6, -2, -14, -14, -14, 3,
    -- filter=25 channel=31
    7, 6, 3, 7, 11, -12, 2, -5, 1,
    -- filter=26 channel=0
    -2, 14, -8, 7, -7, -1, 7, 8, 2,
    -- filter=26 channel=1
    -10, 14, -4, -7, -4, 0, -4, 3, 0,
    -- filter=26 channel=2
    -6, -1, 6, 1, -14, 8, 12, 23, 4,
    -- filter=26 channel=3
    -12, -9, -8, 14, -6, 12, -2, 7, -8,
    -- filter=26 channel=4
    -4, 6, -12, -3, 4, 0, -7, 3, -2,
    -- filter=26 channel=5
    -3, 1, 1, -10, 6, 8, -11, -14, -9,
    -- filter=26 channel=6
    -10, -14, -3, -12, 5, -16, 0, 0, -10,
    -- filter=26 channel=7
    -10, -9, 5, -1, -16, -1, 0, 15, -2,
    -- filter=26 channel=8
    1, -12, -9, 6, -2, -6, 13, 1, -9,
    -- filter=26 channel=9
    9, -11, 1, -16, -7, -17, 0, 3, 6,
    -- filter=26 channel=10
    12, 4, 3, 5, -2, -12, 9, -13, -4,
    -- filter=26 channel=11
    10, 0, 7, 1, -4, -13, 8, -9, 6,
    -- filter=26 channel=12
    -7, -6, -15, 4, -11, 13, 16, 10, 0,
    -- filter=26 channel=13
    -16, 3, -10, -9, 1, -3, 6, -1, 8,
    -- filter=26 channel=14
    11, 0, -5, 14, 2, -11, 10, 2, 12,
    -- filter=26 channel=15
    -3, -5, -1, -11, 10, 6, -3, 2, -11,
    -- filter=26 channel=16
    3, 8, -5, 3, -10, 2, 9, 16, -7,
    -- filter=26 channel=17
    3, 0, -17, 11, -4, 5, 3, 14, -10,
    -- filter=26 channel=18
    -10, 0, 2, -7, 15, -5, -6, 10, -13,
    -- filter=26 channel=19
    12, -5, -12, 0, -10, -8, -15, -14, 11,
    -- filter=26 channel=20
    -10, 1, 4, 5, 5, -1, 2, 3, 7,
    -- filter=26 channel=21
    -5, -3, -3, 6, -16, -13, 8, 0, -3,
    -- filter=26 channel=22
    -10, -14, -12, 8, 11, 6, -14, 1, 9,
    -- filter=26 channel=23
    -4, -18, -6, 6, 14, 1, -2, 5, 18,
    -- filter=26 channel=24
    -7, 3, -9, 12, 7, -2, 4, 16, -2,
    -- filter=26 channel=25
    11, 5, -10, 4, -10, -8, 6, -4, 5,
    -- filter=26 channel=26
    -13, -1, 0, -9, -8, 0, 12, -14, -6,
    -- filter=26 channel=27
    11, -4, -5, 1, -10, 10, 12, 5, -14,
    -- filter=26 channel=28
    12, 5, 9, -13, 11, 3, -10, 4, -9,
    -- filter=26 channel=29
    2, 8, -8, 0, 7, -10, 9, -9, 4,
    -- filter=26 channel=30
    2, 1, 0, 10, -6, -3, -3, 0, -5,
    -- filter=26 channel=31
    6, -13, 11, -10, 14, -8, -3, 2, 2,
    -- filter=27 channel=0
    -14, -9, -1, 8, -3, -4, 3, -4, -6,
    -- filter=27 channel=1
    -6, 0, -12, -1, 12, -6, 13, 8, 8,
    -- filter=27 channel=2
    13, -6, 0, -14, -6, -8, 10, -12, -24,
    -- filter=27 channel=3
    3, -7, -9, 9, 8, -13, -14, 4, -14,
    -- filter=27 channel=4
    10, 26, 19, -5, -5, 8, 17, 6, 5,
    -- filter=27 channel=5
    6, -11, -9, -13, 6, -2, 10, 4, -15,
    -- filter=27 channel=6
    11, -12, -4, 2, -14, -3, 3, 2, -14,
    -- filter=27 channel=7
    -12, 0, 10, -18, -3, -20, 3, -1, 1,
    -- filter=27 channel=8
    12, 3, 13, -11, 17, 10, -10, 1, 12,
    -- filter=27 channel=9
    -11, 7, -5, -14, -16, -13, -2, 1, -16,
    -- filter=27 channel=10
    -5, 5, 7, 5, 2, 0, -1, -10, 3,
    -- filter=27 channel=11
    5, 12, -13, 3, 0, -7, 0, 9, -14,
    -- filter=27 channel=12
    13, -1, -6, -5, 6, 6, -6, -9, 11,
    -- filter=27 channel=13
    -14, 11, 12, 3, 2, 3, -8, 4, -9,
    -- filter=27 channel=14
    25, 10, 7, 9, 15, 6, -6, 11, -8,
    -- filter=27 channel=15
    -14, 0, -9, -5, 11, 0, 3, 9, -2,
    -- filter=27 channel=16
    -14, -9, 13, -4, 5, 8, 10, 8, 11,
    -- filter=27 channel=17
    -3, 13, 0, 6, -8, -16, 13, -4, -7,
    -- filter=27 channel=18
    13, 2, 10, 5, -8, -9, 8, 12, 14,
    -- filter=27 channel=19
    6, 4, 12, 0, 14, -10, 15, 3, 4,
    -- filter=27 channel=20
    8, -10, -9, 5, -19, -11, -12, 0, -17,
    -- filter=27 channel=21
    -16, 10, -13, -14, -11, 1, -5, -8, 7,
    -- filter=27 channel=22
    6, -6, 3, -7, -2, 14, -12, -5, -4,
    -- filter=27 channel=23
    32, 22, -3, 6, 0, 5, 3, 7, 0,
    -- filter=27 channel=24
    -6, -14, 7, -23, -20, -14, -5, -13, -3,
    -- filter=27 channel=25
    0, -1, 2, 9, 1, -7, 11, 8, -1,
    -- filter=27 channel=26
    5, 4, -15, -12, -3, -14, 9, -12, -12,
    -- filter=27 channel=27
    -10, 0, 9, -3, 5, -4, 13, -8, -1,
    -- filter=27 channel=28
    -4, 10, 9, 0, 5, 5, 8, 10, 2,
    -- filter=27 channel=29
    0, 9, 3, -7, -14, -8, 14, 9, -2,
    -- filter=27 channel=30
    13, 5, -2, -3, 7, -6, 3, -10, -6,
    -- filter=27 channel=31
    -12, 11, 6, -8, 2, -14, -9, 8, -13,
    -- filter=28 channel=0
    -5, -5, -6, 6, -14, -1, 0, -2, 13,
    -- filter=28 channel=1
    -2, 4, -6, 10, 6, -9, -7, -6, -6,
    -- filter=28 channel=2
    2, -4, -6, -6, -17, -16, -8, -6, -8,
    -- filter=28 channel=3
    -2, 0, -5, 13, 10, 10, -4, -6, -11,
    -- filter=28 channel=4
    4, 3, 4, -9, 7, -6, 3, 21, 0,
    -- filter=28 channel=5
    -14, 13, 6, -1, -2, 9, 13, -4, 6,
    -- filter=28 channel=6
    -8, 0, 13, 4, -4, -3, -13, -3, -10,
    -- filter=28 channel=7
    -10, 3, 4, -4, 0, 4, -15, 8, 4,
    -- filter=28 channel=8
    7, -9, 10, -1, -2, 14, -2, 13, 0,
    -- filter=28 channel=9
    14, 0, -7, 12, 1, 0, 5, -6, -5,
    -- filter=28 channel=10
    11, 0, 12, -5, 3, -13, 6, -8, -9,
    -- filter=28 channel=11
    1, 0, -2, -1, 0, 12, -3, -6, -10,
    -- filter=28 channel=12
    0, 9, -7, -3, -4, 14, 1, -6, 7,
    -- filter=28 channel=13
    12, -14, -12, 3, 6, 8, 4, 8, 2,
    -- filter=28 channel=14
    1, 15, 4, -1, -4, 12, 4, 16, 16,
    -- filter=28 channel=15
    -9, -7, -14, 13, 13, 8, 1, -11, 14,
    -- filter=28 channel=16
    13, -9, -1, 8, 7, -3, -15, 4, 17,
    -- filter=28 channel=17
    2, 5, -4, -2, -9, -9, -2, -3, 15,
    -- filter=28 channel=18
    -12, 6, 1, 13, 9, 15, -1, -3, 14,
    -- filter=28 channel=19
    8, -8, 15, -2, 7, 14, 7, 21, -4,
    -- filter=28 channel=20
    -10, -12, 9, -4, 2, -8, 1, -3, 6,
    -- filter=28 channel=21
    -3, -11, 2, -10, -8, -8, 11, -10, 10,
    -- filter=28 channel=22
    10, -9, -10, -13, -13, -8, -5, 11, -11,
    -- filter=28 channel=23
    11, -16, -12, -6, 0, 8, -6, 15, 8,
    -- filter=28 channel=24
    -12, 0, 0, -13, -7, -15, -13, 1, 6,
    -- filter=28 channel=25
    0, 4, -3, -1, -8, 3, -9, 11, 9,
    -- filter=28 channel=26
    -10, 16, 1, 0, 4, -3, -7, 7, -5,
    -- filter=28 channel=27
    11, -2, -6, 5, -13, -10, 14, -14, -8,
    -- filter=28 channel=28
    8, 5, -12, -11, -4, -13, -9, -4, 0,
    -- filter=28 channel=29
    13, 14, -6, -2, 3, -5, -2, 1, -1,
    -- filter=28 channel=30
    16, 4, 14, -5, 11, -9, -12, -9, 13,
    -- filter=28 channel=31
    11, 13, 5, -12, 0, -12, -8, 12, 1,
    -- filter=29 channel=0
    -10, 3, -8, 9, 9, 3, 6, 3, 4,
    -- filter=29 channel=1
    0, 0, 1, 10, 0, -14, 12, 0, 7,
    -- filter=29 channel=2
    -21, 16, 31, -29, 10, 13, -8, 9, 18,
    -- filter=29 channel=3
    0, 4, 3, 16, -12, -13, 3, -14, -8,
    -- filter=29 channel=4
    -3, -16, 19, -4, 8, -7, -14, -5, -10,
    -- filter=29 channel=5
    4, 12, 16, -11, -12, -12, -11, -10, 14,
    -- filter=29 channel=6
    2, -14, 0, -14, 9, 0, 14, -7, 6,
    -- filter=29 channel=7
    -16, -1, -4, -10, -7, 12, 12, 1, -6,
    -- filter=29 channel=8
    6, 8, 10, -12, 0, 15, -16, -16, -13,
    -- filter=29 channel=9
    -13, -6, 0, -9, 9, 13, -4, -14, -9,
    -- filter=29 channel=10
    16, -5, -13, -8, 13, 13, -4, 7, -9,
    -- filter=29 channel=11
    12, 6, 8, -4, -11, 8, 13, 0, -2,
    -- filter=29 channel=12
    -19, -11, 5, -7, -10, 4, 6, -12, 14,
    -- filter=29 channel=13
    -7, -16, -1, 7, -13, 6, 10, 8, 1,
    -- filter=29 channel=14
    8, -6, 4, 3, -15, 18, 4, -21, 1,
    -- filter=29 channel=15
    13, 3, -3, 12, 10, -8, -4, -1, -8,
    -- filter=29 channel=16
    14, 1, 8, -13, 13, 15, -4, 11, -3,
    -- filter=29 channel=17
    -3, 9, 4, -17, -12, -4, 8, -18, 11,
    -- filter=29 channel=18
    -12, 11, -12, 12, -5, -6, -14, 10, 7,
    -- filter=29 channel=19
    15, -10, 0, 6, 10, 2, 1, 3, -1,
    -- filter=29 channel=20
    9, 6, 3, -8, -10, -11, -4, 4, 6,
    -- filter=29 channel=21
    8, -15, -8, -3, -5, -7, 3, 5, 3,
    -- filter=29 channel=22
    -5, -12, 2, -9, 1, 2, 2, 11, 5,
    -- filter=29 channel=23
    -20, 4, 25, -18, 14, 26, 0, -9, 20,
    -- filter=29 channel=24
    -11, 8, -3, 0, 8, 13, 2, -17, 14,
    -- filter=29 channel=25
    -14, -13, 1, -11, -14, 2, 7, 0, 0,
    -- filter=29 channel=26
    0, -4, 9, 4, -12, 5, 13, 5, 12,
    -- filter=29 channel=27
    -7, 8, -4, -1, -10, 5, 11, 8, 13,
    -- filter=29 channel=28
    -10, -15, -11, -7, 14, 16, -9, 11, 9,
    -- filter=29 channel=29
    -2, 11, -5, 7, -13, -11, 10, -1, 12,
    -- filter=29 channel=30
    -9, 11, -1, -2, -11, -4, -8, 8, 2,
    -- filter=29 channel=31
    -3, -3, -12, 13, 4, 15, -8, -10, -9,
    -- filter=30 channel=0
    10, -14, 6, -12, -10, 11, -12, -8, 12,
    -- filter=30 channel=1
    -6, 11, -8, 0, 11, 5, -13, -13, 11,
    -- filter=30 channel=2
    18, 20, 24, -3, 16, 13, 5, 16, -1,
    -- filter=30 channel=3
    11, -7, -2, -4, -8, -3, -10, -6, -1,
    -- filter=30 channel=4
    -21, -32, -7, -25, -21, 2, 4, -5, -2,
    -- filter=30 channel=5
    4, 12, -11, 8, 5, 10, -7, -11, -10,
    -- filter=30 channel=6
    -4, 4, 13, 2, 1, 9, -12, 3, 0,
    -- filter=30 channel=7
    5, 17, -1, 0, 9, 16, 17, 10, 4,
    -- filter=30 channel=8
    -14, -2, 6, -4, -25, 0, -13, 5, 0,
    -- filter=30 channel=9
    8, -11, 4, 17, 4, 13, 11, -2, 5,
    -- filter=30 channel=10
    14, 7, 10, -7, -3, -5, 12, 3, 19,
    -- filter=30 channel=11
    -4, -6, -9, -14, 11, 4, -7, 8, -6,
    -- filter=30 channel=12
    -15, -2, 0, -12, -20, 6, 10, 4, 4,
    -- filter=30 channel=13
    -1, 12, 17, 3, 0, 19, 5, 0, 6,
    -- filter=30 channel=14
    -17, -34, -20, -16, -18, -19, 4, -21, 0,
    -- filter=30 channel=15
    12, 15, -9, 1, -12, -2, 13, -5, 3,
    -- filter=30 channel=16
    6, -1, 10, -10, -14, 2, -1, -3, -14,
    -- filter=30 channel=17
    -14, -6, 0, -11, 6, -5, -4, 7, 1,
    -- filter=30 channel=18
    -6, -4, 10, 8, -2, 6, 6, 8, -2,
    -- filter=30 channel=19
    0, -1, -14, -6, -26, 0, 2, -1, -22,
    -- filter=30 channel=20
    -7, 5, -9, 15, -9, 4, 7, 4, 5,
    -- filter=30 channel=21
    19, 19, 25, 12, 14, 17, 0, 14, 0,
    -- filter=30 channel=22
    -7, -19, -4, -12, -18, -17, -5, -12, -16,
    -- filter=30 channel=23
    -30, -20, -8, -22, -37, -5, -18, -23, -5,
    -- filter=30 channel=24
    9, 16, 26, 11, 19, 16, 1, -1, 3,
    -- filter=30 channel=25
    12, -9, -2, -13, 8, -7, -5, 9, -4,
    -- filter=30 channel=26
    8, -3, 11, -3, 5, 0, 2, 20, -2,
    -- filter=30 channel=27
    -13, -8, -7, -8, -15, -10, 5, 11, -10,
    -- filter=30 channel=28
    -9, -17, -6, 8, -6, -2, 4, 0, 4,
    -- filter=30 channel=29
    10, -2, 11, -12, 0, -1, 2, 6, 8,
    -- filter=30 channel=30
    2, 4, -10, 5, -11, -9, 7, -15, 7,
    -- filter=30 channel=31
    -5, 6, -13, -7, -2, 6, 12, 7, 3,
    -- filter=31 channel=0
    -9, -4, 13, -3, 12, -4, -10, -4, 4,
    -- filter=31 channel=1
    -5, -6, 3, -4, -7, 6, 8, -10, -4,
    -- filter=31 channel=2
    7, -5, 10, -4, 0, 6, 2, -10, 12,
    -- filter=31 channel=3
    -2, 6, 9, 3, 10, 12, 0, -8, 12,
    -- filter=31 channel=4
    0, -12, 0, 0, -9, 6, -1, -10, 11,
    -- filter=31 channel=5
    12, 7, 9, 6, -11, 13, 6, -6, -12,
    -- filter=31 channel=6
    3, -7, 4, 1, 14, -10, -11, 0, 6,
    -- filter=31 channel=7
    -9, 0, -2, 6, 2, 5, 12, -9, 2,
    -- filter=31 channel=8
    -4, 8, -7, -14, 7, -3, -14, 4, 5,
    -- filter=31 channel=9
    0, 7, -12, -7, 3, 2, -7, -7, 0,
    -- filter=31 channel=10
    4, -9, 13, -14, -6, -13, 7, 13, -6,
    -- filter=31 channel=11
    -12, 13, 13, 0, -13, 4, -11, 7, -9,
    -- filter=31 channel=12
    -5, -12, -10, 0, -8, 11, 0, -9, -8,
    -- filter=31 channel=13
    -14, -12, -2, -14, 10, -2, 5, 6, -11,
    -- filter=31 channel=14
    13, -11, -12, 8, -3, 6, 9, 0, 14,
    -- filter=31 channel=15
    -4, 9, -14, 13, 8, 4, 9, -2, -1,
    -- filter=31 channel=16
    13, -13, 4, 0, 0, -7, 13, 3, -5,
    -- filter=31 channel=17
    6, 1, 1, -3, -3, 10, 9, -10, 0,
    -- filter=31 channel=18
    -1, 11, -1, 4, -9, 0, -14, 6, -1,
    -- filter=31 channel=19
    1, 11, -10, -4, -11, -7, -13, 14, 11,
    -- filter=31 channel=20
    -8, -5, 3, 0, 12, 6, -8, 9, 7,
    -- filter=31 channel=21
    2, -6, 4, -11, -4, -5, 14, -3, 3,
    -- filter=31 channel=22
    7, 12, -12, -2, 5, -3, -3, -2, 9,
    -- filter=31 channel=23
    -5, 9, -11, 11, 14, -13, 4, 0, 0,
    -- filter=31 channel=24
    -1, 0, -8, -1, -9, -9, 0, -12, -13,
    -- filter=31 channel=25
    -7, 12, -5, -12, -7, -1, 5, 10, 10,
    -- filter=31 channel=26
    1, 2, 0, -5, 11, -2, 4, 0, 1,
    -- filter=31 channel=27
    0, 8, 10, 0, 0, -4, 5, 1, -8,
    -- filter=31 channel=28
    -11, 8, 6, -7, -12, -8, 4, 8, -2,
    -- filter=31 channel=29
    -13, 1, 12, -6, -8, -13, 0, 4, 12,
    -- filter=31 channel=30
    -4, 6, 8, -14, 10, 15, 6, -3, 9,
    -- filter=31 channel=31
    -6, 9, -4, 14, 4, 7, -11, 2, 12,
    -- filter=32 channel=0
    8, -9, -5, 7, 9, -9, -10, -11, -5,
    -- filter=32 channel=1
    10, 6, 9, -9, -3, 8, -11, 7, 13,
    -- filter=32 channel=2
    3, -19, -14, -25, -3, -24, 9, 6, -14,
    -- filter=32 channel=3
    0, -5, -4, 4, -4, -3, -10, 0, 3,
    -- filter=32 channel=4
    19, 18, 11, 13, -1, 29, 2, 3, 32,
    -- filter=32 channel=5
    4, -2, 6, -2, -4, -11, 9, -1, -8,
    -- filter=32 channel=6
    -7, 0, -5, -12, 0, -13, -14, 6, 4,
    -- filter=32 channel=7
    7, -5, 1, -18, -15, -11, -11, -11, -2,
    -- filter=32 channel=8
    -5, 3, -2, -1, 23, 13, 18, 20, 7,
    -- filter=32 channel=9
    -8, -22, 3, -4, 3, -19, -16, -10, 1,
    -- filter=32 channel=10
    5, 7, -18, 4, -13, 7, -9, -9, -15,
    -- filter=32 channel=11
    -9, -1, -6, 13, -9, 3, 7, -1, -11,
    -- filter=32 channel=12
    13, 0, 10, 0, 5, -5, 6, 0, 25,
    -- filter=32 channel=13
    10, 0, -8, -3, -22, 1, -2, -7, -13,
    -- filter=32 channel=14
    13, -3, 12, 15, 6, 21, 22, 21, 30,
    -- filter=32 channel=15
    2, -1, -5, 4, -1, 5, 9, 2, -14,
    -- filter=32 channel=16
    8, 1, -13, 3, 7, -3, -7, 9, 13,
    -- filter=32 channel=17
    -18, -7, 9, -3, -16, 0, -10, 9, 16,
    -- filter=32 channel=18
    -11, -9, 4, 0, -9, 9, -4, -9, -8,
    -- filter=32 channel=19
    0, 0, -4, 0, 2, 11, -2, 12, 11,
    -- filter=32 channel=20
    -11, 2, -7, -2, -8, 3, -1, -2, -1,
    -- filter=32 channel=21
    2, -23, -17, 2, 1, -26, -17, -8, -10,
    -- filter=32 channel=22
    6, 2, 4, -13, 0, 1, 7, 15, -7,
    -- filter=32 channel=23
    17, 5, 14, 2, 9, 24, 13, 28, 36,
    -- filter=32 channel=24
    -17, -27, -14, -11, -3, -2, -19, 6, 4,
    -- filter=32 channel=25
    12, 2, -6, 13, -1, 8, 13, 0, 13,
    -- filter=32 channel=26
    -4, -21, -18, 0, -24, -9, -21, -6, -18,
    -- filter=32 channel=27
    1, -10, 1, 10, 8, -4, -5, -2, -3,
    -- filter=32 channel=28
    1, -1, -11, 9, -14, 15, 9, 3, 0,
    -- filter=32 channel=29
    -2, 0, 9, -5, 12, 8, -3, 6, 3,
    -- filter=32 channel=30
    -17, -4, 2, 0, 9, -2, 0, -6, -7,
    -- filter=32 channel=31
    -6, 2, 13, 14, -1, 11, 0, -6, -9,
    -- filter=33 channel=0
    13, 12, 4, 1, 3, 0, -2, -8, 5,
    -- filter=33 channel=1
    7, 2, -12, 13, -2, -11, 8, 0, 1,
    -- filter=33 channel=2
    9, 15, -13, 14, -12, -14, -2, -14, -4,
    -- filter=33 channel=3
    -5, -16, 10, 7, -11, 9, 15, 7, -12,
    -- filter=33 channel=4
    8, 16, 11, 12, 17, 8, 5, -14, -12,
    -- filter=33 channel=5
    15, 10, 1, 6, 3, -1, -12, 5, 15,
    -- filter=33 channel=6
    6, 5, -3, 3, -12, 6, -4, -11, 5,
    -- filter=33 channel=7
    -1, -9, -2, -1, 8, -5, -4, -21, -10,
    -- filter=33 channel=8
    -2, 1, -3, -5, -3, 4, -18, 3, 3,
    -- filter=33 channel=9
    3, 4, 6, -6, 7, 2, -13, 7, -1,
    -- filter=33 channel=10
    4, 0, -16, -12, 3, 6, -12, -3, 3,
    -- filter=33 channel=11
    7, -1, 5, -9, 7, -12, -8, -6, 10,
    -- filter=33 channel=12
    -2, 18, 10, 5, -9, 4, 1, -19, -16,
    -- filter=33 channel=13
    -6, -1, 2, -8, -14, 5, -1, 0, 1,
    -- filter=33 channel=14
    22, 15, 11, 0, -5, -9, 0, -9, -5,
    -- filter=33 channel=15
    8, -14, -6, -13, -13, -8, -14, 6, 7,
    -- filter=33 channel=16
    12, 0, -12, 14, 6, 8, -10, 2, -7,
    -- filter=33 channel=17
    -12, 5, 0, -8, -16, 10, 5, -12, 8,
    -- filter=33 channel=18
    13, -1, 9, 13, 5, -12, -12, 14, -8,
    -- filter=33 channel=19
    -7, -13, 14, 14, -7, 1, 2, 7, 3,
    -- filter=33 channel=20
    7, 7, -13, -11, -10, 2, 7, -6, 12,
    -- filter=33 channel=21
    -16, 3, -6, 12, 3, 6, -15, 11, 6,
    -- filter=33 channel=22
    -6, 5, 0, 9, 9, -12, -6, 12, -15,
    -- filter=33 channel=23
    22, 12, 21, 10, 14, 23, -21, -29, -16,
    -- filter=33 channel=24
    12, -15, -3, -10, -5, -17, -5, -3, -4,
    -- filter=33 channel=25
    2, -14, 0, -6, -1, -13, -3, 0, -5,
    -- filter=33 channel=26
    4, -4, 4, 13, -11, 9, 0, -7, 6,
    -- filter=33 channel=27
    -6, -6, 10, -13, -11, -8, -5, 8, 8,
    -- filter=33 channel=28
    11, -5, -9, -10, 11, 7, -12, -1, 13,
    -- filter=33 channel=29
    14, 0, -6, 14, 2, 14, 0, 8, -15,
    -- filter=33 channel=30
    -8, 5, -2, -12, -5, -4, -5, 6, -4,
    -- filter=33 channel=31
    -1, 5, -8, 4, 4, 3, -6, 0, 1,
    -- filter=34 channel=0
    -6, -2, 6, 0, 10, -3, -2, 3, 14,
    -- filter=34 channel=1
    14, 3, 10, 0, -10, 3, 9, 2, -8,
    -- filter=34 channel=2
    0, -14, 14, -13, 1, 0, -8, 0, -2,
    -- filter=34 channel=3
    6, 4, 8, 4, -6, 2, -9, 14, -4,
    -- filter=34 channel=4
    13, 0, 14, -6, 0, 0, -3, -10, -11,
    -- filter=34 channel=5
    0, 5, -12, 14, 6, 3, -14, 2, -9,
    -- filter=34 channel=6
    -2, 0, 4, -9, 0, 2, -8, 2, -8,
    -- filter=34 channel=7
    0, 9, 6, 10, 3, 5, 12, -14, 8,
    -- filter=34 channel=8
    -4, 3, 1, 12, -7, -6, -8, 7, -4,
    -- filter=34 channel=9
    -4, -8, 7, -8, 1, -6, 12, -2, -11,
    -- filter=34 channel=10
    0, -6, 2, -13, -2, -4, -1, -7, -5,
    -- filter=34 channel=11
    -1, 3, -2, -1, 14, -13, 9, 2, -3,
    -- filter=34 channel=12
    -5, -12, 0, 5, -7, 10, 3, -5, 0,
    -- filter=34 channel=13
    0, 10, -8, -5, 4, 1, -2, -7, -5,
    -- filter=34 channel=14
    8, -4, 0, -4, 0, 6, 0, 6, 8,
    -- filter=34 channel=15
    -7, 14, -3, 7, 3, -2, -4, -6, 5,
    -- filter=34 channel=16
    -4, -10, 11, -7, 0, 5, 13, 3, 1,
    -- filter=34 channel=17
    3, -8, -4, 11, -14, 8, 7, 5, 11,
    -- filter=34 channel=18
    3, 5, 11, -1, 0, -6, -14, -12, -5,
    -- filter=34 channel=19
    -10, -1, -8, -11, 5, -11, -9, -12, 0,
    -- filter=34 channel=20
    3, 0, 13, -10, -6, 6, 3, 14, 13,
    -- filter=34 channel=21
    5, -13, -9, 7, -13, 10, 2, -10, -8,
    -- filter=34 channel=22
    -14, -14, -4, -5, 10, -5, 14, 1, 1,
    -- filter=34 channel=23
    7, -1, -12, -9, 3, -14, 0, -6, 10,
    -- filter=34 channel=24
    6, -13, 14, -12, -14, 3, -10, -6, 1,
    -- filter=34 channel=25
    1, -14, 0, 12, -1, -11, -2, -1, -3,
    -- filter=34 channel=26
    -2, 13, -9, 2, -6, 0, -7, 3, -13,
    -- filter=34 channel=27
    -9, -14, -10, -7, 11, -10, -4, 1, 0,
    -- filter=34 channel=28
    7, 6, -8, 8, -6, -13, 5, 3, 14,
    -- filter=34 channel=29
    0, -4, -8, -2, 2, 0, -11, 14, 0,
    -- filter=34 channel=30
    -1, -11, 13, 4, -4, -9, 5, 9, 3,
    -- filter=34 channel=31
    -6, 10, 0, 2, 4, -3, -10, -13, -8,
    -- filter=35 channel=0
    2, -9, 12, 8, 1, -2, 11, -8, 9,
    -- filter=35 channel=1
    14, -1, -13, -3, -11, -1, 4, 4, 1,
    -- filter=35 channel=2
    -14, 0, -17, -3, -12, -7, 6, -16, 8,
    -- filter=35 channel=3
    -9, -2, 3, -12, -9, 0, 9, 12, 1,
    -- filter=35 channel=4
    -6, -1, 0, 2, 16, 26, 2, 21, 5,
    -- filter=35 channel=5
    8, -2, 13, -15, 11, -7, -4, 7, -5,
    -- filter=35 channel=6
    13, -7, -6, 7, -9, -5, 1, -1, 17,
    -- filter=35 channel=7
    -9, 1, -13, -3, 5, -13, -3, -13, 9,
    -- filter=35 channel=8
    1, 6, 13, -7, 12, 17, -5, 15, 19,
    -- filter=35 channel=9
    -16, -10, -15, -14, -14, 12, -11, -14, -11,
    -- filter=35 channel=10
    6, 3, -11, 5, -8, -1, 12, -4, 9,
    -- filter=35 channel=11
    7, -10, 12, 12, 9, 9, -5, -9, -6,
    -- filter=35 channel=12
    -3, -8, 16, -13, -8, 2, -9, 9, 6,
    -- filter=35 channel=13
    7, 9, -12, 8, -19, -6, -8, -17, -4,
    -- filter=35 channel=14
    10, 12, 13, 7, 4, 6, -3, 3, 29,
    -- filter=35 channel=15
    0, 14, -4, -8, 6, -3, -13, -3, 8,
    -- filter=35 channel=16
    6, 13, 15, 8, 6, 8, 10, -3, 14,
    -- filter=35 channel=17
    -8, 5, 1, -9, -12, 19, 17, -11, 1,
    -- filter=35 channel=18
    -2, -2, -6, 15, -9, 0, 11, 11, 13,
    -- filter=35 channel=19
    -9, 17, 6, 4, 17, 3, 0, 0, 27,
    -- filter=35 channel=20
    -12, 8, 7, 14, -13, -5, 3, -11, -2,
    -- filter=35 channel=21
    6, 9, -5, -5, 0, -16, -5, -13, -13,
    -- filter=35 channel=22
    -3, 10, 8, 0, 8, -6, 12, -1, 16,
    -- filter=35 channel=23
    -4, 2, -1, 4, 10, -1, -8, 2, 5,
    -- filter=35 channel=24
    -3, -9, 5, -2, 5, -6, 16, -8, -13,
    -- filter=35 channel=25
    10, -9, 12, -11, 14, 8, -1, -8, 13,
    -- filter=35 channel=26
    4, 5, -11, 6, -16, 12, 10, -8, 11,
    -- filter=35 channel=27
    9, -13, 6, 1, -12, 3, -4, -3, -3,
    -- filter=35 channel=28
    0, 11, 0, 4, 11, 8, 14, 11, 9,
    -- filter=35 channel=29
    0, 9, -11, 6, -5, 4, -14, 6, 7,
    -- filter=35 channel=30
    5, -5, -6, -12, -1, -10, 15, 4, 9,
    -- filter=35 channel=31
    9, -3, 4, -1, 0, -13, -10, 12, -11,
    -- filter=36 channel=0
    4, -1, 8, -12, 12, 4, -12, 1, 10,
    -- filter=36 channel=1
    8, -7, -12, 4, -13, -7, -2, -12, 13,
    -- filter=36 channel=2
    -7, 12, -13, 11, -9, 1, -6, -14, -14,
    -- filter=36 channel=3
    -6, 14, 4, -12, -13, 3, -5, -14, -11,
    -- filter=36 channel=4
    3, -12, -12, 6, 13, -2, -4, 8, -3,
    -- filter=36 channel=5
    -11, -9, 0, -10, -8, 6, 14, 1, 7,
    -- filter=36 channel=6
    3, 2, -7, -5, -9, -7, 1, -11, -5,
    -- filter=36 channel=7
    6, 0, 0, 8, 6, -14, -13, -5, 11,
    -- filter=36 channel=8
    -8, -8, 7, -10, 1, -9, -6, 5, 9,
    -- filter=36 channel=9
    -12, 8, 9, 5, -6, -4, -4, -13, 8,
    -- filter=36 channel=10
    11, 7, -8, 1, 8, -11, -12, -4, 14,
    -- filter=36 channel=11
    3, 2, -5, -3, 9, 4, 12, 4, -4,
    -- filter=36 channel=12
    12, 11, 6, -1, -1, -8, 0, 1, -12,
    -- filter=36 channel=13
    -8, -9, 13, 9, -14, -3, 8, -10, 2,
    -- filter=36 channel=14
    3, 7, 13, -2, 1, -15, -13, -12, 1,
    -- filter=36 channel=15
    12, -6, -13, 10, -14, -13, 6, 0, 8,
    -- filter=36 channel=16
    -5, -6, 8, -12, -4, -8, -9, -11, 0,
    -- filter=36 channel=17
    7, 7, -12, -11, -15, -2, -3, 12, 11,
    -- filter=36 channel=18
    -8, 0, -6, -5, -5, 2, 7, 4, 0,
    -- filter=36 channel=19
    10, 8, -2, -9, -10, 4, -1, 1, 8,
    -- filter=36 channel=20
    9, 0, -6, -8, -13, 4, 10, 11, 14,
    -- filter=36 channel=21
    -1, -9, 12, 12, 10, -7, -13, -6, -10,
    -- filter=36 channel=22
    0, -3, -5, 0, -10, -7, 11, 14, -4,
    -- filter=36 channel=23
    -2, 2, 13, -6, -14, 1, 12, -6, 12,
    -- filter=36 channel=24
    4, -8, -8, -15, 7, 2, 1, 7, -5,
    -- filter=36 channel=25
    -10, 9, -8, 6, 0, -4, -2, 11, -11,
    -- filter=36 channel=26
    1, 2, -8, 13, -12, 10, -13, 8, 9,
    -- filter=36 channel=27
    -10, -13, 5, -1, 13, -3, 2, -1, -8,
    -- filter=36 channel=28
    -9, 14, -10, 7, 1, -7, 6, 11, 6,
    -- filter=36 channel=29
    -13, 0, 2, -6, 8, 7, -11, 8, -11,
    -- filter=36 channel=30
    -7, 13, -6, 14, -10, -13, -13, 0, 0,
    -- filter=36 channel=31
    -5, 14, -8, -6, -5, 13, 2, -13, 14,
    -- filter=37 channel=0
    11, -6, -2, 13, -13, -13, -10, -12, -9,
    -- filter=37 channel=1
    4, 6, 9, -4, 2, -8, 10, -1, -13,
    -- filter=37 channel=2
    10, 3, 3, 6, -4, 19, 13, 3, 23,
    -- filter=37 channel=3
    12, 12, -6, 12, 8, 2, 5, -12, -12,
    -- filter=37 channel=4
    6, -5, -10, -12, -14, -13, 5, -20, -3,
    -- filter=37 channel=5
    9, -1, -6, -6, 14, 12, 10, 7, -10,
    -- filter=37 channel=6
    -7, 6, 16, -10, 0, 5, 15, 11, -8,
    -- filter=37 channel=7
    18, 12, -3, 1, 11, 17, -5, -6, 7,
    -- filter=37 channel=8
    -2, 4, -13, -3, -19, 4, -10, -4, 0,
    -- filter=37 channel=9
    12, 16, -6, -6, -11, 11, 13, 0, 14,
    -- filter=37 channel=10
    1, 11, -8, 0, -10, 16, 3, -11, 6,
    -- filter=37 channel=11
    9, -6, -8, -8, 13, 8, -13, 6, 5,
    -- filter=37 channel=12
    -14, -9, 0, 5, -14, -16, -8, -15, -11,
    -- filter=37 channel=13
    -5, 10, 16, 6, 3, -3, 9, 3, 4,
    -- filter=37 channel=14
    -13, -11, 7, -4, -22, -8, 8, -13, -10,
    -- filter=37 channel=15
    -5, 3, -3, -6, 14, -10, 5, 0, 0,
    -- filter=37 channel=16
    14, 2, -1, 11, -2, 12, 16, 7, -4,
    -- filter=37 channel=17
    -1, 6, 11, 19, -2, 0, 19, 3, -4,
    -- filter=37 channel=18
    9, -9, -10, -5, 1, 8, -5, -4, 2,
    -- filter=37 channel=19
    -5, 3, 2, -13, -10, -6, 12, -12, 8,
    -- filter=37 channel=20
    0, 13, 19, -9, -10, 16, 11, 8, 18,
    -- filter=37 channel=21
    -7, 0, 11, 6, -7, 12, -2, 0, -3,
    -- filter=37 channel=22
    12, -14, -1, -3, 2, -13, 0, 11, 0,
    -- filter=37 channel=23
    -8, -14, 6, 0, -27, -4, -16, -15, -11,
    -- filter=37 channel=24
    3, 4, 8, -12, 13, 0, -8, 16, -4,
    -- filter=37 channel=25
    -8, 3, 7, 7, 7, -13, 11, -5, -11,
    -- filter=37 channel=26
    -4, 11, -1, 5, 0, 12, -2, 14, 0,
    -- filter=37 channel=27
    -5, 6, 12, -2, -5, -7, -3, 14, 10,
    -- filter=37 channel=28
    13, 10, -10, -2, -11, 7, 15, 3, -9,
    -- filter=37 channel=29
    -5, -3, 9, 5, -7, 2, -13, 8, -10,
    -- filter=37 channel=30
    -4, 14, -5, -1, 2, 2, 8, -1, -9,
    -- filter=37 channel=31
    -2, -4, -8, -13, -12, -9, 6, -9, 4,
    -- filter=38 channel=0
    0, 2, 2, 0, 13, 2, 14, 3, -3,
    -- filter=38 channel=1
    8, -10, 9, 6, -5, 13, 0, -1, -12,
    -- filter=38 channel=2
    10, -13, 3, -4, -21, 13, -3, -2, 13,
    -- filter=38 channel=3
    -7, 5, 13, -3, 15, 10, 6, 5, -11,
    -- filter=38 channel=4
    6, 2, -1, 1, 9, 1, 0, -6, 12,
    -- filter=38 channel=5
    -10, -9, -8, 3, 14, 11, 4, 10, 10,
    -- filter=38 channel=6
    -7, 0, 11, -13, 3, -12, 10, -6, -13,
    -- filter=38 channel=7
    -6, 7, 16, 10, -8, -7, -5, 4, 8,
    -- filter=38 channel=8
    -10, 1, 8, -8, -8, 0, 0, 8, -1,
    -- filter=38 channel=9
    -9, 1, 6, 3, -15, -5, -9, -4, -1,
    -- filter=38 channel=10
    9, 2, 2, 7, -3, -9, -13, -13, -1,
    -- filter=38 channel=11
    4, 0, 8, 7, 8, 3, 5, 3, -12,
    -- filter=38 channel=12
    13, -10, 0, 9, 0, 5, -11, -15, -12,
    -- filter=38 channel=13
    0, -4, -9, 3, 6, 11, 2, -7, 1,
    -- filter=38 channel=14
    1, 2, 14, 0, 3, -11, 14, -14, 5,
    -- filter=38 channel=15
    -2, 1, 3, 10, 9, 12, 4, -4, -5,
    -- filter=38 channel=16
    7, 4, -9, -2, -14, 4, -3, 7, -3,
    -- filter=38 channel=17
    5, 0, -13, -5, -10, -15, -3, 0, 16,
    -- filter=38 channel=18
    7, 10, 0, 12, 7, 5, 3, -14, 4,
    -- filter=38 channel=19
    5, -10, -9, -8, 8, 12, 6, 15, 7,
    -- filter=38 channel=20
    6, 9, 3, -3, 9, 1, -9, 14, -3,
    -- filter=38 channel=21
    4, -9, -10, 1, -6, -9, -2, -7, -3,
    -- filter=38 channel=22
    10, 1, 3, -4, 7, 11, 7, 6, 1,
    -- filter=38 channel=23
    3, 4, 20, 4, -6, 11, -9, -16, -2,
    -- filter=38 channel=24
    -7, 8, 19, -3, -17, 9, 16, -9, 9,
    -- filter=38 channel=25
    -8, -14, 2, -8, 12, -13, -9, -1, 12,
    -- filter=38 channel=26
    -3, -5, 6, -8, 12, 4, 11, 8, -1,
    -- filter=38 channel=27
    9, 9, 9, -6, 6, -12, -3, -10, -2,
    -- filter=38 channel=28
    5, -5, -3, -5, 5, -12, 5, 0, 0,
    -- filter=38 channel=29
    -2, 2, 0, -9, -5, -7, -6, 1, 13,
    -- filter=38 channel=30
    0, 6, 4, 7, -10, 11, 8, -7, 0,
    -- filter=38 channel=31
    14, 2, 8, -14, -6, -6, 4, -10, -1,
    -- filter=39 channel=0
    8, 2, -2, -11, 8, -9, -3, -10, 3,
    -- filter=39 channel=1
    13, 10, -11, -10, 4, 10, -5, -7, -5,
    -- filter=39 channel=2
    24, 28, 2, 13, 5, 23, -22, -39, -33,
    -- filter=39 channel=3
    4, 0, -3, -13, -3, -6, -1, -4, 11,
    -- filter=39 channel=4
    -10, -11, -13, 10, -2, 13, -12, -7, 8,
    -- filter=39 channel=5
    -6, 2, -3, -2, 12, 8, 12, 0, -6,
    -- filter=39 channel=6
    -9, -3, 8, -3, -8, -4, 0, 4, -6,
    -- filter=39 channel=7
    21, 4, -3, 16, -10, 14, -22, -16, -4,
    -- filter=39 channel=8
    -2, 0, 0, -6, 1, -1, 3, -2, -19,
    -- filter=39 channel=9
    13, 8, 4, 4, 14, 18, -15, -4, -8,
    -- filter=39 channel=10
    -7, -8, 14, -6, 15, -4, -14, -9, -11,
    -- filter=39 channel=11
    14, 5, -3, 13, 5, 15, -13, 0, -13,
    -- filter=39 channel=12
    16, 9, -5, -4, -7, 7, 1, -20, 8,
    -- filter=39 channel=13
    8, 16, -8, 3, -2, -9, 2, 0, -22,
    -- filter=39 channel=14
    3, 11, -6, 1, -7, 6, -11, -24, -7,
    -- filter=39 channel=15
    11, 4, 0, 0, -10, 13, -7, 0, -2,
    -- filter=39 channel=16
    -4, 4, -3, -8, 3, -1, -6, -8, -3,
    -- filter=39 channel=17
    21, 16, -6, -9, -2, 1, -18, -27, -8,
    -- filter=39 channel=18
    -9, -6, 14, 4, 12, 6, -8, -11, -9,
    -- filter=39 channel=19
    0, -1, 3, -6, 17, 17, -8, 2, 7,
    -- filter=39 channel=20
    14, -7, -7, -13, -6, 14, -11, -23, -15,
    -- filter=39 channel=21
    7, 7, -6, -14, -7, 17, -2, -9, 9,
    -- filter=39 channel=22
    -1, 15, -1, 17, 5, -9, 1, 3, 13,
    -- filter=39 channel=23
    -2, 6, 9, 8, 22, 4, 3, -6, 1,
    -- filter=39 channel=24
    11, 21, -1, -11, 3, 15, -12, -21, -21,
    -- filter=39 channel=25
    -13, -2, -9, 2, -9, 2, 0, -11, -9,
    -- filter=39 channel=26
    5, 20, 20, 10, 1, 17, -18, -13, -9,
    -- filter=39 channel=27
    8, 13, 2, 4, 12, 7, -9, 5, 13,
    -- filter=39 channel=28
    0, 12, 4, -7, 14, 11, -7, 9, 0,
    -- filter=39 channel=29
    12, 8, 6, -2, -7, -5, -7, 13, -12,
    -- filter=39 channel=30
    -3, -1, 4, -7, -8, -8, 3, 6, 8,
    -- filter=39 channel=31
    15, -1, 8, -9, -8, 6, 0, 12, 6,
    -- filter=40 channel=0
    11, 4, 7, 7, 6, -4, -12, 0, 13,
    -- filter=40 channel=1
    -9, 5, -6, -3, 2, 0, 5, -14, 0,
    -- filter=40 channel=2
    -1, 17, 2, -8, 0, 5, -21, 9, 16,
    -- filter=40 channel=3
    3, 10, 0, 2, -3, 2, 5, 12, -6,
    -- filter=40 channel=4
    9, -15, 2, 9, -14, -2, -3, -16, -2,
    -- filter=40 channel=5
    -10, 13, 7, -10, 19, 15, 5, -1, -9,
    -- filter=40 channel=6
    -6, 4, 19, -2, 10, -8, 14, 3, 8,
    -- filter=40 channel=7
    12, 12, 25, -17, 4, 1, -8, 16, 14,
    -- filter=40 channel=8
    13, 10, -1, 13, -12, 7, -12, -21, 2,
    -- filter=40 channel=9
    -3, 10, 18, 6, 15, -11, 10, -2, 12,
    -- filter=40 channel=10
    0, 16, 0, 7, 17, 12, -8, 15, 23,
    -- filter=40 channel=11
    -10, 3, 12, 3, 0, 7, 6, 12, 15,
    -- filter=40 channel=12
    13, 0, 8, 1, -8, -19, 3, -15, 5,
    -- filter=40 channel=13
    7, 14, 16, -12, 0, -2, -3, 20, 11,
    -- filter=40 channel=14
    6, 10, -4, -8, -11, -1, -10, 2, -19,
    -- filter=40 channel=15
    -2, -7, -10, 2, -7, -3, -3, 8, 2,
    -- filter=40 channel=16
    -9, 16, 0, -12, 7, -8, 12, 16, -2,
    -- filter=40 channel=17
    -3, 5, -2, -7, 6, 5, 14, 15, 19,
    -- filter=40 channel=18
    -4, -1, -5, -4, 6, 14, -11, -8, 0,
    -- filter=40 channel=19
    9, 12, 14, 0, -11, 4, 1, -5, 2,
    -- filter=40 channel=20
    -11, 3, 0, -10, -4, 4, 3, 10, 13,
    -- filter=40 channel=21
    -15, 13, -4, 0, 18, 0, -8, 22, 19,
    -- filter=40 channel=22
    0, -9, 0, 13, -2, -16, -13, -5, -12,
    -- filter=40 channel=23
    20, 0, 6, -8, -32, -30, -16, -19, -27,
    -- filter=40 channel=24
    -9, -2, 16, -17, 13, 10, -15, 15, 4,
    -- filter=40 channel=25
    13, 0, -12, -10, 7, -2, 9, -10, 6,
    -- filter=40 channel=26
    5, 15, 3, -1, 0, 24, -7, 15, 0,
    -- filter=40 channel=27
    13, 4, 8, -7, 4, 4, -12, -11, 8,
    -- filter=40 channel=28
    3, 12, -2, 9, -1, 8, -9, 6, -8,
    -- filter=40 channel=29
    10, 10, 4, 7, -11, 3, 2, 8, 4,
    -- filter=40 channel=30
    -10, 7, 7, -9, 4, 18, 4, -5, 16,
    -- filter=40 channel=31
    2, 13, 3, -13, -9, 10, 8, 3, 13,
    -- filter=41 channel=0
    2, 3, 7, -6, 10, 2, -10, 8, 13,
    -- filter=41 channel=1
    -4, 12, -10, -15, 7, -1, -10, -1, 12,
    -- filter=41 channel=2
    -16, -11, -27, -7, -11, 8, 21, 6, 22,
    -- filter=41 channel=3
    1, -7, 12, 9, 11, -14, -6, -12, -5,
    -- filter=41 channel=4
    0, -8, 12, -12, -10, 13, 6, -5, 13,
    -- filter=41 channel=5
    -4, -17, -13, -7, 2, -8, 9, -5, 8,
    -- filter=41 channel=6
    -11, 0, -17, 0, -2, 0, 4, -3, 3,
    -- filter=41 channel=7
    -1, -10, 1, -2, 2, -4, 12, 7, -2,
    -- filter=41 channel=8
    -4, -2, 6, -16, 7, -2, 10, 13, 13,
    -- filter=41 channel=9
    -16, -11, -14, -16, -4, -1, 0, 5, 9,
    -- filter=41 channel=10
    -15, 1, -8, -13, 6, -16, -1, 10, -1,
    -- filter=41 channel=11
    -5, -2, 10, -10, 12, 3, 8, -4, -8,
    -- filter=41 channel=12
    -7, 6, 11, -2, 4, 13, 11, 4, 19,
    -- filter=41 channel=13
    -10, -12, -1, -1, 3, 0, -3, 10, 16,
    -- filter=41 channel=14
    13, -4, -3, -11, -7, 13, 0, 3, 1,
    -- filter=41 channel=15
    -7, -7, -2, -6, -12, 2, -10, -14, 12,
    -- filter=41 channel=16
    12, -8, -6, 0, -5, 3, -8, -9, 14,
    -- filter=41 channel=17
    1, -7, 3, 1, -5, 0, 14, 8, 20,
    -- filter=41 channel=18
    8, 2, 2, 10, -3, -10, -9, 5, 11,
    -- filter=41 channel=19
    6, -13, -8, -8, 7, -6, -1, -20, -5,
    -- filter=41 channel=20
    4, -4, -6, -8, -8, -15, 1, 6, 9,
    -- filter=41 channel=21
    1, -19, -16, -12, -16, -11, -1, 13, 10,
    -- filter=41 channel=22
    3, -11, -8, -7, -3, 9, -1, -1, 1,
    -- filter=41 channel=23
    17, 11, 3, -14, -16, 5, -5, 20, 4,
    -- filter=41 channel=24
    -5, -6, -7, 5, 3, -14, 6, 10, 19,
    -- filter=41 channel=25
    9, -2, -7, -9, 14, -7, -3, 1, -15,
    -- filter=41 channel=26
    3, -23, -18, -12, 1, -1, 10, 14, 5,
    -- filter=41 channel=27
    -10, 3, 3, 7, 13, -13, -2, -13, 0,
    -- filter=41 channel=28
    -15, 13, -1, 8, -11, -3, -6, -4, -2,
    -- filter=41 channel=29
    -11, 7, 0, -9, -3, 5, 5, 10, 12,
    -- filter=41 channel=30
    10, -10, 0, -9, 1, 1, -11, -8, -6,
    -- filter=41 channel=31
    -8, 4, 12, 3, -12, 5, -12, -4, -2,
    -- filter=42 channel=0
    3, 7, 10, 13, -12, 7, -7, 6, -6,
    -- filter=42 channel=1
    -13, 6, 1, 15, 3, 1, -13, 8, 0,
    -- filter=42 channel=2
    26, 0, -48, 20, 9, -77, 18, -8, -54,
    -- filter=42 channel=3
    1, -6, -8, 15, 3, 16, 18, -7, -2,
    -- filter=42 channel=4
    4, 9, -11, -9, 10, -31, 21, -11, -9,
    -- filter=42 channel=5
    13, -10, 0, -1, -5, -3, 23, 5, 4,
    -- filter=42 channel=6
    25, -2, 0, 9, -3, 15, 6, 4, 0,
    -- filter=42 channel=7
    14, 4, -30, 8, 4, -42, 24, -7, -18,
    -- filter=42 channel=8
    5, 10, 5, 0, 9, -13, -1, -10, -1,
    -- filter=42 channel=9
    17, 2, -16, 13, 7, -36, 17, -18, -34,
    -- filter=42 channel=10
    14, -7, 14, 16, 3, 5, 8, 14, -7,
    -- filter=42 channel=11
    4, 5, -3, -6, -4, 2, -14, 10, -2,
    -- filter=42 channel=12
    8, 11, -10, 5, 7, 0, 22, -8, 9,
    -- filter=42 channel=13
    -1, 0, -17, 2, 10, -29, 20, 0, -14,
    -- filter=42 channel=14
    9, 7, -15, 17, -4, -30, 18, 4, 2,
    -- filter=42 channel=15
    -13, -12, 2, -7, 9, -3, 0, 0, 14,
    -- filter=42 channel=16
    2, 8, -17, 14, 7, -19, 27, 1, 6,
    -- filter=42 channel=17
    33, 25, -3, 32, 29, 9, 41, 28, 3,
    -- filter=42 channel=18
    1, 0, -4, 6, 1, 12, 12, 0, 0,
    -- filter=42 channel=19
    5, -3, 4, 31, -1, 16, 25, 0, 18,
    -- filter=42 channel=20
    9, 13, -15, 1, 12, -16, 16, -6, -12,
    -- filter=42 channel=21
    19, -5, -21, 7, 1, -5, 15, 12, -24,
    -- filter=42 channel=22
    2, 3, 16, 6, 8, -7, 7, 4, 5,
    -- filter=42 channel=23
    7, -8, -28, 4, -20, -47, 13, -12, -37,
    -- filter=42 channel=24
    13, 14, -16, 30, 3, -34, 13, 3, -13,
    -- filter=42 channel=25
    -11, -1, 1, 2, -12, -6, 12, 14, 5,
    -- filter=42 channel=26
    23, 24, 9, 19, 23, 4, 16, -1, -8,
    -- filter=42 channel=27
    14, 0, -3, -14, 10, -8, 11, -3, 5,
    -- filter=42 channel=28
    16, 4, -4, 16, 10, 9, -9, 6, 14,
    -- filter=42 channel=29
    14, -2, -10, -11, 13, 9, 14, 3, 13,
    -- filter=42 channel=30
    -2, -1, 13, 3, -1, 5, -8, -1, 0,
    -- filter=42 channel=31
    -1, -13, -11, 4, -12, 8, -8, 5, 1,
    -- filter=43 channel=0
    -11, 0, -13, -4, 11, 1, 5, -2, -13,
    -- filter=43 channel=1
    -8, 1, 12, 2, -6, -8, 15, 14, -4,
    -- filter=43 channel=2
    28, 17, 5, 23, -1, -10, 6, 6, -2,
    -- filter=43 channel=3
    3, -11, 0, -19, -7, 8, -8, -4, 7,
    -- filter=43 channel=4
    0, 11, 27, 21, 1, 8, -3, 22, 25,
    -- filter=43 channel=5
    6, -3, -14, -18, -18, -20, -1, -2, 1,
    -- filter=43 channel=6
    0, -20, -13, -6, -28, 5, -2, -24, -16,
    -- filter=43 channel=7
    0, -19, 2, -3, -25, 0, -6, -2, 3,
    -- filter=43 channel=8
    16, 13, 8, 19, 0, 4, 8, 0, 29,
    -- filter=43 channel=9
    -3, -11, 5, 11, 1, -15, 6, -13, -13,
    -- filter=43 channel=10
    -11, -11, -20, 0, 2, 6, -2, -20, 3,
    -- filter=43 channel=11
    -6, 2, -5, 11, 0, -10, 3, 12, 0,
    -- filter=43 channel=12
    2, 16, 23, 15, -8, 2, 15, 14, 14,
    -- filter=43 channel=13
    -3, -12, -6, -3, 0, -3, -1, -16, -8,
    -- filter=43 channel=14
    9, 11, 8, -10, 12, 4, 9, -4, -1,
    -- filter=43 channel=15
    -13, -2, 1, 6, 12, 14, -1, -7, 8,
    -- filter=43 channel=16
    -16, -6, 7, -8, -5, -10, 11, 1, -21,
    -- filter=43 channel=17
    -1, -28, -12, -19, -37, 4, -20, -4, -18,
    -- filter=43 channel=18
    -4, 3, -2, 8, -19, 7, -6, 9, -4,
    -- filter=43 channel=19
    -15, -37, -23, -7, -34, -29, -9, -33, -22,
    -- filter=43 channel=20
    -14, -23, -3, -6, -11, -12, 8, 0, -12,
    -- filter=43 channel=21
    -8, -20, -7, 5, -20, -18, 4, -20, -6,
    -- filter=43 channel=22
    9, -3, -6, 12, -13, 14, -2, 4, 8,
    -- filter=43 channel=23
    33, 21, 34, 31, 25, 34, 34, 13, 24,
    -- filter=43 channel=24
    -10, -5, -3, -4, -12, -19, -10, -1, -29,
    -- filter=43 channel=25
    1, -3, 4, 7, 3, -4, -4, -7, 8,
    -- filter=43 channel=26
    -1, -16, -13, -12, -29, -9, 0, -9, -18,
    -- filter=43 channel=27
    1, 9, 1, -4, 11, 2, -15, 8, -3,
    -- filter=43 channel=28
    6, 1, -5, 1, -23, 16, -7, -3, 13,
    -- filter=43 channel=29
    -8, 7, -3, -9, -5, 8, 5, -3, 2,
    -- filter=43 channel=30
    -22, -24, -22, -25, 0, 1, 1, -3, 0,
    -- filter=43 channel=31
    -6, -1, 3, -2, -15, -1, 5, 9, 10,
    -- filter=44 channel=0
    -6, 4, -8, 8, -2, -12, -8, 10, 9,
    -- filter=44 channel=1
    -1, 4, -10, -1, -13, 2, -6, 13, 0,
    -- filter=44 channel=2
    2, 18, -14, 6, 12, -24, 7, -2, 0,
    -- filter=44 channel=3
    4, -13, -13, 10, -14, 11, -1, 0, 14,
    -- filter=44 channel=4
    -13, -1, 3, -4, -8, -10, -4, -12, -1,
    -- filter=44 channel=5
    -6, -13, 1, 13, -11, -15, 7, -8, 5,
    -- filter=44 channel=6
    11, 1, 8, 7, -7, 2, 6, 0, 10,
    -- filter=44 channel=7
    -4, 6, -12, 11, 0, 2, -8, -8, 0,
    -- filter=44 channel=8
    3, 6, 0, -1, 5, 12, -6, -11, -10,
    -- filter=44 channel=9
    10, 14, 1, 1, -6, -19, 5, 0, -7,
    -- filter=44 channel=10
    -6, -4, -3, 4, 6, -14, -11, 12, 8,
    -- filter=44 channel=11
    -5, -14, 13, 9, 1, 7, 7, 6, -3,
    -- filter=44 channel=12
    -4, 10, -5, -13, 8, -11, -6, -8, 17,
    -- filter=44 channel=13
    5, 0, 9, 8, 12, -12, 2, 5, -3,
    -- filter=44 channel=14
    -5, -6, -4, 3, 0, 5, 8, 10, 18,
    -- filter=44 channel=15
    10, 6, -5, 9, -9, -1, -10, 5, -11,
    -- filter=44 channel=16
    -11, -9, 1, -13, -8, 12, 0, 4, -1,
    -- filter=44 channel=17
    8, -6, 9, -9, 11, -12, 0, 7, 15,
    -- filter=44 channel=18
    0, 1, 9, 13, 10, -11, -11, 0, 14,
    -- filter=44 channel=19
    -1, 0, 11, 7, -6, -1, 0, 9, -8,
    -- filter=44 channel=20
    1, 6, -11, -11, 3, -1, -14, -7, 10,
    -- filter=44 channel=21
    -13, 6, 11, 11, 7, -16, 1, 4, -2,
    -- filter=44 channel=22
    -15, -11, 1, 11, 11, 4, 13, 9, -8,
    -- filter=44 channel=23
    -14, 13, 13, -10, 0, 1, -4, 14, 9,
    -- filter=44 channel=24
    10, -11, 13, 2, -4, -3, -13, -9, -8,
    -- filter=44 channel=25
    -11, 0, 2, 14, -14, 0, 9, 8, -6,
    -- filter=44 channel=26
    4, -10, 3, 5, 7, -9, -11, 1, 3,
    -- filter=44 channel=27
    8, 13, 0, 7, 6, -1, 2, -3, 9,
    -- filter=44 channel=28
    -1, -12, -7, -8, -1, 3, -6, 11, -6,
    -- filter=44 channel=29
    2, 14, -3, -2, 11, -5, -5, -2, -8,
    -- filter=44 channel=30
    7, 5, 13, -6, 11, 8, -2, 14, -4,
    -- filter=44 channel=31
    10, 2, 5, -12, -2, -2, 2, -14, -5,
    -- filter=45 channel=0
    -1, 3, -8, -9, 4, 7, -4, 0, 1,
    -- filter=45 channel=1
    8, -15, 0, 7, 13, 0, 10, -1, 9,
    -- filter=45 channel=2
    25, 15, 31, 8, -17, 7, -33, -25, -7,
    -- filter=45 channel=3
    11, -10, 4, -15, 2, 6, 12, -12, -10,
    -- filter=45 channel=4
    -12, -4, -10, -11, -12, 11, -18, -4, 4,
    -- filter=45 channel=5
    12, -6, 10, -6, 7, 9, -16, 2, 1,
    -- filter=45 channel=6
    -7, 5, 18, -10, 3, 7, -10, -11, 6,
    -- filter=45 channel=7
    25, 9, 4, 3, 17, 16, -10, -19, -6,
    -- filter=45 channel=8
    4, 2, 2, 2, -5, -11, 4, -15, -7,
    -- filter=45 channel=9
    24, 20, -1, 14, -15, -2, -23, -24, -14,
    -- filter=45 channel=10
    19, 15, 16, 8, -10, 15, 4, 4, 10,
    -- filter=45 channel=11
    6, -13, 6, -14, -15, -6, -8, -14, 12,
    -- filter=45 channel=12
    -9, -6, 6, -14, 8, 9, -2, 0, 12,
    -- filter=45 channel=13
    0, 8, 7, 0, -8, 0, -15, 1, -8,
    -- filter=45 channel=14
    2, -18, 0, -2, 4, -1, -18, -3, 2,
    -- filter=45 channel=15
    6, 3, -12, 9, 4, 0, -6, -12, 2,
    -- filter=45 channel=16
    -4, 12, 4, -3, -7, -8, -6, -12, -9,
    -- filter=45 channel=17
    22, 13, 7, 14, -7, -16, -3, -24, 3,
    -- filter=45 channel=18
    -13, -17, 1, 11, 9, 1, -1, -13, 10,
    -- filter=45 channel=19
    -1, -21, -4, -12, 5, -16, -5, -8, 6,
    -- filter=45 channel=20
    11, 4, 0, 11, 15, 2, -3, 0, -1,
    -- filter=45 channel=21
    23, 21, 2, 8, -1, 6, -14, 6, -8,
    -- filter=45 channel=22
    0, -11, -10, -13, -10, 6, 9, 1, 0,
    -- filter=45 channel=23
    -1, 5, 2, -17, -4, -2, -6, 4, -2,
    -- filter=45 channel=24
    19, 18, 22, 11, -5, 1, -3, -8, -18,
    -- filter=45 channel=25
    -3, 5, -4, 0, -6, 10, 7, 13, 7,
    -- filter=45 channel=26
    2, 3, 8, 9, 8, 6, -19, -18, 0,
    -- filter=45 channel=27
    -12, -11, 9, -5, -4, -6, -13, -2, 6,
    -- filter=45 channel=28
    -10, -11, 6, 0, -11, 13, -9, -6, 1,
    -- filter=45 channel=29
    8, 6, -7, 12, 0, 0, 5, 0, -4,
    -- filter=45 channel=30
    -11, -4, 5, -7, -9, 7, -14, -15, 7,
    -- filter=45 channel=31
    12, -13, -2, 4, -15, -14, 14, 13, -13,
    -- filter=46 channel=0
    4, 10, 2, 2, 1, 6, -14, -2, 11,
    -- filter=46 channel=1
    13, 2, -5, 3, -14, 2, -7, 0, 1,
    -- filter=46 channel=2
    35, 16, 11, 5, -10, -5, 3, 0, 20,
    -- filter=46 channel=3
    11, -1, -2, -14, -12, 3, 4, 2, -1,
    -- filter=46 channel=4
    -16, 1, 9, -10, -8, 13, -7, -13, 21,
    -- filter=46 channel=5
    0, 7, -4, -2, -9, -18, 3, 0, 10,
    -- filter=46 channel=6
    0, 5, -11, -6, -7, -15, 10, -11, -3,
    -- filter=46 channel=7
    7, -6, 11, -7, -19, -7, 8, -4, -4,
    -- filter=46 channel=8
    3, 9, -5, 4, -13, -7, 3, 13, 20,
    -- filter=46 channel=9
    0, 8, 18, 0, 4, -7, 6, -5, -3,
    -- filter=46 channel=10
    1, 6, 9, -3, -12, -5, -7, 3, -9,
    -- filter=46 channel=11
    13, -1, -4, 7, 10, 0, 9, 12, 0,
    -- filter=46 channel=12
    0, -10, 10, -10, -1, -8, -1, 7, 8,
    -- filter=46 channel=13
    12, -15, 15, -12, 8, 8, 13, 10, -13,
    -- filter=46 channel=14
    -19, 3, 16, -17, 0, 11, -15, -6, -1,
    -- filter=46 channel=15
    0, 6, -15, 14, 0, 7, -5, 14, 12,
    -- filter=46 channel=16
    -9, -18, 10, -17, -11, 9, 0, 0, 11,
    -- filter=46 channel=17
    10, -16, -17, -22, -3, -10, 2, -1, -2,
    -- filter=46 channel=18
    -5, -12, -11, 5, -19, 0, 2, -10, -13,
    -- filter=46 channel=19
    -8, -22, -23, -13, -10, -16, -22, -12, 0,
    -- filter=46 channel=20
    -1, 10, -12, 4, 3, -15, -15, 10, -15,
    -- filter=46 channel=21
    10, -2, 1, 9, -10, 1, -5, -7, 16,
    -- filter=46 channel=22
    1, -13, 10, 8, 10, 10, 9, 5, 3,
    -- filter=46 channel=23
    -2, -3, 25, 3, 10, -4, 11, 7, 13,
    -- filter=46 channel=24
    21, 6, 16, -6, -10, 9, 2, -13, 4,
    -- filter=46 channel=25
    5, 2, 2, 5, -5, 5, -7, 8, -11,
    -- filter=46 channel=26
    7, 9, 0, 10, -3, -13, -12, -11, 8,
    -- filter=46 channel=27
    -14, 1, 8, 0, 1, 9, 8, -13, -4,
    -- filter=46 channel=28
    -11, -14, 2, -11, -4, -14, 6, -9, -8,
    -- filter=46 channel=29
    4, -7, 8, -4, 5, -5, -8, -4, 6,
    -- filter=46 channel=30
    9, -7, 3, 6, -20, -15, 11, 5, -15,
    -- filter=46 channel=31
    13, -11, 6, 0, -9, -14, -6, 11, 7,
    -- filter=47 channel=0
    9, -9, -11, -2, 10, -8, 7, 8, -10,
    -- filter=47 channel=1
    10, 2, -14, 12, -9, 12, -6, 0, -12,
    -- filter=47 channel=2
    -34, 7, 25, -28, -10, 26, -4, -21, 0,
    -- filter=47 channel=3
    6, -5, 2, 7, 3, -10, 0, 9, 5,
    -- filter=47 channel=4
    4, 0, 3, -19, -7, 0, -15, 5, 6,
    -- filter=47 channel=5
    0, 10, -5, 5, -9, -8, -6, 0, 2,
    -- filter=47 channel=6
    -6, -7, 16, -1, -13, 14, 8, -15, 6,
    -- filter=47 channel=7
    -4, -5, -2, -24, -6, -3, 6, -21, -1,
    -- filter=47 channel=8
    -18, -6, 21, -1, -14, 14, -7, -19, 4,
    -- filter=47 channel=9
    -3, 5, 5, -2, -2, 10, 8, -7, -12,
    -- filter=47 channel=10
    -12, -7, 7, -9, -8, -2, -4, -3, -11,
    -- filter=47 channel=11
    0, -10, 0, -13, 11, 7, 0, 11, 13,
    -- filter=47 channel=12
    -15, 13, 11, -1, 11, 9, 13, -21, -12,
    -- filter=47 channel=13
    -10, 12, 8, 1, -5, 8, -4, -18, 0,
    -- filter=47 channel=14
    -2, 1, 3, 6, -8, 0, -2, -17, 12,
    -- filter=47 channel=15
    -5, 12, 9, 14, 1, 9, 1, 11, -12,
    -- filter=47 channel=16
    1, 17, 18, 9, -8, 12, -6, -3, 9,
    -- filter=47 channel=17
    -14, 5, 17, -14, 6, 25, 18, -20, -6,
    -- filter=47 channel=18
    -12, 0, 13, 5, -9, -12, 6, 12, -7,
    -- filter=47 channel=19
    14, 12, 0, 19, 2, 6, 6, 7, 1,
    -- filter=47 channel=20
    2, -2, 7, 9, 11, -9, 3, 7, 6,
    -- filter=47 channel=21
    -17, -8, 12, 4, 6, 13, -6, 0, 9,
    -- filter=47 channel=22
    -12, 4, 12, 13, 10, -9, 0, -2, -14,
    -- filter=47 channel=23
    -4, -5, 20, -4, 18, 28, -6, -21, 0,
    -- filter=47 channel=24
    -22, 11, -5, -22, 5, 10, -8, -21, 10,
    -- filter=47 channel=25
    9, -14, 4, 1, 8, 5, -5, -2, 0,
    -- filter=47 channel=26
    2, 11, 16, -6, 1, 16, -10, 1, 8,
    -- filter=47 channel=27
    0, 9, -3, -8, 8, 4, 1, 11, -13,
    -- filter=47 channel=28
    0, -13, 16, 6, 6, 16, 12, -10, -2,
    -- filter=47 channel=29
    -6, 8, 4, -8, -9, 7, 0, -13, 6,
    -- filter=47 channel=30
    10, 8, 4, 14, 5, 4, -10, -13, -4,
    -- filter=47 channel=31
    14, 9, 5, 12, 8, 9, -3, -9, -7,
    -- filter=48 channel=0
    4, -3, 10, -8, 8, -5, -7, -10, 5,
    -- filter=48 channel=1
    -11, -12, 7, 11, 13, 0, 14, 0, -7,
    -- filter=48 channel=2
    1, 1, -2, 2, -14, -21, -6, 3, -4,
    -- filter=48 channel=3
    11, -8, 7, 2, 3, 4, 0, -18, 7,
    -- filter=48 channel=4
    -5, 0, 16, 3, 17, 18, 4, 26, 7,
    -- filter=48 channel=5
    0, -10, -21, -10, 6, 3, 0, 7, -16,
    -- filter=48 channel=6
    -17, -8, 11, 7, -21, 0, -16, -16, 4,
    -- filter=48 channel=7
    -16, -8, -12, -7, -7, -19, 11, -22, 5,
    -- filter=48 channel=8
    -7, 26, 4, 8, 9, 28, 8, 22, 12,
    -- filter=48 channel=9
    4, 8, -8, -13, -11, 0, 15, 11, -9,
    -- filter=48 channel=10
    4, -15, -13, 0, 6, -10, -10, 1, -4,
    -- filter=48 channel=11
    0, 2, -2, -5, -11, -12, 8, -12, -2,
    -- filter=48 channel=12
    4, -3, 24, -3, -5, -2, -8, 13, 23,
    -- filter=48 channel=13
    0, 3, -12, -6, 2, -8, 11, 0, 0,
    -- filter=48 channel=14
    9, 21, 2, 17, 19, 25, 10, 3, 14,
    -- filter=48 channel=15
    12, -8, 13, 1, 6, 8, -4, 11, 7,
    -- filter=48 channel=16
    0, 12, 12, 10, -15, 1, 4, 6, -11,
    -- filter=48 channel=17
    -17, -4, -7, -13, -22, 7, 0, 3, -5,
    -- filter=48 channel=18
    -4, 10, -10, -2, -2, -2, -4, 2, 10,
    -- filter=48 channel=19
    -17, 3, 10, -13, 7, -3, -1, 3, 1,
    -- filter=48 channel=20
    -10, -5, 6, 4, 8, -3, 11, -11, -6,
    -- filter=48 channel=21
    -4, -21, -11, -19, 2, -4, 8, -21, -1,
    -- filter=48 channel=22
    -11, -6, -9, 0, -8, 3, -13, 11, 8,
    -- filter=48 channel=23
    2, 8, 14, 17, 12, 18, 24, 7, 36,
    -- filter=48 channel=24
    -23, -15, -8, -15, -6, -19, 5, -14, -22,
    -- filter=48 channel=25
    -11, -5, -10, -9, -10, 13, 7, 6, 1,
    -- filter=48 channel=26
    -11, -25, -15, -16, -27, -24, -12, -15, -10,
    -- filter=48 channel=27
    1, 2, -13, 9, -8, -15, -10, -5, 3,
    -- filter=48 channel=28
    0, -13, 2, 1, 0, -2, 12, -12, 11,
    -- filter=48 channel=29
    1, -4, 11, 13, 0, -2, -1, 12, -6,
    -- filter=48 channel=30
    -2, -6, 6, -19, -13, -9, -2, -14, 1,
    -- filter=48 channel=31
    -9, -11, 3, -15, -14, 5, -1, 1, 13,
    -- filter=49 channel=0
    11, 3, 3, 12, 12, 2, 0, -12, -4,
    -- filter=49 channel=1
    8, 9, 2, -5, -5, -8, 0, 10, -12,
    -- filter=49 channel=2
    -3, -7, -11, -21, -24, -1, -12, 2, 13,
    -- filter=49 channel=3
    -9, 13, -8, -9, -9, 10, -15, -4, 5,
    -- filter=49 channel=4
    21, 5, 27, 13, -5, 7, 6, -4, 7,
    -- filter=49 channel=5
    2, -1, -6, 11, -1, -1, 14, 12, -5,
    -- filter=49 channel=6
    3, 4, -16, -2, -8, -4, 4, -6, 3,
    -- filter=49 channel=7
    13, 6, 8, 0, 0, -6, -16, -13, 1,
    -- filter=49 channel=8
    1, -4, 8, -6, 9, 7, -13, 0, 8,
    -- filter=49 channel=9
    12, 1, -5, -17, 1, -16, 4, 12, -15,
    -- filter=49 channel=10
    3, -5, -17, -17, -1, -8, -7, -3, -4,
    -- filter=49 channel=11
    11, -12, 5, -9, -9, 2, -11, 6, -6,
    -- filter=49 channel=12
    18, 0, 15, 3, -2, 14, -8, 11, -3,
    -- filter=49 channel=13
    -11, 0, -16, -19, -2, 0, 10, 3, 4,
    -- filter=49 channel=14
    10, 8, 5, 4, 0, 0, 8, -3, -5,
    -- filter=49 channel=15
    -12, -1, -13, -12, 4, 12, -13, 12, -14,
    -- filter=49 channel=16
    3, 11, 0, -11, -5, -1, 6, -11, -4,
    -- filter=49 channel=17
    -13, 0, -2, -18, -18, 6, 3, -4, 0,
    -- filter=49 channel=18
    6, 4, -1, -5, 8, 3, 6, 8, 7,
    -- filter=49 channel=19
    7, 13, -10, 10, 1, 10, -7, -14, 13,
    -- filter=49 channel=20
    -12, -4, -2, -6, 3, 5, -7, 3, -12,
    -- filter=49 channel=21
    -13, -19, -10, 0, -3, -4, 7, -5, -16,
    -- filter=49 channel=22
    6, 2, 11, 13, -2, -9, -5, 9, 4,
    -- filter=49 channel=23
    32, 30, 20, 11, -5, -1, 9, -1, 14,
    -- filter=49 channel=24
    9, 8, -15, -9, 2, -3, 2, -13, -13,
    -- filter=49 channel=25
    10, 8, -11, -11, 8, -4, 0, 1, -13,
    -- filter=49 channel=26
    -3, -5, 0, -9, -17, -1, -16, -16, -19,
    -- filter=49 channel=27
    11, -9, -9, -12, 5, -13, 11, -13, 6,
    -- filter=49 channel=28
    -8, 8, 2, -16, -15, 10, -11, 11, -11,
    -- filter=49 channel=29
    1, 6, -7, 3, -5, 9, -9, -3, 10,
    -- filter=49 channel=30
    -5, -12, 5, -13, 10, -2, 6, -9, -14,
    -- filter=49 channel=31
    -6, 11, 1, 4, 3, -5, -15, 6, -4,
    -- filter=50 channel=0
    13, 5, 5, -2, 10, -2, 8, 2, 9,
    -- filter=50 channel=1
    2, -1, -7, -13, -6, -5, 11, 12, -10,
    -- filter=50 channel=2
    -46, -36, -1, 14, 0, 5, 36, 30, 21,
    -- filter=50 channel=3
    -7, 12, 7, -2, 10, 5, 12, 11, 6,
    -- filter=50 channel=4
    -3, 4, -2, -8, -5, 7, 1, 3, 1,
    -- filter=50 channel=5
    4, -10, 0, 3, 9, 6, 1, 6, -11,
    -- filter=50 channel=6
    -5, -11, 4, 2, 7, -12, 20, 16, 7,
    -- filter=50 channel=7
    -35, -17, 0, 2, 0, -9, 27, 11, 2,
    -- filter=50 channel=8
    -17, 4, -15, 2, -16, -3, 1, 1, 12,
    -- filter=50 channel=9
    -21, -2, -6, 12, 12, 8, 0, 5, -8,
    -- filter=50 channel=10
    -11, -19, -18, 0, -10, 6, -4, 15, 16,
    -- filter=50 channel=11
    3, -7, -6, -13, -13, -9, -8, 15, 13,
    -- filter=50 channel=12
    -2, 8, -2, -9, -13, -16, 1, 6, 13,
    -- filter=50 channel=13
    -5, -15, 0, -5, 5, 14, -4, 12, -6,
    -- filter=50 channel=14
    4, 15, 8, -16, 6, -9, 16, 12, -8,
    -- filter=50 channel=15
    8, -10, 12, 3, -3, -6, -11, -4, 3,
    -- filter=50 channel=16
    -19, 6, -13, 13, 6, 5, 9, 6, -8,
    -- filter=50 channel=17
    -24, -28, -17, 8, 8, -14, 14, 0, -9,
    -- filter=50 channel=18
    4, 13, -2, 7, -11, -12, 12, 8, 10,
    -- filter=50 channel=19
    19, -6, 9, -2, -5, -15, -3, -19, -4,
    -- filter=50 channel=20
    2, 2, -1, -5, -14, 0, 17, 7, -12,
    -- filter=50 channel=21
    -21, -8, -6, -2, 2, 16, 21, -3, 16,
    -- filter=50 channel=22
    4, -15, -3, 4, -2, 12, 0, 8, 10,
    -- filter=50 channel=23
    -12, -13, -1, -28, -15, 3, 11, 11, 1,
    -- filter=50 channel=24
    -24, -29, -6, 20, -10, 3, 26, 20, 13,
    -- filter=50 channel=25
    6, 0, 14, 4, 2, 13, -7, 3, 0,
    -- filter=50 channel=26
    0, 0, -11, -11, -1, 13, 24, 4, 15,
    -- filter=50 channel=27
    -2, 14, 14, 8, -10, 3, 11, 15, -10,
    -- filter=50 channel=28
    -7, 2, 14, 0, -11, -2, -1, 11, -4,
    -- filter=50 channel=29
    -1, -11, 2, 6, 5, -11, -11, -4, -3,
    -- filter=50 channel=30
    -10, -4, 3, 4, -5, -2, -6, 7, -11,
    -- filter=50 channel=31
    15, -12, 13, 5, 6, -4, 7, -9, -6,
    -- filter=51 channel=0
    3, -7, 14, 9, 2, -7, 8, -14, 0,
    -- filter=51 channel=1
    -7, 3, 0, 14, 12, -14, -2, 1, -3,
    -- filter=51 channel=2
    15, -13, 4, -11, -18, 1, 27, 11, 36,
    -- filter=51 channel=3
    -5, 1, 13, 11, 10, -3, -4, -3, 0,
    -- filter=51 channel=4
    -3, 2, 10, 0, 1, -7, -14, 2, 12,
    -- filter=51 channel=5
    13, -5, 1, -16, -6, -17, 1, -15, -4,
    -- filter=51 channel=6
    6, -3, -13, -11, -7, 11, -12, 0, 9,
    -- filter=51 channel=7
    16, 4, 13, -14, 2, -8, 14, 16, 9,
    -- filter=51 channel=8
    11, -1, -3, 7, -11, 4, -7, -2, 5,
    -- filter=51 channel=9
    8, -7, -12, 8, -10, 8, 11, 16, 16,
    -- filter=51 channel=10
    1, 0, -10, -10, -1, -14, 11, 12, -3,
    -- filter=51 channel=11
    -7, 14, 14, -11, 12, 5, -9, -13, -6,
    -- filter=51 channel=12
    9, -2, 13, 1, 0, -16, -10, -7, 0,
    -- filter=51 channel=13
    1, 12, 8, -8, 11, 0, 12, 17, 9,
    -- filter=51 channel=14
    1, -2, 14, -3, -12, -14, -12, -8, 0,
    -- filter=51 channel=15
    10, -1, -8, -6, -4, -14, 4, 0, 11,
    -- filter=51 channel=16
    -1, 7, 8, -12, 6, 10, 0, 4, -3,
    -- filter=51 channel=17
    17, 2, 1, -13, 2, -17, -3, -9, -7,
    -- filter=51 channel=18
    1, -10, 4, 3, 7, 2, -10, -14, -8,
    -- filter=51 channel=19
    -6, -5, -5, -3, 0, -9, 4, -17, -2,
    -- filter=51 channel=20
    -6, 3, -4, -12, 0, 7, -6, 14, -3,
    -- filter=51 channel=21
    1, -3, -2, -9, -9, 14, 19, 16, 0,
    -- filter=51 channel=22
    0, 0, 12, -1, -9, -5, -8, -10, -2,
    -- filter=51 channel=23
    15, -12, 5, -18, -30, 2, -2, -10, -2,
    -- filter=51 channel=24
    16, -4, -5, -1, -9, -11, 23, 11, 28,
    -- filter=51 channel=25
    -13, 9, 2, 9, 14, -3, 0, 6, 9,
    -- filter=51 channel=26
    -7, -12, -13, 0, -1, 9, 16, 0, 1,
    -- filter=51 channel=27
    3, -1, 2, 11, 2, 7, 0, 7, -1,
    -- filter=51 channel=28
    -1, -10, -2, 3, 9, -4, -14, 4, 15,
    -- filter=51 channel=29
    -2, 5, 4, -12, -14, 0, 11, 7, -6,
    -- filter=51 channel=30
    -2, -10, 13, 15, -9, -4, -13, 12, -8,
    -- filter=51 channel=31
    -5, -8, -9, -9, 1, 4, -3, 0, -7,
    -- filter=52 channel=0
    14, -10, -4, -13, -9, -3, -7, -7, -12,
    -- filter=52 channel=1
    3, 5, 10, 11, -13, -12, -1, 13, 12,
    -- filter=52 channel=2
    -12, 4, -1, -19, 1, -16, -26, -30, -11,
    -- filter=52 channel=3
    -7, -4, 10, 11, -1, -10, 8, 0, -12,
    -- filter=52 channel=4
    3, 14, 0, 15, 23, 6, 4, 2, -1,
    -- filter=52 channel=5
    5, -3, 4, 0, 14, -4, -11, -11, 15,
    -- filter=52 channel=6
    2, -2, 5, 14, 14, -8, -9, 0, 6,
    -- filter=52 channel=7
    -7, -3, -19, -5, 1, 7, 2, -1, -8,
    -- filter=52 channel=8
    3, 25, -1, 2, 13, -15, 7, 4, 7,
    -- filter=52 channel=9
    -18, 4, -14, 5, 8, -13, -17, 0, 4,
    -- filter=52 channel=10
    -13, -7, -10, 2, -14, 3, 13, -5, 11,
    -- filter=52 channel=11
    6, -7, 3, -12, -2, -11, 0, 3, 0,
    -- filter=52 channel=12
    -4, 13, 10, 16, 23, -2, -3, -8, -14,
    -- filter=52 channel=13
    -6, 4, -12, -13, 4, 9, 8, -2, -5,
    -- filter=52 channel=14
    7, 20, 11, 13, 22, 7, 4, -3, -6,
    -- filter=52 channel=15
    -5, -9, -9, -13, 10, 12, 0, 10, -10,
    -- filter=52 channel=16
    -4, 16, 7, -7, 14, 1, -17, -11, -8,
    -- filter=52 channel=17
    -13, 9, -15, -3, -7, -13, 1, -18, -14,
    -- filter=52 channel=18
    -9, 2, 12, -2, -5, 11, 6, -4, 9,
    -- filter=52 channel=19
    -7, 10, 0, -8, 9, -13, 11, 10, 9,
    -- filter=52 channel=20
    8, -13, -12, 5, 12, 1, -7, -3, -10,
    -- filter=52 channel=21
    4, 1, -14, -15, -10, -1, 9, 0, 0,
    -- filter=52 channel=22
    -2, 15, 9, -8, 18, -5, 14, 7, 2,
    -- filter=52 channel=23
    18, 26, -6, 9, 24, -2, -17, 0, -6,
    -- filter=52 channel=24
    -16, -6, 8, 4, 4, 6, -4, -9, -7,
    -- filter=52 channel=25
    11, 1, 7, 9, 12, -14, 4, -10, -12,
    -- filter=52 channel=26
    -10, 9, 8, 4, 10, -18, -7, -17, -5,
    -- filter=52 channel=27
    2, 9, -1, 0, -3, 13, 13, -1, 3,
    -- filter=52 channel=28
    -13, -3, -2, -12, -4, 12, -8, 6, -3,
    -- filter=52 channel=29
    -8, 3, 14, 13, -6, 6, 8, 5, -12,
    -- filter=52 channel=30
    -6, -6, -13, 5, 11, 2, -7, 12, -5,
    -- filter=52 channel=31
    9, -9, 8, -2, -8, -10, 10, 0, 3,
    -- filter=53 channel=0
    -13, -13, -3, 8, -5, 9, 4, -2, -12,
    -- filter=53 channel=1
    -8, -10, 6, 1, 10, -2, 13, 2, 10,
    -- filter=53 channel=2
    8, 11, -13, 1, -1, 0, -15, -4, 12,
    -- filter=53 channel=3
    -5, -13, -14, 11, 10, 0, 3, 6, -14,
    -- filter=53 channel=4
    -11, -12, -2, -1, -10, 12, 3, -12, 6,
    -- filter=53 channel=5
    -14, 11, 9, -1, 8, -1, 13, 13, -12,
    -- filter=53 channel=6
    1, -12, 12, -4, 10, 14, -11, -4, -4,
    -- filter=53 channel=7
    0, 5, 4, 0, -13, 2, 3, -2, 4,
    -- filter=53 channel=8
    -13, 3, -14, -8, -3, -8, -9, -3, 13,
    -- filter=53 channel=9
    -7, 6, -9, 3, -10, 8, 13, -6, 10,
    -- filter=53 channel=10
    7, 3, -5, 2, -14, 4, -4, -15, -5,
    -- filter=53 channel=11
    -2, -8, 1, -3, 2, 13, 10, 0, 3,
    -- filter=53 channel=12
    -1, 14, 11, -12, 12, 9, -4, 2, 0,
    -- filter=53 channel=13
    -2, 12, -12, 0, 5, -7, 1, 9, 16,
    -- filter=53 channel=14
    -3, 8, 7, 9, -9, -8, -4, -6, 2,
    -- filter=53 channel=15
    4, 0, 9, 6, 1, 8, 11, 5, -7,
    -- filter=53 channel=16
    -3, -8, 14, -8, 12, 2, -10, 3, 16,
    -- filter=53 channel=17
    -5, 0, 7, -13, 0, 6, 14, -10, 13,
    -- filter=53 channel=18
    14, 0, -10, 10, 12, 7, 9, -1, -4,
    -- filter=53 channel=19
    -9, 11, -8, -4, 8, -6, -8, 11, 13,
    -- filter=53 channel=20
    -15, -11, 1, 9, -12, -4, 8, 2, 15,
    -- filter=53 channel=21
    -7, -12, 11, 9, -1, -9, 12, -8, 0,
    -- filter=53 channel=22
    8, -4, 5, 2, -3, -13, 7, 10, 10,
    -- filter=53 channel=23
    -3, 4, -7, 7, 3, -13, 1, -3, 0,
    -- filter=53 channel=24
    10, -7, -14, -2, -8, -4, -15, 6, -2,
    -- filter=53 channel=25
    1, -1, 0, -7, 0, 2, 13, 13, 2,
    -- filter=53 channel=26
    7, 5, 12, 2, -8, 9, 13, -4, -7,
    -- filter=53 channel=27
    7, 14, -12, 5, -3, -2, 8, -3, 12,
    -- filter=53 channel=28
    13, -2, -8, 11, 0, 3, -4, 8, -6,
    -- filter=53 channel=29
    -10, 15, -6, 0, -4, 0, 7, -10, 12,
    -- filter=53 channel=30
    -14, -7, 12, -8, 10, 13, -14, -11, 10,
    -- filter=53 channel=31
    0, -3, -14, 14, -2, -1, -1, 13, -1,
    -- filter=54 channel=0
    8, -12, -2, 5, 7, 7, 10, -10, 10,
    -- filter=54 channel=1
    0, 7, 10, -10, 8, 14, 14, -12, -12,
    -- filter=54 channel=2
    -6, -9, 10, 6, 11, 11, 13, 0, 12,
    -- filter=54 channel=3
    7, 3, -10, -3, 11, -2, 11, 4, 10,
    -- filter=54 channel=4
    0, -2, -7, -8, -6, -4, -14, -1, 7,
    -- filter=54 channel=5
    14, 13, 0, -3, -12, -8, 10, 6, -10,
    -- filter=54 channel=6
    5, -12, -1, -9, -7, -2, 2, 11, 14,
    -- filter=54 channel=7
    -4, 11, -10, -9, -11, 1, -6, -14, 3,
    -- filter=54 channel=8
    -4, 13, 7, -12, 2, -1, 5, 3, 3,
    -- filter=54 channel=9
    -12, -5, 14, -14, -6, -9, -2, 7, 7,
    -- filter=54 channel=10
    -3, 5, 1, -12, -8, -8, -2, -10, -8,
    -- filter=54 channel=11
    13, -10, 14, 2, 9, 6, 0, -6, -7,
    -- filter=54 channel=12
    14, 8, -15, -12, -7, 13, -9, -14, -14,
    -- filter=54 channel=13
    3, -8, 6, 0, 4, -12, 11, -3, -9,
    -- filter=54 channel=14
    -1, -6, 0, -11, 10, -8, -9, 1, 0,
    -- filter=54 channel=15
    1, -2, 7, -1, -13, -5, -12, 2, 2,
    -- filter=54 channel=16
    11, 0, -1, -11, -8, -5, -14, -9, -7,
    -- filter=54 channel=17
    -7, 7, -1, -13, 0, -15, -1, -11, 0,
    -- filter=54 channel=18
    12, 2, 3, 14, -4, 3, -7, 8, -7,
    -- filter=54 channel=19
    -4, -4, -9, -8, -1, 0, 2, -11, -1,
    -- filter=54 channel=20
    3, 14, -8, 3, -10, -7, -6, 5, -11,
    -- filter=54 channel=21
    0, -4, 7, -2, -10, -8, 3, -1, 0,
    -- filter=54 channel=22
    1, 4, 12, 8, 8, 4, 11, -12, -2,
    -- filter=54 channel=23
    9, -15, 2, -14, 13, -3, 0, 9, -12,
    -- filter=54 channel=24
    -15, 6, 3, 0, 9, -14, 12, 6, -8,
    -- filter=54 channel=25
    10, 5, -6, 3, 1, 7, -13, -8, 5,
    -- filter=54 channel=26
    3, 5, -13, -9, 7, 13, -9, -1, 8,
    -- filter=54 channel=27
    -2, 3, 0, -9, 6, 3, 13, 0, 13,
    -- filter=54 channel=28
    3, -12, 0, -4, -13, 10, 7, 13, -11,
    -- filter=54 channel=29
    10, -7, 5, -7, 10, -1, 2, 11, 6,
    -- filter=54 channel=30
    -12, -8, -1, -3, 2, 13, -6, 7, -14,
    -- filter=54 channel=31
    3, 4, -10, -14, -9, 5, 6, -10, 2,
    -- filter=55 channel=0
    1, -10, -6, 2, 0, -1, -3, 12, 8,
    -- filter=55 channel=1
    11, 0, 14, 13, -4, -4, -14, 9, 4,
    -- filter=55 channel=2
    0, -12, -25, 3, 4, -1, -23, -10, -5,
    -- filter=55 channel=3
    6, -10, 3, 8, -6, 4, 8, -9, 10,
    -- filter=55 channel=4
    11, 8, 9, -1, 11, 4, -6, 16, 24,
    -- filter=55 channel=5
    0, 6, 8, -11, -13, 4, 3, 1, 3,
    -- filter=55 channel=6
    10, -11, 11, -15, -19, 8, -16, -8, 9,
    -- filter=55 channel=7
    -1, -17, 2, -15, -24, -2, -16, -10, 0,
    -- filter=55 channel=8
    1, -2, 14, 17, 24, 23, -12, 20, 10,
    -- filter=55 channel=9
    10, -10, -5, -6, -11, -9, 1, 5, -10,
    -- filter=55 channel=10
    7, 7, 3, -15, 6, 0, -14, -11, -14,
    -- filter=55 channel=11
    3, 6, 13, -6, -10, 0, -6, -15, 9,
    -- filter=55 channel=12
    10, 3, 0, 15, 22, 0, -14, 9, 3,
    -- filter=55 channel=13
    -15, 6, -1, -3, -2, -13, -2, -7, 6,
    -- filter=55 channel=14
    -5, 23, 29, 15, 22, 3, -9, 15, 26,
    -- filter=55 channel=15
    -8, 1, -3, 1, -6, -13, -6, 6, -4,
    -- filter=55 channel=16
    -5, -1, -9, -1, -12, 8, -11, -11, -12,
    -- filter=55 channel=17
    -18, 3, -5, 5, -2, 11, -12, -10, 7,
    -- filter=55 channel=18
    5, -12, 4, 14, 8, -8, 9, 0, 14,
    -- filter=55 channel=19
    0, -7, -7, -9, -8, 1, 7, 11, -3,
    -- filter=55 channel=20
    1, -17, -4, 0, -13, 6, 9, -5, 9,
    -- filter=55 channel=21
    -16, -11, -9, 0, -21, -19, 3, -15, 4,
    -- filter=55 channel=22
    10, 11, 5, -10, 12, 9, 15, 6, 9,
    -- filter=55 channel=23
    12, 27, 21, 8, 7, 22, 12, 21, 28,
    -- filter=55 channel=24
    -14, -16, -12, -10, -25, -24, -19, -17, 1,
    -- filter=55 channel=25
    4, 2, -4, -13, -5, -2, 13, 12, -3,
    -- filter=55 channel=26
    0, -21, -13, -17, -5, 2, -13, -9, 6,
    -- filter=55 channel=27
    -15, 1, -9, 6, 8, 12, 1, -14, 0,
    -- filter=55 channel=28
    -2, -7, -5, 1, -4, -1, 11, -14, 14,
    -- filter=55 channel=29
    -5, -10, 10, 10, 11, 13, -7, -9, 11,
    -- filter=55 channel=30
    2, 1, -1, -2, -11, 0, -2, -5, -5,
    -- filter=55 channel=31
    -12, -4, -13, 8, 3, 12, -7, -13, 3,
    -- filter=56 channel=0
    4, 3, 6, 9, 4, -1, 10, 13, -5,
    -- filter=56 channel=1
    0, -1, 0, 9, -14, -4, 10, 1, -7,
    -- filter=56 channel=2
    18, 33, 5, 0, 1, 0, -20, -51, -40,
    -- filter=56 channel=3
    15, 1, 0, -1, 8, 11, 1, 12, 10,
    -- filter=56 channel=4
    -3, -2, 2, -4, 12, 13, 0, -12, 12,
    -- filter=56 channel=5
    -2, 14, -7, -1, 9, -13, -15, 1, 5,
    -- filter=56 channel=6
    13, 13, 9, 9, -7, 4, 18, 5, -11,
    -- filter=56 channel=7
    16, 6, 3, 8, 11, 7, 4, -20, -30,
    -- filter=56 channel=8
    9, 6, -8, -9, 1, -14, -12, -14, -16,
    -- filter=56 channel=9
    13, 10, -3, -12, 3, 7, -20, -5, -23,
    -- filter=56 channel=10
    21, 0, 13, 6, -8, 8, -10, -11, -12,
    -- filter=56 channel=11
    -10, 14, 3, -11, -10, -11, -9, -13, 9,
    -- filter=56 channel=12
    -12, 0, 3, -5, -8, -2, -14, -3, -8,
    -- filter=56 channel=13
    17, 20, 5, -9, -15, -12, -11, -7, -11,
    -- filter=56 channel=14
    -6, -2, 10, -2, -2, 7, 2, -10, 6,
    -- filter=56 channel=15
    13, 0, 0, 3, -14, 6, -9, 0, -7,
    -- filter=56 channel=16
    -8, -7, 6, -13, 10, 5, -3, -9, 8,
    -- filter=56 channel=17
    23, 0, 0, 9, -1, -13, 9, -17, 0,
    -- filter=56 channel=18
    4, 10, -4, 12, -10, -3, 16, -3, 5,
    -- filter=56 channel=19
    3, -10, 3, 15, 0, 11, -6, 16, 16,
    -- filter=56 channel=20
    18, 3, 4, -10, -12, 12, 12, -16, -15,
    -- filter=56 channel=21
    24, 6, 0, 2, -4, -6, -16, -18, 1,
    -- filter=56 channel=22
    -4, -6, 8, 4, -11, 8, 7, 1, 1,
    -- filter=56 channel=23
    10, 8, 13, -12, 18, 14, -19, -16, 0,
    -- filter=56 channel=24
    28, 7, 17, 9, 10, 2, -13, -11, -23,
    -- filter=56 channel=25
    -8, -13, -12, -3, 10, 11, -13, -5, 6,
    -- filter=56 channel=26
    20, 22, 5, 13, 0, 9, -6, -9, -17,
    -- filter=56 channel=27
    -7, -8, 0, 9, 1, -13, 3, 0, -9,
    -- filter=56 channel=28
    9, 12, 10, -5, -15, 7, 13, 1, 2,
    -- filter=56 channel=29
    -11, -5, 10, 11, -3, 0, 2, 5, 0,
    -- filter=56 channel=30
    4, -5, -4, 0, 0, 14, 13, 8, 10,
    -- filter=56 channel=31
    -3, -4, 14, 3, 11, 15, -6, -10, -2,
    -- filter=57 channel=0
    12, 2, 0, 0, -2, 0, -14, 8, -2,
    -- filter=57 channel=1
    1, 7, -9, 5, -4, 12, -11, -1, 2,
    -- filter=57 channel=2
    12, -13, 11, -11, 9, -10, -2, -13, 9,
    -- filter=57 channel=3
    -5, 7, -5, 7, -8, 8, 7, 6, 0,
    -- filter=57 channel=4
    15, -10, 8, 2, 6, 5, 0, -11, 12,
    -- filter=57 channel=5
    2, 1, 14, -1, 3, -7, 7, -4, -1,
    -- filter=57 channel=6
    8, -14, -2, 3, -1, -3, 5, -9, -9,
    -- filter=57 channel=7
    -6, 6, -13, -7, -11, -4, 6, 6, 12,
    -- filter=57 channel=8
    -8, -12, 11, 0, -13, -11, -5, -5, 0,
    -- filter=57 channel=9
    -9, 4, -9, -5, -11, -6, 9, -11, -8,
    -- filter=57 channel=10
    -13, -11, 6, 1, -12, 5, 13, 9, 0,
    -- filter=57 channel=11
    0, 1, 0, 4, -3, -14, 4, 2, -12,
    -- filter=57 channel=12
    -14, 7, -9, 10, 8, -3, -11, 9, 4,
    -- filter=57 channel=13
    -11, -5, -13, -4, 14, -6, -14, 3, -3,
    -- filter=57 channel=14
    -2, 9, -13, -7, 3, 5, 2, -1, 5,
    -- filter=57 channel=15
    12, -6, 2, 14, 10, 0, -8, 9, 1,
    -- filter=57 channel=16
    -13, 11, 14, -12, 10, -13, 9, -14, -5,
    -- filter=57 channel=17
    -12, -6, 4, -8, 10, 12, -5, 9, -12,
    -- filter=57 channel=18
    0, 0, -14, 4, -3, 14, 1, 9, -5,
    -- filter=57 channel=19
    9, -5, -3, -8, 5, -5, 1, -13, 12,
    -- filter=57 channel=20
    -5, -10, -6, -9, 9, -6, 4, -7, 3,
    -- filter=57 channel=21
    0, 7, 1, 5, -9, -5, 9, 9, 12,
    -- filter=57 channel=22
    -8, -5, 0, -7, -6, 1, -12, -5, -11,
    -- filter=57 channel=23
    -6, -12, 10, -10, -5, 5, 7, -2, 6,
    -- filter=57 channel=24
    -10, -5, -5, -1, 0, 8, 6, -10, -8,
    -- filter=57 channel=25
    9, -3, 8, 5, 6, 2, 13, 4, -7,
    -- filter=57 channel=26
    8, -1, 0, 0, -7, 7, 3, 1, -14,
    -- filter=57 channel=27
    5, -11, 14, 10, 2, 12, 0, 4, -11,
    -- filter=57 channel=28
    14, -14, -12, -2, 5, 7, -2, -6, -9,
    -- filter=57 channel=29
    7, -13, -10, 8, 6, 7, 11, 5, 3,
    -- filter=57 channel=30
    1, -8, -12, -4, -2, 3, 11, 6, -13,
    -- filter=57 channel=31
    -3, 2, -12, -3, -2, -9, 3, 0, 2,
    -- filter=58 channel=0
    0, -9, 8, 8, -12, 2, -8, 1, 0,
    -- filter=58 channel=1
    -3, -3, 11, -5, 0, -5, -6, 8, -11,
    -- filter=58 channel=2
    -13, -10, -2, -18, 6, 3, 6, -18, -19,
    -- filter=58 channel=3
    -9, 6, 14, 17, 15, 14, 16, 0, 0,
    -- filter=58 channel=4
    15, 2, 0, -13, -10, 9, 5, -3, -16,
    -- filter=58 channel=5
    4, 4, -9, -11, 17, 3, 12, 9, -9,
    -- filter=58 channel=6
    13, 18, 2, 9, -7, -8, -4, -3, 4,
    -- filter=58 channel=7
    7, 2, -13, -9, 12, -4, 3, -4, -15,
    -- filter=58 channel=8
    -9, 6, -12, -1, 11, 3, 4, -14, 0,
    -- filter=58 channel=9
    12, -12, -6, -13, 17, 12, 4, 0, -19,
    -- filter=58 channel=10
    -1, -13, -8, -11, 15, 3, 3, 17, 4,
    -- filter=58 channel=11
    -13, -2, -5, -7, -1, 10, -5, 10, 3,
    -- filter=58 channel=12
    -4, 4, 11, 12, -3, -5, -4, -6, 9,
    -- filter=58 channel=13
    -2, 8, 2, -7, 2, -6, 8, -14, 0,
    -- filter=58 channel=14
    3, 15, 3, 0, 1, 2, 6, 7, 10,
    -- filter=58 channel=15
    1, -2, -6, 12, 9, -14, -3, -13, -3,
    -- filter=58 channel=16
    0, -1, 14, 1, 14, 3, -9, -3, -6,
    -- filter=58 channel=17
    3, 10, 12, 11, 8, 16, -4, 13, 16,
    -- filter=58 channel=18
    -13, -4, -9, 7, -5, 8, -11, 12, 3,
    -- filter=58 channel=19
    7, 16, 11, 22, -1, -5, 17, 2, 15,
    -- filter=58 channel=20
    15, -5, 1, 8, 13, 4, -9, 0, -14,
    -- filter=58 channel=21
    -6, -2, 12, 13, 16, 0, -5, 10, -7,
    -- filter=58 channel=22
    7, 2, -6, -9, 0, -2, 6, 6, -9,
    -- filter=58 channel=23
    4, -2, -4, -11, -15, -12, 6, -16, -2,
    -- filter=58 channel=24
    14, 11, 0, 6, 16, 5, -13, -16, -6,
    -- filter=58 channel=25
    9, 14, -3, -3, 5, -10, -1, -11, -13,
    -- filter=58 channel=26
    -10, 20, 5, 4, 9, 13, 0, 10, -1,
    -- filter=58 channel=27
    -5, -12, -12, 10, 2, -6, 8, -11, 9,
    -- filter=58 channel=28
    10, 1, 15, 15, 7, 0, -6, 9, 1,
    -- filter=58 channel=29
    6, 10, 8, -8, 5, 14, -2, -6, 15,
    -- filter=58 channel=30
    11, 12, -3, -5, -8, 7, -4, 11, 9,
    -- filter=58 channel=31
    -6, -4, 11, -3, 3, -1, -4, -2, -10,
    -- filter=59 channel=0
    3, -7, 13, -5, 3, 9, 13, 4, 15,
    -- filter=59 channel=1
    -1, 11, 5, -14, 9, -9, -3, 5, -6,
    -- filter=59 channel=2
    12, 19, -19, 14, -10, -32, 14, -3, -29,
    -- filter=59 channel=3
    10, -4, -12, -1, 10, 5, 5, 2, 5,
    -- filter=59 channel=4
    18, 12, 11, -2, 8, -13, 10, -3, -17,
    -- filter=59 channel=5
    1, -12, 8, -4, 7, -9, 0, -14, 9,
    -- filter=59 channel=6
    0, 13, 4, 13, 10, 3, 11, 15, -13,
    -- filter=59 channel=7
    19, 0, -16, 17, -4, -24, 25, -14, 0,
    -- filter=59 channel=8
    0, -8, -1, 7, 6, -16, -5, -5, -6,
    -- filter=59 channel=9
    9, 12, -10, -7, -7, -10, 7, -4, -11,
    -- filter=59 channel=10
    -8, 10, -11, 10, -4, 7, 17, 10, 6,
    -- filter=59 channel=11
    2, 0, -2, -7, -4, -11, -8, 13, 0,
    -- filter=59 channel=12
    -4, 19, 2, 12, 3, -3, 0, 9, -11,
    -- filter=59 channel=13
    1, 13, -2, -8, 12, -18, 4, 10, -20,
    -- filter=59 channel=14
    -12, 17, -18, 0, -3, -15, 7, 5, -11,
    -- filter=59 channel=15
    -3, -7, 3, 12, -14, -2, -4, 0, 3,
    -- filter=59 channel=16
    0, -10, -16, 7, 0, 1, 19, -9, -15,
    -- filter=59 channel=17
    17, 0, 8, 22, -5, -7, 26, 4, 12,
    -- filter=59 channel=18
    14, 15, 5, -12, 0, 15, -8, 0, 1,
    -- filter=59 channel=19
    0, -5, 4, 19, 17, 1, -6, 16, 4,
    -- filter=59 channel=20
    -11, 10, -18, 14, 0, 1, 3, 11, 0,
    -- filter=59 channel=21
    13, -10, 1, 6, -3, -6, 19, -10, -15,
    -- filter=59 channel=22
    -11, -4, 0, -6, 17, 13, 10, 4, -4,
    -- filter=59 channel=23
    7, 0, -17, 2, 4, -22, -3, 5, 2,
    -- filter=59 channel=24
    15, 12, -8, 6, -2, -25, 5, 6, -14,
    -- filter=59 channel=25
    -6, 4, 9, -13, 0, -7, -7, 12, 11,
    -- filter=59 channel=26
    6, -8, 10, 3, 5, -20, -3, 7, 7,
    -- filter=59 channel=27
    -14, -8, -5, 1, -3, -12, 13, 9, 1,
    -- filter=59 channel=28
    2, -2, -8, 0, 18, -7, -8, 17, 17,
    -- filter=59 channel=29
    -10, 10, 2, -5, -11, -9, 3, -13, 0,
    -- filter=59 channel=30
    -9, -13, -6, -10, -1, 5, -7, -10, -7,
    -- filter=59 channel=31
    -9, -13, -8, -15, 6, 7, 11, -5, -5,
    -- filter=60 channel=0
    -2, -6, 12, 7, 3, -5, -9, -2, -12,
    -- filter=60 channel=1
    2, -1, 9, 5, 8, 0, 12, 8, 5,
    -- filter=60 channel=2
    -5, 19, -5, -2, 11, 7, -3, -2, 14,
    -- filter=60 channel=3
    7, 8, -3, 7, 3, 5, -8, -10, 13,
    -- filter=60 channel=4
    -16, -12, -9, -28, -21, 0, -10, -4, -8,
    -- filter=60 channel=5
    17, 0, 1, -1, -8, -1, 0, -11, -1,
    -- filter=60 channel=6
    18, 3, -12, -1, 11, 13, 7, 8, 0,
    -- filter=60 channel=7
    23, 2, 12, 18, 14, 6, 17, 6, -1,
    -- filter=60 channel=8
    -14, -6, 3, -24, -4, 11, -13, -18, 1,
    -- filter=60 channel=9
    11, 17, 5, 14, -5, 10, -6, -13, -10,
    -- filter=60 channel=10
    0, 10, 12, 18, -3, -2, 12, 15, 2,
    -- filter=60 channel=11
    2, 13, -3, 2, 13, 14, 0, 0, -9,
    -- filter=60 channel=12
    -17, 1, -18, -21, 0, 8, -12, -18, 12,
    -- filter=60 channel=13
    12, 18, 18, 0, 13, 1, 3, 2, -2,
    -- filter=60 channel=14
    -20, -14, 2, -21, -15, 6, 0, -15, 4,
    -- filter=60 channel=15
    1, -9, -1, -4, 1, 11, -14, 2, -12,
    -- filter=60 channel=16
    -11, -5, 8, 7, -5, -3, 7, 12, 3,
    -- filter=60 channel=17
    -2, 18, 9, 0, -7, 6, -4, 2, -17,
    -- filter=60 channel=18
    0, -14, 0, 7, -15, -4, -11, -5, -13,
    -- filter=60 channel=19
    9, 3, -17, -1, 2, -9, -13, 4, -1,
    -- filter=60 channel=20
    -8, -5, 12, 0, -1, 3, -3, -7, 14,
    -- filter=60 channel=21
    -4, 22, 0, 21, 2, 6, 16, -7, 5,
    -- filter=60 channel=22
    6, 7, -7, -10, -8, 6, 0, -6, -1,
    -- filter=60 channel=23
    -24, -19, -12, -11, -26, -1, -14, -5, -15,
    -- filter=60 channel=24
    18, 14, -2, 7, 3, -10, -9, -8, 2,
    -- filter=60 channel=25
    12, 5, 7, -4, -3, 12, 9, 4, -8,
    -- filter=60 channel=26
    5, 21, 14, 2, -4, 0, -9, 21, 15,
    -- filter=60 channel=27
    -12, -9, 8, -12, -11, -5, -11, 3, 10,
    -- filter=60 channel=28
    -5, 0, 11, 11, 6, 9, -5, -2, 12,
    -- filter=60 channel=29
    12, -7, -11, -3, -7, -7, 11, 7, -12,
    -- filter=60 channel=30
    14, 9, -10, 12, -7, -1, 12, -5, -10,
    -- filter=60 channel=31
    4, -15, 12, -13, 11, -14, -11, -9, 0,
    -- filter=61 channel=0
    -7, -2, -4, 9, -10, -14, 10, 8, -11,
    -- filter=61 channel=1
    9, 4, 9, 8, 0, 13, 1, -3, 2,
    -- filter=61 channel=2
    -14, -29, 24, -23, -19, 23, -3, -1, 12,
    -- filter=61 channel=3
    -2, -9, -3, 0, -5, 13, -4, 6, 15,
    -- filter=61 channel=4
    6, -7, 13, -19, 1, 11, -7, 6, 13,
    -- filter=61 channel=5
    -5, 13, -5, -9, -2, 5, -7, 12, 0,
    -- filter=61 channel=6
    10, 4, 13, 5, 0, 24, -1, 0, 15,
    -- filter=61 channel=7
    -1, -12, 8, -11, -14, 26, -10, -7, 11,
    -- filter=61 channel=8
    6, -9, -3, 1, 9, 10, -2, 4, -11,
    -- filter=61 channel=9
    -5, -21, 2, 7, -7, 8, -1, -8, 0,
    -- filter=61 channel=10
    1, -13, 0, 12, -19, -4, -10, -5, 18,
    -- filter=61 channel=11
    0, 10, -10, 8, -8, -2, -10, 8, -14,
    -- filter=61 channel=12
    1, 8, 8, -9, -4, 22, 6, 6, -10,
    -- filter=61 channel=13
    -4, 1, 16, 4, -19, 12, 0, -18, -7,
    -- filter=61 channel=14
    -2, 2, -3, -19, 10, 20, 2, 11, -6,
    -- filter=61 channel=15
    1, -9, 12, 0, 1, 14, -2, 8, -2,
    -- filter=61 channel=16
    10, 6, 5, 11, 17, 16, 2, 13, 15,
    -- filter=61 channel=17
    14, 3, 15, 14, -18, 22, 4, 6, 10,
    -- filter=61 channel=18
    -8, 5, -1, 0, -12, 7, -7, -1, -5,
    -- filter=61 channel=19
    -9, 29, 15, -3, 28, 2, 7, -3, 9,
    -- filter=61 channel=20
    0, -4, 10, 8, 5, 14, -8, 10, 2,
    -- filter=61 channel=21
    3, -16, 10, 11, -12, -3, -13, -2, 3,
    -- filter=61 channel=22
    6, -8, -1, -10, -10, 13, -3, -10, -1,
    -- filter=61 channel=23
    4, -4, -7, -21, -12, 18, -20, 6, -4,
    -- filter=61 channel=24
    4, -13, 15, -15, -20, 12, 0, -15, -2,
    -- filter=61 channel=25
    14, -4, 0, -12, 14, 4, 14, 8, -6,
    -- filter=61 channel=26
    -7, -17, 13, 5, -17, 21, 3, -1, 8,
    -- filter=61 channel=27
    13, 3, -11, 12, -11, -7, -6, -10, 7,
    -- filter=61 channel=28
    12, 15, -5, 1, 12, 9, 1, -9, -8,
    -- filter=61 channel=29
    -11, 0, -6, 14, 8, 5, 10, -12, 13,
    -- filter=61 channel=30
    2, 18, 0, -9, 2, -4, 14, 7, 2,
    -- filter=61 channel=31
    -1, 11, 2, 14, 6, -2, -10, 4, 14,
    -- filter=62 channel=0
    -12, 8, 1, 7, -5, -12, 2, 0, 7,
    -- filter=62 channel=1
    -13, 14, -6, -9, 1, 4, -4, 0, -11,
    -- filter=62 channel=2
    -6, -26, 0, 0, -25, 26, -15, -30, 46,
    -- filter=62 channel=3
    13, -7, 13, -9, 10, -10, -9, 2, 6,
    -- filter=62 channel=4
    -3, -5, -3, -16, 3, 15, 5, -20, 8,
    -- filter=62 channel=5
    10, 1, 20, -6, 0, 11, 12, 5, 23,
    -- filter=62 channel=6
    14, 0, -5, 0, 12, 0, -6, 1, 2,
    -- filter=62 channel=7
    16, 3, 0, -2, -23, 19, 0, -5, 24,
    -- filter=62 channel=8
    7, -6, -14, 9, -11, -5, -8, -20, -1,
    -- filter=62 channel=9
    6, 3, 13, 8, 0, 14, -16, -9, 30,
    -- filter=62 channel=10
    18, -4, 0, -7, -9, 7, 8, 0, -6,
    -- filter=62 channel=11
    -10, -5, -5, 6, 16, -3, 2, 7, -5,
    -- filter=62 channel=12
    -13, 8, -9, 5, -20, -5, 0, -22, 21,
    -- filter=62 channel=13
    3, -4, -4, 12, -18, 2, 1, -22, 9,
    -- filter=62 channel=14
    8, -9, -10, 3, -17, 16, 1, -1, 18,
    -- filter=62 channel=15
    0, -6, -11, -10, -5, 12, 2, -10, -12,
    -- filter=62 channel=16
    5, 5, 5, 5, 1, 17, -13, -4, 26,
    -- filter=62 channel=17
    -1, -4, 3, 0, -3, 17, -3, -7, 27,
    -- filter=62 channel=18
    9, -8, 14, 6, -4, 13, 13, 12, -7,
    -- filter=62 channel=19
    6, 4, 8, -9, 25, 11, 12, 17, 26,
    -- filter=62 channel=20
    -7, 2, 14, 4, -17, 0, 2, -16, 8,
    -- filter=62 channel=21
    13, -15, -12, 14, -10, -13, 9, -19, 2,
    -- filter=62 channel=22
    3, 14, 7, 11, -5, 13, 11, -15, 4,
    -- filter=62 channel=23
    -5, -17, 14, -11, -18, 30, -25, -1, 36,
    -- filter=62 channel=24
    -4, -9, 17, 4, -32, 5, 12, -11, 16,
    -- filter=62 channel=25
    6, -8, -11, 13, 4, -1, 1, 4, 0,
    -- filter=62 channel=26
    13, 10, 1, 18, -11, 3, 17, -17, 11,
    -- filter=62 channel=27
    0, 4, -9, 2, 10, -6, 1, 4, 5,
    -- filter=62 channel=28
    -9, 3, -5, -7, -1, 15, 16, 11, 2,
    -- filter=62 channel=29
    -12, 5, 10, 10, 9, 3, 9, -11, -14,
    -- filter=62 channel=30
    -8, 6, 0, -2, -4, -10, 7, -7, -8,
    -- filter=62 channel=31
    -8, 12, -5, -14, -10, 4, 15, -7, 4,
    -- filter=63 channel=0
    -2, 8, 0, -4, -2, 11, -8, -4, 10,
    -- filter=63 channel=1
    7, 9, 9, 9, -9, 9, -14, -11, -13,
    -- filter=63 channel=2
    -13, -10, 11, -12, 14, 9, 11, 16, 5,
    -- filter=63 channel=3
    -2, 2, 13, 7, -11, -9, 9, -3, 14,
    -- filter=63 channel=4
    -11, 5, -9, -7, -15, -5, -11, -7, -15,
    -- filter=63 channel=5
    -9, -10, 0, -15, -2, -4, -11, -5, -6,
    -- filter=63 channel=6
    10, -8, 0, -2, 6, -3, -5, -5, 7,
    -- filter=63 channel=7
    -8, 10, -6, 12, -11, 4, -2, 9, 0,
    -- filter=63 channel=8
    -12, -4, -11, -8, 7, -8, -15, -6, -7,
    -- filter=63 channel=9
    4, 12, -3, -12, -2, -11, 0, 9, 0,
    -- filter=63 channel=10
    -7, -9, 13, 9, 5, -3, 1, 6, -13,
    -- filter=63 channel=11
    -1, 0, -4, -6, 14, -2, 12, -8, 11,
    -- filter=63 channel=12
    -6, -14, -14, 7, 6, 2, -6, 7, -7,
    -- filter=63 channel=13
    10, 13, 0, 9, 9, 12, -13, 3, 0,
    -- filter=63 channel=14
    7, -6, -15, 5, 0, 9, 13, 11, -4,
    -- filter=63 channel=15
    0, -12, 4, 3, -10, 12, 11, 0, -9,
    -- filter=63 channel=16
    5, -7, 12, -5, -3, -7, -9, -2, 12,
    -- filter=63 channel=17
    4, -15, -13, -1, 10, -11, 5, 1, -7,
    -- filter=63 channel=18
    13, 1, 0, -1, 0, 12, 14, 7, -4,
    -- filter=63 channel=19
    0, -3, 6, 0, 13, 0, 5, -2, -15,
    -- filter=63 channel=20
    -14, -14, 0, -12, -14, 14, 14, -2, 11,
    -- filter=63 channel=21
    -9, 11, 2, -3, 1, -11, -12, 7, 6,
    -- filter=63 channel=22
    12, -1, -4, 5, 8, -8, 7, 2, 8,
    -- filter=63 channel=23
    10, 0, -9, -10, 6, -5, -13, 0, 3,
    -- filter=63 channel=24
    -11, -1, 11, 8, -9, -9, 6, 16, -10,
    -- filter=63 channel=25
    10, -14, -10, 0, 9, -4, 7, -14, -10,
    -- filter=63 channel=26
    -7, 9, -12, 11, 0, 7, -7, 6, 11,
    -- filter=63 channel=27
    10, -12, -7, 9, 2, -8, 0, 0, -13,
    -- filter=63 channel=28
    10, 3, 4, 4, 8, -12, -5, -13, -10,
    -- filter=63 channel=29
    3, -7, 11, 10, -13, 11, 3, 1, -2,
    -- filter=63 channel=30
    -2, -10, 4, 14, 0, 14, 3, -1, -11,
    -- filter=63 channel=31
    -12, -7, 14, -8, 3, 5, -13, 14, 5,

    -- ifmap
    -- channel=0
    29, 34, 33, 34, 34, 29, 30, 27, 
    4, 19, 32, 6, 27, 0, 22, 19, 
    0, 52, 0, 0, 14, 0, 0, 28, 
    0, 17, 21, 0, 13, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 
    22, 0, 0, 0, 0, 0, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 0, 
    22, 1, 3, 0, 0, 0, 6, 0, 
    
    -- channel=2
    89, 110, 240, 245, 154, 270, 122, 0, 
    384, 307, 519, 472, 421, 615, 314, 0, 
    1060, 795, 1031, 1021, 676, 852, 410, 63, 
    1322, 978, 1009, 1146, 794, 957, 453, 243, 
    1575, 1390, 1052, 926, 808, 517, 383, 305, 
    1548, 1771, 1794, 1114, 909, 847, 1041, 971, 
    1368, 1752, 1682, 953, 993, 1140, 1332, 1260, 
    1141, 1140, 970, 857, 1029, 1126, 1356, 1220, 
    
    -- channel=3
    79, 54, 67, 60, 61, 57, 48, 59, 
    89, 45, 92, 22, 99, 44, 14, 54, 
    150, 59, 86, 48, 111, 64, 27, 51, 
    178, 49, 103, 54, 109, 19, 39, 31, 
    186, 59, 56, 51, 47, 21, 71, 55, 
    179, 136, 20, 37, 26, 62, 52, 41, 
    163, 111, 30, 69, 77, 84, 98, 100, 
    161, 83, 72, 57, 74, 75, 91, 54, 
    
    -- channel=4
    561, 575, 606, 559, 528, 399, 473, 484, 
    539, 612, 643, 573, 457, 415, 410, 483, 
    483, 676, 682, 515, 462, 422, 328, 360, 
    501, 660, 713, 631, 565, 541, 380, 419, 
    487, 462, 660, 662, 580, 537, 444, 504, 
    531, 598, 487, 402, 345, 208, 227, 302, 
    369, 644, 501, 202, 90, 0, 0, 31, 
    59, 345, 238, 87, 94, 90, 125, 82, 
    
    -- channel=5
    66, 0, 17, 0, 37, 21, 0, 0, 
    108, 11, 48, 0, 102, 59, 0, 0, 
    241, 0, 127, 0, 104, 81, 0, 0, 
    303, 0, 130, 29, 112, 44, 35, 0, 
    337, 0, 82, 24, 38, 6, 52, 0, 
    326, 191, 28, 87, 25, 115, 119, 70, 
    289, 253, 0, 96, 130, 137, 164, 128, 
    204, 206, 103, 122, 140, 150, 192, 67, 
    
    -- channel=6
    31, 27, 7, 97, 29, 74, 60, 154, 
    63, 55, 71, 160, 74, 177, 125, 152, 
    157, 253, 175, 248, 178, 249, 130, 157, 
    217, 290, 35, 263, 201, 260, 119, 207, 
    245, 319, 192, 156, 218, 166, 58, 227, 
    199, 270, 414, 193, 228, 119, 122, 380, 
    155, 184, 418, 212, 176, 198, 217, 453, 
    207, 186, 295, 159, 162, 209, 230, 429, 
    
    -- channel=7
    54, 54, 123, 139, 90, 157, 93, 21, 
    210, 145, 250, 244, 256, 404, 221, 19, 
    639, 445, 553, 545, 382, 515, 256, 116, 
    821, 573, 542, 625, 456, 570, 279, 182, 
    958, 809, 651, 566, 489, 331, 262, 233, 
    985, 1034, 1122, 778, 682, 693, 783, 782, 
    986, 1140, 1106, 778, 838, 936, 1078, 1089, 
    989, 936, 818, 755, 873, 930, 1121, 1078, 
    
    -- channel=8
    352, 397, 427, 427, 356, 319, 324, 312, 
    335, 452, 474, 423, 325, 312, 294, 300, 
    385, 487, 495, 456, 388, 359, 284, 255, 
    397, 498, 502, 513, 434, 374, 304, 310, 
    384, 471, 464, 456, 437, 362, 306, 365, 
    407, 535, 474, 397, 358, 210, 237, 279, 
    260, 521, 432, 204, 110, 56, 82, 88, 
    93, 239, 213, 72, 77, 94, 108, 109, 
    
    -- channel=9
    17, 2, 73, 61, 46, 90, 7, 0, 
    101, 72, 199, 173, 177, 311, 122, 0, 
    451, 299, 463, 424, 295, 399, 152, 0, 
    588, 392, 504, 510, 352, 465, 182, 84, 
    762, 596, 457, 424, 320, 257, 155, 101, 
    773, 782, 825, 519, 434, 393, 490, 447, 
    692, 840, 815, 493, 501, 571, 668, 631, 
    621, 614, 519, 450, 531, 571, 699, 622, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 40, 0, 145, 83, 0, 
    213, 167, 172, 174, 67, 169, 101, 33, 
    288, 228, 107, 238, 119, 207, 103, 66, 
    379, 258, 130, 181, 128, 133, 78, 43, 
    355, 254, 418, 315, 303, 163, 222, 230, 
    357, 344, 486, 325, 270, 308, 341, 395, 
    370, 346, 411, 280, 275, 313, 373, 429, 
    
    -- channel=11
    66, 67, 68, 57, 65, 46, 56, 41, 
    15, 13, 18, 7, 3, 0, 10, 0, 
    22, 29, 16, 0, 23, 0, 0, 1, 
    0, 5, 3, 0, 21, 0, 0, 0, 
    0, 13, 0, 0, 0, 7, 25, 3, 
    46, 19, 21, 23, 42, 32, 36, 23, 
    43, 14, 6, 8, 8, 15, 18, 8, 
    20, 8, 17, 18, 32, 40, 37, 44, 
    
    -- channel=12
    373, 395, 428, 436, 337, 316, 297, 317, 
    364, 446, 467, 429, 299, 344, 280, 288, 
    414, 479, 516, 495, 338, 387, 272, 219, 
    441, 467, 491, 516, 354, 411, 268, 309, 
    475, 454, 444, 456, 381, 360, 280, 342, 
    451, 478, 550, 353, 318, 184, 209, 249, 
    231, 493, 490, 136, 79, 45, 72, 146, 
    45, 224, 155, 50, 64, 69, 101, 127, 
    
    -- channel=13
    68, 54, 91, 82, 41, 106, 43, 25, 
    144, 104, 140, 156, 144, 222, 127, 2, 
    378, 254, 323, 350, 215, 290, 163, 80, 
    486, 360, 314, 367, 242, 325, 169, 136, 
    563, 495, 403, 358, 275, 152, 158, 140, 
    543, 607, 622, 418, 410, 418, 463, 491, 
    542, 602, 575, 448, 479, 534, 625, 620, 
    516, 468, 462, 418, 487, 519, 619, 590, 
    
    -- channel=14
    590, 603, 688, 630, 518, 488, 470, 514, 
    562, 675, 717, 602, 525, 502, 403, 494, 
    566, 725, 776, 627, 579, 559, 363, 363, 
    576, 656, 768, 705, 585, 560, 407, 454, 
    593, 540, 636, 597, 549, 520, 447, 528, 
    587, 750, 652, 533, 351, 240, 278, 357, 
    332, 715, 471, 144, 66, 28, 52, 103, 
    54, 253, 122, 35, 56, 46, 99, 69, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 
    25, 0, 0, 0, 0, 0, 0, 0, 
    18, 33, 11, 10, 12, 26, 22, 16, 
    
    -- channel=16
    223, 134, 195, 151, 165, 166, 109, 101, 
    322, 210, 291, 167, 265, 224, 105, 112, 
    452, 239, 337, 258, 333, 285, 104, 106, 
    528, 187, 367, 265, 342, 268, 155, 116, 
    571, 308, 323, 280, 228, 148, 204, 171, 
    558, 525, 365, 295, 170, 215, 243, 248, 
    454, 510, 280, 177, 208, 224, 276, 263, 
    355, 330, 107, 162, 227, 239, 294, 214, 
    
    -- channel=17
    236, 206, 228, 359, 199, 291, 236, 304, 
    383, 321, 387, 443, 180, 454, 353, 312, 
    631, 608, 563, 632, 411, 571, 359, 292, 
    771, 756, 388, 667, 419, 581, 329, 392, 
    827, 769, 569, 539, 567, 394, 243, 464, 
    745, 722, 963, 515, 617, 399, 460, 726, 
    538, 649, 1011, 514, 480, 504, 590, 880, 
    534, 569, 701, 436, 477, 528, 641, 821, 
    
    -- channel=18
    107, 97, 101, 115, 86, 76, 88, 88, 
    91, 92, 84, 68, 50, 74, 69, 82, 
    107, 124, 84, 79, 29, 90, 59, 85, 
    81, 106, 63, 84, 60, 89, 77, 106, 
    100, 63, 78, 31, 84, 65, 75, 104, 
    86, 55, 94, 44, 59, 1, 15, 69, 
    53, 45, 61, 10, 5, 11, 5, 95, 
    83, 25, 24, 27, 36, 37, 48, 64, 
    
    -- channel=19
    407, 229, 318, 113, 268, 143, 189, 229, 
    421, 344, 316, 112, 356, 149, 144, 267, 
    545, 377, 404, 69, 407, 176, 101, 172, 
    593, 169, 495, 68, 342, 114, 177, 140, 
    651, 161, 215, 241, 159, 126, 257, 198, 
    665, 277, 0, 54, 0, 123, 126, 70, 
    446, 350, 0, 12, 38, 48, 58, 48, 
    329, 104, 31, 37, 68, 58, 122, 0, 
    
    -- channel=20
    45, 16, 60, 56, 48, 99, 47, 0, 
    138, 79, 92, 91, 120, 212, 79, 22, 
    315, 200, 256, 225, 203, 275, 107, 69, 
    372, 233, 259, 289, 206, 284, 136, 92, 
    455, 332, 303, 272, 224, 135, 143, 115, 
    486, 482, 499, 350, 327, 372, 391, 392, 
    490, 522, 482, 373, 410, 441, 528, 509, 
    495, 443, 374, 381, 434, 439, 546, 486, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 0, 
    32, 0, 0, 18, 58, 160, 53, 0, 
    280, 127, 218, 238, 134, 231, 79, 0, 
    411, 229, 205, 274, 181, 258, 87, 50, 
    531, 426, 283, 267, 195, 57, 43, 11, 
    532, 564, 609, 385, 362, 437, 475, 487, 
    541, 577, 575, 493, 544, 604, 686, 702, 
    599, 510, 437, 477, 569, 595, 727, 680, 
    
    -- channel=22
    107, 115, 130, 151, 116, 109, 116, 126, 
    116, 123, 153, 177, 98, 133, 126, 127, 
    122, 184, 165, 151, 75, 149, 112, 131, 
    141, 201, 169, 192, 128, 166, 106, 126, 
    117, 133, 161, 173, 168, 182, 85, 153, 
    116, 110, 205, 115, 126, 58, 53, 138, 
    55, 158, 220, 43, 20, 0, 0, 121, 
    50, 121, 115, 49, 64, 56, 74, 105, 
    
    -- channel=23
    621, 678, 736, 677, 619, 493, 512, 508, 
    601, 716, 789, 693, 557, 552, 447, 486, 
    634, 898, 946, 784, 584, 568, 439, 294, 
    647, 830, 987, 924, 787, 730, 509, 483, 
    756, 727, 845, 882, 709, 704, 526, 569, 
    786, 968, 779, 630, 495, 233, 288, 339, 
    526, 985, 770, 308, 119, 29, 47, 30, 
    85, 443, 337, 141, 184, 201, 252, 147, 
    
    -- channel=24
    94, 81, 133, 131, 57, 132, 44, 6, 
    213, 148, 227, 244, 228, 368, 169, 0, 
    632, 445, 611, 583, 346, 510, 242, 30, 
    809, 577, 569, 659, 423, 549, 245, 156, 
    992, 830, 610, 551, 454, 260, 222, 166, 
    980, 1024, 1083, 658, 587, 587, 666, 648, 
    870, 1027, 1001, 650, 702, 798, 919, 890, 
    787, 740, 693, 612, 715, 770, 931, 855, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 2, 1, 
    0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    24, 13, 26, 89, 22, 97, 64, 67, 
    149, 52, 142, 157, 119, 286, 193, 35, 
    478, 357, 340, 406, 255, 358, 224, 137, 
    611, 480, 284, 440, 303, 378, 231, 142, 
    668, 569, 417, 351, 391, 221, 160, 162, 
    652, 666, 766, 585, 498, 409, 486, 515, 
    660, 726, 850, 557, 532, 603, 689, 766, 
    709, 668, 607, 507, 565, 619, 743, 821, 
    
    -- channel=27
    48, 47, 54, 40, 48, 11, 35, 37, 
    60, 51, 50, 19, 19, 0, 31, 43, 
    0, 58, 51, 0, 17, 0, 0, 16, 
    0, 22, 66, 2, 8, 0, 12, 8, 
    0, 0, 26, 33, 0, 17, 32, 35, 
    23, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=28
    22, 12, 14, 61, 17, 55, 43, 81, 
    54, 18, 7, 64, 0, 71, 77, 86, 
    73, 115, 41, 111, 4, 99, 66, 74, 
    57, 126, 0, 100, 15, 105, 22, 108, 
    47, 99, 75, 63, 98, 45, 14, 131, 
    2, 0, 125, 29, 120, 42, 32, 181, 
    0, 0, 133, 7, 10, 0, 0, 177, 
    0, 0, 54, 0, 0, 6, 10, 158, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 0, 0, 0, 24, 
    0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=30
    20, 26, 28, 48, 50, 52, 52, 49, 
    65, 56, 35, 80, 83, 48, 71, 53, 
    24, 83, 22, 60, 118, 67, 80, 84, 
    23, 100, 38, 59, 105, 84, 89, 57, 
    22, 99, 88, 81, 59, 98, 84, 52, 
    13, 88, 135, 97, 143, 126, 87, 118, 
    93, 34, 200, 133, 118, 98, 109, 112, 
    102, 66, 154, 95, 86, 114, 87, 127, 
    
    -- channel=31
    4, 0, 0, 2, 0, 0, 0, 0, 
    18, 25, 1, 12, 9, 6, 0, 0, 
    40, 26, 33, 9, 7, 20, 0, 0, 
    6, 0, 0, 0, 4, 0, 0, 10, 
    12, 0, 24, 12, 11, 0, 0, 0, 
    0, 0, 50, 0, 0, 5, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end inmem_package;
