library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    0, 0, 0, 0, 76, 58, 135, 292, 0, 193, 0, 0, 0, 0, 136, 171, 555, 457, 0, 0, 0, 0, 0, 0, 0, 0, 0, 180, 277, 241, 0, 0, 0, 222, 0, 182, 0, 0, 0, 0, 0, 0, 0, 0, 0, 94, 0, 0, 0, 0, 0, 0, 0, 0, 549, 859, 586, 1015, 424, 401, 734, 430, 487, 168, 0, 0, 0, 0, 0, 289, 103, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 107, 0, 0, 0, 0, 24, 151, 0, 0, 563, 481, 428, 279, 396, 178, 764, 593, 729, 0, 0, 304, 0, 0, 0, 307, 0, 0, 328, 84, 216, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 315, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 79, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 157, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 267, 76, 0, 143, 45, 257, 0, 29, 303, 0, 0, 0, 0, 38, 185, 0, 0, 0, 0, 0, 64, 68, 0, 61, 0, 172, 8, 13, 24, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 190, 358, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 217, 519, 0, 305, 319, 0, 0, 0, 0, 0, 0, 0, 0, 164, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 200, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 0, 0, 0, 0, 0, 0, 0, 0, 159, 207, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 130, 128, 11, 0, 0, 0, 0, 0, 0, 0, 40, 66, 0, 0, 0, 0, 375, 668, 0, 65, 0, 0, 0, 37, 0, 0, 0, 332, 421, 406, 36, 391, 188, 0, 0, 0, 804, 589, 385, 712, 697, 736, 518, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 384, 157, 283, 0, 0, 90, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 83, 30, 0, 0, 0, 0, 0, 0, 0, 0, 93, 0, 164, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 81, 315, 292, 0, 0, 0, 79, 242, 276, 0, 81, 61, 15, 136, 124, 383, 320, 97, 357, 94, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 34, 165, 268, 562, 307, 233, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 285, 143, 0, 436, 187, 221, 0, 0, 186, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 302, 386, 347, 442, 521, 360, 18, 166, 19, 234, 238, 448, 183, 317, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 285, 213, 143, 243, 387, 417, 256, 80, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 52, 0, 279, 0, 0, 0, 0, 359, 0, 0, 172, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 164, 0, 0, 31, 0, 0, 0, 0,
    others => 0);
end ifmap_package;
