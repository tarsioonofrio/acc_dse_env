library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 14, 7, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 8, 25, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 11, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 16, 13, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 13, 11, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 12, 29, 6, 0, 0, 0, 0, 0, 0, 0, 17, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 22, 34, 21, 0, 0, 0, 0, 0, 0, 0, 7, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 30, 29, 35, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 37, 36, 39, 43, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 30, 36, 38, 40, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 28, 27, 30, 24, 7, 12, 13, 0, 0, 0, 0, 0, 0, 11, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 16, 25, 18, 19, 17, 3, 20, 57, 52, 11, 0, 6, 3, 20, 33, 27, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 31, 37, 21, 23, 26, 11, 15, 46, 69, 55, 17, 13, 17, 26, 22, 20, 15, 4, 0, 0, 4, 10, 20, 31, 26, 24, 24, 19, 16, 21, 34, 
    0, 42, 49, 37, 38, 38, 19, 25, 46, 35, 32, 32, 12, 13, 15, 11, 22, 28, 18, 15, 31, 39, 39, 43, 51, 58, 61, 59, 58, 57, 61, 60, 
    3, 47, 37, 42, 39, 28, 19, 33, 39, 36, 44, 31, 29, 31, 31, 30, 32, 37, 37, 39, 48, 51, 54, 58, 63, 70, 71, 67, 66, 66, 70, 69, 
    29, 74, 45, 31, 41, 30, 15, 31, 35, 41, 41, 42, 44, 45, 45, 43, 43, 44, 46, 50, 53, 59, 63, 67, 71, 73, 70, 68, 73, 80, 86, 80, 
    35, 89, 64, 39, 34, 30, 32, 42, 45, 36, 37, 51, 51, 50, 49, 47, 46, 47, 50, 53, 59, 67, 73, 74, 72, 71, 67, 71, 85, 93, 89, 85, 
    35, 92, 77, 59, 38, 25, 46, 61, 51, 34, 43, 51, 56, 52, 47, 47, 49, 52, 55, 60, 64, 68, 73, 77, 79, 73, 73, 82, 91, 90, 85, 78, 
    34, 92, 83, 73, 58, 31, 35, 61, 45, 37, 49, 55, 57, 59, 53, 47, 47, 51, 58, 62, 67, 74, 74, 73, 75, 78, 84, 88, 92, 91, 75, 61, 
    39, 92, 83, 80, 73, 51, 29, 38, 43, 32, 41, 48, 55, 59, 59, 57, 55, 57, 60, 64, 69, 70, 71, 71, 74, 81, 89, 100, 107, 91, 63, 51, 
    35, 94, 80, 79, 78, 67, 50, 41, 35, 41, 40, 41, 43, 45, 51, 52, 52, 57, 66, 72, 71, 69, 68, 67, 70, 81, 96, 105, 97, 87, 67, 51, 
    33, 88, 74, 72, 74, 68, 57, 49, 43, 45, 43, 45, 46, 43, 38, 35, 38, 47, 57, 65, 70, 68, 61, 58, 63, 74, 86, 93, 90, 80, 67, 57, 
    0, 5, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 11, 4, 2, 0, 
    
    -- channel=2
    293, 198, 206, 190, 181, 196, 201, 193, 194, 201, 203, 195, 194, 204, 212, 211, 208, 206, 204, 194, 180, 177, 179, 184, 181, 174, 176, 181, 183, 177, 170, 55, 
    354, 289, 306, 290, 279, 292, 295, 290, 288, 286, 290, 283, 282, 299, 311, 312, 306, 293, 279, 268, 253, 249, 255, 262, 266, 260, 251, 255, 264, 257, 247, 108, 
    355, 292, 313, 295, 282, 297, 296, 291, 291, 293, 290, 258, 243, 282, 306, 301, 292, 260, 243, 228, 202, 180, 192, 222, 235, 261, 266, 260, 265, 262, 250, 104, 
    357, 291, 304, 298, 287, 303, 302, 294, 297, 307, 338, 253, 166, 233, 285, 262, 247, 238, 220, 199, 150, 114, 101, 124, 160, 192, 242, 267, 268, 259, 254, 107, 
    346, 276, 288, 295, 293, 304, 308, 296, 301, 315, 381, 333, 173, 200, 243, 234, 193, 194, 222, 188, 132, 101, 77, 85, 99, 119, 167, 250, 275, 253, 242, 104, 
    323, 211, 256, 327, 315, 303, 307, 300, 299, 311, 336, 311, 226, 182, 152, 160, 157, 160, 213, 189, 125, 105, 104, 109, 104, 78, 96, 194, 276, 264, 234, 98, 
    283, 115, 146, 312, 331, 301, 308, 311, 298, 291, 284, 265, 237, 173, 103, 117, 131, 123, 200, 229, 136, 82, 116, 147, 121, 80, 85, 130, 239, 278, 241, 93, 
    253, 39, 97, 229, 267, 284, 307, 308, 293, 238, 229, 248, 230, 153, 87, 113, 138, 118, 163, 257, 206, 91, 96, 145, 139, 103, 80, 97, 185, 280, 260, 88, 
    278, 0, 94, 199, 173, 241, 300, 317, 283, 160, 89, 189, 199, 125, 77, 96, 129, 120, 139, 228, 241, 133, 78, 95, 131, 124, 91, 68, 114, 251, 294, 96, 
    301, 47, 114, 169, 135, 209, 273, 352, 347, 171, 47, 116, 159, 91, 86, 79, 107, 95, 130, 237, 216, 130, 80, 69, 120, 126, 104, 77, 67, 164, 278, 125, 
    286, 70, 181, 152, 117, 191, 245, 307, 411, 243, 83, 120, 163, 72, 78, 98, 85, 73, 140, 281, 195, 101, 85, 66, 135, 148, 103, 84, 59, 97, 194, 119, 
    271, 57, 209, 163, 118, 191, 246, 220, 331, 296, 125, 177, 218, 97, 45, 105, 106, 36, 147, 314, 188, 77, 83, 75, 134, 159, 132, 100, 75, 77, 125, 76, 
    263, 45, 210, 130, 111, 223, 267, 196, 262, 282, 152, 198, 263, 142, 36, 90, 128, 53, 148, 303, 162, 70, 74, 91, 123, 148, 155, 128, 94, 89, 110, 44, 
    264, 56, 216, 73, 46, 230, 287, 204, 234, 271, 212, 220, 218, 174, 95, 101, 106, 69, 174, 282, 143, 72, 71, 73, 104, 122, 148, 149, 103, 103, 143, 48, 
    282, 64, 205, 62, 0, 168, 272, 201, 204, 245, 267, 243, 100, 98, 133, 145, 120, 77, 182, 277, 156, 78, 94, 91, 118, 145, 145, 155, 125, 131, 185, 72, 
    304, 65, 178, 87, 0, 88, 226, 181, 175, 254, 296, 281, 130, 63, 140, 148, 143, 126, 200, 255, 188, 117, 73, 74, 115, 162, 160, 158, 160, 182, 225, 80, 
    325, 52, 146, 117, 0, 30, 203, 166, 121, 203, 287, 225, 176, 133, 145, 147, 142, 159, 188, 227, 241, 207, 98, 78, 116, 163, 177, 162, 179, 222, 239, 78, 
    358, 53, 114, 125, 20, 0, 161, 192, 96, 126, 188, 191, 179, 145, 158, 121, 106, 189, 175, 123, 180, 222, 132, 87, 131, 158, 194, 205, 207, 241, 248, 87, 
    390, 91, 106, 124, 58, 0, 106, 193, 136, 108, 62, 159, 207, 157, 197, 98, 31, 180, 205, 134, 124, 107, 112, 114, 133, 158, 191, 242, 235, 246, 256, 95, 
    412, 143, 113, 133, 89, 2, 69, 164, 93, 103, 81, 120, 208, 183, 215, 106, 0, 91, 201, 186, 150, 90, 94, 125, 147, 179, 206, 254, 240, 250, 257, 96, 
    411, 193, 114, 141, 105, 22, 98, 216, 78, 0, 21, 91, 135, 166, 173, 91, 6, 17, 77, 119, 121, 106, 81, 77, 99, 121, 168, 200, 183, 182, 191, 60, 
    379, 215, 100, 133, 100, 18, 130, 272, 168, 0, 0, 55, 138, 161, 155, 122, 61, 44, 51, 44, 62, 69, 72, 59, 47, 55, 88, 108, 101, 92, 94, 0, 
    322, 225, 125, 125, 94, 36, 161, 269, 176, 62, 0, 38, 128, 142, 131, 126, 83, 52, 57, 53, 49, 41, 46, 45, 33, 25, 33, 45, 36, 25, 24, 0, 
    224, 158, 183, 166, 105, 113, 225, 244, 116, 26, 0, 35, 64, 62, 58, 59, 53, 37, 36, 43, 43, 33, 29, 26, 25, 18, 11, 16, 12, 9, 9, 0, 
    151, 25, 130, 199, 128, 155, 274, 198, 38, 0, 10, 27, 31, 23, 22, 30, 33, 26, 25, 29, 29, 20, 16, 20, 18, 15, 6, 6, 1, 2, 4, 0, 
    151, 0, 35, 132, 159, 209, 268, 116, 0, 0, 41, 24, 20, 18, 20, 26, 28, 26, 24, 25, 21, 17, 9, 10, 14, 13, 14, 21, 17, 8, 11, 0, 
    162, 0, 0, 41, 119, 264, 267, 43, 0, 1, 32, 33, 15, 6, 23, 29, 26, 23, 22, 21, 14, 16, 23, 14, 0, 0, 10, 26, 25, 9, 15, 0, 
    162, 0, 0, 0, 41, 201, 291, 48, 0, 37, 30, 30, 23, 0, 6, 20, 27, 29, 23, 17, 12, 3, 13, 16, 3, 0, 3, 13, 5, 0, 15, 0, 
    154, 0, 0, 0, 0, 76, 206, 115, 0, 55, 54, 52, 43, 21, 6, 5, 16, 17, 16, 10, 6, 2, 1, 10, 17, 13, 7, 0, 0, 0, 1, 0, 
    171, 0, 0, 0, 0, 7, 64, 81, 28, 29, 47, 56, 56, 54, 41, 30, 34, 28, 18, 2, 0, 0, 0, 15, 40, 46, 11, 0, 0, 0, 0, 0, 
    180, 0, 0, 0, 0, 0, 12, 30, 26, 13, 32, 35, 33, 39, 46, 64, 73, 65, 56, 29, 0, 0, 4, 33, 67, 75, 36, 0, 0, 0, 0, 0, 
    218, 87, 85, 94, 95, 97, 95, 101, 98, 87, 97, 100, 96, 95, 88, 107, 133, 146, 153, 140, 109, 102, 105, 122, 161, 176, 159, 104, 60, 72, 79, 19, 
    
    -- channel=3
    0, 2, 6, 5, 4, 4, 6, 6, 3, 4, 5, 4, 3, 6, 6, 7, 8, 7, 6, 5, 3, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    0, 137, 137, 154, 161, 147, 148, 154, 151, 147, 140, 145, 148, 151, 156, 159, 160, 155, 145, 145, 146, 138, 132, 131, 137, 142, 137, 133, 133, 134, 128, 188, 
    0, 90, 82, 108, 122, 103, 109, 116, 120, 113, 102, 103, 106, 108, 117, 124, 131, 126, 104, 90, 75, 61, 51, 52, 72, 86, 102, 105, 106, 112, 107, 235, 
    0, 95, 85, 112, 124, 108, 113, 119, 123, 118, 112, 125, 146, 127, 119, 124, 127, 118, 97, 59, 64, 58, 40, 22, 17, 29, 52, 85, 101, 111, 109, 244, 
    0, 107, 99, 122, 126, 108, 108, 121, 116, 102, 82, 145, 235, 154, 104, 101, 86, 77, 45, 44, 69, 85, 77, 51, 42, 9, 18, 39, 69, 95, 106, 246, 
    0, 95, 81, 95, 118, 106, 108, 121, 115, 87, 0, 62, 190, 126, 55, 49, 49, 45, 0, 0, 34, 64, 79, 76, 55, 46, 4, 0, 14, 77, 107, 254, 
    0, 69, 26, 0, 64, 109, 116, 127, 122, 100, 0, 29, 143, 127, 102, 71, 70, 22, 0, 0, 26, 45, 45, 43, 45, 79, 38, 0, 0, 37, 102, 259, 
    0, 136, 35, 0, 6, 101, 116, 121, 125, 116, 78, 75, 83, 127, 162, 78, 37, 6, 0, 0, 31, 83, 50, 2, 34, 75, 67, 0, 0, 0, 82, 265, 
    0, 219, 86, 0, 22, 106, 114, 111, 127, 135, 132, 66, 44, 110, 142, 49, 2, 11, 0, 0, 0, 114, 74, 5, 22, 60, 67, 27, 0, 0, 40, 267, 
    0, 239, 69, 0, 85, 127, 105, 96, 111, 237, 240, 96, 27, 105, 132, 61, 2, 14, 0, 0, 0, 106, 119, 69, 34, 47, 67, 72, 0, 0, 0, 232, 
    0, 201, 0, 0, 141, 144, 90, 5, 0, 182, 255, 92, 46, 128, 144, 88, 42, 25, 9, 0, 0, 100, 145, 123, 36, 23, 60, 88, 63, 0, 0, 174, 
    0, 103, 0, 0, 166, 165, 126, 0, 0, 0, 187, 103, 75, 160, 145, 106, 67, 83, 0, 0, 0, 106, 126, 120, 12, 6, 43, 83, 103, 18, 0, 132, 
    0, 62, 0, 0, 168, 156, 157, 29, 0, 0, 111, 51, 13, 177, 181, 118, 87, 138, 0, 0, 0, 108, 126, 106, 0, 0, 26, 55, 84, 61, 7, 132, 
    0, 83, 0, 1, 142, 95, 129, 177, 0, 0, 77, 11, 0, 148, 232, 124, 69, 159, 0, 0, 14, 139, 127, 83, 1, 0, 0, 21, 65, 62, 69, 167, 
    0, 85, 0, 76, 150, 42, 70, 196, 3, 0, 25, 0, 0, 72, 162, 106, 67, 143, 0, 0, 35, 146, 126, 92, 42, 0, 0, 4, 53, 57, 74, 191, 
    0, 68, 0, 140, 197, 27, 13, 181, 69, 0, 0, 0, 68, 107, 72, 55, 68, 111, 0, 0, 32, 119, 102, 67, 14, 0, 0, 0, 44, 62, 49, 217, 
    0, 71, 0, 119, 236, 61, 0, 144, 89, 0, 0, 0, 93, 97, 29, 3, 46, 83, 0, 0, 29, 97, 102, 96, 17, 0, 0, 0, 37, 57, 49, 245, 
    0, 91, 0, 57, 235, 85, 0, 63, 135, 0, 0, 0, 27, 79, 25, 16, 29, 38, 0, 0, 0, 0, 98, 97, 0, 0, 0, 0, 52, 55, 76, 275, 
    0, 97, 0, 7, 202, 135, 0, 0, 160, 47, 0, 0, 0, 81, 45, 60, 50, 0, 6, 93, 2, 0, 57, 59, 4, 0, 0, 10, 56, 63, 94, 288, 
    0, 76, 3, 0, 143, 183, 0, 0, 75, 93, 103, 20, 0, 51, 0, 108, 114, 0, 0, 134, 60, 22, 56, 51, 0, 0, 0, 14, 71, 90, 104, 290, 
    0, 32, 26, 0, 87, 190, 22, 0, 29, 87, 129, 0, 0, 0, 0, 136, 200, 0, 0, 0, 22, 57, 25, 1, 0, 0, 0, 13, 89, 104, 96, 277, 
    0, 0, 50, 5, 61, 168, 21, 0, 102, 204, 213, 77, 22, 0, 0, 118, 233, 129, 25, 15, 11, 33, 29, 0, 0, 0, 0, 0, 53, 53, 43, 216, 
    0, 0, 58, 16, 69, 172, 0, 0, 79, 295, 234, 96, 0, 0, 0, 0, 89, 89, 67, 67, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 158, 
    0, 0, 0, 0, 81, 181, 0, 0, 0, 159, 173, 0, 0, 0, 0, 0, 0, 0, 8, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 121, 
    0, 0, 0, 0, 20, 82, 0, 0, 19, 118, 115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 120, 
    0, 0, 0, 0, 0, 0, 0, 0, 115, 160, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 162, 
    0, 0, 0, 0, 0, 0, 0, 16, 216, 119, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 180, 
    0, 0, 0, 0, 0, 0, 0, 110, 250, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 145, 
    0, 0, 0, 0, 0, 0, 0, 79, 182, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 102, 
    0, 0, 0, 0, 0, 0, 0, 0, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 73, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 70, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    
    -- channel=5
    93, 90, 98, 95, 89, 93, 93, 92, 89, 88, 94, 94, 93, 95, 95, 95, 94, 92, 93, 89, 83, 81, 79, 83, 82, 80, 77, 75, 74, 71, 67, 7, 
    69, 18, 27, 21, 20, 28, 27, 24, 23, 24, 23, 22, 21, 22, 23, 23, 23, 21, 14, 6, 1, 0, 3, 8, 12, 18, 15, 13, 15, 13, 10, 0, 
    69, 18, 28, 25, 22, 28, 27, 23, 23, 29, 46, 38, 9, 11, 23, 23, 24, 9, 0, 4, 0, 0, 0, 0, 0, 0, 13, 16, 16, 16, 14, 0, 
    73, 24, 27, 25, 25, 30, 28, 22, 24, 34, 88, 72, 0, 5, 20, 8, 0, 0, 13, 17, 15, 4, 0, 0, 0, 0, 0, 7, 17, 14, 12, 0, 
    73, 16, 18, 23, 21, 26, 24, 20, 21, 30, 69, 51, 3, 0, 0, 0, 0, 0, 17, 39, 30, 19, 5, 5, 11, 0, 0, 0, 18, 14, 8, 0, 
    68, 0, 0, 20, 28, 23, 25, 23, 23, 26, 34, 0, 0, 0, 0, 0, 0, 0, 50, 56, 19, 0, 0, 10, 1, 0, 0, 0, 15, 21, 11, 0, 
    69, 0, 0, 3, 21, 21, 26, 29, 28, 22, 11, 8, 14, 5, 0, 10, 18, 10, 39, 60, 25, 0, 0, 0, 0, 0, 0, 0, 8, 19, 10, 0, 
    88, 0, 0, 54, 16, 11, 26, 31, 36, 13, 0, 34, 49, 18, 0, 0, 12, 0, 8, 35, 29, 0, 0, 0, 0, 0, 0, 0, 0, 25, 18, 0, 
    112, 0, 27, 69, 22, 4, 24, 62, 95, 49, 7, 31, 51, 8, 0, 0, 0, 0, 0, 33, 27, 0, 0, 0, 0, 0, 0, 0, 0, 6, 24, 0, 
    104, 0, 66, 54, 0, 0, 16, 80, 139, 84, 27, 55, 41, 0, 0, 0, 0, 0, 0, 65, 64, 11, 0, 0, 9, 8, 0, 0, 0, 0, 7, 0, 
    94, 0, 52, 46, 0, 0, 9, 41, 92, 59, 0, 14, 38, 0, 0, 0, 0, 0, 11, 115, 75, 10, 0, 0, 3, 15, 1, 0, 0, 0, 2, 0, 
    85, 0, 57, 21, 0, 0, 16, 10, 55, 12, 0, 8, 68, 12, 0, 0, 6, 0, 27, 128, 54, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    80, 0, 72, 0, 0, 0, 18, 0, 53, 39, 0, 28, 68, 28, 0, 0, 11, 0, 49, 116, 24, 0, 0, 0, 0, 0, 1, 6, 0, 0, 0, 0, 
    85, 0, 83, 0, 0, 0, 16, 0, 29, 43, 33, 65, 59, 4, 0, 10, 1, 0, 42, 102, 6, 0, 0, 0, 0, 2, 10, 17, 4, 0, 0, 0, 
    100, 2, 72, 0, 0, 0, 20, 0, 20, 45, 75, 105, 19, 0, 0, 0, 0, 0, 30, 75, 13, 0, 0, 0, 4, 22, 29, 23, 0, 0, 11, 0, 
    117, 2, 59, 7, 0, 0, 29, 0, 0, 48, 97, 62, 0, 0, 0, 0, 0, 0, 40, 65, 8, 0, 0, 0, 0, 7, 9, 0, 0, 4, 21, 0, 
    135, 0, 44, 22, 0, 0, 36, 25, 0, 20, 31, 0, 0, 0, 0, 0, 0, 4, 17, 0, 5, 19, 0, 0, 0, 3, 4, 0, 0, 14, 22, 0, 
    149, 6, 33, 23, 0, 0, 23, 31, 0, 0, 0, 0, 0, 0, 13, 1, 0, 24, 24, 0, 0, 0, 0, 0, 0, 0, 7, 21, 28, 32, 27, 0, 
    149, 9, 25, 24, 0, 0, 10, 27, 0, 11, 0, 0, 18, 21, 68, 29, 0, 11, 26, 16, 16, 0, 0, 0, 3, 17, 29, 42, 30, 25, 16, 0, 
    143, 19, 13, 21, 0, 0, 2, 50, 0, 0, 0, 15, 26, 46, 72, 23, 0, 0, 0, 0, 0, 0, 0, 0, 16, 25, 40, 41, 12, 5, 6, 0, 
    138, 33, 5, 21, 0, 0, 7, 114, 73, 0, 0, 9, 55, 62, 70, 25, 0, 0, 0, 0, 0, 0, 0, 2, 4, 7, 0, 1, 0, 0, 0, 0, 
    137, 44, 1, 17, 0, 0, 34, 134, 96, 50, 28, 18, 61, 62, 33, 0, 0, 0, 0, 0, 0, 0, 10, 23, 21, 8, 1, 0, 0, 0, 0, 0, 
    110, 36, 10, 22, 7, 0, 83, 142, 72, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 12, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    70, 0, 0, 27, 0, 11, 118, 120, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    65, 0, 0, 0, 0, 26, 101, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 9, 0, 
    71, 0, 0, 0, 0, 64, 110, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 10, 0, 
    69, 0, 0, 0, 0, 65, 102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    67, 0, 0, 0, 0, 30, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 18, 3, 0, 0, 0, 0, 
    76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 10, 1, 0, 0, 0, 0, 13, 36, 30, 0, 0, 0, 0, 0, 
    71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 9, 3, 0, 0, 0, 0, 28, 38, 18, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=7
    0, 23, 24, 22, 23, 26, 25, 26, 26, 27, 26, 23, 21, 25, 28, 28, 31, 32, 30, 27, 24, 21, 19, 20, 19, 21, 20, 20, 21, 23, 23, 12, 
    0, 8, 7, 5, 8, 8, 8, 10, 10, 11, 6, 4, 5, 7, 11, 13, 15, 15, 9, 4, 0, 0, 0, 0, 0, 0, 2, 7, 8, 10, 11, 4, 
    0, 10, 8, 7, 11, 8, 8, 9, 10, 11, 8, 5, 5, 7, 12, 11, 6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 8, 9, 3, 
    0, 11, 7, 6, 10, 9, 8, 8, 9, 9, 15, 2, 3, 7, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 6, 2, 
    0, 4, 0, 0, 7, 9, 8, 10, 11, 8, 3, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 3, 9, 9, 11, 12, 8, 0, 0, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 5, 11, 12, 12, 11, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 1, 12, 12, 10, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 1, 10, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 3, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 2, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 7, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=8
    0, 30, 32, 41, 37, 30, 34, 35, 35, 31, 31, 35, 31, 28, 29, 27, 29, 29, 30, 37, 41, 38, 35, 30, 33, 32, 30, 24, 23, 26, 27, 74, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 9, 12, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 76, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 17, 0, 0, 0, 0, 19, 15, 16, 29, 31, 17, 0, 0, 0, 0, 0, 0, 0, 1, 79, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 80, 20, 0, 11, 13, 6, 6, 44, 73, 86, 68, 46, 22, 0, 0, 0, 0, 0, 0, 80, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 91, 48, 15, 4, 3, 0, 25, 64, 106, 122, 124, 95, 69, 61, 10, 0, 0, 0, 1, 82, 
    0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 66, 62, 42, 19, 37, 36, 23, 70, 128, 135, 119, 102, 110, 88, 53, 0, 0, 0, 6, 83, 
    0, 76, 3, 0, 0, 0, 0, 0, 0, 0, 5, 3, 35, 81, 95, 69, 63, 65, 33, 63, 133, 138, 102, 93, 95, 98, 76, 15, 0, 0, 1, 86, 
    14, 129, 50, 0, 0, 0, 0, 0, 1, 35, 24, 17, 59, 109, 123, 90, 70, 78, 50, 27, 94, 140, 110, 73, 69, 88, 76, 49, 0, 0, 0, 92, 
    38, 177, 96, 55, 46, 12, 0, 0, 35, 113, 123, 82, 98, 126, 130, 92, 72, 78, 48, 0, 58, 132, 127, 87, 69, 77, 83, 66, 17, 0, 0, 88, 
    45, 190, 133, 100, 102, 34, 13, 0, 76, 186, 215, 121, 119, 145, 129, 114, 79, 75, 36, 4, 69, 133, 155, 120, 71, 77, 89, 84, 53, 0, 0, 68, 
    52, 177, 142, 128, 126, 54, 25, 15, 29, 147, 208, 152, 128, 172, 138, 116, 93, 94, 24, 8, 120, 163, 160, 123, 75, 74, 91, 91, 80, 26, 0, 41, 
    65, 178, 106, 152, 138, 58, 23, 39, 0, 97, 172, 122, 109, 192, 169, 115, 113, 117, 36, 26, 142, 184, 149, 120, 75, 63, 92, 92, 91, 62, 18, 41, 
    66, 176, 106, 176, 128, 37, 9, 54, 8, 44, 115, 100, 109, 197, 209, 137, 116, 136, 56, 38, 150, 194, 143, 112, 75, 57, 63, 88, 99, 81, 46, 70, 
    63, 180, 118, 196, 141, 22, 0, 51, 28, 18, 80, 122, 133, 181, 190, 147, 131, 132, 65, 50, 167, 180, 145, 120, 84, 69, 67, 90, 106, 88, 44, 92, 
    58, 190, 125, 207, 195, 38, 1, 51, 39, 28, 66, 133, 214, 177, 159, 140, 125, 114, 65, 57, 152, 181, 149, 116, 78, 72, 77, 83, 101, 69, 29, 103, 
    53, 207, 135, 204, 240, 94, 36, 66, 75, 28, 64, 133, 206, 174, 124, 102, 101, 100, 47, 52, 130, 162, 137, 119, 83, 62, 76, 71, 59, 37, 22, 99, 
    54, 229, 161, 202, 252, 152, 53, 94, 110, 38, 62, 80, 123, 148, 87, 97, 90, 69, 64, 61, 49, 98, 151, 113, 65, 39, 43, 50, 31, 23, 16, 100, 
    47, 247, 191, 200, 245, 202, 72, 103, 133, 105, 54, 48, 79, 97, 86, 120, 104, 57, 76, 61, 56, 77, 98, 79, 43, 21, 10, 29, 33, 20, 14, 111, 
    23, 244, 209, 202, 234, 231, 105, 88, 135, 129, 108, 49, 69, 79, 84, 154, 154, 55, 67, 111, 113, 69, 59, 62, 26, 26, 7, 13, 31, 17, 16, 106, 
    0, 214, 212, 197, 219, 233, 137, 92, 164, 153, 125, 61, 37, 72, 107, 182, 200, 94, 52, 86, 87, 75, 57, 32, 35, 23, 10, 8, 25, 17, 16, 95, 
    0, 182, 207, 186, 211, 224, 136, 94, 210, 227, 161, 125, 86, 137, 155, 200, 233, 158, 83, 69, 55, 68, 69, 62, 73, 56, 60, 48, 61, 59, 55, 101, 
    0, 159, 211, 187, 205, 209, 120, 120, 244, 326, 272, 194, 150, 157, 161, 192, 212, 170, 122, 94, 91, 93, 105, 120, 120, 116, 107, 105, 122, 123, 113, 141, 
    0, 127, 198, 191, 206, 214, 148, 155, 241, 338, 307, 181, 131, 128, 131, 140, 157, 148, 133, 140, 132, 130, 134, 144, 154, 160, 159, 165, 169, 173, 174, 169, 
    42, 116, 148, 167, 209, 187, 152, 188, 288, 295, 232, 178, 132, 126, 129, 128, 145, 154, 142, 143, 147, 155, 155, 158, 165, 178, 182, 180, 183, 187, 181, 179, 
    86, 153, 120, 129, 175, 144, 151, 232, 310, 252, 208, 167, 150, 152, 146, 145, 145, 149, 150, 151, 156, 163, 168, 170, 179, 187, 191, 191, 194, 189, 192, 215, 
    110, 203, 147, 108, 123, 127, 158, 273, 292, 230, 179, 162, 162, 158, 151, 148, 150, 152, 154, 160, 164, 172, 181, 188, 193, 188, 190, 187, 193, 208, 225, 232, 
    105, 220, 178, 135, 108, 95, 159, 296, 284, 217, 163, 160, 165, 163, 152, 149, 152, 157, 161, 163, 176, 182, 184, 192, 194, 191, 183, 183, 209, 230, 211, 203, 
    101, 220, 196, 170, 139, 84, 120, 278, 269, 186, 163, 158, 171, 174, 163, 155, 152, 155, 161, 170, 180, 182, 182, 188, 192, 192, 189, 212, 222, 211, 171, 175, 
    108, 226, 199, 186, 168, 123, 90, 201, 224, 162, 150, 152, 161, 177, 176, 162, 156, 163, 172, 177, 181, 189, 184, 174, 176, 192, 217, 233, 229, 217, 164, 150, 
    106, 225, 194, 189, 181, 161, 120, 137, 192, 147, 134, 140, 146, 155, 159, 160, 161, 170, 176, 190, 199, 190, 179, 169, 172, 194, 236, 258, 258, 216, 173, 130, 
    89, 222, 194, 182, 183, 175, 162, 142, 160, 150, 133, 133, 134, 139, 139, 133, 134, 151, 172, 196, 204, 188, 178, 164, 165, 190, 235, 266, 246, 200, 181, 133, 
    24, 118, 105, 94, 98, 96, 90, 83, 79, 82, 73, 72, 76, 74, 68, 59, 60, 71, 83, 96, 107, 103, 93, 84, 81, 91, 110, 135, 133, 112, 96, 82, 
    
    -- channel=9
    19, 4, 5, 10, 8, 2, 3, 4, 1, 0, 0, 11, 5, 0, 0, 0, 0, 0, 0, 11, 23, 26, 23, 19, 18, 18, 15, 8, 3, 6, 16, 58, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 81, 74, 36, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 103, 115, 108, 101, 82, 46, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 74, 96, 99, 82, 69, 72, 82, 73, 26, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 72, 93, 86, 71, 71, 77, 60, 37, 41, 52, 47, 52, 25, 0, 0, 0, 0, 
    98, 67, 63, 35, 0, 0, 0, 0, 0, 0, 0, 0, 7, 46, 51, 64, 73, 71, 50, 17, 14, 35, 38, 28, 22, 47, 68, 50, 0, 0, 0, 0, 
    136, 122, 128, 108, 0, 0, 0, 0, 0, 43, 52, 45, 54, 46, 38, 53, 58, 47, 36, 19, 11, 27, 56, 55, 42, 59, 84, 83, 29, 0, 0, 0, 
    120, 105, 157, 116, 0, 0, 0, 0, 6, 81, 89, 76, 59, 34, 39, 60, 72, 55, 38, 60, 88, 69, 63, 67, 70, 76, 78, 79, 66, 8, 0, 0, 
    136, 81, 125, 93, 0, 0, 0, 0, 0, 0, 0, 9, 46, 49, 44, 58, 72, 67, 61, 104, 128, 79, 51, 38, 48, 72, 78, 82, 82, 68, 0, 0, 
    139, 88, 114, 65, 0, 0, 0, 0, 0, 0, 0, 0, 23, 58, 61, 53, 79, 97, 87, 118, 102, 41, 26, 25, 53, 54, 57, 79, 95, 94, 48, 8, 
    139, 93, 136, 75, 0, 0, 0, 0, 0, 0, 0, 0, 36, 56, 60, 64, 69, 84, 98, 124, 67, 22, 24, 34, 59, 52, 49, 73, 98, 88, 47, 25, 
    141, 97, 148, 101, 0, 0, 0, 0, 0, 0, 0, 47, 59, 14, 8, 54, 69, 55, 74, 108, 59, 36, 58, 76, 85, 82, 79, 92, 95, 61, 10, 12, 
    145, 104, 137, 98, 42, 0, 0, 0, 0, 12, 32, 106, 105, 32, 0, 7, 34, 43, 59, 72, 41, 31, 42, 51, 63, 81, 91, 79, 47, 4, 0, 0, 
    149, 111, 131, 105, 98, 60, 0, 0, 0, 5, 19, 30, 11, 0, 0, 0, 1, 15, 37, 32, 0, 26, 58, 55, 56, 64, 58, 28, 0, 0, 0, 0, 
    163, 126, 133, 112, 114, 87, 58, 19, 12, 0, 2, 0, 0, 0, 0, 16, 33, 34, 10, 0, 0, 0, 25, 35, 38, 42, 30, 5, 0, 0, 0, 0, 
    160, 129, 144, 119, 110, 108, 89, 53, 40, 38, 17, 0, 0, 3, 37, 80, 71, 43, 32, 9, 0, 0, 0, 0, 20, 35, 15, 0, 0, 0, 0, 0, 
    131, 99, 130, 118, 103, 109, 109, 69, 37, 68, 63, 11, 21, 33, 72, 127, 103, 49, 11, 19, 68, 50, 0, 11, 67, 74, 30, 0, 0, 0, 0, 0, 
    99, 70, 103, 101, 95, 102, 122, 137, 98, 47, 34, 39, 50, 53, 101, 125, 119, 74, 0, 0, 0, 6, 28, 62, 90, 73, 5, 0, 0, 0, 0, 0, 
    88, 69, 89, 86, 83, 74, 98, 165, 228, 200, 128, 138, 168, 163, 168, 132, 123, 132, 74, 14, 10, 52, 125, 165, 180, 136, 58, 12, 0, 0, 0, 6, 
    125, 114, 100, 93, 92, 85, 115, 176, 194, 222, 230, 193, 164, 147, 98, 60, 69, 84, 103, 126, 161, 192, 209, 234, 244, 216, 178, 141, 123, 132, 145, 104, 
    167, 135, 100, 112, 116, 122, 162, 200, 137, 76, 89, 97, 80, 63, 35, 34, 67, 101, 128, 174, 229, 250, 247, 243, 247, 257, 255, 239, 233, 239, 255, 177, 
    226, 157, 86, 103, 102, 91, 134, 158, 88, 49, 42, 96, 152, 159, 154, 158, 173, 193, 208, 224, 240, 247, 254, 261, 269, 280, 285, 277, 268, 273, 286, 196, 
    294, 261, 159, 108, 94, 79, 114, 113, 54, 41, 108, 201, 234, 241, 235, 233, 237, 238, 241, 253, 265, 270, 275, 287, 297, 295, 287, 287, 292, 303, 320, 230, 
    310, 316, 258, 169, 104, 109, 148, 106, 55, 84, 188, 243, 247, 241, 236, 235, 238, 245, 255, 268, 283, 293, 304, 305, 296, 278, 265, 277, 306, 326, 332, 225, 
    302, 314, 293, 246, 166, 133, 144, 107, 83, 163, 238, 247, 250, 243, 236, 239, 246, 256, 266, 277, 287, 290, 292, 296, 289, 273, 277, 303, 328, 318, 282, 159, 
    299, 315, 309, 291, 247, 165, 105, 78, 103, 191, 246, 253, 256, 262, 258, 247, 242, 251, 265, 274, 286, 291, 286, 277, 277, 294, 321, 344, 332, 274, 227, 138, 
    310, 322, 315, 307, 285, 226, 116, 58, 106, 186, 214, 233, 246, 254, 264, 264, 264, 271, 276, 279, 282, 285, 286, 279, 285, 316, 353, 368, 334, 280, 247, 170, 
    299, 313, 308, 308, 294, 269, 213, 141, 152, 216, 221, 223, 218, 216, 224, 238, 255, 272, 286, 295, 294, 284, 276, 280, 297, 329, 358, 349, 317, 297, 282, 184, 
    282, 291, 295, 296, 288, 271, 253, 228, 220, 236, 245, 246, 236, 223, 205, 196, 207, 227, 251, 271, 275, 270, 266, 272, 285, 296, 300, 294, 285, 276, 285, 189, 
    120, 65, 79, 88, 84, 78, 68, 68, 74, 81, 91, 91, 87, 91, 85, 71, 58, 50, 44, 39, 38, 50, 66, 66, 55, 31, 11, 18, 50, 82, 98, 68, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    59, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    88, 11, 19, 11, 0, 0, 0, 0, 0, 7, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    111, 14, 43, 45, 0, 0, 0, 0, 0, 65, 38, 0, 15, 15, 0, 0, 0, 0, 0, 0, 41, 3, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    124, 9, 61, 56, 0, 0, 0, 0, 0, 38, 22, 0, 16, 31, 0, 0, 0, 0, 0, 0, 59, 19, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    130, 4, 65, 70, 0, 0, 0, 0, 0, 5, 0, 0, 0, 45, 0, 0, 0, 0, 0, 26, 67, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    130, 0, 68, 91, 0, 0, 0, 0, 0, 0, 0, 0, 11, 39, 11, 0, 0, 0, 0, 42, 61, 15, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    127, 9, 71, 92, 0, 0, 0, 0, 0, 0, 0, 37, 60, 23, 10, 0, 0, 0, 0, 22, 49, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    130, 28, 74, 89, 41, 0, 0, 0, 0, 0, 0, 35, 58, 29, 0, 0, 0, 0, 0, 0, 5, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    138, 56, 80, 91, 77, 0, 0, 0, 0, 0, 0, 25, 21, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    138, 81, 92, 98, 95, 20, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    121, 85, 92, 99, 96, 45, 0, 36, 10, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    86, 82, 78, 82, 89, 60, 10, 52, 58, 0, 0, 0, 0, 0, 9, 48, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    52, 86, 65, 67, 81, 58, 5, 59, 114, 68, 1, 0, 16, 18, 53, 78, 48, 5, 0, 0, 0, 0, 0, 1, 11, 10, 0, 0, 0, 0, 0, 0, 
    45, 110, 77, 64, 79, 57, 3, 72, 120, 110, 76, 26, 50, 79, 92, 95, 79, 39, 25, 10, 9, 21, 36, 52, 73, 67, 62, 48, 36, 27, 35, 31, 
    61, 129, 109, 86, 88, 60, 14, 94, 132, 131, 87, 84, 82, 96, 95, 93, 96, 76, 61, 50, 65, 82, 92, 103, 115, 122, 124, 120, 119, 115, 120, 89, 
    98, 139, 113, 114, 104, 45, 49, 119, 136, 126, 105, 82, 88, 95, 90, 92, 95, 92, 94, 96, 108, 117, 120, 131, 136, 144, 145, 145, 146, 143, 148, 113, 
    130, 153, 118, 107, 116, 50, 72, 130, 129, 99, 92, 93, 101, 105, 100, 100, 105, 110, 111, 116, 125, 134, 136, 140, 151, 152, 152, 152, 157, 156, 166, 130, 
    145, 165, 135, 115, 100, 63, 108, 147, 114, 84, 95, 118, 118, 116, 113, 110, 108, 109, 114, 120, 132, 143, 150, 153, 155, 156, 156, 157, 173, 178, 178, 142, 
    153, 176, 151, 131, 103, 70, 151, 167, 92, 80, 109, 119, 129, 119, 110, 112, 112, 116, 121, 129, 143, 147, 158, 167, 169, 161, 158, 170, 188, 186, 180, 141, 
    153, 180, 166, 149, 127, 95, 140, 183, 74, 94, 116, 124, 129, 123, 118, 113, 115, 121, 132, 139, 148, 157, 160, 164, 163, 165, 168, 186, 194, 192, 159, 122, 
    159, 178, 171, 168, 148, 123, 122, 147, 91, 95, 109, 121, 132, 129, 127, 121, 122, 128, 134, 141, 150, 152, 155, 155, 157, 166, 181, 203, 208, 181, 129, 105, 
    155, 181, 165, 171, 159, 139, 123, 123, 90, 99, 104, 115, 119, 122, 125, 121, 122, 131, 141, 151, 149, 145, 145, 141, 148, 167, 197, 209, 192, 164, 137, 92, 
    148, 174, 156, 161, 157, 145, 123, 115, 104, 101, 101, 114, 113, 116, 108, 103, 113, 126, 137, 150, 149, 140, 135, 127, 144, 166, 194, 200, 181, 156, 144, 89, 
    51, 85, 75, 77, 74, 69, 57, 46, 46, 41, 39, 44, 42, 45, 44, 37, 37, 45, 56, 70, 70, 61, 59, 55, 64, 79, 97, 101, 90, 70, 70, 33, 
    
    -- channel=11
    155, 255, 251, 258, 263, 258, 260, 262, 262, 262, 252, 250, 259, 267, 270, 270, 267, 261, 256, 255, 252, 244, 241, 238, 239, 240, 235, 233, 230, 227, 219, 197, 
    51, 148, 138, 144, 153, 152, 159, 162, 163, 160, 149, 145, 151, 157, 159, 161, 163, 163, 155, 142, 124, 111, 103, 106, 118, 127, 141, 145, 143, 147, 148, 173, 
    58, 155, 143, 142, 149, 153, 163, 164, 167, 164, 153, 165, 186, 169, 155, 160, 160, 157, 132, 101, 102, 101, 96, 77, 74, 84, 100, 131, 148, 155, 155, 180, 
    60, 160, 157, 156, 154, 154, 159, 164, 161, 157, 153, 205, 260, 192, 149, 142, 124, 83, 67, 97, 135, 143, 134, 116, 91, 78, 95, 107, 130, 148, 153, 178, 
    53, 150, 142, 143, 150, 152, 153, 158, 156, 151, 130, 146, 184, 153, 110, 67, 39, 53, 64, 104, 135, 153, 164, 147, 133, 127, 99, 72, 93, 132, 152, 180, 
    31, 118, 93, 67, 124, 159, 160, 161, 165, 157, 88, 83, 109, 116, 104, 82, 91, 99, 71, 91, 138, 147, 125, 124, 135, 136, 102, 73, 63, 107, 147, 180, 
    28, 123, 81, 54, 115, 163, 162, 160, 164, 167, 135, 110, 111, 154, 179, 145, 131, 119, 78, 78, 134, 153, 122, 101, 110, 123, 109, 76, 53, 76, 128, 180, 
    50, 204, 130, 101, 166, 172, 159, 158, 158, 167, 153, 118, 139, 180, 183, 134, 109, 107, 73, 44, 80, 149, 140, 92, 84, 99, 116, 100, 55, 48, 108, 187, 
    53, 229, 178, 157, 211, 195, 161, 146, 166, 239, 261, 199, 153, 168, 153, 118, 93, 98, 58, 11, 57, 144, 152, 128, 103, 110, 125, 126, 86, 43, 64, 165, 
    39, 213, 145, 183, 223, 197, 151, 121, 131, 267, 284, 190, 134, 159, 150, 136, 115, 89, 78, 33, 93, 174, 186, 169, 113, 114, 137, 137, 111, 53, 40, 124, 
    13, 175, 101, 157, 222, 208, 157, 84, 4, 66, 175, 141, 131, 173, 179, 138, 129, 126, 85, 47, 150, 204, 173, 150, 100, 101, 125, 138, 134, 94, 57, 109, 
    27, 146, 57, 137, 221, 201, 177, 86, 0, 0, 120, 92, 103, 197, 210, 164, 141, 164, 109, 46, 153, 174, 149, 125, 87, 92, 111, 124, 132, 127, 102, 127, 
    27, 146, 59, 146, 189, 141, 161, 157, 42, 15, 92, 91, 118, 205, 245, 189, 155, 175, 106, 36, 139, 166, 147, 121, 90, 76, 81, 104, 136, 139, 139, 158, 
    34, 164, 78, 158, 172, 115, 133, 174, 84, 37, 99, 125, 148, 167, 180, 163, 154, 166, 73, 39, 141, 168, 151, 145, 116, 95, 105, 116, 144, 149, 149, 171, 
    34, 164, 89, 177, 196, 132, 119, 178, 119, 82, 98, 137, 195, 169, 118, 132, 124, 133, 74, 46, 120, 167, 162, 128, 102, 96, 107, 118, 136, 137, 138, 184, 
    27, 166, 99, 175, 225, 163, 111, 184, 172, 107, 54, 117, 146, 134, 97, 78, 100, 128, 83, 62, 124, 136, 143, 135, 99, 75, 82, 94, 107, 122, 143, 196, 
    16, 175, 116, 159, 228, 175, 89, 148, 189, 122, 23, 9, 52, 83, 86, 88, 103, 113, 122, 103, 48, 66, 152, 142, 73, 44, 45, 74, 119, 140, 160, 200, 
    3, 178, 130, 138, 210, 180, 95, 105, 199, 155, 77, 25, 48, 119, 121, 141, 140, 112, 117, 123, 84, 83, 84, 71, 51, 38, 63, 101, 149, 158, 158, 196, 
    0, 163, 139, 132, 195, 203, 104, 70, 145, 147, 149, 103, 77, 132, 122, 182, 187, 98, 104, 179, 153, 109, 75, 62, 64, 84, 120, 139, 162, 160, 157, 198, 
    0, 132, 151, 135, 171, 202, 123, 68, 138, 175, 139, 82, 63, 89, 126, 211, 212, 129, 84, 80, 76, 72, 65, 60, 53, 91, 115, 140, 161, 156, 148, 192, 
    0, 105, 164, 138, 157, 190, 117, 84, 186, 253, 230, 144, 150, 162, 166, 208, 236, 182, 119, 63, 35, 57, 76, 92, 78, 83, 90, 106, 117, 120, 114, 165, 
    0, 84, 167, 144, 151, 176, 114, 102, 258, 332, 325, 248, 154, 108, 92, 104, 137, 142, 116, 107, 104, 111, 123, 118, 109, 94, 74, 81, 102, 101, 93, 156, 
    0, 35, 106, 130, 161, 207, 165, 132, 203, 261, 216, 90, 9, 0, 0, 0, 8, 43, 83, 106, 112, 106, 94, 83, 79, 76, 78, 81, 90, 92, 92, 158, 
    0, 0, 15, 59, 143, 178, 118, 146, 188, 150, 84, 39, 20, 18, 19, 23, 48, 67, 75, 72, 73, 79, 74, 68, 72, 82, 90, 87, 91, 92, 89, 159, 
    0, 35, 2, 6, 65, 105, 89, 161, 177, 123, 73, 85, 87, 88, 88, 81, 78, 78, 75, 74, 74, 76, 80, 82, 88, 101, 104, 98, 96, 92, 101, 197, 
    9, 105, 44, 2, 33, 56, 97, 173, 178, 104, 74, 81, 87, 80, 73, 75, 80, 83, 85, 87, 85, 87, 95, 102, 97, 88, 80, 72, 77, 107, 131, 212, 
    0, 110, 79, 33, 28, 3, 50, 180, 202, 116, 91, 80, 80, 86, 76, 74, 80, 86, 87, 86, 86, 87, 82, 79, 80, 73, 59, 58, 91, 113, 86, 154, 
    0, 102, 90, 73, 36, 0, 0, 128, 184, 101, 87, 81, 93, 102, 94, 83, 72, 69, 71, 78, 78, 71, 67, 67, 72, 74, 80, 91, 93, 63, 31, 113, 
    0, 114, 86, 76, 64, 0, 0, 40, 98, 75, 64, 58, 77, 98, 103, 94, 80, 81, 86, 82, 83, 83, 75, 65, 67, 90, 111, 109, 95, 88, 60, 116, 
    0, 108, 83, 69, 78, 52, 2, 42, 73, 69, 50, 43, 50, 54, 67, 79, 87, 92, 95, 104, 111, 99, 82, 76, 83, 105, 126, 146, 138, 118, 71, 124, 
    0, 102, 87, 71, 74, 87, 76, 75, 83, 83, 64, 53, 48, 43, 48, 40, 37, 55, 80, 106, 117, 104, 95, 85, 76, 90, 115, 132, 117, 96, 74, 130, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 
    
    -- channel=12
    117, 162, 171, 173, 165, 160, 164, 163, 160, 158, 161, 166, 166, 169, 169, 168, 163, 157, 156, 158, 156, 151, 150, 148, 148, 141, 136, 133, 129, 121, 110, 63, 
    122, 128, 137, 144, 139, 138, 144, 142, 141, 136, 133, 141, 145, 145, 143, 140, 136, 131, 129, 125, 119, 111, 111, 113, 120, 121, 120, 113, 108, 99, 89, 47, 
    121, 123, 131, 140, 135, 139, 147, 145, 143, 142, 151, 163, 154, 142, 143, 145, 145, 135, 116, 102, 92, 81, 75, 77, 86, 95, 112, 115, 113, 107, 98, 52, 
    124, 130, 136, 146, 140, 144, 150, 148, 143, 147, 185, 234, 207, 154, 145, 144, 126, 102, 87, 99, 117, 116, 99, 76, 62, 63, 78, 101, 116, 114, 105, 57, 
    128, 136, 141, 149, 142, 140, 143, 142, 137, 140, 181, 259, 226, 146, 115, 96, 62, 41, 65, 131, 155, 158, 144, 121, 102, 82, 69, 75, 103, 116, 108, 57, 
    120, 109, 91, 114, 140, 142, 142, 141, 138, 135, 132, 157, 128, 105, 67, 34, 33, 47, 95, 157, 171, 160, 142, 130, 120, 100, 49, 40, 80, 119, 117, 64, 
    110, 83, 24, 53, 127, 149, 144, 147, 148, 142, 125, 122, 120, 129, 107, 78, 86, 80, 102, 169, 197, 160, 121, 116, 120, 89, 46, 30, 52, 101, 116, 65, 
    138, 112, 51, 95, 148, 150, 141, 148, 160, 152, 121, 123, 155, 176, 140, 99, 102, 92, 86, 138, 192, 172, 120, 100, 95, 70, 45, 23, 29, 77, 113, 70, 
    192, 163, 113, 181, 205, 161, 144, 168, 215, 231, 182, 167, 207, 203, 144, 92, 81, 75, 61, 87, 154, 175, 139, 98, 77, 78, 67, 44, 12, 39, 99, 75, 
    214, 201, 187, 246, 231, 170, 140, 174, 292, 371, 315, 250, 235, 198, 147, 106, 83, 61, 42, 88, 182, 200, 174, 126, 98, 97, 88, 71, 28, 11, 55, 55, 
    209, 189, 213, 274, 242, 170, 135, 128, 240, 336, 306, 237, 246, 214, 163, 128, 97, 61, 45, 136, 250, 239, 196, 128, 96, 111, 105, 82, 51, 21, 33, 26, 
    216, 169, 210, 266, 252, 185, 153, 96, 125, 217, 242, 209, 258, 259, 192, 146, 120, 93, 60, 184, 292, 236, 175, 104, 82, 102, 109, 99, 79, 57, 46, 16, 
    216, 160, 209, 261, 224, 172, 163, 115, 89, 180, 195, 186, 258, 306, 238, 175, 154, 131, 96, 210, 279, 208, 150, 94, 82, 84, 95, 98, 100, 86, 77, 26, 
    221, 174, 237, 266, 172, 132, 158, 130, 78, 150, 190, 231, 286, 305, 251, 202, 168, 131, 103, 221, 262, 203, 150, 105, 85, 80, 95, 118, 127, 106, 97, 47, 
    235, 199, 256, 272, 165, 127, 156, 141, 85, 133, 197, 300, 304, 245, 193, 188, 171, 125, 100, 203, 244, 197, 157, 123, 100, 106, 124, 141, 138, 108, 100, 62, 
    250, 227, 268, 280, 198, 140, 170, 167, 116, 143, 210, 315, 315, 221, 158, 149, 130, 112, 114, 184, 212, 190, 151, 96, 68, 91, 116, 124, 117, 101, 109, 77, 
    267, 256, 275, 294, 241, 149, 174, 196, 147, 118, 155, 200, 176, 130, 125, 117, 111, 120, 130, 150, 151, 171, 159, 111, 67, 68, 89, 100, 102, 112, 135, 85, 
    280, 282, 281, 294, 263, 153, 152, 204, 203, 133, 128, 111, 117, 120, 125, 135, 112, 138, 165, 130, 69, 105, 110, 54, 18, 27, 61, 103, 128, 144, 147, 85, 
    271, 289, 283, 288, 274, 186, 143, 190, 208, 178, 132, 82, 130, 156, 181, 203, 133, 123, 178, 172, 137, 110, 48, 14, 24, 54, 89, 132, 152, 151, 137, 81, 
    241, 283, 278, 280, 275, 210, 146, 182, 196, 177, 150, 95, 129, 157, 218, 260, 177, 113, 129, 130, 117, 73, 18, 13, 36, 95, 136, 167, 165, 148, 135, 81, 
    199, 279, 281, 276, 268, 212, 156, 234, 292, 226, 148, 115, 170, 212, 287, 304, 231, 155, 108, 48, 22, 12, 19, 31, 48, 94, 126, 158, 153, 134, 127, 73, 
    158, 283, 291, 277, 263, 199, 158, 278, 413, 393, 299, 234, 249, 277, 295, 280, 233, 179, 134, 77, 40, 52, 79, 99, 113, 115, 127, 135, 131, 117, 111, 66, 
    114, 260, 286, 286, 275, 233, 231, 356, 434, 398, 294, 203, 152, 148, 141, 135, 118, 94, 92, 84, 94, 102, 104, 106, 110, 108, 111, 119, 125, 114, 108, 74, 
    60, 161, 210, 265, 278, 263, 302, 410, 404, 301, 161, 75, 67, 66, 60, 61, 65, 72, 81, 78, 86, 94, 95, 95, 100, 109, 113, 116, 116, 109, 111, 77, 
    52, 95, 118, 190, 235, 236, 314, 406, 340, 200, 94, 86, 95, 96, 93, 88, 84, 81, 77, 75, 81, 89, 93, 101, 114, 128, 132, 130, 128, 125, 134, 103, 
    76, 110, 97, 128, 179, 233, 356, 386, 258, 110, 80, 100, 101, 96, 89, 85, 81, 79, 80, 85, 93, 103, 112, 122, 130, 134, 128, 126, 136, 152, 174, 143, 
    80, 112, 96, 95, 125, 211, 362, 355, 198, 92, 97, 103, 104, 89, 83, 87, 89, 91, 93, 100, 104, 109, 124, 131, 125, 108, 99, 110, 143, 167, 170, 121, 
    76, 110, 101, 99, 102, 154, 285, 303, 161, 107, 106, 106, 110, 102, 91, 87, 87, 92, 98, 104, 106, 102, 102, 107, 108, 101, 106, 129, 153, 136, 102, 69, 
    82, 111, 101, 103, 101, 100, 161, 188, 109, 80, 89, 100, 117, 119, 112, 100, 91, 93, 100, 105, 105, 99, 97, 94, 99, 117, 141, 159, 139, 89, 56, 57, 
    96, 121, 99, 101, 102, 93, 87, 98, 58, 57, 53, 65, 83, 95, 104, 105, 112, 121, 128, 128, 118, 103, 92, 90, 114, 158, 191, 187, 144, 102, 67, 53, 
    89, 118, 98, 99, 99, 101, 91, 85, 68, 56, 51, 56, 54, 53, 56, 68, 89, 111, 132, 150, 141, 114, 98, 101, 137, 184, 216, 193, 134, 89, 69, 43, 
    21, 42, 29, 26, 23, 26, 24, 16, 12, 0, 0, 2, 0, 0, 0, 0, 0, 16, 39, 56, 51, 36, 31, 31, 51, 79, 94, 74, 36, 10, 14, 2, 
    
    -- channel=13
    162, 129, 139, 135, 125, 127, 127, 125, 121, 117, 125, 133, 136, 134, 131, 127, 119, 114, 118, 118, 112, 112, 113, 116, 113, 107, 104, 103, 97, 84, 74, 0, 
    182, 105, 119, 117, 111, 117, 116, 112, 106, 103, 109, 120, 122, 117, 111, 107, 98, 92, 87, 83, 81, 81, 91, 97, 101, 105, 97, 88, 81, 69, 58, 0, 
    177, 97, 114, 117, 111, 117, 118, 112, 109, 112, 138, 146, 113, 104, 110, 109, 106, 85, 69, 77, 67, 59, 54, 65, 77, 88, 103, 95, 86, 76, 66, 0, 
    179, 100, 116, 120, 114, 120, 121, 113, 112, 124, 203, 215, 117, 98, 111, 101, 76, 62, 86, 101, 103, 92, 76, 60, 51, 67, 73, 91, 97, 85, 71, 0, 
    179, 100, 117, 128, 115, 116, 115, 109, 107, 120, 203, 217, 136, 83, 70, 60, 45, 45, 100, 150, 152, 138, 111, 92, 90, 54, 51, 80, 107, 97, 77, 0, 
    169, 60, 61, 125, 132, 114, 114, 109, 107, 109, 142, 137, 73, 58, 28, 23, 26, 56, 145, 195, 166, 133, 116, 119, 98, 54, 21, 45, 106, 116, 88, 0, 
    169, 17, 7, 93, 133, 118, 113, 116, 111, 100, 92, 98, 110, 95, 52, 62, 78, 76, 144, 214, 186, 117, 99, 113, 95, 46, 8, 30, 86, 120, 97, 0, 
    202, 20, 38, 147, 138, 112, 111, 120, 128, 99, 72, 125, 164, 139, 80, 75, 93, 79, 108, 185, 199, 126, 85, 88, 83, 47, 19, 1, 50, 116, 112, 0, 
    260, 75, 115, 206, 163, 109, 110, 160, 229, 185, 122, 156, 205, 158, 90, 70, 76, 56, 64, 156, 191, 139, 98, 73, 68, 65, 46, 12, 4, 73, 117, 0, 
    286, 125, 214, 246, 157, 108, 100, 199, 343, 321, 220, 230, 229, 153, 103, 78, 64, 42, 44, 173, 228, 173, 119, 74, 92, 93, 63, 32, 0, 32, 88, 0, 
    282, 145, 245, 271, 161, 107, 91, 155, 316, 354, 235, 223, 247, 168, 115, 92, 77, 17, 68, 251, 268, 192, 130, 71, 94, 111, 87, 47, 12, 17, 62, 0, 
    275, 133, 268, 261, 166, 126, 109, 87, 222, 273, 193, 212, 291, 208, 124, 108, 99, 35, 96, 304, 279, 176, 107, 60, 84, 108, 91, 76, 52, 43, 46, 0, 
    270, 132, 284, 231, 133, 136, 131, 59, 152, 237, 176, 218, 299, 256, 145, 128, 130, 62, 141, 315, 257, 135, 87, 58, 76, 90, 98, 98, 81, 71, 56, 0, 
    278, 154, 306, 204, 85, 115, 143, 63, 99, 193, 207, 259, 297, 246, 178, 167, 138, 63, 153, 310, 230, 137, 104, 70, 71, 87, 106, 123, 109, 81, 71, 0, 
    303, 184, 308, 202, 67, 110, 155, 77, 84, 166, 255, 341, 264, 178, 159, 156, 134, 84, 150, 274, 223, 141, 99, 80, 91, 115, 137, 147, 112, 82, 89, 0, 
    334, 205, 306, 238, 89, 105, 174, 117, 85, 155, 289, 329, 241, 167, 136, 135, 110, 86, 160, 240, 193, 150, 110, 55, 59, 107, 127, 125, 98, 92, 99, 0, 
    370, 223, 298, 275, 132, 96, 190, 181, 88, 129, 201, 218, 149, 89, 113, 103, 96, 121, 146, 128, 150, 174, 102, 49, 59, 89, 112, 109, 98, 108, 110, 0, 
    398, 245, 288, 287, 172, 87, 179, 209, 137, 110, 123, 126, 133, 98, 127, 109, 85, 153, 158, 95, 85, 99, 60, 20, 19, 63, 99, 122, 127, 130, 118, 0, 
    404, 256, 276, 284, 206, 97, 153, 212, 170, 150, 87, 90, 146, 146, 209, 164, 75, 142, 176, 128, 111, 75, 16, 0, 47, 89, 123, 146, 132, 121, 102, 0, 
    386, 270, 260, 272, 228, 119, 142, 229, 179, 119, 83, 110, 152, 192, 263, 208, 96, 103, 123, 104, 75, 31, 0, 14, 71, 119, 157, 162, 124, 103, 96, 0, 
    357, 289, 252, 267, 228, 119, 155, 319, 289, 159, 81, 119, 199, 246, 305, 257, 142, 103, 81, 19, 8, 3, 20, 48, 72, 108, 125, 133, 105, 86, 83, 0, 
    329, 313, 258, 265, 223, 121, 197, 391, 394, 283, 202, 177, 247, 287, 290, 243, 162, 115, 86, 50, 35, 53, 78, 102, 115, 114, 123, 126, 102, 87, 91, 0, 
    270, 304, 278, 280, 243, 175, 285, 440, 420, 276, 151, 154, 161, 162, 151, 133, 101, 78, 68, 65, 89, 103, 109, 111, 113, 114, 117, 122, 116, 106, 103, 0, 
    185, 206, 239, 293, 250, 231, 374, 450, 340, 172, 71, 52, 80, 83, 75, 78, 70, 69, 78, 82, 94, 98, 101, 107, 115, 122, 121, 120, 114, 107, 111, 0, 
    147, 116, 166, 240, 231, 265, 396, 397, 213, 83, 55, 78, 99, 98, 94, 93, 91, 82, 79, 84, 91, 96, 101, 114, 132, 135, 132, 129, 125, 132, 151, 2, 
    155, 93, 120, 176, 200, 310, 430, 323, 111, 42, 74, 107, 103, 96, 94, 90, 84, 80, 84, 91, 101, 113, 122, 130, 132, 131, 124, 130, 151, 169, 178, 16, 
    163, 88, 95, 121, 167, 317, 439, 252, 63, 52, 98, 109, 106, 86, 86, 94, 94, 95, 99, 107, 111, 115, 132, 138, 123, 103, 103, 139, 166, 163, 160, 8, 
    164, 92, 94, 105, 133, 256, 363, 210, 47, 85, 106, 118, 111, 96, 91, 88, 94, 102, 111, 114, 111, 110, 113, 112, 106, 103, 126, 152, 152, 118, 108, 0, 
    173, 91, 98, 109, 112, 159, 230, 135, 46, 68, 91, 116, 125, 116, 105, 100, 104, 108, 111, 113, 110, 101, 99, 103, 115, 137, 162, 161, 126, 57, 67, 0, 
    183, 99, 101, 111, 108, 107, 127, 88, 28, 50, 66, 83, 93, 101, 106, 111, 124, 132, 140, 133, 111, 96, 92, 105, 145, 192, 205, 164, 100, 63, 74, 0, 
    184, 100, 100, 109, 106, 99, 89, 85, 53, 47, 61, 69, 67, 65, 62, 81, 112, 132, 150, 150, 122, 103, 95, 118, 175, 222, 217, 153, 86, 70, 65, 0, 
    85, 52, 50, 53, 47, 43, 35, 31, 24, 13, 20, 22, 21, 19, 13, 16, 30, 49, 70, 73, 56, 46, 45, 62, 92, 118, 113, 69, 31, 27, 28, 0, 
    
    -- channel=14
    61, 63, 64, 58, 57, 61, 61, 60, 60, 64, 59, 58, 64, 66, 71, 72, 68, 65, 62, 56, 50, 49, 49, 52, 48, 45, 46, 49, 48, 43, 37, 0, 
    151, 175, 181, 176, 174, 176, 178, 175, 174, 171, 168, 172, 180, 185, 191, 191, 181, 172, 165, 161, 150, 148, 149, 151, 152, 147, 145, 147, 147, 139, 128, 21, 
    151, 171, 179, 177, 176, 180, 180, 178, 177, 172, 167, 156, 165, 180, 184, 180, 174, 156, 150, 130, 111, 100, 108, 124, 132, 151, 149, 146, 146, 141, 130, 20, 
    149, 166, 174, 179, 180, 186, 184, 182, 182, 183, 192, 151, 144, 162, 170, 162, 160, 149, 120, 92, 71, 54, 49, 59, 81, 103, 132, 144, 146, 142, 136, 23, 
    140, 162, 173, 183, 183, 187, 188, 183, 185, 190, 230, 225, 162, 145, 152, 148, 117, 100, 95, 87, 74, 59, 39, 39, 38, 52, 90, 128, 142, 137, 134, 24, 
    127, 133, 169, 189, 181, 183, 187, 182, 182, 190, 219, 226, 167, 115, 91, 84, 57, 58, 94, 99, 88, 82, 72, 60, 47, 40, 39, 90, 134, 137, 132, 25, 
    98, 76, 94, 156, 175, 181, 188, 186, 180, 178, 173, 168, 139, 89, 48, 42, 39, 45, 99, 126, 99, 83, 84, 82, 70, 38, 23, 43, 110, 140, 134, 25, 
    73, 32, 34, 91, 150, 177, 186, 183, 175, 147, 147, 136, 123, 95, 60, 58, 58, 48, 86, 153, 133, 80, 73, 89, 77, 42, 18, 16, 75, 136, 135, 22, 
    94, 19, 37, 89, 123, 162, 179, 183, 159, 107, 80, 118, 128, 109, 69, 60, 61, 54, 70, 128, 140, 98, 62, 61, 65, 48, 21, 1, 32, 116, 143, 21, 
    124, 65, 66, 121, 125, 154, 165, 204, 198, 151, 94, 126, 134, 105, 76, 47, 55, 38, 54, 101, 117, 108, 66, 52, 59, 52, 39, 11, 2, 62, 130, 29, 
    127, 100, 120, 141, 129, 148, 146, 195, 276, 227, 152, 147, 147, 95, 84, 63, 44, 22, 53, 113, 118, 117, 87, 64, 69, 69, 46, 25, 0, 16, 80, 24, 
    119, 100, 148, 151, 137, 152, 148, 146, 237, 229, 167, 175, 174, 109, 82, 78, 52, 6, 61, 146, 151, 124, 96, 61, 68, 82, 62, 39, 11, 8, 39, 0, 
    116, 89, 140, 140, 148, 165, 165, 116, 167, 195, 155, 162, 199, 145, 87, 83, 79, 24, 74, 168, 158, 114, 83, 58, 59, 77, 76, 53, 33, 29, 36, 0, 
    114, 89, 145, 115, 108, 160, 174, 120, 144, 172, 149, 151, 197, 187, 127, 96, 87, 53, 98, 169, 146, 106, 66, 45, 49, 54, 66, 67, 52, 54, 65, 0, 
    124, 98, 159, 104, 54, 124, 158, 120, 122, 141, 167, 170, 150, 167, 141, 123, 100, 60, 105, 174, 146, 98, 81, 60, 58, 60, 69, 86, 78, 81, 90, 0, 
    138, 107, 161, 116, 35, 83, 127, 116, 106, 149, 180, 225, 176, 125, 131, 121, 105, 76, 116, 162, 155, 109, 74, 52, 58, 77, 85, 101, 103, 99, 109, 10, 
    152, 112, 155, 140, 53, 58, 123, 111, 92, 129, 186, 219, 183, 122, 111, 92, 94, 90, 108, 158, 181, 134, 75, 57, 55, 77, 93, 93, 101, 113, 130, 20, 
    177, 119, 146, 155, 81, 41, 114, 124, 80, 87, 140, 151, 121, 101, 91, 66, 75, 102, 102, 103, 119, 137, 100, 53, 50, 60, 91, 97, 109, 138, 152, 28, 
    203, 140, 146, 156, 104, 37, 92, 132, 110, 80, 59, 105, 103, 103, 107, 62, 48, 114, 117, 80, 69, 84, 69, 31, 32, 46, 86, 119, 137, 154, 157, 30, 
    219, 160, 151, 158, 122, 53, 72, 111, 88, 101, 61, 76, 114, 111, 132, 96, 35, 77, 128, 121, 100, 52, 26, 24, 31, 72, 103, 145, 156, 160, 154, 33, 
    216, 170, 154, 160, 134, 75, 88, 125, 71, 35, 43, 45, 74, 101, 145, 122, 53, 40, 63, 82, 65, 26, 0, 0, 14, 55, 90, 128, 126, 120, 118, 18, 
    190, 172, 147, 156, 134, 76, 101, 166, 154, 60, 20, 64, 102, 140, 173, 152, 100, 63, 34, 10, 0, 0, 0, 0, 0, 18, 48, 68, 64, 56, 51, 0, 
    154, 178, 147, 149, 129, 75, 118, 204, 229, 163, 109, 99, 124, 142, 145, 133, 94, 55, 27, 3, 0, 0, 1, 8, 5, 3, 12, 19, 15, 6, 1, 0, 
    95, 135, 158, 155, 135, 130, 174, 231, 217, 173, 102, 52, 47, 46, 44, 41, 28, 10, 3, 4, 4, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    30, 33, 102, 154, 137, 158, 212, 231, 180, 114, 35, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 20, 98, 126, 157, 221, 203, 127, 47, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 7, 10, 3, 0, 4, 0, 
    32, 0, 0, 22, 82, 180, 227, 160, 70, 13, 6, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 3, 4, 14, 34, 0, 
    34, 0, 0, 0, 24, 151, 238, 128, 50, 17, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 12, 17, 27, 0, 
    27, 0, 0, 0, 0, 65, 177, 123, 33, 22, 14, 13, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39, 0, 0, 0, 0, 0, 57, 66, 10, 0, 2, 10, 18, 18, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 0, 
    51, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 1, 8, 17, 24, 24, 22, 11, 0, 0, 0, 0, 20, 45, 43, 12, 0, 0, 0, 0, 
    91, 37, 29, 34, 33, 32, 28, 27, 22, 10, 12, 15, 14, 14, 15, 26, 45, 61, 76, 77, 59, 43, 38, 50, 82, 113, 117, 80, 33, 16, 9, 0, 
    
    -- channel=15
    45, 26, 30, 27, 23, 26, 27, 25, 25, 25, 27, 30, 28, 27, 31, 29, 26, 27, 27, 25, 23, 23, 22, 23, 22, 21, 23, 23, 22, 20, 16, 0, 
    129, 123, 134, 136, 129, 127, 128, 127, 124, 124, 127, 132, 133, 132, 135, 137, 134, 129, 125, 119, 113, 112, 112, 116, 117, 113, 110, 111, 112, 104, 95, 36, 
    125, 118, 129, 137, 135, 132, 130, 129, 129, 124, 123, 128, 130, 132, 138, 140, 134, 122, 105, 100, 92, 90, 97, 104, 114, 117, 113, 110, 110, 103, 93, 35, 
    127, 121, 129, 138, 136, 136, 133, 131, 130, 130, 138, 131, 109, 119, 134, 133, 127, 106, 97, 86, 68, 52, 49, 67, 75, 96, 109, 110, 108, 104, 97, 36, 
    130, 127, 126, 134, 134, 137, 136, 133, 133, 135, 166, 157, 105, 106, 119, 111, 95, 97, 91, 77, 58, 47, 37, 30, 44, 51, 70, 98, 108, 104, 99, 41, 
    122, 114, 117, 130, 131, 132, 136, 133, 132, 130, 134, 174, 137, 96, 80, 84, 72, 57, 69, 77, 64, 57, 47, 49, 41, 32, 39, 73, 105, 109, 99, 41, 
    109, 68, 74, 124, 131, 128, 135, 136, 132, 129, 118, 122, 117, 86, 47, 36, 36, 32, 66, 88, 68, 54, 62, 64, 51, 39, 22, 37, 88, 114, 104, 43, 
    92, 37, 22, 81, 114, 124, 133, 138, 137, 125, 106, 103, 102, 77, 44, 36, 41, 31, 55, 102, 96, 60, 56, 64, 63, 37, 25, 24, 61, 108, 108, 40, 
    96, 20, 33, 70, 87, 114, 131, 133, 138, 102, 81, 93, 95, 77, 50, 42, 51, 46, 41, 90, 123, 81, 47, 52, 59, 44, 21, 14, 36, 93, 112, 38, 
    128, 35, 41, 89, 89, 102, 123, 149, 160, 119, 58, 76, 101, 85, 63, 44, 39, 38, 45, 77, 103, 87, 59, 37, 44, 47, 34, 18, 10, 56, 110, 46, 
    123, 65, 76, 95, 94, 100, 108, 141, 186, 165, 114, 106, 118, 83, 71, 47, 38, 28, 37, 92, 99, 78, 65, 42, 53, 50, 36, 29, 17, 22, 73, 45, 
    121, 46, 101, 112, 98, 100, 109, 86, 170, 193, 136, 121, 138, 92, 57, 65, 41, 20, 40, 111, 108, 75, 71, 47, 52, 65, 46, 33, 23, 18, 37, 24, 
    121, 39, 103, 111, 104, 114, 124, 86, 109, 159, 118, 130, 152, 115, 56, 59, 62, 26, 38, 115, 118, 76, 65, 46, 45, 55, 56, 45, 35, 27, 34, 6, 
    124, 45, 102, 87, 86, 123, 132, 97, 88, 133, 121, 115, 136, 131, 78, 60, 64, 49, 51, 120, 108, 70, 53, 41, 39, 45, 57, 52, 41, 37, 46, 5, 
    130, 52, 111, 88, 48, 90, 126, 95, 73, 114, 125, 126, 103, 114, 109, 88, 62, 48, 65, 121, 103, 76, 59, 37, 39, 45, 47, 58, 52, 45, 67, 19, 
    143, 62, 112, 96, 35, 57, 111, 90, 64, 88, 133, 156, 92, 73, 87, 88, 82, 57, 58, 115, 114, 72, 54, 48, 48, 61, 61, 64, 65, 70, 83, 31, 
    151, 71, 111, 105, 43, 38, 96, 89, 46, 87, 124, 137, 140, 85, 79, 81, 68, 62, 78, 104, 111, 103, 60, 33, 35, 56, 66, 67, 81, 92, 98, 38, 
    159, 76, 103, 110, 63, 17, 87, 102, 63, 49, 92, 105, 106, 84, 74, 62, 53, 80, 69, 71, 103, 113, 65, 45, 43, 51, 69, 81, 89, 101, 108, 42, 
    169, 88, 93, 103, 78, 23, 57, 112, 87, 45, 52, 85, 93, 73, 78, 53, 29, 75, 95, 66, 39, 51, 64, 41, 36, 42, 58, 94, 98, 108, 112, 47, 
    170, 104, 93, 101, 89, 39, 40, 88, 92, 79, 38, 50, 91, 88, 106, 73, 16, 53, 101, 89, 62, 38, 33, 33, 39, 57, 70, 106, 115, 117, 114, 45, 
    166, 121, 93, 105, 97, 54, 45, 94, 57, 38, 59, 43, 79, 92, 100, 90, 43, 20, 57, 67, 66, 43, 14, 18, 25, 61, 86, 105, 104, 100, 96, 32, 
    150, 127, 93, 104, 94, 52, 61, 129, 118, 28, 16, 39, 61, 80, 104, 102, 70, 41, 22, 17, 16, 12, 9, 0, 2, 25, 45, 59, 58, 45, 46, 0, 
    119, 118, 94, 99, 91, 55, 71, 127, 147, 118, 38, 36, 74, 91, 103, 100, 75, 52, 41, 13, 0, 0, 0, 3, 1, 0, 5, 6, 3, 0, 0, 0, 
    68, 91, 102, 103, 96, 76, 96, 143, 137, 94, 63, 39, 38, 45, 45, 44, 36, 15, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 10, 72, 105, 88, 100, 140, 157, 107, 62, 29, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 64, 91, 103, 147, 130, 68, 31, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 0, 0, 7, 69, 113, 148, 99, 37, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 0, 0, 0, 12, 97, 150, 89, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 0, 0, 0, 0, 28, 119, 84, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 0, 0, 0, 0, 0, 26, 58, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 6, 4, 0, 0, 0, 0, 0, 0, 11, 7, 0, 0, 0, 0, 0, 
    47, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 20, 25, 28, 24, 12, 5, 1, 9, 28, 41, 44, 20, 0, 0, 0, 0, 
    
    
    others => 0);
end gold_package;
