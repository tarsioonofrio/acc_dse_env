library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -- layer=3
    -4623, -5437, -262, 4537, 8565, -5190, 9754, -9573, 3234, -3646,

    -- weights
    -- layer=3 filter=0 channel=0
    -3, -46, 2, 17, -5, 0, 4, -54, -39, -8, 1, -14, -13, 5, 13, 17, 39, -13, -28, -11, 15, 0, 6, -2, -43, 9, -17, 0, -9, 5, -49, -65, 7, 3, 6, -8, -9, -7, -27, 9, 5, 28, -11, 2, 34, 0, 5, -5, -20, 15, 45, -35, -38, 28, -11, -10, -10, -6, 0, -10, -24, -39, -6, -1, -3, 1, -16, 3, 12, 5, 33, -6, -3, 3, 4, -12, 0, 14, 2, -5, 39, 15, 8, 6, 2, -21, -13, -12, 27, -79, -7, -13, -9, -8, 24, -5, -25, 8, -4, 4, 4, 30, -16, -17, -44, -3, 21, -7, -44, -11, 7, -46, 21, -7, 2, 3, 13, -35, 22, 43, -4, -36, 10, -7, -9, 16, -25, 4, -13, -22, -17, 12, -2, -4, -31, -1, -26, -3, -1, -10, -15, -23, 0, -70, -12, -6, 5, 34, -16, 3, -12, -4, -26, 0, -7, 12, -10, -14, 56, -14, -41, 21, -1, 24, -11, 2, -11, -6, -16, -29, -27, -15, 112, 6, 3, -7, 10, 4, -54, -11, 5, -40, -38, 8, 25, -26, 8, 18, 40, 30, 5, -26, -48, 6, 16, -31, -9, -3, 2, -14, -6, 5, 16, 8, 42, -24, 15, -11, -9, -1, -4, 32, -51, -40, 57, -30, 33, 19, -33, 6, 5, -3, -48, -10, 3, 27, -5, -63, 11, -39, -11, -1, 11, -18, 12, -39, -9, -12, -35, 10, -27, 5, -2, 3, 13, -9, -24, -14, -7, 9, -11, -8, -57, 2, 39, -3, -23, -11, 8, -13, -8, -35, 4, -45, -13, -35, -1, -4, -30, 7, 25, 13, 11, -27, -1, -11, 4, 7, 0, 13, 2, 8, 27, 8, -9, 44, -57, -2, 2, 6, 1, 8, -8, 2, 19, -25, 7, -6, -20, 22, -36, 8, 10, -9, -5, 20, -12, -7, -6, 2, -11, 4, -1, -6, -6, 8, -9, 26, -10, -16, -10, -14, 17, -40, 9, -9, 11, 10, 13, 10, 10, 1, -5, 16, -7, -7, 47, 27, -7, -28, 8, 3, 3, 23, -12, -20, -35, -8, 5, 2, 13, -12, -24, -7, 5, -64, -9, 8, -3, -18, -20, -13, -16, 0, 34, 5, 7, -30, 30, -7, 13, -5, -4, 5, 1, -8, 53, 12, 1, -13, -9, 1, -31, 2, 4, 0, 37, 4, -9, 3, 19, 7, 5, -6, -11, 6, -1, -20, -28, -36, -6, -39, 38, -24, -22, 4, -24, -3, -19, 0, 0, 8, 0, 8, 28, -19, -16, 10, -56, 15, -4, -26, -18, 13, 18, -25, 24, -12, 51, 12, 3, -1, -17, -6, -8, 4, 12, -22, 37, -18, 8, -3, -11, -11, -20, -2, 12, -5, -9, 2, 21, -20, 0, -3, 1, -7, -20, 8, -49, -7, -4, 5, 28, -2, -12, 0, -78, -29, -31, -8, 22, 6, 2, -9, -31, 3, 15, -5, 3, 7, -4, 33, -15, -81, 7, -19, 4, -4, -53, -7, 0, 26, 0, 13, -20, 3, 11, 0, -1, -3, -21, -18, -29, 4, 13, 2, -12, 10, 1, 22, 0, 8, 20, 49, -11, 11, 4, -41, -7, -37, -14, -8, -5, -18, -21, -11, 30, -24, 10, -22, -24, -4, 16, -8, 3, 31, 21, 0, -5, -18, -8, -2, -19, -60, 6, -3, -2, -4, -5, 0, 0, -23, 30, 1, 17, 27, -10, 14, 5, -2, -16, -17, -11, -47, -26, -1, -4, -26, -15, -10, 11, 24, 21, 4, -3, 2, 28, -9, 11, 10, 5, -3, 37, -16, -8, 0, -16, -37, -8, 3, -1, 11, 4, 19, 6, 6, 0, 2, 9, 5, 33, -60, -22, 9, 4, 7, 26, 31, 3, -4, -29, -35, -32, 10, 18, -24, 25, -11, -23, -12, -21, -23, 21, -4, -9, 10, -28, -46, 6, -35, -6, 13, -20, -14, 0, 5, 7, -6, -9, -20, -7, -38, -13, 7, -7, 10, 36, -6, 54, -1, -2, -11, -4, 35, 16, 8, 10, 11, -27, -12, -28, 1, -3, 7, -24, -28, -11, -1, 12, -4, 7, -3, -64, -3, -48, 16, -15, 15, -18, 7, -7, 28, 54, -10, -5, 9, -11, -8, 13, 11, 15, 13, -6, -32, 11, -1, -50, 20, 5, 18, 7, -26, 0, -18, -16, 12, 0, -33, 10, 6, -14, 9, -10, 9, 31, -9, -22, -15, 9, 0, 8, 1, -35, 11, -53, 13, 30, 27, -48, 21, -71, 2, 20, -1, 32, -32, 9, -32, -12, 7, 1, -8, 0, 10, 52, 8, 29, 44, -16, -42, 30, -7, -12, -3, -6, -14, -28, 30, -44, 23, 41, -18, -24, -3, -37, 20, -42, -4, 16, 3, -11, -34, 0, -16, 0, -10, -13, -5, -6, 0, -33, 16, 21, 32, 62, 0, -29, -16, 9, 6, -13, 26, -40, 32, 14, -8, -1, 20, 6, -28, -3, -2, 9, -8, -8, -2, -3, 3, -26, 21, 15, -35, 9, -14, -10, 4, -3, -9, -8, 15, -28, 0, 7, -25, 4, 9, 0, -12, -57, -27, -6, -36, -14, 4, -9, -1, 5, 0, -5, 16, 11, -7, 10, -11, -4, 14, 0, -4, -31, -25, 2, -47, -7, -17, -2, -31, -14, -105, 18, 6, -7, -12, 0, 21, -4, -4, -4, 1, -2, 10, 28, -27, -9, 5, -17, -1, -27, -15, -39, 0, 7, -3, -7, 16, 39, -12, 15, 28, 23, -51, -50, 5, -12, -3, 39, 27, -6, -21, 27, 4, 2, -3, 16, -9, -26, -14, -15, 1, -6, 32, -21, 8, 8, -6, 12, -20, 23, 9, -74, 0, 4, 3, 10, 7, -33, 10, 71, -23, -22, -45, 9, 12, -5, 28, -14, 5, -14, -13, -37, -7, 26, 8, -15, -12, 0, -10, 31, -5, -8, -68, -20, 9, -24, 10, -13, 32, 15, -16, 7, 10, 9, 0, 15, 32, -10, 5, -8, 11, -20, -15, -41, -5, 15, -3, 10, 13, -11, 3, -29, 18, 14, -11, 32, -15, 24, 3, 11, 10, -29, 5, -26, -13, -4, 23, 20, 30, -12, -1, -4, 0, -23, -27, -1, -5, 15, -21, -30, -50, -23, -3, -8, 3, 31, -8, -37, -21, -54, 10, 4, 5, 2, -8, -3, -4, -29, 55, -5, 7, -7, 82, 5, -5, -23, 6, 3, -1, -5, 0, 14, -15, 3, -16, 19, 9, 17, 1, 30, -15, 3, -2, -13, 1, 11, -37, -19, 29, 8, 0, 3, -7, 6, -1, -38, 19, -43, 1, -42, -29, 2, 1, -10, -9, -10, -11, 25, 14, -19, 17, 8, -1, -47, 14, 1, -24, 33, -29, -7, -18, 2, 10, 28, -45, 10, 6, -13, 4, 6, 3, 0, -49, 4, 23, 8, 11, 18, -30, 4, 13, 11, 18, -1, 31, 29, 33, 6, -37, 13, -15, 17, 8, -13, -11, -12, -14, 26, -22, 23, -7, -15, -23, -25, -4, 21, 2, 34, 16, -15, -1, 13, -5, 11, 7, 28, 3, 30, 8, -16, -3, -2, 9, 77, 35, -3, -35, 23, 10, 5, -2, 2, -1, -9, 14, -16, 0, 0, -5, -25, 14, -2, 10, 7, 0, -13, -8, -15, 2, -25, 2, 12, -9, 14, 6, -15, 11, -22, -4, -1, -2, -13, 38, 5, -6, 2, 20, -28, -10, -27, -7, -5, 4, -7, 3, 11, -10, 12, -32, -44, -32, 11, 21, -3, 22, -17, -69, 22, -24, 11, -26, -10, 16, -1, -1, 13, -5, -9, 24, 20, 11, -1, -38, 7, 8, -49, 4, -46, 5, -6, 27, -8, -14, -35, -43, -17, 9, -13, -3, 13, -4, -6, 33, 32, -30, -6, 34, -6, 8, -54, -4, -30, -17, -25, -16, -14, -19, 10, 0, 26, 1, -21, -14, -7, -21, 10, 36, -2, -11, 49, 24, -4, -2, -14, 22, -2, -19, 18, 5, -19, -10, -9, 23, -7, -20, -41, -29, 41, 16, 0, 0, -18, 25, 17, 2, 24, 15, -60, 32, -28, 11, 1, -14, -38, -71, 0, -4, 3, 7, 8, 4, 9, 35, -17, 17, -26, -20, 12, 18, -2, 5, 2, 30, 3, -64, 46, -10, 7, -4, -60, 8, 12, 17, 18, 2, -11, 7, -11, -2, 12, -4, 1, -3, -1, 35, 10, -5, 15, 12, -7, -18, 5, -6, -20, -31, -3, 36, 1, 2, -11, 8, 7, -77, 23, -13, 8, 14, 25, 31, 5, -7, -28, -33, -18, -47, -5, -5, 33, -9, -36, 0, -68, 6, -10, 20, -31, -10, 19, -13, -18, -22, -19, 6, 17, 1, -25, -6, 3, 8, -10, -11, -11, -13, 17, -21, -1, -3, -25, 5, 5, -25, -3, -2, -15, 33, 0, -7, -7, 43, -20, -13, 23, -3, -55, 0, -4, 5, -4, 9, 0, 7, -5, -14, -43, -36, -31, 36, -10, 3, -6, 8, 9, 35, 68, 10, -32, -10, -15, 0, -14, -8, 37, 2, -8, 7, -18, 0, 30, -3, -16, 14, 30, -24, -14, -23, -34, -31, 19, 17, 5, 9, 19, 5, 32, 4, 4, 17, -24, 30, -15, -7, -10, -10, 30, 18, 10, -26, -16, 26, -41, -8, -22, 0, 32, -8, 6, -18, 0, -18, 17, 42, -1, 11, 0, -5, -36, 28, -14, -30, -45, 29, 3, -51, 30, -5, -8, -11, -58, -8, -17, 67, 4, 18, -10, 0, 5, 17, -25, -10, -7, -9, 8, -14, 0, 27, -16, 22, -21, 12, 4, 0, 16, -2, -6, 11, 48, -10, -43, 34, -8, -3, 30, 17, 23, 4, 30, -43, -1, 8, 9, -1, 11, 2, 15, -6, -11, -4, 40, -7, 20, -9, 48, 0, 40, 17, 1, 4, 11, 37, 30, 37, -17, -12, 5, 0, 17, 7, -7, -31, 43, -6, -4, -9, 3, -6, -15, 3, -4, 0, -9, -22, -5, 2, 8, -39, -2, -5, -6, -6, -14, -16, -5, 0, 9, 31, 2, -12, -40, -48, -27, 21, -5, -18, 33, 20, 10, 14, 5, 6, -14, 13, 2, -18, 25, 9, -25, -1, -41, -23, -9, -8, 29, 6, -21, -19, 17, 27, -58, -8, -11, 42, 28, 1, 12, 15, 50, -37, 6, -29, 47, 28, 9, 10, 17, 9, 42, 32, -6, 3, -3, 24, 3, -2, 9, -12, -2, 1, 21, -8, -38, -10, 4, 26, 3, 0, 30, 2, 23, 14, 7, 6, 22, 1, -11, 4, -8, -5, -13, 2, 21, 2, -24, 1, 2, -9, 13, 0, 7, -1, 5, -35, 40, -12, -6, -46, 0, -28, -18, -31, -12, 13, 47, 2, 36, 8, 0, 9, -26, -8, 26, -16, -31, -16, -15, -40, 11, -19, -50, -14, -2, -13, -17, -36, -25, -2, 24, -25, -15, -6, -33, -1, 33, 19, 6, -17, 20, 15, 8, 47, 1, -5, 7, 24, -32, -26, -30, 17, 6, 7, -36, -10, 8, -8, 71, 14, -14, 37, 15, -23, -23, -2, -20, -14, -16, -12, -10, 14, 8, -18, 7, 27, 18, 12, -27, -14, -14, 13, -24, 9, 25, -5, 23, -9, 0, 14, -6, 9, -15, -3, 34, -4, 17, 7, 4, -3, 27, 51, -7, 4, -5, -13, 9, -10, -14, -14, 67, 0, 13, -9, -17, -8, 5, 5, -4, -9, 14, -6, 5, -24, -8, -19, -27, 10, -6, -1, 2, -21, -11, 3, 19, 6, -27, -5, 0, -4, 5, 8, 8, 2, 22, 6, -4, -46, 9, 7, 30, -7, -6, -15, 5, -4, 1, 8, 25, 23, -62, 27, -3, -17, -1, -17, 18, -1, -25, -22, 17, 15, 7, -13, 17, -7, 40, -4, -4, 55, -5, 2, 19, -10, 19, -25, 23, 11, -2, -2, -46, 46, 2, -5, 0, 2, 32, 27, 0, -21, 18, 11, 6, 4, 6, -3, 0, -24, -14, -3, 7, -31, 12, -12, 11, -7, -22, 26, 19, 2, -127, 7, -12, -22, 8, -5, -1, -11, 18, -21, -5, 16, 22, 6, -7, -37, -12, 12, -8, 23, -9, -1, -14, 0, 0, 0, -14, 6, -13, -6, 3, -10, 21, 12, 17, -28, -9, -6, -2, 0, 29, -12, 10, -31, 1, 6, 7, -14, -20, -5, -25, 16, -14, -16, 8, -33, 27, -7, -37, 0, 14, -6, -9, -29, -12, 17, 18, -29, -49, -6, -55, 5, 12, 19, 10, -14, -3, 18, 1, -2, -4, -8, 8, -8, -23, 20, -9, 58, -6, 29, -4, -6, 2, 14, 73, 9, 5, -14, 32, 5, -12, 8, 3, 43, 50, -11, 1, -33, -8, -14, -2, 36, 15, 8, -35, -9, -4, -17, -22, -12, -15, 7, 0, -25, 14, -25, 13, -7, -23, -23, -38, 20, 16, 1, 14, 29, -5, 1, 1, -7, -7, 0, -8, -10, -16, 15, 12, 8, -44, -2, -21, -32, 12, -6, 5, 21, 21, -22, -6, 11, -12, -3, 8, 10, 3, -68, 59, 11, -2, 35, 28, -4, 1, -2, -8, -12, 25, 10, 10, -2, 6, -7, -2, 12, -6, 11, 12, -12, -9, 29, 0, 24, 6, 24, 40, -68, 26, 41, 3, -1, 0, -25, 0, -12, -89, -21, 48, -54, -16, -2, 22, -16, -11, -12, -39, -17, -27, 1, -31, 5, 32, 14, 4, -4, -12, 41, -98, 22, -36, -2, 5, 10, -53, -28, -5, 8, 0, 32, 11, 2, 18, -10, -62, 28, -6, 7, -4, 17, -40, 12, 12, 13, -12, 31, -8, 0, -70, -8, 3, -28, 10, -1, 0, 8, -15, -14, -11, 0, 11, 13, 3, -25, 2, -3, -14, -2, 7, -9, -12, -9, -20, -10, 9, 13, 20, -8, 0, -1, -29, 7, -23, -22, 3, -39, 11, -31, -60, -51, -40, 31, 25, -17, 6, -11, 24, 2, 15, 6, -16, -8, -7, 9, -32, -16, -27, -7, -3, -2, -21, 16, -17, -14, 17, -23, -45, -6, 16, 2, -20, -51, -19, -28, -8, 43, -14, 3, -4, -3, -33, 0, -74, 10, 14, 8, 14, -1, -8, 7, -23, 4, -17, 10, -21, 13, 0, 11, 0, -8, 7, 17, 35, 0,
    -- layer=3 filter=0 channel=1
    18, 4, -1, -14, -3, -18, -12, 19, -12, 37, -11, 1, 23, 30, -21, 30, -11, 4, -2, -3, -16, 20, 13, 4, -1, -29, -18, 1, 6, -37, -3, -5, 6, 9, 6, 9, -5, 7, 54, 11, 25, -26, 3, -10, 19, -4, -12, -9, 24, -41, 14, 25, -1, -18, 5, -23, -13, 8, -4, -26, -10, 21, -5, 0, -16, -3, -55, 0, 6, 7, 13, -2, -3, 2, -13, -11, 12, 12, -5, 8, -12, -39, 0, 15, -10, 17, 8, -5, 14, 15, 3, -54, -11, -7, -24, -12, 14, 0, -12, -20, 9, 5, -34, -1, -37, -11, 10, -6, 19, 13, -71, 6, -5, 0, -37, 17, 7, -8, -11, -18, -9, 22, -20, 5, -10, -41, -21, 3, 5, 6, -9, -12, 8, -10, -8, 1, 10, 13, -9, -9, 2, -34, 11, 46, 1, -27, -5, -11, 39, 4, -7, -8, 5, -26, 6, 4, -2, 1, 19, 3, 4, 9, 14, 7, -10, 35, 15, -5, 0, -42, -23, 13, -49, -7, -24, 4, -9, 0, -16, -9, 11, 24, -12, -33, 0, -13, 0, -6, -18, 58, -10, 27, 38, -13, 17, -9, -7, 7, 4, 8, 5, -6, -48, -2, 0, -16, 32, -10, -1, 12, -18, -24, 49, 33, -16, -7, 4, 5, 17, 4, -8, 8, 39, -24, -15, -42, 25, -22, -7, -4, -7, 6, 57, 9, -10, 7, 22, -24, 18, -62, -19, -6, -10, -1, 54, -11, 24, -40, 11, -1, -4, -5, -21, -20, 7, -3, -6, -50, -16, 7, -9, -16, -6, -10, 1, -2, 0, 2, 10, -16, -17, 7, -28, 3, -8, -5, 36, 2, 3, -6, -1, 40, -7, -15, -9, -42, -23, 31, 4, 1, 14, 11, 2, -6, -13, -8, -16, 6, -23, 32, 6, 27, -19, -13, 8, -6, -12, -40, 44, -6, -7, -1, -5, 13, -3, -25, -14, -10, 8, -28, -16, 6, 1, -63, 0, -5, 8, -4, -11, 1, -4, -3, -16, 2, 12, -9, -32, -32, -4, 19, -3, -8, 11, 1, 21, 11, 12, -14, 11, -14, 13, -18, 0, -17, 8, -2, -6, 1, -31, -3, 0, -2, -9, -6, -30, 15, -19, 25, 15, -6, -6, -10, 0, 10, -25, 10, -13, -9, -8, 1, -5, -19, 1, 14, 10, -29, 6, -11, -9, 0, 13, 2, -5, -33, -11, -11, 2, -20, -40, -37, 8, 0, 0, -34, -31, 0, 47, 5, -3, 26, 12, 0, -2, -3, -12, 3, 2, -3, 26, 3, -4, -23, -11, -5, 9, -16, 24, 7, -33, 0, -9, 6, 3, -10, 15, -2, -2, 17, -31, 9, 6, 6, 8, -12, 14, 51, -14, 19, 28, -4, 5, -3, -7, 11, 7, 4, 25, 4, 0, 5, 40, 8, -38, -7, -51, 14, 12, -49, 34, -29, 13, 38, -21, -9, -16, -2, -27, -11, 24, 23, -8, 10, 23, 3, 2, -18, 2, 0, -35, 1, -39, 0, -12, 4, -38, -41, -40, -6, -7, -7, -40, 7, -10, 7, 11, -3, -19, -9, 2, -28, 1, -9, 26, -53, -3, 8, 2, -4, -16, -12, 32, -1, -7, -4, -20, 8, -13, 17, -43, -14, 43, 21, 13, 4, 21, -28, -25, -8, 14, -4, -6, 15, 6, 22, 8, 10, 4, -19, 5, 8, 13, 7, -36, -38, 5, -7, 9, -53, -18, 13, 22, -27, 8, -24, 38, -21, -6, 7, 29, 8, -4, 27, 0, 13, -1, -10, 7, -1, -2, 2, 7, -3, -10, 21, 8, 9, -10, -29, -17, 13, 5, 6, 33, -15, -1, -8, 10, -1, 3, 12, 14, 16, 36, 14, -4, -8, -4, -33, 10, -2, -7, 12, 16, 19, -21, -19, -40, -7, -4, 12, 0, 5, -35, 23, 0, -10, 14, 17, -25, 9, 22, 12, -23, -27, 0, 3, 13, -14, -41, 18, 5, 15, 17, 6, -12, 3, 22, -10, -31, -10, 2, -6, 0, 36, -1, -20, -12, 33, 0, 12, -16, 2, -27, 7, 12, -18, -9, -11, -9, -8, -35, 2, 31, 21, 20, 10, -8, 0, 6, 2, -9, 1, 10, -17, -1, -10, -48, -3, 8, 3, 6, -14, -4, -24, -2, -8, 12, 14, -12, -31, -11, 33, -12, -2, -9, -28, 16, 15, 13, 0, 7, 10, 29, 4, -49, 4, 34, -10, 21, 0, 24, -5, 10, -29, 3, 39, 20, 0, 2, -10, -15, 14, 35, -14, -21, 33, -5, -7, -28, -72, 1, -27, -8, -9, -15, 22, -14, -55, -23, -5, -36, -34, 7, 8, -4, 9, 3, -38, -11, -15, 11, -6, -13, -6, 18, 5, 8, 4, 36, -63, -12, 42, -12, 36, -13, 32, 31, 7, -8, 12, -81, -14, -15, 23, 22, -5, -13, -20, -4, -12, -1, 14, -9, -32, -5, 38, -5, -52, -46, -18, 3, 3, -12, 10, 3, 0, -34, 49, -19, 15, 17, -3, 19, -5, -7, 10, 10, -1, 37, 49, 15, 2, 3, -19, -4, 7, 13, -11, -9, -24, 3, 1, 12, 0, -33, 61, 27, -2, -69, -53, 9, 7, -4, 42, 10, 1, -9, -3, 27, -77, -11, -5, -1, -18, -13, -19, -1, 25, -25, 11, -9, -34, -20, 24, 1, -6, -78, 0, 7, -35, 3, 18, 11, -3, 35, -10, 16, 9, 45, -27, -25, 3, 24, -6, -2, -24, 6, 19, -2, -16, -14, -3, -12, 33, -5, 22, -1, -20, 30, -4, -4, -11, 3, 11, 16, 19, -7, 0, -7, -18, -32, -64, -8, -39, 14, -26, 20, -3, 4, 8, 12, -18, 1, 6, -13, 12, -51, -2, -9, -46, -3, -8, -22, -4, -3, 9, -10, -6, -34, -9, -1, 1, -21, -6, -33, 3, 11, 10, 10, 38, -52, 4, -19, -36, 0, -17, 11, -6, 7, 34, 25, -10, 32, 16, 7, 16, 9, -7, -3, -7, 40, -22, -15, 40, -13, -15, 14, 2, -19, 40, 7, 34, 20, 10, -13, 34, 16, 0, -38, 0, -36, 8, -11, 37, -27, -64, 12, 31, -2, 1, -4, 13, -30, 7, -31, 4, 18, -5, 32, 4, -1, 3, -2, 19, 46, -15, -15, 12, -1, -9, -17, 3, 28, -10, 8, 13, -14, 35, -12, 10, -20, 3, 7, -6, 0, 1, -34, -6, 50, -3, -15, 15, -18, 25, 33, -14, 41, 33, -20, 29, 5, -16, 0, -42, 0, -1, 4, -2, -12, 20, 10, -13, -13, 27, 17, 72, -31, -28, -6, -2, -7, -7, 11, 34, 5, -68, -26, 12, -16, 10, -64, -1, -9, 41, 35, 13, -11, -2, -20, 4, 39, 20, 1, 4, -83, 28, 1, 7, -22, -16, 5, 1, 5, -9, -36, -7, -1, 10, -1, -22, -12, -29, -20, 5, 47, 2, 12, -41, 39, 0, 2, -3, -61, -2, -53, 11, 20, -18, 36, -3, 38, -10, 2, 14, 33, -47, -24, 2, -15, -26, 25, -84, -2, 0, 2, 9, 0, -18, 0, -9, 0, 1, 9, -37, 6, -34, 0, 7, -3, 0, -1, 20, -16, 6, -8, 15, -42, -33, 12, -17, 27, 13, -20, 9, 0, 3, -1, -4, -9, 12, -10, -7, -49, 5, -3, -99, -9, 17, -11, -29, -1, 12, -6, 28, 9, 4, 38, 8, -24, 11, 0, -12, 20, 14, 7, 44, -63, 26, -30, -27, 13, 2, 49, -87, -17, -22, -2, 0, 9, 18, -2, 8, 19, -6, -14, -4, -20, -13, -57, 40, 11, -16, -17, -7, -24, 30, 12, 15, -45, 33, -10, -1, 2, 4, -36, 7, -38, -24, 4, -20, 34, -49, 4, -2, -11, 1, -27, 7, -13, -3, -16, 48, 0, -2, 3, -11, -9, -4, -40, 34, -8, 7, 25, 1, -4, -6, 15, -49, 27, 1, 9, 13, 6, 11, 3, -36, 0, -17, -13, 2, 5, 3, 24, -7, 31, -20, -15, -4, -36, 8, -16, -11, 26, 26, -44, -17, 0, -27, 9, -44, 1, -8, -3, 1, 1, 20, -11, 7, -6, 25, 1, -8, -5, -16, 36, 9, 0, -7, -10, -40, 10, -27, 19, -16, -4, -51, -38, 14, -9, 30, -27, -23, 4, -14, -4, -10, -16, -11, 3, -1, -58, -31, 2, 7, -34, -34, 0, 38, -10, -9, -27, -64, 5, 2, -8, 8, 9, 8, -14, 61, -53, -18, -3, 4, 1, 14, -9, 16, -23, -15, -35, 2, -46, 0, 24, -6, 14, -7, -10, 46, 48, -54, -8, -1, -5, 12, -33, -12, 28, 15, 27, -96, -18, 0, 0, -22, -10, 6, 0, -32, 7, -26, 4, -8, 37, 9, 20, -22, 0, -2, -4, 3, -5, -10, -6, 35, -25, 9, -5, -2, -33, -1, -1, 13, -5, 12, -17, 2, -56, -5, 12, -27, 24, -5, 5, 5, -20, -3, 0, 38, -7, -3, 10, -6, 22, -9, -30, 3, 13, -10, 2, 14, -58, -17, -19, -20, -10, -56, 11, -49, -4, -4, 5, 1, -17, 11, 6, -7, 2, 3, 6, 9, 4, -6, -31, -28, -24, -9, 0, -2, 18, 11, -39, -4, -31, 22, -14, -80, 2, 4, -40, -5, -36, 21, -2, 19, -1, 59, 6, 0, -10, 11, -5, 29, -29, 1, -57, -24, -5, 18, 16, 6, -5, -21, 31, 38, -34, -32, -35, 36, -11, -10, 25, -24, 11, 10, 24, -24, -2, -10, 0, 19, 2, -13, -5, -57, 11, 1, -29, 27, 39, -3, -21, 15, -70, -71, 34, 0, -2, 31, -38, -13, -22, 54, 10, 20, -27, -15, 9, 1, -5, -6, 10, -9, -53, 38, 1, -13, -36, -7, -34, 3, -16, -1, -11, -6, 30, 6, -16, 24, -8, -7, 30, -4, -2, 15, -25, -63, -5, 3, 1, -2, 7, -13, 9, -12, 21, -4, -5, -6, -2, -9, -5, -34, -5, -1, -30, 15, 1, 6, -15, -27, -14, -7, 41, 3, -9, 25, -12, -29, -9, -17, -10, 0, -83, -22, 22, 7, -19, 15, 59, 4, 53, 3, -20, -28, -1, -22, 5, -5, -2, -19, 10, 22, 51, 59, -15, -5, -2, -1, 1, -6, 14, 17, 1, 43, -72, -28, 7, 9, 5, 11, -38, -83, 8, -7, -10, 1, -5, 0, 0, -23, 0, -25, 18, -10, 28, -13, -7, -25, 6, -8, -73, -1, -27, -2, -16, -10, -30, 14, -19, -4, 2, -5, 3, -28, -44, 10, 18, -1, -60, 0, -19, -8, -5, 12, 0, 17, 16, -1, -62, 44, 6, -3, -22, 41, 18, -23, -14, -33, -37, 22, -1, -2, -18, -12, -20, -11, 17, 7, 7, 42, 24, -6, -11, 0, 44, -6, -4, -24, -54, -4, -78, -74, -19, -14, -68, -2, 6, -6, 8, 6, -67, -33, 9, 1, 3, -2, 14, -49, -21, -24, 8, 21, -9, 12, -30, -12, 12, 3, -14, 0, 46, -25, -10, 0, -18, 3, -6, -60, 3, 1, 22, 21, 4, 24, -13, -48, 6, 12, -18, -13, -4, 0, 8, 31, -25, 6, -32, 1, -61, 11, 14, -14, 52, -30, 9, -1, 6, -39, 10, -24, -72, -12, 0, -8, -2, 13, 11, -3, -21, 29, -16, 41, -33, 0, 35, 29, -23, -5, -6, 21, 17, -5, -1, 46, 4, 45, -18, 8, -9, 25, -45, -80, -9, 12, -59, -4, -12, -13, 2, 3, -27, 26, -1, -14, -30, 10, 0, 8, 3, 12, 23, -37, -8, 4, -1, 1, 5, 21, 8, 16, 22, 14, -2, 16, 23, 43, 3, -14, -2, -9, -2, -88, -13, -14, 55, -14, 17, -1, 17, 0, 1, 19, -30, -13, 15, 17, 17, 16, 68, -9, 43, 8, -11, 0, 0, -24, 13, -26, 6, -13, -18, -11, 7, -8, -19, 7, 13, -20, 8, -7, 2, 16, -41, 15, 1, -20, 6, -66, -20, 25, 41, -7, -1, 68, 11, -6, 18, 1, -12, 15, -28, -77, -11, 9, 2, 3, -3, 2, 1, 24, -45, 11, 8, -3, -10, 6, -19, -12, 23, 8, 4, 1, -40, 16, 29, -16, 17, 28, 21, -13, 15, -14, -9, -38, 29, -18, 0, 12, -33, 10, 19, 8, 14, -10, 35, -29, -54, -5, 15, -11, 8, 42, 25, 26, -38, 45, -9, -24, -42, -12, 29, 1, 4, 22, -4, 34, 0, 6, 11, -13, 2, -11, 18, 9, 45, -7, -36, -54, -26, -5, -29, -7, -49, -6, -35, 13, 51, -25, 19, 0, 14, 0, 11, 21, 1, -7, 22, -21, 3, -2, -4, -25, 6, -7, -10, -7, 2, -20, -24, -2, 8, -34, -7, 4, -7, -16, -12, -5, 30, 19, 54, -21, -13, -51, -9, 4, -61, -23, -4, 3, 1, 13, 0, -6, -9, 45, -21, -20, 1, 24, -17, -7, -19, 6, -10, -28, -24, -40, -15, 29, -5, -5, -32, -9, 10, 10, -50, -37, -3, -34, -18, 2, -3, -12, 9, -1, -1, 34, -7, 6, 20, 18, -3, -42, -7, -9, 7, 13, 5, -21, -11, -64, -9, -6, 2, 14, -56, -60, 7, -3, 20, 27, -9, 3, -6, -13, -19, -19, 10, -15, 55, -4, 23, 1, -23, -1, 12, 15, -60, 5, -6, 24, -38, -1, 39, 2, 59, 46, -5, 2, 3, -21, 23, 15, -6, -34, -49, -35, 4, 0, -3, -7, 40, -26, -9, -3, -6, 23, 31, -55, 4, 6, -27, -40, 5, 0, 25, -2, -12, -35, 5, -1, 1, 13, 28, 3, 0, 21, 4, -12, -2, -27, 6, 8, -10, 42, -14, 12, -74, 4, -17, 4, -10, -7, 29, -9, 9, 20, 30, 4, -22, -7, 0, -4, 0, 7, 54, -29, 19, -44, -47, 7, 4, -2, -62, -2, 10, 19, 20, -5, 16, 29, -47, -4, -43, -9, 26, 26, 7, -18, -25, 18, -23, -25, -19, 12, 4, 1, -7, 65, 2, 33, 2, 42, -10, -28, -11, -4, 29, 7, -19, -3, -16, 13, 7, 12, 28, 12, -8, -9, 11, 23, 69, 11, 59, 4, 5, -3, -39, 41, -3, 0,
    -- layer=3 filter=0 channel=2
    -22, 14, -3, 11, -7, 35, -8, 0, 6, 3, 9, -1, 3, -6, -7, 14, -7, 14, -38, 22, -22, 4, -7, -25, 21, 36, 40, -21, -3, 23, 0, 15, -1, 14, -17, 0, -1, -5, 2, -23, -3, 2, 23, 19, 25, -24, -13, -4, 20, -3, -44, -13, -16, 10, 3, -17, 8, 8, -8, -23, 0, 11, 5, 17, 8, 5, -3, 8, -19, -10, -12, 8, 0, 7, -24, -12, -7, -11, -10, 1, -27, -20, 7, -31, -11, -4, -17, -37, -23, -43, 24, -27, -5, -10, -12, 0, -7, -2, 46, -3, 45, -28, -4, 4, 8, -10, -5, 6, -1, 0, 25, 3, -8, 5, 42, -20, 5, -43, -25, -25, 26, 27, -33, -12, 18, -10, 17, -1, -14, 19, 0, 3, -2, 6, -12, -5, -14, 14, 9, 7, 9, 18, -15, -4, -1, -22, -1, -42, -36, -1, 9, -2, -2, 10, -5, -3, -9, -5, -21, 0, 5, -7, -25, 42, -9, 17, 7, 13, -9, 10, -112, -4, -32, -4, -28, -14, -15, -9, 1, -7, 13, -40, 12, 10, -34, 8, -7, -12, -38, 25, 18, -12, 41, 9, -10, -30, 2, 6, 27, -9, -34, 1, -16, 6, -17, 6, -5, -7, -26, -5, -30, -19, 38, 11, 57, 13, -16, -17, -13, 10, 0, -15, 0, -13, -5, 22, 26, 23, -9, 26, -5, 5, 4, -34, -4, 40, 5, 31, -2, -35, -13, 3, 9, 8, 10, -3, 18, 18, 3, 25, 24, 5, 22, 10, -23, 11, -8, 13, 10, 13, 11, 8, -7, 0, -31, -40, 13, 0, 23, -8, -10, -9, 27, 9, -2, 14, 13, 3, -7, 1, 9, -19, -5, -10, -5, 2, 10, -7, -3, 9, -21, 0, -13, 14, -28, 6, -6, -38, 21, -17, 31, 5, -6, -2, -6, 8, -6, -10, -3, -6, 3, -21, -23, -5, 13, 1, 25, 7, 0, -37, -54, -6, -8, -41, -20, -9, 12, -15, 13, 10, -27, -41, 9, -37, -8, -6, -38, -7, 8, 42, 6, -12, 8, 20, 12, -34, -3, -14, -2, 1, -17, 27, 1, 7, 37, 13, -6, 5, 0, -23, 18, 23, -22, 9, -3, 14, -8, 28, 12, 7, -4, -24, 2, 10, -33, -3, -41, -7, 36, 11, -1, -6, -31, -30, -3, 49, -15, 6, 2, -3, -25, 6, -6, -29, 0, -6, -7, -7, -28, 5, 9, 45, -21, 10, -12, -7, -5, -6, 8, -39, -6, 8, 6, 10, 26, 7, 5, 4, 7, -20, 5, -5, 0, -4, 0, 31, 7, 2, 31, -8, 2, 5, 19, 0, 33, 7, -5, -8, 23, 5, -3, -24, 0, -20, 33, 18, -23, -7, 15, -24, 35, -15, -12, -13, -3, -5, 7, 9, 11, 0, -11, -4, 34, -19, 5, -10, 2, -18, 17, -13, 68, -26, -5, 12, -15, 7, -27, 8, 10, -24, 0, -17, -36, -18, 1, -6, -3, 1, 7, 0, 11, 23, -14, -21, 52, -16, -27, 10, -7, 5, 37, -37, 27, 5, -28, 26, -1, -4, 4, -24, 57, 6, 3, -24, 0, -12, -3, 20, -2, 1, 29, -22, -5, -18, 0, -23, -16, 26, 38, 8, -1, -12, 14, 9, 12, -20, 21, 26, 3, 0, 6, 2, 17, 0, -6, -2, -18, 33, -11, 0, 14, -13, -4, 7, -25, 15, -29, 1, -27, 5, -24, -11, -14, 5, 9, 22, 5, -57, -13, 5, -4, -32, -19, -21, -6, -18, 5, 13, 16, -13, -4, -6, 8, 3, -2, -9, -23, 6, -5, -8, 9, 8, -64, 48, 4, -12, 11, -15, -7, -17, 5, -33, -3, -4, 5, -7, -27, -24, 0, -13, 4, -8, 31, -29, -4, 17, 7, 5, -36, 6, -13, -6, -3, 6, 18, 12, 31, 7, 9, -29, -12, -55, 0, 37, -3, -4, -3, 0, -26, 16, -9, 26, 8, 32, 0, -1, -6, -1, -1, -10, 12, 8, 5, -4, -42, -18, -10, 16, 4, 14, -2, -10, -77, -5, -9, 1, -6, 4, 20, -11, 13, -15, -5, 18, 37, -4, -4, 6, 2, 6, -17, 14, -51, -31, 30, 6, -12, -4, 7, 0, -44, 6, 10, -3, 57, -26, 13, -23, -5, -18, -3, 53, -7, 2, 43, -55, 20, -11, 3, -11, -9, 0, 15, 8, 16, -12, 0, 62, 20, -9, -7, -5, -67, -12, 63, -31, 20, 13, -16, -27, -11, 7, -8, 8, -23, -2, 4, -6, 2, -3, 1, -15, 13, -3, -1, -69, 23, -25, 14, 34, 32, -20, 16, 0, 2, 6, -13, 23, 0, 21, -38, 0, 0, 0, 11, 11, 20, -19, -4, 10, 4, -58, 10, 29, -6, -10, 23, -33, -5, 2, 36, 35, 0, -25, -6, -6, -14, 42, 48, 6, -12, 16, -11, 11, 28, -1, 9, 16, 0, -30, 7, 0, -15, 14, 10, -2, -14, -39, -1, 0, -20, 27, 16, 12, -5, -7, -4, 19, -1, 3, -20, -25, 16, 34, 13, 4, 3, 16, 9, 36, -11, 6, -36, 0, -12, 21, -1, -15, 22, 38, -6, 2, 39, 26, -3, 26, -15, 9, -55, 27, -4, -36, -16, 24, 5, 39, -12, -23, -56, -17, -13, -2, 11, 25, -10, -12, 4, -7, -11, 9, -23, -10, -1, 0, -15, -1, 3, -27, 0, 5, 27, 0, -32, 13, 39, -26, -6, -25, -37, -9, 26, -9, 10, -15, 11, -33, -8, 10, -11, 11, -12, 5, -52, 10, 53, -11, -18, 10, 1, -22, 18, -6, 5, -3, 7, 12, -32, 0, -38, 8, 0, -2, 3, 0, -15, 2, 12, -6, -8, 28, -5, 15, -6, -17, 4, 0, 7, -43, 2, -7, 21, 9, -17, 1, 18, 2, -48, 9, -6, 6, 31, -44, 7, 19, 4, 0, -30, 31, 24, 28, 6, -52, 40, 35, 2, -4, 0, 4, 21, -12, -36, 3, 13, -7, 35, 9, 8, -7, -55, -48, -9, -17, -17, 5, 5, 5, -25, -3, 3, 5, -2, 6, 2, 13, -3, -2, -14, 31, 10, -2, -27, 10, 8, -32, 0, -10, -14, 34, -1, 5, 10, 0, 40, -42, -49, -8, -23, 17, -12, -3, 7, 42, 25, -7, 5, -19, 9, -31, 1, -12, -6, 9, 29, -21, -6, -2, -26, 39, 26, 97, -12, 17, 16, 28, -17, -15, 1, 22, -5, -59, -63, 50, -15, 22, 31, -39, 10, -2, -7, -1, 4, -2, -8, -44, -14, -16, 24, -7, 18, 15, -8, 5, 3, -22, 5, 6, -11, -14, -1, -29, 9, 0, 3, 0, -40, -33, 0, -30, -2, 8, 0, 8, -23, -4, 18, 31, -1, 10, 2, 25, 0, 13, -1, -7, -41, -24, -3, 9, 0, -28, 0, 18, 0, 10, -2, 16, 3, 8, 51, -17, 2, -15, -7, -13, -1, -42, -1, -15, -23, -1, -72, 8, -69, -6, -19, 20, 8, 0, -9, -2, -23, 44, -27, 12, -40, -39, -28, -11, 14, 14, -36, -42, -3, -1, -49, -44, -9, 7, -19, 5, 11, 22, -4, 10, -11, -16, 5, -29, 9, 53, -110, 11, -20, 8, -15, 8, 13, -38, 0, -5, 18, -8, 25, -10, -15, 29, 27, 14, -17, 4, 4, 12, -13, 0, -25, -1, 28, 13, -1, -7, 11, 3, 16, -5, 2, -11, 0, -26, 14, -15, 6, -2, 26, 0, 22, 27, -28, 3, 38, 44, -5, 6, 36, -3, -31, -35, 13, 6, 9, 69, -9, -4, 16, 2, 30, -36, -81, -13, 26, -6, -20, 36, -8, 9, -35, 0, -3, 6, -6, -8, -41, 16, 0, -10, -1, 0, -13, -8, 2, -4, -26, -38, 75, -4, -25, 8, 0, 11, 32, -10, 0, -10, -36, 8, -12, -14, -28, -2, 11, 1, -36, -2, 7, -2, -15, 18, -14, -17, -29, -36, 10, 2, 5, -13, -6, 61, -5, -2, 12, 5, 4, 14, -21, 6, 45, 28, 17, 13, -4, 15, 0, -37, -8, 8, -14, 3, 3, -5, -26, -12, 9, 0, -16, 6, -77, -29, 5, 0, 15, 5, -36, 10, -52, 5, -14, -26, 1, -7, -13, -6, 21, -22, 2, -5, 29, -11, 19, -22, -21, -16, 28, 23, -1, -13, 21, 38, -2, 9, -8, 10, -85, -13, 10, -27, -27, 7, 4, 74, 9, -53, 50, 11, -16, -5, -13, -34, -4, 2, 34, 19, 0, 15, -3, -26, -28, -17, -62, 0, -15, -27, 15, 15, -20, 4, -10, 4, 6, -27, 20, -6, -48, 45, 21, -6, -2, 17, -58, 20, 0, -19, 27, 5, -3, -9, 20, -14, 22, 21, -1, 8, -9, -17, -19, 15, -10, 42, -29, -38, -24, 10, 17, 6, -11, -7, 10, 3, 17, 0, -5, 4, -5, -7, -18, -39, -28, -13, -14, 0, -7, 0, -66, -9, 32, 5, -5, 6, -3, 12, 12, -10, 6, -23, 25, 25, 10, -59, -5, 49, 55, -6, 23, 13, -12, 16, -7, -45, -12, -13, -11, -15, -11, -47, -2, -15, 14, 22, 0, 7, 2, -9, 35, -39, -11, 0, 40, 37, 4, -4, -38, 2, 12, -15, 21, -18, 4, -43, -6, 9, -10, -28, 10, -13, 8, -45, 18, 3, 9, 10, 24, 15, 48, 8, -20, -3, 6, -37, 34, 5, 24, -8, -14, 4, 2, -12, 27, -14, -17, -32, -4, -39, -2, 45, 4, 11, -89, 5, 2, 4, 8, -45, -2, -50, -21, -3, 37, 16, 23, -6, -16, 38, 24, 16, 7, -73, 9, -27, 13, -40, -4, 1, -16, -8, 6, 12, 27, 11, 38, 55, 11, -4, -9, -1, -12, 7, -8, -20, -39, 15, 8, -32, -17, -30, 13, 7, -13, 6, 41, 8, 5, 18, 5, 10, 39, -3, -10, -4, 20, 10, 0, 2, 31, -1, -5, -9, -8, 0, 55, 0, 11, -45, 0, 32, -3, -31, -26, -4, 17, -39, -8, 3, 58, 40, -12, -5, 2, -12, -21, 20, -20, 15, -12, 5, -36, 6, 7, -6, -4, -5, 5, -6, -4, -10, 0, -34, -55, -61, 56, -33, -19, 0, 0, 16, 9, -24, 9, 4, 38, 35, -6, -16, -27, 13, 63, 59, -5, 7, 3, -27, 25, -28, -1, 21, 54, 15, -6, -8, -52, 9, 17, -12, 12, 11, 10, 3, -20, -9, 0, 3, 2, 12, -5, -7, 12, 2, -12, 38, 33, -3, 0, 5, 35, 7, -25, -8, 1, -14, -11, 7, -24, 28, -1, 20, -9, -9, -11, -13, -6, -9, 11, 17, 21, 15, -3, 6, -5, 0, 7, -50, 10, -22, -48, 35, 2, 0, 18, 6, -59, -23, -13, 45, 29, 18, 51, 16, 6, 10, 12, -33, -10, -24, 0, 17, 27, 0, 8, -24, -8, 3, -3, -8, -30, 8, -11, -1, 9, -15, -10, -5, -11, -8, -38, 29, -42, 35, 39, 9, -7, -7, -1, -1, -31, 6, -1, -5, 10, -1, -5, 9, -16, -34, -10, 12, -7, 2, -11, -27, 6, 46, 0, -6, 37, -13, -44, -13, -46, -3, -36, -30, -35, 26, 5, 28, 59, -21, 0, 11, -20, -9, -2, 12, -1, -12, 0, -23, 10, -39, -6, -49, -1, 1, -2, 16, -7, -7, -4, -10, -2, 1, 8, 2, -11, 23, 29, 18, -3, -12, 14, -1, -20, 41, -21, 3, 22, -35, -9, -8, -25, 24, 1, -3, 3, 0, 0, 28, 7, -39, -17, -12, -8, -25, 35, -22, -13, 25, -18, -3, 18, -26, -15, -9, 42, -24, -31, 62, -54, -33, -17, -8, -8, 8, -21, -26, -53, -21, 5, 0, -8, -13, 9, -44, -29, 50, -10, -20, -28, 6, 2, -27, 14, 19, 1, -6, -36, 22, 1, -10, 18, 13, -30, 8, -3, 7, 0, 31, 37, -8, 11, 27, -20, 13, 36, -1, 0, -6, -20, -9, 7, 5, -6, -12, -5, 1, -30, 20, -5, 25, 6, 26, -11, -5, 19, 0, 13, 10, 21, -7, 19, -8, -9, -4, 19, -3, -13, -57, 21, 31, -13, 12, -14, -12, -12, -15, 3, -20, -1, 8, -9, 6, 0, -12, -4, 0, -32, -9, -37, 16, -16, 36, -7, -10, 16, -4, -75, 11, 5, 34, 5, -49, 18, 27, 17, -1, -39, 0, -9, -1, 3, -7, -26, 30, -15, 15, -5, -10, -18, -11, -31, -28, 7, 34, 21, 5, 48, 9, -15, -10, 10, 44, -52, 49, -46, -28, 10, 4, -22, 27, 0, -22, -31, -24, 7, 7, 5, 24, -7, -22, -27, 2, 10, -7, 17, -34, -50, 50, -13, 21, -7, 25, -8, -12, -39, 46, 4, 1, -22, 9, 4, -16, 41, -32, -6, -8, -11, -3, -13, 10, -15, -3, 22, 14, -34, -16, 8, -27, 6, -17, 0, 15, -9, 15, 15, 38, -11, -4, -11, 0, 7, -26, 3, 11, 8, 39, -12, -8, 16, 31, -6, -9, 22, -48, 4, 0, 32, 43, -18, -15, -11, 9, 3, 4, 0, 5, 2, -32, 1, -13, -42, -46, 22, -16, -6, 16, -14, -15, -13, 4, 22, -8, -3, 44, 4, -9, -19, -21, -38, -7, 27, -10, 24, -38, 2, -12, 4, 9, -21, -60, -40, 25, -49, 7, 28, 7, -2, 7, 24, 13, -5, 5, 42, 2, 0, -10, 9, -5, -24, 19, -12, -4, 7, -6, -10, -6, 5, -23, 0, 1, 14, 0, 0, -10, -7, -10, 12, 1, -14, 10, -37, -2, 22, 29, -2, 15, -9, -15, 1, -8, -21, -51, -8, -13, 17, 1, 38, 3, -1, 5, -15, 10, 10, -10, 7, -36, 17, -9, -11, 14, -14, -10, 5, 15, 13, -9, 35, -29, -12, 0, -35, -6, -24, -70, 13, -4, 7, -29, -36, 0, 19, 3, -47, 14, -6, 22, -8, 2, 11, 42, 30, -3, 10, -17, -4, -39, -12, -4, 6, 28, 8, 38, -11, -3, -39, 5, -11, -23, -1, 2, 28, -6, 32, -10, 3, 10, 25, 4, -12, 30, -56, 28, -5, 6, 22, 2, 36, 7,
    -- layer=3 filter=0 channel=3
    11, -5, 11, -32, -4, -25, 1, 9, -5, 27, 14, -7, -25, 29, 14, -14, 26, -6, 44, -40, 18, -2, -21, 0, 30, -9, -12, 9, 2, 35, 5, -1, 1, 0, 10, 7, -9, -18, 6, -15, -67, -51, -3, 12, -22, -2, 5, 10, -5, -30, 28, 10, -30, 4, 8, 1, 32, -1, 10, 13, -27, -4, -9, -18, -36, -9, -11, 4, -13, 1, -7, 5, 11, 1, -17, 14, -6, 9, 2, 12, 14, 4, -1, 0, 3, -13, 8, -13, 35, -6, 4, -39, 5, -13, 12, 2, -15, -5, 6, 9, 23, 10, -2, 0, -23, 16, -38, -14, -8, 0, 2, 20, -13, 3, -13, 23, -21, 38, 3, -19, 17, -13, -4, -7, -4, -19, 14, -18, 0, 4, -40, -29, -7, -3, -5, -1, -6, -8, 9, -9, -12, -36, -2, -3, -12, 17, -25, 16, -39, 0, -40, 6, 11, -34, 2, 7, 7, 3, 2, -5, -51, 12, 1, -31, 3, 5, -20, -22, -1, 7, 26, -10, -9, -2, -10, 6, 13, 11, 29, 2, 10, 20, -35, -8, 33, -37, -4, 8, 6, -27, 20, -1, 23, -21, 9, 19, 6, -25, 35, 0, 16, -9, -25, 0, 23, 5, 5, -11, 26, 2, -40, -6, -37, 16, -49, 17, 15, -17, 45, -4, 22, 5, -7, -18, -12, -37, 39, 5, 3, -10, 9, -13, 14, 0, 3, 28, -2, -7, 7, 4, 20, -10, 5, -1, 0, 1, 26, -24, -55, -20, -1, -1, -22, 15, 0, 3, 11, 41, -14, -6, -10, 38, -19, 52, 23, 8, -5, 3, -19, 30, -2, -18, 15, -24, 17, 38, -43, -29, 16, 11, -3, 5, -18, 7, -3, -24, 23, -3, 10, -2, 5, 10, -6, -9, 42, 5, -27, -12, 20, 5, -51, -4, 14, 0, 4, 19, 43, 22, 20, 2, -8, -4, -2, -6, 13, -3, -3, 19, 8, 5, 32, -3, -18, 21, 24, 5, -4, -10, -9, 8, 3, 41, -14, 9, 3, 9, -25, -16, 4, -8, 11, -8, 6, -29, 29, 18, 2, 12, -7, -29, -20, 7, 18, -7, 23, -31, 2, 0, 6, -2, -25, -9, 20, -2, -9, -5, -1, 0, -11, 2, -11, 29, 8, 19, -7, -29, 52, 0, -1, 3, -13, 7, 3, -14, -10, 34, 9, -65, -7, -8, -29, 4, -12, 8, -4, 0, 3, 21, 17, -2, 2, 2, -3, 8, 20, 0, -19, 0, 0, -17, 4, 7, 14, 6, 14, 19, 9, -15, -27, -30, -5, 5, 2, 1, -14, 7, -46, 16, -10, 3, 39, -6, 31, 4, -9, -6, -5, 24, 19, 1, 21, 0, 3, -7, 0, -13, 19, 29, -11, 11, -26, 8, -8, 1, -28, -1, -25, 23, -19, 0, 3, 8, 3, 0, -11, 0, -21, 4, 35, 12, -31, 2, 25, 6, -17, 4, -9, 4, 8, 4, 1, -29, -43, -13, 6, 7, 10, 0, 6, -26, -1, 5, 11, -16, 24, -30, 19, 11, 19, -5, -25, -22, -17, -23, -50, -50, -34, 8, 17, 15, -23, 9, -16, 9, 5, -43, -16, 7, -22, 11, -44, 10, -2, 3, 10, 14, 3, 20, -15, -12, -13, -55, -11, -5, -22, 5, 0, -34, -13, 16, -3, 2, 6, -34, 2, 1, -18, 3, 1, -6, 36, 30, -48, 2, 30, -8, 61, 8, 9, -5, -9, -33, 14, -59, 9, 5, 4, 42, -1, 5, 0, 0, -11, -6, 12, 1, 11, 5, -79, 36, 7, -7, -21, -11, 6, 9, -13, 19, -14, -34, 3, -12, -40, -17, -4, 39, -9, -9, 9, 8, 36, -11, -2, 7, -7, -25, -13, 2, 0, 3, 19, -8, -31, 17, 19, -3, -32, 2, 14, -12, 7, -2, -38, -15, 11, 1, -36, 22, -37, 39, 12, -16, -43, -7, 47, 1, 17, -57, -26, 13, 6, 60, -10, -12, -1, -1, -16, -13, 9, -16, -3, 0, -4, -8, 22, 25, -10, 38, 6, -1, -21, -8, 21, 8, 19, -2, 6, -3, 42, 10, 9, -15, 10, 35, -60, -43, -4, 8, -4, 0, -24, -15, 30, -7, -16, 0, 6, 0, -36, 9, -15, 4, -3, 0, -39, -6, -7, -19, 0, -2, -20, -61, -32, 29, -11, 14, -49, -16, 7, -7, 0, 0, -33, -28, -11, -21, 0, -49, -7, -13, 0, 12, 53, -13, -18, 4, 3, 7, -9, 12, 18, 7, -8, -2, 31, -22, 9, -1, 16, -19, 8, 58, -3, 8, 10, -11, 4, 37, 2, 12, 0, 6, -13, 1, -22, -9, 29, -16, 26, 34, -27, -3, -6, -1, -13, -9, 0, 0, 13, -9, -3, -23, 7, -5, -4, -2, -1, 15, -6, 11, -3, -5, -38, -29, 2, -9, 28, 12, -43, -19, -61, -6, 6, -34, 0, -13, 0, -11, 13, 10, -10, -7, -5, -8, -5, -4, -3, 26, -27, -46, 3, -30, 5, 8, -1, 18, 9, -2, -35, -14, -5, -7, -17, -26, 12, 0, 4, -28, 43, 0, 2, -17, 17, 10, -52, -10, -7, -3, 31, 7, 6, -12, 1, -7, 6, 17, -9, -13, 9, 6, -7, 11, -5, -16, -4, 23, 0, 1, -5, -36, 7, -11, 3, -9, -18, -13, 20, -4, -24, 10, -26, 14, 16, 6, 33, 0, 8, 12, -2, 3, -7, 5, -28, -9, -12, -33, -11, -7, -23, -4, -6, 7, -8, 23, -46, -51, -12, -3, -27, 37, 4, -4, 20, -3, 21, 23, -5, 1, 4, 6, -27, 10, 1, 11, -11, -13, 2, 5, -16, 12, -5, -20, 8, 7, 21, -1, 10, -4, 10, -2, -26, 20, -4, -9, -6, -6, -9, -20, 5, 4, 3, -2, -12, 3, -10, 6, -6, 4, -5, -4, -63, 4, 16, -26, 0, -29, -74, 6, 40, 5, 38, -7, -1, -19, -10, -2, 2, -2, 2, 25, 16, -1, 16, -31, -8, -17, -21, 5, 13, -85, -10, 15, -10, -8, -20, 8, -27, -7, -4, -10, 15, 14, -12, -43, -4, -27, -14, -29, -11, 9, -19, -2, -9, 12, -3, 16, 24, -9, -5, -7, 10, 2, 20, -10, 35, -12, 16, 7, -21, -8, 18, 1, 24, 13, -55, 39, -4, 37, 0, 31, -3, -15, 18, -8, -11, -3, 17, -19, -17, -76, -7, -18, 17, -10, 21, 10, -24, -34, 17, -2, 15, -26, -2, 2, 25, 22, 7, -7, 6, 6, 8, -8, -9, -46, -10, -34, -31, -33, 24, -30, -2, 5, 22, -38, -33, 17, 33, -20, 0, -49, -7, -13, 7, -7, -3, 19, 11, 8, 23, -10, 5, 43, -8, -15, 0, -30, 3, -8, -13, -5, -9, -37, -4, -3, -31, 4, -5, -22, -7, -2, -7, -9, -31, -4, 15, -40, -7, -19, -34, -72, 2, -6, -1, -5, -17, -1, -59, 10, 9, 24, 10, -5, 45, 26, 35, 35, 31, -6, -3, 7, -28, -23, 0, 7, -11, 36, 10, -7, -15, -27, 18, -4, 6, 27, 10, 28, -7, -16, 3, -9, -9, 8, -12, -12, 6, -24, 15, -3, 4, -21, 15, -17, 16, -12, 12, 5, -7, 35, 9, 2, -2, -5, 58, 11, 29, -11, -25, -5, 10, -8, 7, 0, 0, -10, -38, 0, -48, -8, 41, -8, 18, -10, -5, 11, -2, -27, 35, -27, 31, 16, -1, -4, -38, 36, -13, -8, -9, -19, 31, -14, -4, 10, -8, 0, 0, -38, 9, -16, 14, 45, -7, 0, 18, -8, -5, -67, 9, 15, 7, -15, 10, -9, -25, -8, 27, 0, 5, -18, -5, -20, -2, -8, -11, -9, 2, -9, -1, -19, 4, 1, 16, 18, -2, 15, 20, 8, -5, -7, 6, -16, 24, 15, 5, -22, -4, -4, -15, 20, -66, 0, -56, -1, 11, 16, -2, 34, -14, -16, -4, 19, 4, -3, 14, -6, -17, 29, -6, -4, 20, -22, -15, 0, -65, -23, 14, -4, -3, 14, -1, 31, -4, 19, 6, 10, -3, -2, -12, 0, 10, 14, -26, -8, 30, -13, 29, 4, -6, -3, 0, -50, -23, 33, 0, 34, 8, 7, -1, -7, 7, -18, -9, 16, -6, 3, 0, 13, -12, -16, 1, -18, 5, 5, -14, 0, 28, -7, 0, -23, -2, 14, -26, 7, -1, -34, 3, 15, 3, 2, -11, 27, 10, 22, 10, 5, -22, 7, 3, 0, -37, -28, -19, -22, -2, 33, 6, 14, 24, 3, 12, 3, -9, 6, 4, -2, 1, -45, -30, 22, -11, -15, -32, -12, -20, 3, 2, 0, 68, 11, 7, 11, -17, -2, -8, 1, -32, -7, -53, 0, -10, 8, 6, 7, 24, 5, -10, -21, -23, -10, 6, 9, -12, -9, -9, -24, -9, -2, 39, 0, 19, 18, 6, 43, -19, 17, 3, -6, 9, -6, 2, -20, 33, -11, -16, -6, -10, 9, -5, -5, -24, -2, 5, -28, -30, -7, -29, 17, 2, -17, -10, 32, -16, -2, 0, -34, 10, 25, -6, -11, -2, 2, -24, -28, 44, -2, 6, 45, -2, 7, 4, 4, -62, -30, 9, -4, -5, -35, -27, -6, 10, 10, 11, -8, -16, 1, -16, 13, 3, 1, 1, 5, 5, -2, -2, -22, 30, 12, 16, 5, 0, 28, -36, 2, -22, 0, 47, 30, -7, -7, 12, -29, -23, 9, -21, -8, -36, -11, -30, -22, -10, -11, -2, -4, 14, -38, 73, -14, 3, 10, -55, 13, -16, 42, -8, -9, 30, 3, -1, 1, 25, -41, 1, -28, -20, -8, 0, 3, 22, 8, 0, -4, -14, -14, -5, -7, -34, -32, -15, -31, 12, 9, 38, 6, 1, -10, 0, 12, -46, -13, -7, 3, 0, -10, -13, -1, 0, 11, -6, -11, -5, -40, 2, 6, -33, -26, -10, -15, 1, 8, -5, 6, 22, -23, 17, 31, 1, 0, -42, 22, -5, -3, -1, 7, 0, 36, 23, -4, 3, 21, -14, 2, -8, 7, -1, -18, 10, 0, 15, 9, 3, -2, 40, 0, 13, -3, 19, 40, -16, -2, 12, 10, 37, 10, 16, -12, 12, 3, -56, -24, -27, -5, -4, -15, 3, -59, -10, -14, -22, -29, 11, 13, -12, -12, 28, 41, -16, -6, 0, 19, 0, 0, -9, 31, -15, 17, -14, 4, -24, -3, 4, 8, -7, -2, 11, -11, 7, 0, -17, 1, -25, -22, -6, 4, 6, -14, -5, 27, -7, 11, 29, -4, -7, 0, 30, -12, -27, 8, -5, 36, -30, -48, 2, -15, -7, 8, -29, 5, 8, -2, -30, -22, -4, -7, -9, -13, 6, -8, -23, 19, -17, 17, 21, -27, 11, 0, 32, -3, 8, -16, 9, -17, 11, 17, 5, -1, 20, 3, 28, -2, 7, 14, -18, 21, -19, -43, -9, -21, -6, 0, -11, 1, 15, -13, -2, 12, 17, 11, 20, -6, -22, -10, 14, -1, 10, 34, -36, 21, -9, 5, -2, 31, 15, 3, 39, -3, -14, -23, 0, 2, -5, -4, -11, 15, 0, -4, 16, 7, -10, -77, -15, -1, 7, 30, 24, -6, 29, -5, 3, -10, -46, -5, -2, 18, 4, 9, 2, -11, 31, -19, 0, 0, 9, 6, -33, 1, 6, -25, 33, 28, 3, 10, -25, 12, -31, 2, 9, -30, 3, -17, 4, -10, -5, -29, -9, 21, 12, -34, 1, -5, 7, -11, 2, -2, -10, 8, -11, 0, 31, 8, -5, -2, 0, -11, -7, -4, -11, 7, -6, 34, 1, 24, -19, 16, 43, -27, -6, 0, -14, -19, -2, 16, -9, -14, 9, 14, -26, 8, -15, 9, -17, -14, -5, -13, -69, 9, 39, 0, 12, -32, 15, 0, -42, -4, 38, 9, -106, 14, -6, 24, -26, -4, -5, 7, 43, -28, 3, 11, 28, -9, -36, 5, 0, 9, -3, -17, -6, 7, 1, -8, 2, -9, -8, -2, 8, -4, 11, -4, 14, -8, -10, 0, 26, -1, 24, -37, 22, -21, 2, 5, 4, -7, -16, -40, 28, -22, 3, -1, 10, 2, 16, -14, -1, -4, 3, -8, -22, -20, -18, -13, -13, 22, -1, 42, -33, 22, -29, 44, -28, 30, 7, 10, -1, -7, 32, -59, 9, 9, 8, -35, -8, -17, 0, 2, -16, -20, 6, -19, 21, 27, -14, 14, 7, 9, 18, 2, 15, -3, 10, -15, 20, -17, -11, -4, -4, -14, 29, 0, -5, -13, -6, -21, -38, 20, 0, 5, -23, -5, -23, 32, -11, 34, -32, -10, -23, 9, 2, 11, -24, 7, -16, 13, 6, -2, 3, -9, -26, 4, -24, 3, 4, -12, -39, 7, 43, 20, -9, -6, 13, -20, 11, -11, -15, 1, 0, -42, 35, 20, -12, 0, 0, 0, -8, 3, 21, -5, 0, -1, 3, -8, -20, 17, 34, 10, 4, 6, 24, -8, 2, 5, -8, -3, -22, -25, -2, -11, -22, 6, 5, 0, -11, 20, 9, -1, 23, 0, -10, -18, 0, -3, 11, 35, -9, 5, -36, -8, 9, 0, 1, -7, 17, -16, -4, -26, 17, 27, 2, 5, -2, -10, 8, 23, -9, 25, -5, 36, 1, -14, 15, 8, 12, -15, -29, -36, -36, 8, -44, -8, 38, -13, -31, 4, 9, -11, -7, -17, 17, -33, 18, -25, -4, -15, -14, -5, 8, -36, 0, -13, 7, -6, -13, 10, 8, -9, -9, 4, -3, 31, -3, 14, -19, 0, 4, -7, 12, 32, -20, 32, -49, 9, 25, 12, 3, 19, -7, -7, -25, 13, -15, 13, -11, -13, -33, 4, -6, -17, 14, 3, 14, -8, 6, 8, -14, 1, -27, 8, 9, 10, -11, 12, 11, -31, -55, 9, 9, -7, -4, 27, -20, -2, -53, 21, 36, -30, 21, -27, 2, -9, -5, 2, 23, -59, 15, -16, -6, 43, 39, -8, -2, -11, -45, -10, -6, -11, 28, -4, -49, 5, -11, -4, -15, 6, 8, -4, -2, -19, 1, -25, 10, -4, -1, 6, 0, 12, 17, 16, 3, -11, -6, 10, -33, 4, -16, 4, 5, -35, -11, 4, 6, 13, -3, -8, -13, 1, -14, -4,
    -- layer=3 filter=0 channel=4
    1, -39, -8, 1, -4, 31, 4, -30, -59, -2, -3, -2, 7, -15, 3, 27, -14, -1, -1, 28, 31, -15, 17, -6, -8, 4, -10, 11, -2, -32, 15, 14, 7, -6, 3, -7, -5, -13, -16, 12, 3, 26, -11, -27, 0, 2, 1, 3, 2, -20, 7, 12, 9, 23, 4, -14, -32, -15, 7, 12, 38, -26, -5, 6, 23, -10, 39, 15, -6, -13, 6, -5, 7, -7, -1, -8, -6, -35, 0, -13, -69, 0, -1, -23, 10, -35, -6, 36, -54, 46, -39, 14, 0, -5, -11, -38, 18, -5, -39, -13, -30, -15, 17, -14, 28, -22, 11, -6, 38, 29, 12, -13, -1, 0, 5, -37, -32, -26, 22, -17, 16, 11, -13, 11, -7, -6, 23, -40, 3, 1, -12, -31, -11, -12, -21, -7, -7, 1, 2, -2, -10, 7, -10, 35, -3, -59, -19, -13, -11, 6, 47, 3, -17, 9, -6, -4, 24, 6, 17, 11, 31, 5, 31, 26, -2, -20, -12, 9, 1, -39, -41, 1, 42, 10, -37, -5, -43, -12, -3, 4, -4, 14, 10, -15, -13, -43, 5, -7, 33, 37, 5, 1, -90, 22, -9, 50, -12, 1, 5, 7, -11, -35, 6, -2, -12, 16, -38, -18, -4, -6, 11, 6, 4, -15, 13, -14, 11, -39, 7, 10, -8, 3, -48, -8, 7, -18, 7, 44, -8, 6, 0, 1, -54, -18, 34, -2, 7, -3, -76, 15, -9, 8, -1, -12, -10, 5, 12, -27, -22, -1, -6, -14, 13, 48, 11, 7, -7, -37, 8, -12, 9, 26, -3, -6, 4, -4, 10, -13, -3, -8, 20, 19, -67, 0, -26, -9, -6, -22, 6, 16, 5, 22, 20, -32, 4, 22, -3, 3, 10, -3, -10, -35, 8, 4, 19, 1, 24, 11, -27, -13, -28, -11, -15, 6, -2, 66, -25, 43, 31, -7, 9, -63, -18, 6, -12, 14, -4, 14, 7, 45, -9, 8, -9, 35, -23, -15, 11, -29, -12, -13, 22, -63, -16, -5, 3, 6, -10, 22, 6, -44, 9, 2, 6, -12, -27, -5, -23, -11, -5, 7, 0, -47, 1, -9, -56, -3, 14, -21, 32, -14, 33, -16, -23, 4, 54, -44, 0, -30, -15, -11, -35, 11, -18, 2, 20, -31, -4, 41, 12, 2, -15, 27, 30, 25, -10, 3, -48, 5, 6, 10, -1, -1, 22, 9, 4, -5, -6, 21, -10, -8, 12, -35, -19, -15, -33, 7, -5, -1, -13, -20, 5, 0, -4, 3, 37, 1, -11, 27, -11, 18, 12, -22, -4, -13, -12, -23, -4, -11, -38, -1, -13, 2, 3, -1, -10, -3, -7, 4, -9, -34, 2, 3, -7, 37, -4, 24, 16, -1, -20, 20, -12, -52, -5, -1, -28, -3, 27, -16, 0, 12, 7, -42, 8, -10, -14, 2, -57, 16, 20, -12, -35, -7, 6, 2, -3, -6, -11, -8, 1, -19, -1, -11, 42, 32, -7, 13, 4, 5, -14, -38, 8, -7, 13, 0, -52, 18, 7, 7, -17, 1, 20, 9, 8, -42, 18, 12, 13, -5, 13, 0, -36, -17, -67, 37, -8, -40, 0, 40, -21, 32, 21, 7, 2, -14, 52, -55, 42, -55, -13, -11, -39, 21, 39, -11, -8, 34, 22, 24, -9, -60, -11, 1, -13, 33, -7, 5, 1, -1, 10, 2, -13, -2, 13, 11, 6, -33, -25, -1, -14, 5, 12, 22, -63, 6, 24, -24, 6, -14, -27, 10, -4, -4, 10, 15, -12, 15, -8, -10, 40, 7, 0, -8, 8, -19, 4, 9, 24, -51, 2, -7, 5, -6, 17, 11, 4, -14, 7, -10, -7, -8, -32, 20, -19, 5, -6, -17, 31, 4, 13, 7, -3, 6, -33, -32, -40, -22, 27, -7, 25, 7, 45, 30, -4, -13, -62, -13, -41, -5, -48, -21, -1, 1, 29, -12, -29, 7, 5, 8, 46, -13, -14, -40, 8, 1, 1, 1, -55, -7, 58, -4, -3, 5, 5, -19, 4, 39, 5, -74, 8, -32, -11, 8, -1, 7, -3, -23, -3, 3, -39, 10, 29, 2, 2, -8, -12, -5, 12, 1, -13, 5, -1, 21, -56, -17, -26, -11, 31, 2, -28, 0, 49, -6, 8, -47, 10, 15, -34, 11, 9, 38, -8, 18, -3, -18, 11, 17, 3, -39, 9, 2, -10, -8, 26, -22, 3, 7, -16, -37, -1, -8, -13, -5, -8, 3, -3, 45, 5, -43, 18, -1, 15, -6, -37, 12, 6, 33, 3, -33, 16, 2, 0, 14, 4, 5, -6, 5, -11, -32, -14, -7, -53, 43, -4, -2, 7, 3, 0, 42, 6, -23, -12, 52, 21, 5, 21, 7, -36, -3, -68, 20, -17, 38, -3, -2, -11, -25, 11, -13, 9, 4, -3, 30, 17, -15, -16, 0, -60, 4, 23, -5, 20, -58, -16, -10, 37, -19, 0, 25, 26, 41, -4, 3, 8, -28, -7, -7, 20, 21, 54, -28, -8, 11, -13, 14, -3, -4, -18, 0, 6, -4, -16, 9, -1, 4, -11, -10, 9, 35, 18, -1, 4, 17, -28, 7, 13, -20, 4, -3, -24, 16, 4, -6, -3, 34, -16, -1, -10, 8, -22, 14, -6, 0, -12, 1, -6, 4, -1, 53, -9, -7, -7, -2, -3, -10, 18, 0, -20, 3, 7, -11, 19, 4, -35, -4, -11, 5, -8, 33, -18, 5, -3, 6, 27, -21, -28, -18, -39, -33, -63, -18, -35, -3, 0, -41, -23, -18, 3, -18, 6, -22, 9, -7, 16, -7, -50, 4, 8, 8, -12, -2, 14, 3, -7, -18, 35, 45, 10, 0, 23, -11, -10, -3, 3, 4, 10, 14, -35, -5, 20, -5, 35, -1, 18, -13, 0, -6, -16, -6, -51, -12, 3, 9, 32, 14, -12, -8, -67, -3, -11, 4, -9, -33, -4, -30, 12, -3, 2, -4, -33, -63, -61, 71, 37, 3, -12, 1, -6, 8, 0, -14, 18, -7, 12, -63, 21, -9, 20, 4, -40, 45, 3, 5, -7, -9, 36, -23, -11, -8, -21, 8, 4, 40, 4, 10, 42, 8, 1, 18, -4, -13, -31, -46, -14, 25, -26, 38, -42, 21, 9, -7, 26, 4, -32, 28, -11, 2, -21, -8, -1, 9, 0, -15, -11, -7, -32, 1, -13, 1, 10, -14, 13, 7, -7, -9, 10, 3, 8, 9, 7, -27, 36, -2, 0, 34, -106, -8, 66, 21, 0, -69, 16, 72, -10, 3, 2, -14, 7, 7, -9, -4, -6, -9, 17, -43, -19, -48, 14, 6, -6, -15, -7, 7, -10, 12, 19, 4, -9, -37, 9, 40, 0, 11, 10, -19, -32, 0, -12, -1, -23, 0, -65, 0, 0, -7, -3, -17, 5, -15, 25, -6, -10, -68, -12, -10, -32, 11, -2, 5, -2, -12, -10, 2, 0, -5, -43, 19, -11, -15, -14, 13, 17, 1, 17, 9, 37, 24, -10, -2, 14, -9, 16, -10, -60, 4, -22, 13, -27, -1, -4, 21, -4, 7, -33, -10, -1, 19, 29, 0, 13, -12, -58, -27, 2, -22, -69, -54, -2, 5, -47, -5, 7, 0, -5, -2, -3, 18, 2, 12, 0, -12, 36, 24, 0, 9, 32, 14, -9, -64, -7, 6, 49, -6, -26, -6, -5, -47, 37, -8, 1, 8, -11, 1, 9, 27, -29, -8, -29, 5, 28, 0, -28, -8, -32, -10, 3, 8, -29, -11, 0, 32, -7, -5, 19, -4, -12, 5, -21, -11, -42, -24, 7, -15, -25, -1, -50, 35, 5, -1, 24, -37, 17, -5, 6, 1, 0, 98, 16, 11, -17, -41, -2, 30, 0, 9, -24, 6, 0, 20, -2, -6, -69, 37, 2, -23, 5, 9, 18, -4, 12, 6, -11, -31, -8, -83, 13, -13, 2, -12, 7, -10, 1, -57, 26, -40, -1, -11, -27, -59, -17, -2, 48, 38, -11, 6, -14, -6, 0, -14, 25, -19, 2, -15, 4, -2, -24, 25, 12, -19, 2, -9, 14, -5, 36, 12, 9, 23, -8, 18, 8, -11, 14, -4, -11, 10, -5, -15, 8, 0, 15, -34, 41, -9, -7, -3, -24, -42, -14, -7, -7, 15, -42, -6, -15, -13, -10, 31, 21, 12, 0, 11, 36, 18, 1, 15, -62, 0, -44, 12, -16, 3, -26, -21, -13, 2, -43, -13, 0, 16, 5, 3, -55, 4, -8, -2, 0, -4, -9, 7, 21, 6, 52, -3, -9, -27, -18, 26, 20, 7, 1, -20, 29, 10, -44, -18, 0, -11, -11, -5, -25, -17, 45, 21, -8, 9, 25, -25, 25, -8, -27, 2, 22, -29, -1, -7, 2, 0, 49, -20, 0, -7, 37, 22, -10, 6, 20, -3, 31, -8, 4, 9, -4, -3, -5, 9, 3, -64, 16, 24, 6, 5, 6, 0, 1, -6, 11, -10, 3, 10, -31, 9, -4, 0, -17, -26, 20, 22, 2, -6, 9, -15, -17, 4, -8, 3, 36, 0, -40, 9, -29, -2, 0, -24, -29, -32, -6, -32, -6, -25, -4, -1, -31, 0, 0, 25, 14, -42, -4, -6, 4, 0, -27, 16, -1, 5, -9, -47, 2, 12, 7, -13, -40, 48, 16, -11, -29, 27, 0, 23, 30, 10, 13, 5, 37, -9, 12, -12, -18, 32, -3, -22, -2, -4, 42, 20, -8, 26, 13, -40, 0, -8, 15, -7, -5, -17, -2, -26, 15, -38, 5, 47, -4, -9, -19, -7, 20, 8, -82, 0, -13, 35, 8, 11, 4, 19, -21, 19, -3, 4, 15, -38, -17, -11, -17, -14, -16, -46, -33, -9, 28, 5, -18, -9, -17, -16, -3, -2, 13, 3, -5, 0, 12, -4, -3, 4, 5, 42, 17, 14, 16, -20, 22, 0, -3, 11, -23, 13, -31, -3, 10, 1, 1, 33, 5, -1, 0, -44, -26, 21, 6, 7, 20, 8, 12, 39, 4, 14, -1, 24, 0, 3, -18, 17, -4, 35, -2, 0, 12, -13, -1, 37, 6, 21, 5, -37, -55, 73, -8, 11, -7, 6, -5, 35, -5, -3, -10, 19, -3, -5, -44, 2, -7, -10, -27, 2, -10, -24, -24, -9, 66, -6, 25, 23, 4, -16, 0, -17, -22, 17, -12, -6, 2, -2, -44, -19, -8, -4, 26, -21, 4, -3, -39, 0, -35, -8, 9, 0, 2, -1, 28, 9, 5, 2, 11, 3, -21, 6, 58, 8, 9, -21, 8, 1, 30, -1, -33, -3, 9, 26, -9, -32, 16, 26, -9, 16, 4, -1, -33, 2, -78, -1, 48, 5, 21, -11, 16, -3, 4, -43, -24, -3, 26, -20, -11, 26, 7, -11, -19, -56, -13, 21, -16, -22, -9, -7, 14, 0, -38, 37, -27, -6, -13, -66, -38, -1, 36, -1, -40, 2, 30, 1, -2, 4, -8, 35, -22, -5, 41, -10, 12, 19, -2, -22, 62, -1, -7, 15, -3, 2, -8, -12, 28, 19, 19, 19, -14, 42, 7, -1, 31, 7, 15, -60, -10, 24, 18, -17, -5, 5, 6, -10, 41, 2, -7, 8, -2, -23, 1, -26, 16, 2, -39, -1, -2, -2, 19, 13, 0, -47, 21, 1, 6, -48, -56, -2, -1, -37, 43, -22, 36, 0, -1, 21, 5, -21, 9, 3, 16, 28, 3, 7, 7, -44, -11, -36, 10, 66, 43, -19, -1, 3, -4, -14, 37, 19, -6, -27, 0, -39, 15, 4, 11, -9, -13, 16, 11, -20, -28, 8, -42, 2, 7, 1, 7, 6, 5, -6, -5, -26, -7, -16, 6, 6, -40, 30, -9, 35, -1, 0, 0, -12, 0, 26, 11, -26, -3, -10, -54, 0, 0, -5, 45, -11, 12, -19, -39, -1, -18, 0, -61, 3, -18, 26, -5, 8, -13, 7, -23, 19, -16, -50, 6, -58, 13, 64, 50, -7, 13, -35, -26, -47, -12, 8, -13, -30, 0, 2, -42, 0, -8, -36, -5, -2, 4, -12, 18, -10, -8, 19, 23, 7, -13, -8, -7, 6, 3, 4, 0, 3, -36, -9, 11, 7, -26, 62, 27, -4, 4, 34, -2, 9, -9, 18, 59, 3, -40, 8, 33, -1, -11, -9, 0, -5, 2, -107, -45, -35, 19, -43, 11, -40, -14, -18, 5, 2, -26, -56, -55, -6, 6, -18, 30, -10, -30, -26, -20, -2, 23, 18, 3, 0, -2, -4, 43, -11, 11, 18, -20, -46, -9, 47, 13, -12, 12, -3, 5, 14, 13, 1, 56, -42, -4, 44, -2, -8, -15, 4, 6, 31, 27, 8, -3, 0, 0, -3, -3, 8, -5, -27, 10, -1, -14, -62, -13, -7, 9, 16, -4, -1, -32, -17, -6, 17, -8, 44, 1, 11, -1, 3, -14, -19, 36, 0, -59, 7, -14, -13, -11, 17, -38, 12, 19, -10, 19, -26, -18, 16, 9, -14, 17, 17, 6, -1, -3, 5, -7, 3, -20, -15, 13, 12, -9, 30, 0, 22, 0, 10, 17, 32, 2, 9, 14, -5, 9, -12, 22, -9, 1, -65, 1, -10, -8, -3, -20, 4, -27, 40, -25, -4, 5, -21, 9, 9, -43, -18, 6, 4, -2, -10, -47, 2, -3, 23, -14, -12, 0, 11, -6, 57, -6, 39, -3, 20, -53, -13, 0, -13, 42, 17, -5, 24, 0, 21, 2, -20, -38, -6, -34, -26, -1, -1, 20, 7, 22, 3, 37, -7, -25, 3, 8, -16, 25, 0, 2, -32, 24, -15, -4, 38, 33, 26, -8, 9, 4, 0, -64, -13, -5, -13, -2, -28, -3, -12, -11, -21, 25, -9, 24, -4, 28, -3, 21, -1, 9, -2, -5, -5, -3, -15, 25, -12, -44, -61, 26, 33, -17, 15, 5, -19, -2, 0, 13, 8, 37, -10, 0, -9, 7, 5, 5, 19, -35, -1, 10, -6, -4, -36, 28, 2, -27, 1, 0, -15, -14, 35, 2, -11, 1, -14, -41, -2, 30, -2, -5, -7, 50, -2, 9, 3, -25, 0, -21, 8, -68, -6, 14, 0, -10, 1, 11, -14, -8, 28, -5, 1, 35, -38, -3, 5, -9, 0, 34, 40, 16, -5, 20, -10, -15, 17, 0, 9, -8, 7, 32, 25, -15, 24, -43, -17, -4, 1, 9, -2, 7, 0,
    -- layer=3 filter=0 channel=5
    -6, 30, 0, -28, -16, -13, -12, -17, -6, 1, -9, 7, -27, 43, 37, -65, 4, 13, 34, 2, 4, -9, -13, 18, 10, -15, -21, 3, 6, -28, 25, 8, 2, 1, -1, -11, -1, -1, -8, 57, -27, 13, -11, -16, -2, -37, 16, -7, -13, -22, 32, 6, 45, -53, -13, 2, -74, 10, -9, -4, -16, 38, 9, -3, 34, 0, 28, 21, -12, 11, 1, 34, -5, 3, -44, 39, -9, 6, -4, 13, -64, -13, -9, 33, 7, 22, -10, 14, 1, -20, 3, 32, 0, 31, -23, -2, -1, -8, -2, -6, -18, 3, 6, -21, -28, 8, -21, 5, -33, 11, -6, 4, 31, -3, -22, -18, -29, 7, 28, -36, -4, -6, -7, 0, 16, -28, -14, -2, 8, 21, -4, -11, 10, 9, 39, -7, 31, -7, -9, -9, -11, 32, -23, 25, -11, 46, -10, -23, -17, -9, -1, 0, -13, 12, -11, 0, 6, 3, -44, 14, -20, -23, -1, -57, -9, 33, 15, 4, 1, 12, 20, -11, -33, 0, -42, -3, 22, 4, -8, -11, -4, -22, 36, -19, -9, 17, -4, -17, -40, 15, -1, 33, 32, 1, -25, -11, 3, 7, -27, -1, -29, 7, 20, -7, 15, -19, 6, -8, -4, 5, 45, 23, -16, 4, 21, 4, -42, 30, -28, -9, 2, 4, 35, 43, 15, 45, -63, 18, -3, 24, 9, 10, 32, 8, -4, -1, -8, 17, 27, 2, 7, 6, -18, 9, -37, 2, 20, 0, 24, 8, -18, 12, 17, 28, -33, -3, -4, 17, -3, 3, 8, -29, -1, 1, 24, 29, -1, -5, 19, 37, 13, -23, 20, 0, 19, -17, -51, -30, 19, 22, -14, -56, 25, -22, 6, -32, -13, -31, -1, 1, -12, -10, 9, -12, 14, 3, -24, -5, 23, 13, -2, -16, -6, -2, 7, -11, 16, 25, -27, -18, 12, 12, -38, -10, 2, 4, 58, -3, 7, 18, -44, -3, 22, 29, -12, 0, -18, 15, -11, 10, -26, 45, -6, -15, 4, -4, -13, 7, -5, 34, -7, -10, 8, 31, 35, 16, 0, 56, -11, 9, -5, 25, 0, 3, 16, -20, -23, -4, -26, -7, -18, -3, -33, -6, -19, 41, 4, 19, -2, -2, 21, -32, 22, -2, 58, -46, -29, -66, 6, -6, 13, -3, 15, 0, 8, -9, 9, 15, 6, 3, -10, -9, 15, 22, 10, 12, 4, 20, -7, 30, 3, 12, -11, 42, 8, 1, 22, 4, 6, 7, 3, -4, 8, 12, -53, -1, -3, -21, 39, 11, 0, 26, 12, -8, 1, 19, -29, 2, -10, -7, -1, 7, -49, 5, 32, -10, -11, -28, -41, 5, -14, 11, -8, -4, -41, -49, -13, 35, 13, -10, 33, 35, -7, 8, 24, -1, -23, -24, 20, 0, 18, 36, -43, -20, 23, -4, -16, 26, -9, 27, -12, -12, -4, 30, 7, 9, 40, 4, 9, 15, 1, 30, -1, 53, -1, 12, 3, -10, -13, -9, 30, 19, 22, -17, 4, 11, -6, -7, 10, 11, 17, 6, 28, -17, -32, -20, 12, 4, -11, -54, -11, 0, 19, -21, -6, 23, 5, -34, 9, 23, -30, -10, -6, -4, -13, 13, 20, -18, 32, 7, 9, -26, -3, -21, -19, 0, -12, -9, 4, -23, -6, 30, -15, -9, -8, -3, -9, -24, 5, -12, 0, 6, 6, 32, 20, -12, -17, -83, 6, 9, 1, -18, 27, 35, -7, -4, 9, -36, -3, 12, -12, -4, 14, -17, 6, -3, 6, -2, 20, 4, -21, -5, 0, 10, -7, 3, 25, 7, -4, -27, 0, -8, -13, 12, -12, -13, 12, 35, -4, 2, 16, 13, 10, -24, -11, 15, 4, 16, -24, 2, 16, 0, 9, -45, -18, -7, -39, -3, -20, 1, 6, 28, -9, 46, -7, -5, 39, 29, 22, -30, 10, 40, 13, 27, -42, -7, -5, 30, -31, -51, 8, -12, -43, -48, 0, 7, -9, -5, -26, 27, 17, 3, -10, 2, 20, -15, 11, -1, -18, 18, -45, 8, 25, 0, 3, -2, 0, -13, -13, -10, -19, -10, -19, -28, 38, 15, 0, 16, 5, 14, -14, 0, -68, -4, 18, 5, 22, -9, 38, 3, 11, 1, -2, 32, -32, -36, 30, -5, 6, -66, -5, -40, -29, 6, 12, -17, -18, 26, 5, 9, 3, -8, -1, -23, -3, 21, 38, 32, 0, -3, 4, -10, 18, 30, 31, -14, -24, -16, 36, -27, 6, -5, -25, -4, -12, 37, -15, 34, -14, 33, -2, -11, 1, 3, -32, -36, 7, 16, -5, 19, 24, 22, -16, -2, 9, 6, 7, -38, 23, -3, -41, -51, -6, -8, 2, -9, 21, -5, -22, 8, -9, 3, -4, -4, -24, 0, -33, 1, 13, 0, 17, 3, 19, 6, -2, 3, 18, -40, -23, 16, 30, -27, 2, -5, -15, -12, 3, 19, -16, -15, 2, 11, 5, -10, -10, 7, 14, 22, 15, -3, 3, 13, -3, 16, 7, -3, -13, 6, -4, 0, 14, -58, -10, -26, 9, 6, 6, 18, -10, -20, 6, 12, 6, 3, 21, 45, 3, -2, 4, 0, 0, 8, -7, -47, 3, -40, 11, 11, -1, 6, -12, -9, -8, 8, 8, 24, 32, 6, 0, 19, 2, -27, -48, 14, 13, -11, 16, -21, 4, -22, -11, -11, 11, 0, -7, 4, 7, 8, -29, -9, 12, 2, 3, 21, -33, 20, 33, -67, -32, 28, -14, 12, 7, -29, -4, -21, -8, -8, 9, -67, -3, -5, -25, -3, -13, -65, -18, 13, -15, -15, 10, 18, 0, 20, -15, 8, -74, 3, -14, 0, -21, -11, 5, -6, 6, -8, -4, 6, -10, 26, -27, -19, 9, -18, 0, 4, -7, 0, 6, -2, -33, 1, -10, 1, 2, -9, -40, -12, -7, 62, 15, -16, -1, -2, -8, 2, -20, 19, -13, -7, 22, -5, -28, -33, 4, 5, -17, -3, 26, 45, -11, -13, -1, 18, 28, -23, 2, -13, 20, -2, -25, 1, 7, -18, 7, 1, -25, 4, 59, -2, 12, -4, -8, -37, 0, 14, -12, -2, 4, 3, -5, -28, -7, -15, 3, 22, 36, 8, 1, -8, -16, -4, 3, -26, 8, -33, 1, -17, 5, -13, -36, 24, -3, -8, -6, 8, -6, -29, 17, 22, 0, -8, -14, 19, 11, -9, 19, 38, 0, -34, 35, 5, -12, -9, 22, -14, -12, -18, 20, -9, -5, -15, 0, 0, 20, 5, 0, -6, -3, -34, -2, 15, 12, -12, -33, -37, -17, -15, 1, -4, 11, 11, -12, -14, 18, -31, 0, -36, -7, -47, 31, 7, -3, -15, -35, -28, 5, -16, -4, 4, -11, -17, -14, 5, -33, -5, 4, -1, 20, 21, 10, -22, 12, 8, -1, -28, 8, 5, -1, -42, -10, 3, 25, 16, -31, 15, 11, -15, -46, -44, 20, -23, -9, -18, 23, 6, 36, -19, 4, -15, 3, 4, 49, 9, -25, 17, -14, -2, -10, -42, -6, -30, 2, -48, 16, -12, -26, -10, -9, 6, 26, -1, -7, 4, -16, 22, -2, 2, 3, 0, -13, -7, 5, -6, -12, 0, 4, 11, 1, 34, -23, -21, 54, 12, -8, 1, 14, 12, -2, -9, -47, -5, -16, -20, 28, 0, 28, 7, -14, -2, -6, 9, -15, 10, -5, 2, -39, 7, -7, 3, -9, 4, 5, 2, 7, 1, -8, -14, -29, -35, 8, 18, -44, 3, -39, -25, 25, -26, -55, -8, -1, -14, -16, -7, 0, 17, -46, 8, -9, -32, 36, 0, -5, -1, -24, -23, 38, -10, -13, -2, -7, -11, 19, -5, -24, -1, 30, 0, -4, 16, 10, -22, -3, -65, 10, 8, -19, -11, -4, 3, 6, 35, 16, 24, -9, 0, -6, 7, -16, 24, 19, 20, -13, -8, -24, 9, -73, -18, 25, -1, -16, 10, 8, 3, 7, -14, -1, 0, -22, 1, -10, -8, -34, -8, 13, -37, 13, 9, -16, 8, 0, 8, 32, -12, 29, -63, 26, 0, 1, 19, -1, -9, 9, 7, -7, -18, 10, 0, 9, -6, 7, 13, 10, -16, 8, -10, 10, 2, -12, 13, 20, -9, -25, -13, 0, 10, 23, -3, 9, -2, -10, 9, -9, 3, 4, 5, -7, 20, -18, 9, -6, -38, -11, -10, 13, -1, 10, 20, -6, 3, 0, 10, 0, -7, -15, 30, 7, -8, 19, 3, -52, 20, -10, -11, -51, -6, -10, -20, 25, 15, 5, 19, 2, -17, -26, -9, 7, 10, 12, -52, -12, 29, 14, 10, -8, -2, -8, 9, -3, -42, 8, -15, 6, -5, -16, -26, -34, -40, -10, 35, -33, -5, -10, 0, -39, 9, -9, 4, -8, 4, -7, 0, 39, 8, -5, -23, -11, -24, -49, 1, 10, -1, 1, 25, 6, 5, 11, 9, -73, 2, -15, -15, 6, -43, 0, -14, 4, 2, -26, -39, -12, -3, 5, 0, 21, 5, 0, 2, -44, 3, -5, 25, -22, -27, -3, 26, 7, 3, -65, 10, -8, -9, -2, 11, -57, 26, 2, 2, 11, 5, -6, -33, -27, 0, 30, -19, 6, -23, -7, 0, -26, -33, 11, -9, 46, -19, 31, -14, 10, 0, -2, 3, 34, -24, 0, -16, -5, -37, 9, -4, 8, -5, -3, -11, 20, 11, 1, 13, 29, -6, -26, 11, 14, -4, 18, -7, 12, 33, -4, 16, 3, 9, 26, 25, -26, -8, -47, 13, -10, 9, 3, 36, -12, 2, 3, -6, -13, 3, -17, -1, 5, -19, -4, -6, 15, 23, -12, 0, -64, -12, 10, -4, -28, 15, -9, -6, 0, 14, 9, 14, 3, -1, -3, -1, -26, -5, 4, -43, -9, 23, -23, 70, -16, -3, 7, 47, 22, -11, 23, -33, -2, 18, -24, 0, 0, -42, -34, 29, -11, -4, -42, -5, -3, -45, -5, -18, 45, 23, 8, -6, 0, -5, -11, -2, 1, 11, 0, 2, 11, -7, 8, -13, -14, 28, -8, -40, 10, -40, -1, -13, -24, -13, 17, -14, -10, 10, -43, -17, -11, -10, -16, -1, 4, -3, -17, 20, 3, 11, -9, 3, 12, -5, -9, -22, 0, -17, -15, 12, -19, 9, 12, -11, -27, -10, -8, -21, 13, 2, 9, 14, 55, 14, -2, -16, 0, 9, -11, -38, -6, 2, -7, 10, 1, 6, -43, -12, 37, -1, -3, -17, 2, 8, 73, -10, -36, 2, -16, -14, -23, -43, -3, -8, 3, -2, 5, 17, -36, 1, 26, 0, -3, 6, -28, 8, 6, 5, 2, -26, -32, 8, 16, -23, 9, 0, -4, -25, -37, 24, 17, -7, -2, -14, 8, -1, 21, -5, 33, 34, 23, -2, 8, -4, 20, -8, 5, -5, -13, 6, -30, 2, 37, -33, -5, 6, -17, -2, 15, 8, 7, -9, 13, -47, -21, 1, -6, 8, -9, -10, 34, -1, 1, 15, -10, -1, -12, -1, 25, 1, 1, 6, -1, -42, 5, -16, -6, 6, -3, 11, -20, 21, -14, 6, -18, -4, 2, 54, -1, -2, -29, -58, 49, -13, 9, 9, -4, 7, -12, 0, -12, -1, -11, -8, 16, 0, -8, 21, -9, -21, -12, 3, 7, -29, 1, 34, 0, -9, -20, -8, -4, 2, -5, 0, -50, -15, 11, -7, -3, 29, 0, 7, -8, 23, 10, -36, -8, -71, 7, -5, -3, -6, 1, -53, -7, -9, 3, -42, 4, 0, 10, -7, 5, -6, -16, 24, 10, -13, -12, -30, -1, 31, 2, 1, -31, 17, -4, 17, 12, -4, 5, -15, -25, 4, -49, -24, -5, 3, -38, -55, 11, 1, -12, 3, -7, 25, 6, -2, 20, -14, 30, 4, 32, -42, -7, 5, -13, -6, 7, -9, 28, 28, 30, -19, -47, -67, 24, 2, 0, -39, -7, -31, -11, 5, -13, -17, -4, 4, -14, -9, -5, 10, -5, 4, 11, -33, 8, 9, -9, -2, -29, 22, -18, 10, -2, -6, -7, -5, -5, 1, -23, 1, 0, -8, 28, 9, -1, -38, -5, -15, 7, 3, -9, -7, -39, -4, -2, 2, -11, 4, 10, -7, -19, -7, 5, 23, -22, -22, -6, 35, 2, -25, -40, -16, 11, 12, -6, -34, 4, -50, -11, -8, 19, -11, 6, 20, -11, 0, -22, 4, 6, -13, 4, -6, -49, -6, -6, -1, 43, -10, -22, 5, 36, -8, -11, -11, -2, 14, 7, -4, -27, -53, -8, -55, 6, 8, -5, 46, 26, 14, -15, -1, -12, -11, -48, 4, -10, -19, -32, 14, 11, 14, 2, 27, -17, 0, 1, -1, 43, 7, 3, 5, 9, 16, 10, -36, -15, -16, 19, -55, 12, -18, -85, 5, -21, -27, -13, 16, 23, 9, 4, -18, -73, -11, -11, -11, 10, -20, 6, 27, -21, -4, 2, -4, 7, -27, 5, -6, -11, -20, -33, -5, 35, -6, 6, 49, -11, 12, -3, -11, -44, -17, -17, 11, 0, 21, 39, 10, 6, -49, -19, 19, 1, -58, -39, 9, 36, -46, -13, -2, -18, 0, -11, 5, 9, 12, -1, 3, -8, 11, -81, 24, 2, 1, 10, 11, -11, -37, 0, -1, -40, -2, -17, -17, -8, -33, 9, -15, -2, -7, 5, 25, 7, -11, 13, 15, 12, 3, 0, 34, -10, 6, -6, 6, -3, -13, 9, 0, -17, -29, 16, -1, -2, -10, -2, -2, -60, -27, -3, 11, -24, 20, -9, 3, -5, 13, -8, 0, -2, -3, -4, -9, 22, -7, -7, -4, 10, 9, 8, -5, 28, 9, -1, -8, -12, 0, 23, 9, -41, -1, -19, -8, -2, -28, -4, 3, -5, -7, -3, -11, -27, -1, 10, 7, -4, 9, 0, -2, -23, -12, -9, 27, -33, 0, 18, 3, 10, -4, 1, -17, -75, 3, -73, -23, -30, -10, 0, 10, 31, -8, -19, -33, -29, -6, -1, 0, -3, -12, 46, -3, 25, -45, 12, 15, 13, -5, -15, 2, 37, -10, -21, -2, -8, 15, 3, -5, -29, -31, 6, 5, 2, 0, -11, -8, 16, 6, -5, 1, 50, 1, -32, -5, 6, 3, -23, 9, -16, 21, 21, 16, -14, -3, 5, 22, -6, -11,
    -- layer=3 filter=0 channel=6
    23, 26, 9, -6, -5, 62, -6, 13, -23, -3, -1, 1, 13, 3, 20, 34, -13, 16, 2, -26, -56, -14, -35, 25, 33, -42, -4, -8, -5, 11, 15, -10, -1, -6, 5, -12, -9, -10, 13, 10, 7, 2, -4, -7, -47, -18, 3, 0, 2, -15, -10, -2, 16, 1, 0, -18, -5, -16, -5, -3, 10, 2, -3, 8, 0, 1, 18, -4, -3, 1, -38, 1, 2, 5, -11, -72, 8, 0, -5, 7, 12, 11, 5, 17, 8, -28, 5, -30, -29, -37, -19, 13, 0, -12, 6, 22, 3, 16, 23, -4, -22, 5, -19, 6, -47, 21, 19, 0, 23, -13, 23, -16, -68, 14, -18, 26, -32, 10, 3, 37, 5, 12, -2, 10, -6, 31, -11, 22, 9, 0, 16, -8, -2, -9, -2, 5, 57, 5, 0, 2, -11, 1, 9, 11, -2, 5, 9, 13, 32, 11, -3, 0, 2, 7, 0, 4, -20, -10, -49, 1, 14, 4, -46, -39, 4, -19, -8, -7, 0, 11, -19, -2, -36, -12, -6, 1, -10, -8, 2, 4, 10, 2, -34, -19, 39, -25, 1, -49, 0, -12, -45, 7, 9, 6, -22, -31, 4, -5, -32, -1, -1, -61, -20, -1, -18, -20, 1, -3, 16, 5, -19, 11, 19, -6, -29, -19, 8, 7, 7, -2, -50, -2, 57, 15, 7, 16, -43, 5, 3, 24, -14, 4, 33, 3, -2, 12, 29, -30, 11, 3, 7, 9, -14, 5, 32, -28, 1, 15, -14, -4, -8, 1, 9, -19, -41, 1, -52, -7, -3, -19, -23, -5, -12, 2, -12, 37, 6, 0, -7, -52, -14, 41, -64, 27, -11, -59, 29, 0, -45, 5, -4, -8, 9, 30, 8, -14, -6, 19, -3, -1, -7, 3, -9, 4, 4, 33, 17, 16, -43, 11, 0, 23, -14, 0, 1, 0, -55, 10, 8, 3, -3, 28, 16, -1, -4, -60, -41, 11, -3, 3, -26, 11, 38, -7, 0, -4, -31, 0, -12, 3, -9, -13, 10, 59, -4, -5, -54, 14, 5, 14, -5, 0, 1, -72, 3, 39, 22, -10, 8, -36, 31, 0, 15, -1, -1, -6, -9, -34, -2, -16, 1, -7, -8, -12, -4, -48, 2, -23, 12, -10, -4, 0, -36, 49, -6, 41, -41, 25, -69, 5, 10, -19, -58, 5, 3, -17, -2, 17, -10, -3, -7, -10, 20, 13, -10, -14, 10, -17, 22, -30, -8, 8, 10, -17, 31, -7, 15, 8, 0, 19, 7, 4, -15, 5, -17, -13, 45, -17, -18, -33, -15, 25, -5, 0, -13, -42, -48, -8, 4, -1, -23, 2, -17, -6, -56, 5, 2, -60, -25, -21, -22, -6, -3, -7, -56, 21, -2, -3, 2, 3, 39, 30, -7, -10, -4, -3, -43, 5, -29, -1, -57, -11, -34, 0, 16, 10, -5, 55, -33, -28, -10, 23, 12, 18, 25, -2, 5, -14, -31, 34, 8, 0, -9, -58, -15, 8, -9, 0, 53, -6, -2, -23, 8, 21, -13, 44, 6, 0, 0, -4, 15, 21, 34, 4, 12, 12, -8, -1, -8, -32, 22, -12, -7, -33, -2, -31, -20, 7, 14, 0, 11, 56, 5, 1, -12, 37, -5, 11, -4, -11, -69, -65, -6, -19, 2, -42, 3, -71, -13, 11, 5, 11, 12, -12, -2, 10, 11, 7, 2, 3, -13, -17, 12, 39, -12, -33, 0, 18, 2, -9, -15, 14, 4, 51, -27, -71, 0, -30, -13, -5, -10, -8, 20, -10, 4, 1, -5, 1, -12, -9, -10, -8, -26, -38, 10, -8, -55, 11, -4, 21, 11, 5, 24, -2, -2, -7, 7, -38, -11, -25, 1, -21, 38, -41, -7, -29, -31, -73, -8, 2, -3, 31, 18, 30, -40, -6, -33, 0, -23, 6, -14, -55, 15, -35, 12, -10, 35, 12, -5, 7, -11, 29, 22, 5, 15, 6, -14, -27, 22, -13, 5, 40, 16, -7, -1, 9, 30, -3, 3, 21, -12, -6, -10, -25, -4, -18, 11, -21, -44, -30, 25, 11, -27, -3, 4, -59, -6, -11, 27, 11, -15, 1, 44, 8, 35, -33, -2, 18, -17, -12, 0, -48, -10, 18, 11, -7, -6, -3, -22, -7, 14, -11, 3, 5, -29, -6, 2, -5, 2, -40, -13, 24, 46, -22, 15, 37, -19, -16, 7, -3, 6, 7, -38, -4, 5, 4, -57, 44, 5, 2, 17, -3, -23, 7, -4, -72, -46, -41, 3, 35, -14, 7, -30, -2, -15, -55, -2, -17, 19, 26, -7, -12, -11, 1, 12, -30, 3, 5, 10, -18, -8, 7, 23, 9, 20, 8, 41, -60, -7, -30, -17, -32, -11, -8, -20, -19, 32, -6, -20, -37, -11, 15, 4, -20, 29, -15, 1, -13, 5, 0, 5, -17, 12, -20, 1, -13, 1, -18, -13, 5, -83, 57, 3, 3, -62, -29, 5, 13, 35, -35, 9, -7, 0, -23, 1, 4, -14, -36, -54, -9, -6, 18, -36, -23, 0, -4, -16, -8, 18, 21, 25, -7, -6, -16, 19, -6, 11, -12, 25, 16, 8, 0, -34, 0, 31, -19, -11, 3, -7, -23, 0, -9, 31, -72, -4, -21, 10, 10, -23, 31, 11, 5, 2, 11, 3, -38, -12, -35, 8, -8, -8, -4, 10, -50, 10, -1, 23, -4, 33, 24, -41, -38, -10, 1, -6, -12, -17, 6, 43, -6, -28, 5, 28, 0, 45, -2, -20, 16, 4, 24, 10, -4, 5, -47, 16, 42, -12, -7, -20, 72, -10, 0, 17, 3, -6, 30, -8, -13, 4, -3, 6, 4, 7, 43, 23, 19, -1, -9, -28, -13, -3, 53, -8, -6, -15, -3, 23, 2, -8, -6, 49, -47, 6, -13, -3, -1, 3, 37, -17, 0, 23, 0, -70, -13, 13, -7, -5, -5, 2, -36, -15, 7, -2, -15, 10, -28, -20, 0, -42, -7, -24, 8, -78, 5, 11, -2, -25, 3, -16, -20, 8, 5, 33, 46, 11, 9, -2, -2, 8, -74, -24, -19, 6, -58, -6, 0, 31, -2, -4, -2, -15, 23, 2, -4, 45, -24, -2, -15, -4, 7, 5, 6, -14, -3, 23, -22, 10, 29, 0, -14, -3, 4, -21, 13, 47, -4, -10, 50, 5, 9, -6, -17, -22, 0, 81, -38, -12, -56, -4, 23, 16, -20, -1, -12, 10, 4, 45, -41, -61, 5, -24, 4, 1, -50, 10, 0, -56, -43, 41, 8, 36, -24, 2, 44, 37, -37, 9, -3, 6, 17, -11, -4, 4, 14, 81, -31, 22, 42, -47, 3, -4, 3, -8, -44, -33, 44, 29, 5, 4, -59, -8, 0, 10, 10, 18, 49, -3, 22, 35, 8, -31, 10, -7, -13, -17, 34, 1, 3, 4, -17, 10, -47, -6, 2, -8, 25, 5, -44, 11, 42, -3, 4, 10, -11, 57, -14, -7, 17, 49, 47, 6, 1, 4, 26, -13, 42, -79, 14, -25, -13, -7, -14, -87, 31, -38, -12, 7, -3, -80, -17, -107, 25, 11, -46, -7, 44, -26, -9, -8, 4, 18, 45, -2, 40, 27, -46, -7, -13, -17, 3, -15, 33, 4, 0, -5, -32, 20, 18, -10, 13, -12, 17, -31, -8, 7, -1, -8, 31, -4, 8, -19, -1, -51, -2, 23, 44, -40, -13, 3, 3, 2, -1, -15, -92, -81, 1, 99, 0, -41, -10, -16, -8, -65, 3, 10, -6, -12, 27, -30, -61, 4, -61, -78, 41, 0, 10, -6, -69, 24, -25, 1, -9, 23, -12, -39, 32, 1, 0, -55, -18, 1, 6, 0, 4, -38, -65, 1, -41, 54, -1, 18, 8, -20, 0, 48, -3, -45, -4, -14, 4, -5, -35, 6, 16, -6, -4, 21, -60, 6, 0, 1, -46, -14, -3, 50, 3, 10, 4, 40, 51, -32, -46, -34, -7, 7, 4, 63, 2, -28, -17, 7, -39, 12, -60, -11, 3, 10, 41, 34, 30, -5, -4, 61, -3, -11, -28, 27, 6, 13, 64, -26, -13, -3, 8, -12, -52, 0, 8, 6, 4, 31, -31, 9, -5, 1, -14, 3, 4, 20, -32, -6, 6, -5, 22, -29, -23, -13, -4, 1, 4, 24, 3, 9, -10, 0, -12, -32, 14, -8, -34, -6, 29, 0, -9, -3, -5, 14, -17, 0, 3, 16, 5, -5, 9, -74, 2, -9, -68, -5, 5, 10, 31, -11, -28, 2, -7, 11, -70, -32, -15, 3, -31, -9, -8, 17, -67, 8, -9, 0, 15, 14, -9, -26, 19, -30, 11, -34, 0, -37, 30, -1, -3, 44, 0, -45, 52, -40, -6, 5, 38, -18, 6, -73, 1, -1, -5, -85, 47, -6, 54, -60, 1, -6, -7, -9, 4, 0, 4, -10, -14, 2, -37, 0, 16, -5, 16, -50, 23, 20, -2, -10, -6, -3, 17, -7, -13, 9, 4, -25, 6, 7, -7, -19, 39, -2, 0, -4, 18, 1, 24, -9, 1, -8, -8, -17, -2, -29, -15, 35, -5, -6, 22, 7, -11, 1, 52, 13, -39, -26, 12, 38, 46, 10, 25, -12, -49, -2, -15, 0, 8, -3, 15, -11, 0, -27, 19, 19, 5, 31, 0, 44, -84, 0, -44, 66, -3, 15, 19, 7, -9, 18, -25, 10, 1, 4, -16, -8, -24, 0, 23, 7, 3, -26, -39, -12, -12, 16, -21, 6, 22, -26, 6, -2, -2, 0, -1, -10, -1, 13, -30, -13, -8, 11, 23, 12, -6, -41, -11, 5, -55, 0, -11, -13, -6, -16, 40, -8, -10, 28, 13, -22, 1, 36, 6, -6, 40, -21, -9, -34, -27, -16, -14, 0, -9, -14, 26, 18, -34, -9, 1, -20, -12, 8, -1, -7, -28, -57, 23, -9, -6, -13, 27, 1, -14, -10, 32, -13, 21, 18, -19, -6, -40, -3, 2, 5, 30, 31, -17, 1, -28, -38, -4, 71, 27, -8, -13, -41, -5, 3, 1, 29, 12, -14, 10, 8, -12, 22, 8, 2, -9, -8, 7, 5, 21, -27, -35, 14, -38, -12, -3, -42, 0, 7, -1, -56, -45, -6, 5, -25, 1, 8, 3, -56, 7, 14, -4, 56, 0, -35, 7, 31, 35, 42, -17, 7, -33, 20, -16, 39, -3, 15, 36, 32, 50, -5, 6, -21, 19, 3, 4, 22, -14, -21, -19, -2, -3, -13, 20, -13, 15, 7, 0, 26, 35, 3, 2, -18, -4, 12, 35, 11, 10, -54, 14, -45, -3, 16, -28, 32, 0, 4, -6, 6, -7, -16, -27, -89, 10, 20, -5, -56, -11, -18, -3, -22, -11, -10, -35, -15, 25, 17, 29, -2, -6, -37, 27, -77, -29, -13, 3, -14, -19, -10, 12, 26, -12, 1, -30, 9, 18, 2, 3, 13, 2, -1, -5, -4, -52, 17, -10, -37, 13, 4, 6, 31, 11, -23, 10, -8, 19, -11, 20, 34, -39, -9, 26, -3, 4, -10, 2, -8, -15, -12, 14, -14, 14, -3, -5, -32, -11, -12, 23, -19, -63, -31, 13, -24, -1, 12, 11, -37, 1, -59, -30, -8, 3, 17, -25, -7, 18, -5, 2, 6, 9, -8, -6, -6, 18, 7, 3, -20, 21, -25, 6, 10, 4, -7, -23, -27, 23, -1, -1, 27, 9, 5, -11, 0, 13, 11, 10, -1, 12, -35, 3, -4, -5, -61, -13, 11, 7, 5, -15, -11, 0, -3, 36, 2, 0, -22, 5, 6, 6, 16, -24, 11, 20, -19, 8, -13, -45, -8, -4, -49, -5, 11, 4, -3, 24, -12, -27, 1, -3, -18, -40, 9, 13, -6, -11, 0, 25, -26, -26, -64, 42, -5, -11, 14, -13, -7, -4, -8, 2, 12, -48, 22, 5, -9, 6, -39, 7, -11, 0, -6, 38, -12, 1, 14, 7, -8, -32, -16, -38, -18, -33, 6, -2, 13, 2, -5, 53, 3, 6, -20, 37, -8, -16, 22, 7, 0, -2, -11, -13, -13, 22, -12, 26, 3, 6, -4, 10, 41, -14, 0, -3, -1, -32, 6, 1, 28, 10, -48, -9, 16, -31, -40, -2, -16, -2, -1, 10, 6, 6, -6, -14, -15, -14, -15, 10, -11, 4, 2, -10, 1, 7, 28, -29, -12, 10, 6, 12, -8, -24, -2, -11, 0, -4, -2, 7, -6, 4, 20, 1, 22, 43, -10, 0, 36, -12, -3, -1, 5, 7, 11, -36, 14, -37, -7, 0, 0, -19, 24, 14, -4, 1, 17, -72, 1, 1, 1, -44, -3, 0, 2, -5, -13, -1, 12, 37, -30, 2, 27, -17, 2, 1, 4, -8, -13, 3, -7, -28, -23, 9, -3, 1, -40, -33, 24, -3, -44, 13, 6, -29, -11, -9, 10, 0, -46, 61, 0, -8, 31, 25, 9, 13, 18, 10, 11, 7, -11, -1, -4, 15, -2, -11, 17, -10, 0, -8, 17, -38, -5, -4, -20, -19, 5, 7, 13, -36, 6, -13, -13, -54, -20, 21, -3, 5, -16, -12, -27, 11, 0, -42, -15, -26, -21, 3, -5, 18, -9, 39, -13, 0, 41, -10, 34, 26, -9, -11, -6, -4, -11, -5, 16, 40, 10, 10, 5, -5, -2, -25, -2, 5, 2, 9, -12, 40, -35, -29, -33, -47, -12, -6, 22, -38, -3, 6, 20, 4, 0, -13, -11, 23, -19, -12, 0, 9, 26, 9, -21, 20, 3, 1, -14, -13, 22, -4, -23, -59, 15, -17, 36, 0, -6, -23, 25, 52, 5, -5, -18, -15, -9, -15, 12, 7, 55, 14, 2, -5, 5, 27, 37, 12, -10, -16, -8, -30, 9, 4, -46, 13, -9, -86, -11, -12, 50, 11, -68, 16, 12, 0, 2, -32, -16, 6, -10, -8, -9, 35, 2, -12, -25, 1, -36, -2, -14, 4, 37, 10, 10, -3, -23, -10, -19, -2, 0, -31, -24, 10, -3, 5, 4, 32, -30, 17, -4, 0, 33, -10, -19, 30, -17, 10, -13, 19, -5, 1, -4, -8, 50, -49, 12, -40, 11, 36, 13, 30, 44, -7, 33, -22, 33, -2, 4, -44, 32, -53, -9, -34, 4, -9, 16, -37, 12, 31, 5, 10, -2, 10, -20, 9, 19, -14, -16, -23, -12, -3, -41, -22, -8, 2, 16, -20, -23, -1,
    -- layer=3 filter=0 channel=7
    -4, -24, 14, -13, 3, -29, 3, 21, 38, -10, 9, 2, 5, -33, 3, -21, 6, -4, 29, 1, -24, -17, 9, 0, -11, 24, 0, -56, 6, -24, -12, 26, -11, 8, 3, -9, 5, 13, -8, 5, 43, -34, -14, 0, -39, 41, -6, 8, 0, 18, -31, -15, -6, 3, -10, -28, -22, -1, 8, -24, 16, 4, 0, -7, 65, 2, -15, -5, -11, 6, -39, 6, 10, -8, 41, 38, 9, 15, 5, -5, 31, 4, 7, 1, 0, 26, 9, 13, -24, 26, -13, 18, -10, -23, 19, 17, -1, 4, -28, -8, -1, -12, 0, -17, -1, -4, -15, -4, -17, -6, 7, 25, -17, -3, 24, 16, 10, -11, 21, 21, -48, -31, -20, -8, 3, 23, -18, -19, 10, -33, 5, 32, 11, 0, 0, -3, -35, 45, 2, -10, -13, 30, 1, -12, -5, 6, 15, 8, 7, 2, -13, -6, 1, 0, -4, -7, -27, -3, -9, -5, 24, -35, 36, -23, 16, -19, 2, -2, 2, 30, 7, 4, 7, -4, 43, 0, 0, 11, 5, -10, -7, 19, -14, -27, -24, -9, -3, -4, 4, -64, 3, 0, -6, 21, 18, -11, 3, -8, 21, 0, 16, 24, -11, -13, -12, -5, 10, 6, -37, 6, 0, -9, 9, 10, -32, -3, 2, 13, -10, -5, -35, 1, 13, -41, 4, 32, -18, -45, -5, -22, -12, 1, -20, 8, -36, -36, 9, -19, 0, 33, -1, 10, -16, -4, -4, 21, -30, 20, 7, -13, -10, -2, 20, -27, -2, -4, 4, -6, 11, 0, -13, -22, -13, -4, -32, -55, 12, -4, -23, 23, 30, -22, 39, -12, 9, -32, 0, 7, 0, -8, -23, -66, -29, 5, 9, 10, 11, 9, -2, -8, 2, 22, 0, -6, -36, -3, -11, -19, 35, -81, 44, -13, -13, 2, 18, 1, -26, 0, -63, 0, 1, -21, -13, 14, -6, 11, 17, -48, 7, -14, 62, 3, 8, -12, 7, -8, -31, 33, -7, -10, 18, 4, 6, -48, -3, -1, 61, 12, -9, -42, -13, 3, -6, 41, -58, -21, -48, -47, -7, 22, -10, -25, -27, -3, -42, 17, 62, 18, -24, 18, 23, 5, 4, 5, 6, 0, -46, 18, -9, 0, -40, 37, -1, -40, -22, -14, 7, -12, 50, -11, 2, -27, -27, -17, -1, 10, -1, 9, -10, 14, 18, 11, 8, 24, -2, -9, -13, 15, -20, 32, 10, -7, -56, -27, -11, 4, -26, -9, 9, -32, 0, -5, -2, -10, -40, -25, -27, -40, -8, 3, -16, -37, -9, 11, -12, 9, -2, -1, 16, -7, 13, -4, -4, -1, 2, -9, -6, 66, -49, 0, -1, -15, 1, 25, -41, -7, 7, 25, -7, -18, -51, -6, 8, -12, 30, -1, 10, -17, -2, 3, 29, -23, -1, 21, -23, 0, 42, -36, -65, 34, 24, 0, -6, -38, 8, -2, 7, 18, 17, -46, -12, 23, 8, 15, 12, -26, -8, -1, -9, 19, -10, -37, -34, 21, 10, 32, -27, -16, -6, 0, 9, 37, -38, 23, 0, -7, 13, -4, 11, 28, 0, -24, -35, -28, -6, 22, -6, -8, -8, 33, 35, -65, 3, -4, -65, 24, 10, 8, -9, -1, 6, 33, -24, -2, 0, 0, -20, -24, -29, -19, -13, -55, 45, 44, 2, -11, -4, -3, -1, -9, -1, -13, 30, -21, -46, -1, -30, 54, -10, 0, 14, 14, -1, 40, 1, 32, 3, -30, -19, 6, -10, -24, -37, -24, -11, 1, 3, 3, 6, -10, 2, -3, -58, 0, 9, -11, 30, 4, 6, 21, 11, -1, 25, 3, -1, 25, 2, 7, -8, 20, -37, 21, 3, 38, 8, -1, 26, 56, -4, 0, 9, 0, 5, -6, -41, 19, 34, 17, 36, -1, -15, 0, 40, -21, 49, -1, -6, -40, 30, 18, 14, -28, -25, -4, 46, 0, -6, -34, -12, 1, 0, 24, -7, 1, -6, -6, -5, -9, -39, -10, 1, 9, -5, 10, -9, -10, -10, -13, -10, 32, 35, -6, 5, 2, 0, -3, 1, -9, -10, -8, -4, -1, -6, -53, -14, -14, 15, -5, -7, -10, -2, 33, 22, -8, 14, -1, 23, -7, 8, 6, -29, 9, 0, 76, -47, 8, 32, -7, 1, -3, 17, 34, 22, -6, -17, -23, 20, 22, -8, -9, -33, -11, 0, 47, -34, -5, -29, 17, -13, 15, -39, 5, -33, -40, -32, 21, 30, -19, -28, -3, 22, 2, -29, -5, 23, -13, -14, -19, -40, 20, -2, -21, 10, 9, 37, 68, -35, 15, -24, -3, -5, 0, -39, -1, -13, 1, -5, -1, -4, -25, 27, -1, -21, -5, 5, 14, -8, -3, -50, 39, -3, 7, -20, -13, 8, 5, -2, 16, 7, 2, 0, -5, 23, 14, 20, -6, 2, 26, -66, 5, -6, -20, 43, -29, -79, 17, -7, -16, 9, 36, 0, -8, -20, -10, -7, -3, 1, -28, 5, 1, 27, -39, 20, 10, -7, 8, -12, 11, -19, 8, 31, -8, -7, -9, 7, -4, 10, -10, -16, 7, 5, 28, 6, 6, -3, 4, -2, -9, -14, 39, -5, 0, -34, -8, -7, 15, -7, 5, 34, 17, -8, 17, 2, -25, 14, -6, -12, 3, 13, 42, 3, 13, 37, 25, -23, -1, 10, 23, -4, -13, 36, 1, -71, 23, -17, -2, 0, 3, -44, 22, -1, 8, 17, -14, -40, -9, 2, -62, 4, -7, -6, -2, -17, 40, -3, -6, -10, 30, -15, -68, 8, 9, 32, 4, -19, -6, -4, 10, -8, -6, 27, -3, -2, -5, -62, -7, 32, 9, 67, 1, 17, -23, 6, -4, 3, 4, -32, 3, 1, 15, -41, -11, -9, 21, 9, -7, -21, 20, 5, 14, -31, 0, 29, 3, -8, 2, 12, -15, -13, -77, -17, -29, 12, 28, -6, -6, 3, -30, 0, 0, -1, -3, 0, 19, 0, -16, 13, 5, -39, -17, -13, 0, -22, -81, -24, 18, 36, 2, 26, 27, 15, 11, 38, 71, 21, 6, -6, -8, -20, 8, 8, 21, 4, -10, -34, 49, 2, -24, 0, -7, 44, 45, 33, 39, 27, -2, 10, 7, -11, -5, -19, 0, -24, 11, -55, 14, 40, -5, -4, 0, 40, -14, -10, -2, -76, -42, 0, 12, 6, -67, 14, 20, -19, 37, -10, 3, -28, 17, 5, 32, -3, -18, -17, -52, -15, 7, -28, 33, -55, 20, 13, -56, -10, -13, -69, -10, 4, -4, -17, -11, 9, 0, -13, 25, -38, 4, -10, -4, -30, 24, -6, 8, -2, 60, 19, -6, -10, 11, 6, 50, -8, 8, -12, 34, 26, 6, 12, -1, -2, -14, -45, -2, -12, -6, 9, -95, -13, -5, 3, -7, -1, 92, 3, -10, 20, 1, 9, 6, 9, -2, 2, -24, -4, 6, -46, 2, -12, 24, -71, 27, -16, 2, 24, -4, -11, -23, -29, 29, -1, 20, 47, 0, 27, -43, -39, -18, 19, -1, 24, 17, 39, -7, 15, -9, 20, -75, 13, 12, 17, -18, -5, 2, -1, -1, 43, 4, 9, 6, -24, 1, 23, -79, -4, 2, 13, -1, -24, 6, 2, -26, 37, -29, -25, 12, -17, 12, -5, -22, 0, 6, -38, 11, -85, 1, -33, -36, 5, -31, -17, 19, 5, 13, -16, -2, -13, -7, -7, 12, 26, -4, -10, 1, 16, -9, -8, -73, -47, 0, -39, -44, -7, 5, -57, -1, -8, -10, -22, 32, -30, -16, 10, 0, -22, 5, 32, -64, -26, 5, 38, -40, -77, 10, 1, -15, -7, 9, -30, 19, -9, -67, -39, -14, 15, 0, 5, -7, 18, 7, 15, 23, -23, 26, -5, 35, -1, -13, 59, 45, 3, 30, 6, 14, -19, 4, -52, -11, -8, 2, -19, -13, -13, 23, -19, -48, 5, -11, -73, 52, 27, -22, -29, -56, 0, -16, 2, -19, 3, 32, 16, 10, -8, -18, -35, 1, -63, -19, 8, -1, 4, -30, -27, -2, -25, -23, -5, 6, 8, -48, 0, -32, 9, 28, -2, 8, 5, 6, -11, -6, -2, -17, -25, 16, 7, -1, -15, 31, 5, 5, 11, -5, 12, -11, 14, 36, -1, -33, 28, -8, -3, -38, -9, -35, 3, -28, 21, -4, -26, 18, -16, 14, -15, -5, -3, -1, 17, -5, -11, 3, -8, -9, 66, -18, 0, 24, -11, -32, 11, -22, -8, 9, -7, 9, -3, 8, -29, -25, 0, 9, -16, -14, -12, -8, -31, -4, 13, -4, -54, 12, 10, 1, -16, -12, 29, 6, 23, 24, 7, -50, -26, -49, 18, 48, -7, 0, -9, 0, 5, -44, 11, -81, -20, -45, -5, 1, -36, 8, -19, 17, 3, 4, -1, 13, -11, 15, 5, -31, 55, 16, 20, 0, -39, -2, 15, -29, 0, 2, 11, 2, -35, 1, -20, -18, 37, -41, -13, 28, 4, -7, -3, 0, -15, 9, 26, -5, 12, -7, 32, -1, -8, -5, -3, -3, 14, 2, 3, -25, 3, -13, 0, -5, -70, 4, 15, -55, -2, 11, 13, -23, -17, 2, 7, -12, -1, -17, 12, -10, 7, 12, -1, 13, -52, -11, 13, 52, -71, -74, -24, -14, -40, -10, -44, -5, -6, 44, -3, 35, -40, -4, -8, 3, -7, 1, 26, -6, 1, 2, 13, 12, -16, 7, -16, -1, -4, -1, 19, 12, 29, -39, -24, 7, -2, -9, -19, 17, 16, 1, 17, 54, -4, 50, 4, -29, -9, -22, -41, -13, -5, -3, 25, -12, -31, 9, 19, -6, 8, -46, -28, -11, 20, 2, 11, 39, 14, -58, 0, 28, -8, 14, -8, 11, 4, -13, -2, -1, 44, -12, 25, -10, 27, 39, 49, -75, -14, 5, 9, -92, -15, -19, 19, -44, 6, -2, 44, 3, 9, -41, 14, 7, -1, 5, 66, 10, 2, -18, 0, 7, 23, 19, 1, 1, -42, -7, 4, -31, 1, 7, -81, 26, -10, 18, -17, -38, -4, 28, -35, 29, 1, -3, 4, 3, 7, 20, -8, -2, 69, -2, 20, 16, -41, -8, 6, 2, -24, -13, 10, 9, 15, 7, -53, 0, -50, -30, -29, -32, 5, -62, 13, -8, 19, 11, 0, -32, -17, -23, 10, -50, -22, -8, -11, 1, -49, 9, 33, -65, -17, 10, 9, 3, 28, -5, 7, -26, -36, -49, 20, -11, 52, 11, -5, -23, -7, 0, 11, 0, 32, -19, -12, 20, 17, 25, -13, 21, -10, -7, -4, 14, -41, 2, -22, -6, 31, 10, -25, 2, 26, -9, 4, -23, -21, -13, 20, -26, 3, -2, 12, 19, 5, 15, 34, -8, 37, 24, -11, 0, -38, 3, -10, -13, -36, -16, 2, -47, -8, -7, -2, -10, 51, 12, 12, 50, 12, 15, 70, 42, 26, -11, 8, 16, 12, 15, 0, -64, 6, 40, 7, 6, 1, -6, 0, 23, 36, 16, 20, -25, -11, 14, 43, 1, -5, 0, 16, 19, 17, -16, 6, -40, -22, 0, 39, -16, -9, 4, -1, -11, 0, -16, -8, 19, 0, -10, -52, 10, 5, 4, 16, 0, -19, -11, -14, -15, 16, -38, -30, -13, -33, -1, 7, 20, 21, -40, -5, -10, -13, 13, 14, -11, -29, -3, -12, 5, 46, -54, 58, 8, 11, 29, -5, -13, -6, 0, 8, -36, -47, 24, 4, 23, -15, -13, 2, 10, -12, -40, -53, 2, -1, 47, -30, -5, -71, 36, -14, 5, 45, 1, -1, 4, -25, -50, 12, 5, -12, -1, 10, -5, 1, 23, -6, -60, 9, -21, -46, -17, 12, -13, 14, -15, 6, 34, -13, -5, -12, 6, -7, -6, -31, -2, 9, 2, 9, -7, -60, -30, 69, 11, 32, -11, -2, 20, -37, -28, -53, -15, 32, -13, 22, -3, -6, 0, -28, -4, -5, -4, -70, -4, 1, 15, -24, 11, -24, 0, -13, -2, -8, 12, -2, -3, -5, -40, 40, -16, -9, 1, -3, -4, -4, 22, -6, -10, 3, 10, -14, 7, 3, 16, 5, -42, -12, 19, -6, -7, -9, 8, -4, 0, -2, 1, 30, -7, 11, 17, -8, -12, -7, 13, 17, 13, 40, -44, 7, -3, 35, 19, -24, -17, -1, -4, -16, -13, -9, -11, -6, 4, -7, 32, 8, -3, 12, -39, 31, 4, 25, -5, -56, -8, 0, 40, 0, -39, -16, 27, -23, -3, -12, -10, -21, 18, -15, -47, -27, 56, -1, 36, 8, -12, -10, -33, 9, -3, 17, -6, -1, 26, 36, 5, 4, 15, 5, -66, -9, -51, -6, -29, 2, -12, 41, 0, 0, -13, -33, -26, 4, 3, -8, -25, -10, -24, 50, 5, -2, -5, 49, -5, -47, -35, 21, -11, 19, -57, 1, -6, 9, -31, -9, 41, 17, -9, 5, 6, -8, 39, 8, -2, -7, -23, -2, 14, 28, -26, -7, 10, -10, 51, 4, -29, -9, -7, 0, -17, 47, 4, 31, 14, 13, 9, 11, -7, -1, 0, -18, -31, -7, 42, -16, 0, -9, 13, 24, 4, 32, 27, 0, 10, -11, -16, 6, 2, -8, -13, -1, 28, -12, -16, 0, -2, -1, -33, 37, 16, -23, 44, -22, -14, -50, 28, 0, -4, -24, 0, 38, -22, -2, -15, 16, -1, -48, -14, -18, 0, 1, 22, 53, 1, 37, -33, 31, 5, 17, -20, -33, 23, -20, 7, -10, 8, -12, -56, 0, -26, -12, -20, 10, -16, -45, 2, -84, -29, -17, 6, -2, -20, -19, 32, 6, -21, 14, -31, -3, 2, -12, 9, -23, 24, -2, -11, -5, -13, -1, -4, 29, 21, 11, -9, -18, 26, -8, -11, -11, -15, -15, -10, 44, 2, -20, 9, -4, 9, -32, 0, -13, -42, 10, -19, 4, -43, -7, -13, 19, 8, -41, 3, -42, -50, -48, -10, 0, -13, -18, 4, 4, 1, -40, 2, 19, -44, -4, 17, 2, -6, -24, 42, 40, 17, 37, -51, -10, 8, -49, 3, 0, 9, -12, -15, 15, 25, -6, 41, -14, 37, 6, 6, -32, -9, 18, -25, 10, 9, -72, -19, 42, 7, 39, 11, -23, -22, -16, -107, -38, -41, -10, 8, -13, 20, 80, -18,
    -- layer=3 filter=0 channel=8
    -25, -18, 0, 2, 2, -78, -13, -14, 10, 33, -8, 9, -38, -40, -23, -33, -27, -15, -61, -1, 9, -6, 8, -35, -25, 28, 9, 5, 10, -3, -39, 34, -12, 0, -7, 0, 8, -2, -31, 2, -4, -5, -15, 19, -14, 23, 4, 4, -39, 17, -24, -11, -45, 1, -6, -20, 2, -11, 4, -6, 29, -19, 3, -14, -36, 10, 27, 31, -10, -18, 9, 6, 6, 13, 3, -44, -2, -17, 9, -7, -25, 32, -8, -8, 4, 17, 2, 26, -22, 12, -34, 25, 5, 0, 8, 4, 8, -18, -68, -1, -54, 0, 2, 8, 47, -11, 27, -10, 23, -1, 7, -35, 24, 10, 20, -30, 4, 0, -27, 32, -19, 30, -44, 5, 5, -28, -34, 9, -6, 0, 11, 15, 1, -8, 11, 8, 10, 3, 10, 11, 0, -35, 32, 23, 11, -47, -24, -5, 21, -2, 10, -7, 3, -7, 1, 0, 19, -12, -18, -13, 30, 10, 10, -8, 5, -19, -5, 2, 1, -4, 19, -12, -18, 0, 51, -1, -12, -1, 32, 5, -14, 6, -12, -21, -24, 34, 4, 14, -4, -40, 4, -34, -1, 33, -1, 4, -1, 6, -40, -4, 30, 15, -13, -8, -48, 34, 12, 3, -5, -10, -9, 10, -1, -25, -44, 37, -2, -68, 3, -7, 23, -2, -17, -22, -7, 13, 11, -12, 1, -19, 4, -4, -28, 23, -3, -2, 0, 6, -10, 27, 23, -9, 3, -10, -28, 3, -98, 10, 17, -2, 6, 0, -43, -23, 19, -7, 3, -34, -6, 4, 11, -21, -2, -8, 17, -36, -13, -6, -2, -27, -1, -35, -15, -19, -40, 8, -28, -7, -1, 2, -28, 0, 10, -45, 6, 7, 37, 15, -6, 5, 0, -15, -12, -5, -20, -3, 11, -2, -2, 10, 23, -6, -1, -2, -4, 0, -21, -48, -1, 7, -9, -25, 15, 10, -3, -26, -1, 0, -5, 10, -15, -14, 8, -24, 0, -1, 50, 28, -12, -5, 10, -25, 14, 3, -9, 10, -8, 0, -3, 7, 2, -10, -7, 7, 14, -21, 8, -12, 4, -10, -7, -7, 2, 0, -28, 14, -18, 10, -3, 4, 7, 3, 32, -1, -11, -9, -15, -19, 4, 2, 2, -9, 7, 6, -29, 35, -42, 15, -38, -11, -15, 17, 22, -7, 0, -25, 0, 17, -1, 9, 8, -7, -31, 2, -3, -1, 0, 9, 19, 13, -13, -23, 7, -10, -16, 12, 0, 0, 0, -29, -10, 13, -13, -8, 2, -14, -11, 39, -26, 32, 0, 7, 1, -11, -1, 14, -7, 4, -20, 9, 3, -2, -7, -15, 4, -6, -12, -66, -24, -6, 8, -7, -15, 7, 15, 3, 0, -50, 1, -11, -24, 5, 7, -4, 0, 11, -6, -4, 6, 0, -56, -44, 7, 16, 10, -4, 3, -55, -15, 10, 27, -12, -11, -3, 33, 3, -4, -7, -18, -25, -7, 0, 0, 12, -3, -46, 6, 0, -49, -6, 0, -6, 35, -11, -33, 7, 12, 0, 19, -12, -31, -4, -43, 0, 9, -12, -1, -5, -14, 18, 4, 7, 12, 20, -5, 8, 5, -9, -6, -61, -43, -22, 10, -11, -22, -31, -12, 6, -44, -7, 0, 0, -16, -10, 3, 30, 0, 26, 37, 5, -14, 20, -11, 15, -2, 0, 7, -7, 0, -3, -26, 4, 6, -18, -3, 25, 14, -5, -3, -7, -16, 6, 31, -25, 8, 17, -5, -24, -1, 1, -12, -14, 22, -3, -6, 6, -34, 8, -8, 5, -1, -15, 24, 31, 10, -3, 14, -10, 4, -9, 0, -10, -54, -58, 5, -10, -5, 26, 14, 20, -23, -8, -27, -1, -6, -13, 21, -10, 4, -18, -51, -38, -5, 35, -10, -25, -15, 5, 17, 0, 18, -33, 6, 3, -1, 0, -12, -32, 27, 22, -20, 40, 2, 26, 10, 0, -17, 9, 3, 0, 0, -60, 21, 8, 3, -4, 2, -10, -18, 11, 8, 4, -6, 8, 0, 20, 1, -36, 40, -46, 0, -2, 3, -9, 19, 4, -5, 8, -32, 10, 27, -8, 6, 32, -36, -11, -1, 16, 3, -5, 1, -34, -29, 0, -6, -3, 12, -8, -26, 7, -1, -2, -10, -73, 4, 10, -66, 6, 9, 19, 5, 1, 22, -25, -4, 13, 16, 21, 12, 9, 7, -1, -11, 12, 25, -9, -47, -59, 4, -1, -26, -12, 15, 6, -10, -44, -9, 12, 3, 19, -31, -6, -6, -14, -18, 8, -19, 32, 16, 11, -8, 10, 0, -11, -30, -4, -3, -7, 16, -34, -41, 17, 53, -9, 5, -8, -66, 40, 12, 25, 17, -3, -28, -8, -42, 26, -19, -23, -1, -24, -7, -12, 7, 8, -41, -3, -30, -31, -5, -5, 5, -19, -48, 37, -74, 0, 5, -4, 9, -6, -4, 18, 1, 23, -5, 10, -8, -13, 10, 47, 10, -7, -10, -8, 8, 0, 6, 11, 25, -5, -21, 56, 3, -2, 11, -10, -15, -18, -14, 5, -4, 11, -7, 5, -20, 3, -5, 23, 14, -39, 8, -39, -16, 0, 34, -108, -1, 12, 35, -17, 0, -9, 8, -13, 2, 5, 12, 0, 46, 30, 7, 7, 0, -42, -9, 0, 17, 51, 18, -38, 0, 0, -4, -18, 0, -21, -44, -36, -6, 5, -18, 7, 34, -28, 11, 0, 9, -13, -4, 9, -38, -14, 13, 31, -33, 37, 41, 47, -14, 23, -18, -6, -15, 10, 3, -5, -13, -14, 12, 14, 3, -1, -27, 5, 33, 26, -16, -3, -15, -15, 11, 2, 0, 0, -19, 12, -15, -10, -50, -7, 17, -2, -11, 0, 10, -13, -50, -18, 16, 7, 0, 3, 9, -14, 2, -8, 1, -4, 20, -14, -24, -10, 21, -8, -1, -8, 28, 8, -6, -17, -18, -8, 18, 20, -10, -8, 24, 12, 3, -56, -20, 36, -16, -28, 2, 7, 20, -1, -5, 12, -8, -17, -20, 4, -44, 4, 4, -9, 21, 25, 5, 16, -22, 13, -41, -59, -62, -9, 32, -15, -10, -44, -3, -5, 0, -33, 5, -40, -7, 5, -44, 13, 24, -31, 31, -4, 25, 29, 30, 0, -8, 5, -64, -17, -44, 23, 35, 26, -9, 5, -29, -27, -53, 10, 45, -34, -11, -13, -8, 13, 5, -8, 9, -3, 8, 7, -62, -46, -13, -28, -32, 21, -2, -15, 60, -21, -2, 3, -5, 21, -54, 25, 2, -5, -13, 17, -2, 2, -2, -28, 7, 2, 21, 23, 48, 1, 11, 4, 16, 12, -12, 3, -10, -1, -12, 13, -5, 15, 0, -7, -1, 11, -5, -6, -23, 13, 2, -23, 27, -11, -24, -28, 3, -21, 67, -14, -1, 12, -14, -1, 1, -41, -4, 10, -59, 9, -1, 10, 2, -16, -9, -18, -1, -7, 40, 22, 5, 4, 27, 5, -1, 2, 23, 8, 6, 59, -25, -12, -19, -2, 16, 2, 20, 12, -13, 5, -1, -6, 38, 26, 20, 20, 2, 37, 16, -25, -18, -15, 3, -4, -46, -9, -6, 0, 3, 5, -9, -8, 44, -14, -7, 14, 10, -10, 6, 18, -13, 22, -5, -22, -41, -15, 13, 19, 37, 4, 23, -3, -12, -8, -25, 3, 59, -27, 16, 39, 17, 27, 5, 17, -8, -14, -15, 18, 65, -18, -15, 4, -50, -2, 13, -9, 17, 3, -4, -29, -19, 10, 28, -3, 7, 15, 3, -46, -2, -16, 13, 65, 25, 9, 0, -7, -25, -16, 26, -27, -17, 0, -1, -50, 6, 6, 17, 10, -5, -1, 42, -39, 3, 33, 31, -37, 7, -8, 4, -2, 0, -16, 2, -14, 19, -18, 1, -41, 5, 3, -28, -15, 27, -10, 28, -4, -47, 76, 31, -3, -36, 5, -55, -29, -33, 14, 2, 33, -24, 5, 20, 5, -4, -12, 19, 32, 1, 3, 1, 11, 11, -3, -6, -32, 5, -12, -65, 40, 22, -61, -7, 0, -25, -14, -1, -6, -19, 2, -28, -4, -11, -6, 5, -7, -12, 33, -5, 1, 12, -20, -11, -15, -48, -36, -10, -29, 12, -1, 35, 12, -14, 5, -5, -4, 6, -25, 5, 7, 3, -11, 11, 9, 10, -14, -37, -10, -6, -22, 7, -11, -9, -8, 0, -15, 55, -20, -7, 0, -16, -31, -21, 8, 3, 5, -27, -6, -1, -24, -10, 0, 11, -38, 0, 2, 17, -19, 3, 14, 21, 17, -17, -14, -22, 8, 15, 46, 18, 1, -31, 0, 14, 7, -17, -18, -14, -4, 39, -2, -33, 9, 12, 47, 29, 27, -11, -45, 32, -12, -13, -9, -8, -3, -4, 24, 18, -9, -1, 1, 46, -7, 24, 19, 2, -5, 0, -34, -19, -21, -6, -54, 44, 37, -11, -3, 50, -8, 4, 10, 4, -3, -11, 0, 71, -11, 45, 42, 20, 5, -4, -3, 6, 1, -21, -38, -48, -20, 24, -11, -11, -1, 7, -12, -7, -10, 9, -61, 0, -32, 14, 15, 0, 26, -16, -2, 7, 5, 33, 53, 19, -41, 0, 0, -44, 2, 36, 36, 1, -17, -45, -50, -35, -8, 8, 11, 26, 35, -36, -21, -31, -2, -15, 42, -17, 9, -5, -20, -16, 2, -6, 1, 9, -31, 0, -19, 7, -12, -8, -1, -16, -31, 3, -12, -43, 40, 18, -3, -15, 5, -51, -9, -49, -45, 42, -23, 0, -2, 4, -5, 4, -20, 11, -48, -3, -10, 9, 10, 0, 28, 13, -23, -8, -13, -36, 10, 0, -26, -9, -20, 49, 39, -19, 0, -35, -7, 21, 17, -13, 60, 0, -10, -25, 7, 0, 4, -14, 11, 0, 0, -18, 2, -59, 23, -47, 0, -51, -4, 2, 0, 3, -36, -19, -58, -65, 21, -2, -36, -5, 10, 10, 10, -27, -3, -2, -30, -10, 7, 15, -79, 0, 11, -31, -3, -5, 0, 19, 34, -20, -15, -3, -9, -74, -33, 1, 4, 2, 4, -10, -17, -20, -19, 26, -12, 1, -6, -9, -33, 0, -9, 11, -8, 6, -25, -7, -21, -60, -16, -6, -11, -33, -13, -10, -20, -10, -8, 5, 53, -64, 4, -28, 16, 29, -68, 31, 6, 0, -10, -53, -33, 1, 0, -5, -2, 12, 5, 49, 9, -9, 53, 16, -12, -5, -18, -74, -37, 4, 38, 3, 24, -10, 13, -29, 5, 13, 56, 4, 2, -18, 4, 19, -11, -20, 17, -16, 2, -14, -73, -13, 4, -4, 4, 18, -6, 59, -10, -37, 8, 9, 11, -12, -14, -1, 0, 41, -11, -26, -30, 8, -51, 19, -39, 12, 1, -30, 29, -9, -6, -9, -6, 58, 4, -5, 9, -4, -1, 35, 43, -7, 4, 0, 4, 14, 12, -24, 19, -49, -55, -70, -27, 1, 10, 33, 4, -34, 3, -17, 12, 2, -2, 8, -76, 7, -14, -14, 1, -23, -5, -33, -37, 37, -46, -37, -7, -15, -1, -49, 8, -16, -9, -69, 27, -11, 0, -3, -10, -30, -5, 4, -41, 6, -12, 0, 2, 7, 27, 16, 28, 1, -7, 41, -24, -4, 17, -27, 6, 5, 14, 48, -13, 19, 1, -25, 4, 27, 16, -2, -7, -51, -62, -13, 0, -9, -16, 2, 3, 0, 11, -6, 4, -67, 21, 14, 24, 5, 6, 10, -9, -5, -5, -15, 39, -6, -11, 13, 9, 0, 7, -4, 33, 8, 9, -17, -5, 52, -26, -10, 8, -8, -13, 6, -9, 0, 5, -5, 47, -4, 1, -10, 15, 8, -37, 3, 24, 3, -14, -18, -21, 67, 5, 3, -11, 25, 20, 1, -3, -38, -5, -44, -1, 10, -3, -51, -16, 5, -11, 29, 31, 41, -51, -33, 0, 15, -2, 3, 20, -35, 7, 1, -11, -2, -8, 0, 1, -68, 6, 7, -3, 29, -30, 13, 0, -17, -6, 59, 36, -19, 9, -9, 8, -41, -38, 0, -4, 29, 31, -8, -18, 34, 11, -4, 24, 8, -7, 36, -12, 26, 0, -46, -41, 26, 31, -4, -55, 7, 3, -10, -12, -39, -15, 48, -1, -27, -1, 1, 6, -6, -7, -9, -4, 9, -7, -68, -23, -3, -3, -8, 2, -8, 34, 29, 66, 59, 13, 9, 3, -3, 6, 29, -2, 18, -9, -11, 36, -17, 10, -35, 4, 38, 79, 38, -26, -5, -2, 11, -29, 28, 9, 62, -11, -72, -80, -17, 0, -5, -6, -3, 13, -5, 3, 28, -29, -20, -58, -16, -51, 81, -41, -15, -6, 21, 4, -6, -18, 25, 12, -19, 35, -12, 10, 37, -38, -46, 7, 47, 40, 5, -29, 0, 9, -12, 24, -16, 0, 8, 8, 2, 5, -1, -71, 24, -8, -24, 15, -8, 3, 37, -34, -10, 17, -18, 47, -6, -20, -25, 27, 2, -9, -12, 17, -5, 8, 7, -3, -85, 31, 57, -53, 27, 21, 3, 1, -10, 0, -8, -49, -70, -3, -4, -17, -8, -7, 10, 18, -30, 4, 6, -81, -51, -7, -36, -11, -7, 14, -47, -45, -12, -2, -4, -39, 3, -7, -5, -5, 15, 2, -5, -36, 6, 4, 13, -44, -48, -1, 83, -30, 13, -15, 5, 54, 13, -8, 15, 23, -46, -3, 11, 11, -29, 4, 10, 10, -32, 36, 35, 12, 38, 10, -42, -7, -9, 35, -16, 0, 1, -78, -17, -10, -2, -18, -12, -18, 0, 23, 6, -41, -5, 2, 22, 8, 19, -31, -20, 8, -1, 1, -7, -4, 1, -30, 10, 21, -5, 0, -56, -4, 10, 52, -6, -3, 9, -4, 26, -8, -52, -11, 22, 25, -9, -41, 8, -5, -14, -23, 20, -13, -30, 2, 33, 13, -47, -11, -39, -3, -6, -23, -10, 1, 1, -25, 10, 6, -17, -4, 5, 30, 17, 58, 17, -28, 1, -9, 29, 0, 43, 28, 18, -5, 24, -11, -20, 5, -42, 16, 3, 33, -12, -34, 22, -19, -34, -2, 4, -3, 0, 11, 29, -2, -6, -18, -6, 11, -5, -41, 9, -13, -7, -25, 18, -48, -40, 20, 8, -34, -10, 10, 18, 5, -6, -5, 23, -5, -5, 4, -15, 0, 4, -41, -81, 11,
    -- layer=3 filter=0 channel=9
    -9, 20, -8, 45, 15, -5, -5, 2, 19, -85, -5, 11, 28, -34, -26, -14, -22, -7, -3, 15, -1, -7, -2, -3, -8, -6, -45, 44, 7, 2, -36, -53, 9, -12, 0, -13, -12, -10, -15, -39, -20, 5, 34, 15, 8, 35, 19, -7, -6, 32, -39, 6, -4, 13, -12, -3, 42, 4, 10, 14, -10, 2, 0, -43, -58, -4, -34, -56, -6, -22, -17, -7, -6, -12, 39, 28, -12, 12, 1, -11, -30, 7, 12, 28, 10, 19, 9, 1, 11, 38, 34, 18, -10, 4, -8, -8, -9, -2, 34, 3, 19, 26, -22, 8, 5, -1, -1, -1, -20, 6, -13, 12, 14, 10, 16, -9, 23, 29, -34, -12, 14, 10, 46, -14, -12, -5, -5, 31, 0, -64, 23, -32, -6, 4, -6, 7, -25, -21, 0, -9, -13, -3, 42, -60, -14, 47, 29, -4, 4, -6, 23, -3, 10, 30, 12, -4, 0, 9, 12, -8, -53, -21, -35, 19, -7, 21, 6, 5, 5, 13, -30, -16, 1, 1, 29, -7, 0, -13, 2, -10, 0, -45, 35, 4, 27, -3, -11, -12, -19, 9, -26, 16, -13, -46, -24, 18, -3, 1, 30, -11, 7, -3, 16, -13, 16, 7, -16, -3, -5, 5, -11, 3, -35, 12, -7, -25, 13, 40, -76, 4, 6, 6, -7, 32, -4, -18, -29, 0, -8, -22, -13, 8, -50, 27, 13, -14, -20, 7, -15, -26, 18, 9, -10, 4, -25, 15, -14, 35, 24, 3, -15, 9, -34, -27, 10, 0, 52, 6, 0, 4, 10, -24, -16, 30, -12, 24, 7, -11, -32, -37, -52, -46, 15, 5, 12, 26, 2, -24, -3, -8, -2, -16, -23, 20, 1, -21, -5, -37, -6, -14, -23, -11, -9, 3, -13, 22, -27, 17, -24, -16, 13, -4, 20, -6, 0, -30, 45, -2, 1, 28, -16, -63, 32, 6, 12, -15, -17, -25, -2, -10, -25, -6, -38, 0, 6, 7, -31, -3, -9, -9, -8, 2, 9, -7, -2, 9, -31, -8, 7, 24, 0, 44, -12, -24, -28, -1, 75, -9, 1, -2, 0, 43, 4, 0, 31, -4, 9, 4, 20, 17, 3, -11, 31, 8, -35, -15, 32, -4, 12, 10, 28, -11, -2, -30, 15, 7, 33, -31, 4, -1, 4, -23, -10, -10, 8, -22, -12, -7, -7, 13, 16, -7, 0, 18, 0, 1, 9, -22, 38, 11, -8, 11, -8, 21, 43, 6, -10, -5, -5, 60, 0, 10, 19, -5, 13, -3, -27, 11, 30, 5, 3, 13, 2, -6, -4, -2, -67, -2, -22, 1, -21, -10, 30, -10, -12, 4, -2, -15, 24, -28, -11, -31, 13, -24, 24, -43, 3, -23, 13, 21, 0, 26, -1, 11, 20, 2, 29, -12, -4, -13, -24, -9, -27, 6, -6, 2, -1, -2, 34, 17, -12, -24, -20, 8, -63, 0, 1, 3, 3, 26, -9, -11, 0, -10, -3, 14, -4, 6, 17, 37, 3, 1, -11, -13, 6, -23, 39, -5, 9, -20, -29, 34, -19, 17, 17, 19, 2, -9, 5, -12, 0, -9, 0, -16, 6, 18, 11, -88, 22, 9, -34, -26, -13, -18, 8, -7, -49, -55, 27, 0, 9, 41, -10, -3, 5, -7, -44, 0, -10, 19, 15, -74, 25, -14, 7, -6, -5, -6, 1, 4, -31, -2, -13, 0, -20, -9, 13, 11, 20, -10, 0, 13, -14, 0, -22, 45, -11, 9, 19, -7, -2, -28, -29, 6, 6, -46, -53, -6, -10, -23, 6, 14, -5, 11, -13, -2, 0, 62, -14, 40, -11, 13, -63, -87, -2, -33, 2, -14, -8, -26, -34, 39, -3, -28, -4, -11, -15, 24, -14, 13, 30, 3, 33, -1, 10, -5, 22, -23, 4, 8, -44, 26, 14, 2, -7, 9, 32, -5, 19, -2, -2, -5, 42, -40, -63, 2, -13, 5, 26, 17, -9, -87, -2, -30, 12, 7, -36, -13, -15, -23, 2, -12, -2, -27, -29, 22, -8, 27, 11, 29, 23, -2, -19, -2, 8, 80, -14, 1, 32, -8, 10, -16, -16, 0, 10, 4, 0, -41, -2, -1, 13, -33, -34, -3, -33, -4, -2, -6, 37, 4, -39, -5, 12, -53, -20, -34, 31, -59, -5, 25, -16, -51, 31, 36, -23, 11, 4, 4, -6, 6, 40, -14, 6, 21, -18, 7, 22, -22, -19, 6, 22, -8, -103, 10, 52, 6, -30, 6, -5, -8, 0, -12, 13, 5, -19, 41, 2, 24, 15, -52, 7, -9, 9, 10, -49, 23, 23, -2, 17, 11, -2, -28, -26, 4, 13, 10, -18, 16, -43, -8, 4, 13, -24, 2, 27, -6, 13, 3, 6, -8, -2, -3, 0, -52, -30, 1, -11, 52, 2, -3, -31, -32, 5, -28, 10, 4, 33, 5, 14, -23, 53, -37, 0, -16, 2, -9, -5, -14, -44, -8, 10, -6, -10, -21, -12, -9, -9, -17, -14, 42, -15, -35, -16, -18, 0, 7, 23, -20, 12, -55, -45, -7, -7, 1, -18, 8, 9, -1, 1, 5, 7, 13, 20, -13, 12, 9, -6, 1, 1, -39, 9, -10, -47, 9, 0, -34, 6, -1, -74, -61, -11, 0, -3, 39, 2, 30, 19, 8, 12, 10, -2, -9, 32, -12, -20, -6, -2, -2, 27, -3, -36, -7, 26, -2, -36, -3, -43, -12, 25, -10, -2, 1, -28, 16, 16, 40, 0, -6, 35, -38, 37, -4, -4, -19, -36, 29, -3, -30, -22, -7, 9, -3, 19, 7, -29, -7, -11, 5, 0, 17, -12, -10, -8, -23, -35, -15, 9, -2, 24, 0, -29, -12, 0, -5, 45, 1, 23, -2, 12, 31, -23, 8, 2, 25, 10, -4, -2, 16, -7, 0, 9, 9, -46, -7, 3, 8, 8, 9, 6, 2, 36, -3, -2, -19, -1, -2, 8, 0, -18, 20, 17, -57, -7, -12, -5, 3, -22, 1, 44, -12, -17, 7, -5, 9, -88, -12, -60, 4, -23, -27, 38, 5, -29, 17, -7, -15, 23, -5, 16, 3, 10, -41, -14, 11, 11, 17, -13, -27, -3, -2, 11, -8, -14, -8, -16, -63, -80, -46, 4, -4, 6, -6, -3, -1, -7, 43, 28, -60, -21, 0, 33, -18, -12, 1, 8, -23, 0, 18, 0, -25, -16, -4, 3, 1, 7, -9, 0, -49, -52, -19, 13, 0, -37, 3, -38, 7, -41, -25, -18, 25, 58, -31, -11, -22, -40, -62, 0, -7, -9, -3, 3, 13, -3, 20, -56, 25, 38, 15, 1, 13, 21, -13, 7, 14, -3, -8, 5, 18, -4, 0, 34, 4, 1, 15, 0, -27, -2, 31, -50, 8, 2, -47, -8, 8, 53, 32, -1, -1, -4, 17, -14, 39, -9, 15, -8, -2, -2, -3, 8, 45, 2, -10, -24, -33, -32, 5, 1, 14, -47, 4, 0, -14, 10, -14, 2, -55, -18, -3, -13, -13, -3, 9, -70, -27, 8, -31, 2, 11, 30, 19, 21, 19, 26, -2, -18, 11, 13, -7, -6, 33, -3, -27, 1, -19, -4, 22, 7, -8, 7, -1, 18, -40, 8, 0, 0, -28, 29, -9, 10, 4, 57, 1, -13, -6, -43, 3, -4, 6, -8, -4, 15, 7, 39, 2, -49, 71, -3, -32, 0, 2, 10, 0, 5, 10, -4, -15, -59, 3, -53, 0, -8, 9, -30, -11, 5, 34, 7, -2, 46, 25, -2, 6, 16, -4, 26, 18, 18, 8, -9, 0, 7, -9, 13, -18, 42, 14, -8, 4, 9, -8, 38, 4, -25, -4, 45, 0, 36, 19, -5, 7, 4, -8, -10, 1, 48, 11, -7, 18, -6, -26, -21, 29, -18, 6, 1, 5, 29, 25, -16, -9, 62, -21, -15, -27, -31, 0, -9, 7, -16, -7, -5, -15, 0, -28, 12, -7, 52, 57, -31, -4, 17, -10, -1, -15, 11, 17, -14, -7, -29, -15, 1, 0, -24, 33, -21, -14, 0, -6, -1, -9, -5, -3, 4, -22, -38, -6, -8, -15, 9, -28, -37, 15, 0, 9, 3, 0, -11, -4, 11, 12, 20, 16, -3, 56, -31, 27, 9, 5, -7, -3, 55, 32, -28, 20, 7, 18, -6, -2, 4, 20, 2, -28, 11, 7, -6, 4, 19, 20, 12, 7, 21, 33, -7, -12, -6, 17, 6, 10, 5, -11, 34, -2, 1, 9, -16, 14, 11, -32, -14, 11, -40, 22, -3, -10, 5, 16, -3, 5, 2, -33, 14, -3, 22, 2, -24, 13, 53, 3, 15, 8, -38, -33, -45, 3, 8, 18, 39, 30, 10, -13, -9, -2, 42, -6, 0, 5, -10, -1, 6, -41, -26, 64, -9, 2, 15, 4, -3, -22, 16, -2, -2, -18, -1, -14, 5, -8, 38, -14, -5, -10, 47, 10, -6, -26, 0, -10, -27, -1, 26, 1, -13, 15, 24, 9, 13, -29, -1, 0, -18, -31, -3, 5, -49, 3, -24, -9, 15, 3, -11, -8, 4, 21, 1, -13, 2, 2, -1, 25, 12, 5, 1, 2, 1, -15, -22, 25, -13, 0, 9, -5, -17, 27, -18, 12, 2, -45, -11, 15, -6, 4, -9, 16, 31, 39, -28, -24, 0, -35, 25, 0, -2, -7, -31, -4, -26, 1, 1, -56, 7, -4, 11, 7, -1, 26, 16, -2, 14, 21, -8, -36, -11, 6, 23, 5, -20, -18, -17, 10, -16, -10, -15, 4, 12, -1, -6, -10, 37, 38, -4, 1, -8, -79, -15, 10, -19, -10, 1, 4, 20, 32, 8, -15, 44, 6, -52, 3, 16, -7, 38, -20, -24, -39, 23, 4, -8, -46, -43, 0, -8, 1, -22, 14, 9, -9, 0, -43, -2, 8, -13, -76, 11, -41, 3, -1, 7, -68, 26, 0, 17, 22, -6, -10, -46, 7, 12, 30, -51, -37, -13, 19, 4, -4, -42, 9, 0, -22, -68, -57, 0, 2, -49, -9, 5, -33, 0, -9, 24, -9, 7, 3, 0, -43, 6, -2, 73, 19, -57, 14, -6, -2, -28, -47, -7, 13, -53, -2, 8, 0, 23, -11, -27, 13, 6, -6, -22, 17, 0, 32, -68, -14, -24, 1, 0, 31, 16, 20, 11, 9, 13, 8, -15, 0, -21, 52, -3, 44, -16, -47, -9, 4, -27, -2, -23, -4, -10, 10, -10, 4, -44, 32, 0, -53, -50, -46, 10, 3, -35, 1, -20, -9, 8, 2, -43, -12, 17, -12, 56, -30, 9, 14, -7, 22, 9, -4, 8, -46, 3, -8, -75, 0, 19, 8, 12, 8, 5, -6, 4, 18, -29, -16, 1, -44, -4, 20, -4, -32, 35, 20, 17, -40, -19, -3, 6, 0, -59, 2, -16, 36, 15, 0, -3, 0, -47, 8, -60, 10, -37, 33, -20, -14, -13, 22, -51, 0, -32, 3, -42, -6, -8, 10, -12, 38, -25, -36, -7, 4, 0, -6, -35, 27, -3, -20, -1, -40, -17, -25, -35, 15, 10, -1, -19, -51, 31, 6, 39, -30, 13, -13, -19, -19, 35, 1, -7, 6, -4, 15, 8, 26, -22, 35, 27, -24, 6, -10, -51, 9, 21, -41, 20, -4, 10, -54, -5, -7, 5, 24, -18, 11, 85, -15, 5, -12, -16, -13, -7, 6, 15, 2, 1, -3, -10, 7, 17, 0, 8, -13, -44, -31, 7, -6, 1, -2, 32, 24, 4, -20, -14, -64, -18, -6, -2, 42, 32, 2, -4, -11, 72, 10, 11, -3, 7, 6, -2, -26, 6, 0, 6, -17, 3, -29, -1, 8, -51, -32, 9, 11, 8, -21, 8, 30, 46, 12, -2, -11, 2, 14, -7, -27, -9, -4, -47, 14, -9, -13, -33, 0, -4, -8, -9, 7, 2, -5, -8, -3, -42, -6, -41, 3, -35, 11, 3, 18, -44, 22, -2, -8, -9, 11, 59, 5, -5, 15, -7, 14, 2, -6, 25, 6, 31, 29, -9, -2, -2, 5, -7, 2, 0, -13, -32, 5, -10, 0, 4, -7, -4, -52, -7, -6, -9, 3, -16, -12, 23, -10, -16, -10, 6, -19, -8, 2, 4, -3, 28, -14, -46, -5, -34, -2, -18, 5, 6, 2, 10, -1, -45, -3, -20, 20, 1, 20, -4, 1, 1, -36, 16, -8, -7, -22, -7, 4, -16, 4, -4, -6, -3, -4, 4, 4, -25, -6, -44, -7, 4, -6, -43, -31, -7, 63, -11, -37, -21, 1, -10, -3, 12, 22, -11, 38, 0, -4, -15, -6, -14, -4, 3, -25, -30, -15, 20, 3, -31, -14, -49, 6, -2, 12, -13, 0, -32, -13, 47, -13, -27, 10, -8, -69, -10, 7, 8, 2, 2, 17, 0, 0, 25, 13, 28, -20, 7, -5, 17, 13, 37, 50, -8, 9, -31, -11, 24, 0, 7, 17, 3, 22, -1, -28, 1, -45, 9, 6, 7, 1, -12, -8, 0, -17, -1, 9, 0, -57, -19, -44, -39, -2, 15, -1, 10, -5, 35, 20, 36, -20, 4, -45, -30, -2, -9, 67, 17, -64, -2, -26, -2, 10, -14, -42, -6, -1, 20, 9, -6, -8, -15, -42, 0, -31, -13, -6, 10, -18, -5, 13, -5, -10, -2, 27, 50, 41, -10, 10, -7, -21, 11, -39, -13, -19, -7, 0, -20, -19, -7, 1, -15, 7, 52, -13, -1, 37, -12, -5, -42, 3, -21, -6, -44, 42, 11, 11, -10, 6, -7, -9, 7, 22, 27, 29, 11, -1, 13, 19, -7, 7, -15, -7, 34, 3, 12, -10, -4, -22, 2, 21, -6, 45, -63, 18, -9, 1, 24, -8, -5, 17, 9, 5, -40, -6, 0, 0, 0, -7, 0, 21, -3, 1, -1, -19, 9, 3, -44, 22, -21, -13, -18, -2, 5, -10, 16, 3, 9, 5, 0, -7, -24, 7, -1, 34, -23, 17, 54, -16, -1, -81, 2, 39, -7, 9, -22, -5, -26, 23, -5, -12, -6, -34, -28, -11, -10, -5, -17, -55, 2, -29, -35, 36, -1, -67, -3, 0, 0, -8, 17, -4, -9, 19, -25, -32, -4, -29, -6, -12, 47, 10, -34, -15, -53, 2, -27, -13, -46, -4, -21, 9, -42, -17, 26, -44, 24, -7, 13, -11, -40, -74, 3, -6,

    others => 0);
end iwght_package;
