library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    68, 68, 63, 65, 63, 66, 66, 68, 65, 67, 57, 53, 46, 46, 45, 
    55, 64, 67, 68, 69, 63, 54, 65, 61, 39, 19, 22, 40, 50, 46, 
    66, 66, 72, 67, 80, 134, 56, 33, 20, 58, 56, 18, 10, 33, 45, 
    2, 28, 68, 69, 64, 51, 49, 22, 21, 94, 43, 56, 19, 0, 44, 
    19, 63, 52, 80, 59, 51, 58, 21, 21, 47, 60, 19, 20, 0, 17, 
    78, 103, 50, 114, 178, 101, 67, 31, 0, 99, 85, 28, 41, 8, 0, 
    57, 102, 65, 44, 103, 104, 127, 51, 19, 124, 70, 27, 29, 40, 18, 
    85, 76, 27, 36, 77, 163, 77, 82, 34, 120, 77, 36, 44, 60, 24, 
    102, 121, 44, 70, 64, 94, 61, 54, 38, 60, 114, 20, 33, 36, 55, 
    133, 130, 45, 79, 63, 29, 48, 62, 54, 73, 12, 0, 9, 54, 59, 
    144, 124, 59, 124, 31, 39, 109, 109, 25, 0, 0, 0, 24, 60, 57, 
    140, 125, 72, 190, 185, 80, 76, 71, 39, 32, 30, 36, 36, 42, 37, 
    29, 115, 112, 205, 57, 26, 26, 24, 24, 24, 26, 34, 46, 47, 38, 
    29, 27, 149, 130, 42, 32, 21, 26, 26, 31, 42, 54, 35, 54, 75, 
    28, 30, 50, 79, 38, 50, 47, 24, 29, 31, 35, 29, 44, 54, 6, 
    
    -- channel=2
    1, 0, 0, 0, 0, 0, 0, 0, 0, 11, 24, 19, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 9, 40, 14, 0, 14, 47, 23, 0, 
    34, 46, 0, 0, 0, 68, 50, 68, 11, 0, 0, 0, 0, 42, 2, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 15, 0, 14, 14, 5, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 25, 
    11, 0, 0, 27, 108, 27, 0, 0, 0, 0, 0, 21, 0, 0, 0, 
    0, 0, 60, 0, 9, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 42, 7, 0, 1, 19, 6, 0, 0, 
    0, 0, 0, 0, 0, 82, 38, 0, 0, 8, 77, 54, 35, 0, 0, 
    3, 0, 0, 0, 3, 0, 0, 0, 0, 43, 30, 23, 0, 0, 2, 
    14, 0, 3, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 43, 49, 
    96, 35, 0, 0, 82, 142, 102, 103, 47, 13, 0, 3, 0, 0, 0, 
    0, 78, 20, 0, 108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 72, 60, 15, 0, 0, 0, 0, 0, 0, 18, 5, 0, 22, 
    0, 0, 15, 107, 32, 37, 22, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 
    4, 3, 0, 0, 0, 54, 5, 0, 0, 20, 34, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 12, 5, 0, 0, 0, 0, 0, 
    23, 45, 0, 4, 9, 24, 18, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 14, 0, 14, 52, 13, 0, 0, 0, 12, 4, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 4, 0, 0, 0, 0, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 6, 15, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 8, 45, 14, 0, 0, 0, 19, 34, 26, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 34, 20, 11, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 8, 17, 16, 7, 16, 18, 20, 0, 
    7, 15, 0, 0, 0, 0, 8, 16, 28, 0, 8, 8, 18, 14, 3, 
    34, 33, 0, 0, 27, 0, 1, 9, 24, 11, 14, 14, 21, 15, 13, 
    28, 43, 0, 0, 0, 0, 7, 0, 21, 23, 16, 23, 24, 20, 21, 
    26, 33, 2, 0, 0, 13, 18, 18, 15, 22, 12, 30, 26, 23, 0, 
    36, 44, 37, 9, 0, 11, 11, 17, 5, 0, 26, 17, 26, 0, 0, 
    34, 47, 38, 33, 28, 1, 0, 15, 35, 2, 6, 16, 11, 0, 0, 
    37, 31, 40, 37, 5, 27, 27, 32, 23, 16, 46, 46, 54, 31, 22, 
    109, 45, 24, 30, 59, 81, 92, 92, 91, 85, 97, 103, 114, 116, 114, 
    129, 105, 32, 54, 75, 96, 98, 97, 99, 105, 111, 117, 115, 110, 121, 
    137, 116, 95, 69, 78, 101, 100, 103, 101, 110, 122, 129, 122, 137, 142, 
    135, 131, 113, 109, 100, 111, 105, 97, 99, 111, 122, 119, 116, 140, 128, 
    
    -- channel=5
    55, 63, 62, 60, 56, 58, 65, 67, 57, 53, 57, 60, 58, 50, 46, 
    55, 62, 65, 64, 61, 45, 47, 64, 57, 11, 0, 0, 16, 46, 52, 
    55, 76, 62, 62, 57, 46, 23, 0, 0, 0, 0, 0, 0, 7, 47, 
    0, 4, 46, 60, 50, 33, 6, 3, 0, 11, 6, 0, 0, 0, 28, 
    0, 0, 41, 54, 52, 31, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 47, 27, 20, 29, 2, 0, 0, 4, 13, 0, 0, 0, 0, 
    0, 0, 28, 46, 21, 11, 22, 11, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 25, 10, 43, 39, 3, 7, 4, 0, 0, 0, 11, 19, 
    0, 0, 0, 0, 6, 0, 0, 0, 2, 0, 0, 12, 0, 1, 28, 
    2, 0, 0, 0, 0, 26, 5, 0, 0, 36, 19, 0, 5, 34, 47, 
    0, 0, 0, 0, 0, 0, 27, 30, 17, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 20, 35, 20, 6, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 23, 12, 23, 0, 9, 9, 0, 0, 
    64, 11, 0, 0, 21, 11, 7, 9, 4, 7, 21, 17, 13, 14, 0, 
    70, 16, 0, 0, 0, 6, 0, 16, 5, 31, 17, 12, 21, 23, 12, 
    71, 14, 0, 0, 0, 0, 28, 8, 25, 23, 23, 20, 13, 30, 8, 
    65, 45, 15, 0, 4, 45, 2, 0, 5, 0, 5, 13, 28, 3, 0, 
    68, 64, 40, 13, 0, 0, 0, 9, 15, 0, 18, 0, 0, 0, 0, 
    41, 54, 43, 38, 53, 5, 12, 39, 15, 6, 0, 30, 18, 0, 0, 
    55, 51, 37, 71, 65, 97, 79, 66, 61, 36, 80, 96, 88, 59, 67, 
    115, 70, 70, 48, 65, 78, 82, 85, 104, 113, 121, 125, 133, 131, 139, 
    142, 100, 66, 49, 92, 116, 117, 109, 116, 127, 138, 146, 142, 148, 156, 
    160, 135, 112, 54, 110, 120, 118, 120, 125, 134, 140, 146, 144, 172, 143, 
    152, 150, 113, 97, 108, 118, 122, 119, 126, 130, 138, 135, 155, 164, 148, 
    
    -- channel=7
    40, 42, 46, 45, 43, 41, 47, 49, 43, 27, 22, 26, 36, 41, 37, 
    44, 44, 43, 45, 40, 63, 53, 34, 17, 18, 25, 20, 16, 20, 32, 
    23, 12, 45, 49, 42, 12, 51, 20, 10, 3, 27, 27, 22, 0, 22, 
    41, 4, 41, 42, 46, 27, 31, 22, 13, 0, 55, 14, 25, 13, 0, 
    58, 15, 56, 9, 53, 54, 56, 45, 15, 0, 40, 42, 14, 21, 0, 
    55, 37, 73, 44, 14, 64, 79, 38, 36, 0, 64, 48, 2, 19, 23, 
    71, 47, 37, 52, 0, 45, 32, 60, 33, 0, 64, 40, 15, 12, 29, 
    74, 52, 42, 35, 0, 0, 69, 29, 36, 0, 56, 39, 0, 12, 43, 
    76, 37, 78, 18, 44, 18, 40, 26, 11, 36, 0, 33, 0, 23, 33, 
    57, 42, 72, 5, 30, 32, 29, 38, 30, 11, 21, 0, 0, 20, 37, 
    7, 46, 67, 1, 110, 28, 0, 25, 41, 20, 0, 0, 0, 0, 0, 
    0, 16, 47, 13, 57, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 23, 42, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 43, 11, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 5, 2, 3, 0, 0, 1, 7, 
    0, 0, 0, 0, 0, 0, 31, 0, 24, 0, 10, 1, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 61, 32, 3, 0, 8, 20, 28, 0, 0, 
    87, 0, 0, 0, 8, 0, 0, 34, 4, 0, 53, 0, 41, 23, 0, 
    120, 0, 49, 0, 0, 19, 43, 48, 12, 0, 1, 64, 0, 40, 0, 
    114, 0, 74, 9, 0, 45, 26, 38, 45, 0, 68, 94, 0, 30, 31, 
    131, 0, 13, 54, 0, 0, 0, 56, 59, 0, 93, 53, 0, 0, 22, 
    90, 10, 55, 20, 0, 0, 103, 3, 44, 0, 50, 56, 0, 0, 23, 
    70, 0, 135, 0, 40, 0, 26, 0, 0, 9, 0, 82, 0, 0, 0, 
    3, 0, 114, 0, 42, 33, 0, 0, 10, 12, 67, 11, 0, 0, 11, 
    0, 0, 99, 0, 107, 25, 0, 5, 91, 54, 0, 0, 0, 0, 20, 
    0, 0, 47, 0, 99, 101, 0, 0, 19, 0, 0, 0, 0, 0, 3, 
    12, 0, 0, 0, 194, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 0, 0, 37, 57, 0, 12, 0, 0, 0, 0, 0, 6, 0, 0, 
    36, 0, 0, 0, 14, 0, 0, 2, 0, 0, 3, 0, 0, 0, 58, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 0, 0, 4, 4, 2, 2, 0, 0, 
    0, 4, 0, 0, 0, 41, 0, 0, 0, 62, 30, 21, 1, 0, 5, 
    0, 29, 0, 0, 0, 8, 15, 0, 6, 73, 13, 20, 0, 0, 31, 
    5, 73, 0, 39, 58, 63, 34, 0, 0, 60, 43, 0, 12, 0, 5, 
    27, 73, 0, 7, 103, 59, 37, 17, 0, 107, 34, 0, 26, 3, 0, 
    27, 66, 7, 0, 78, 61, 67, 24, 0, 128, 22, 0, 18, 25, 1, 
    43, 72, 17, 0, 48, 106, 32, 39, 0, 97, 24, 0, 29, 31, 3, 
    62, 99, 0, 55, 1, 58, 17, 14, 33, 34, 22, 0, 15, 25, 12, 
    73, 93, 6, 99, 16, 15, 52, 51, 24, 6, 0, 0, 24, 27, 0, 
    105, 84, 20, 136, 40, 30, 89, 71, 1, 0, 3, 17, 36, 37, 10, 
    109, 98, 58, 170, 57, 8, 50, 46, 20, 28, 34, 45, 47, 51, 38, 
    35, 93, 100, 110, 0, 37, 38, 35, 30, 32, 44, 48, 52, 52, 60, 
    34, 46, 125, 52, 8, 47, 33, 36, 41, 45, 48, 50, 44, 56, 57, 
    37, 50, 53, 56, 19, 36, 38, 37, 49, 51, 40, 46, 73, 65, 22, 
    
    -- channel=10
    11, 13, 5, 7, 9, 0, 10, 14, 9, 20, 27, 18, 6, 4, 10, 
    2, 0, 5, 12, 2, 0, 0, 14, 53, 0, 0, 0, 0, 6, 7, 
    40, 38, 5, 8, 9, 57, 24, 0, 0, 0, 0, 0, 7, 0, 7, 
    0, 0, 0, 0, 4, 0, 0, 0, 3, 0, 13, 4, 9, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 28, 16, 0, 0, 0, 0, 0, 14, 12, 0, 0, 0, 
    0, 21, 0, 26, 8, 0, 14, 0, 5, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 69, 32, 0, 0, 14, 0, 0, 10, 6, 
    0, 0, 0, 0, 0, 29, 0, 0, 0, 8, 0, 59, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 50, 72, 0, 0, 0, 13, 
    0, 0, 8, 0, 0, 0, 0, 49, 31, 0, 0, 0, 0, 0, 0, 
    14, 2, 0, 0, 93, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 23, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 101, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 
    0, 0, 0, 17, 4, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    50, 54, 54, 57, 56, 54, 53, 53, 50, 41, 36, 37, 46, 44, 41, 
    53, 52, 55, 58, 59, 91, 61, 43, 28, 42, 53, 33, 24, 33, 44, 
    31, 38, 52, 56, 52, 56, 45, 28, 21, 64, 69, 69, 45, 17, 40, 
    58, 46, 53, 55, 52, 58, 68, 46, 45, 45, 79, 38, 38, 14, 23, 
    104, 94, 71, 73, 142, 109, 87, 51, 31, 43, 88, 58, 46, 38, 7, 
    90, 105, 81, 28, 66, 83, 104, 71, 50, 55, 103, 58, 45, 53, 36, 
    102, 95, 52, 46, 49, 83, 104, 93, 61, 72, 95, 55, 44, 52, 53, 
    106, 120, 74, 70, 52, 91, 112, 60, 57, 66, 86, 53, 38, 51, 57, 
    127, 116, 80, 70, 59, 52, 57, 55, 63, 67, 21, 38, 22, 50, 55, 
    119, 116, 99, 78, 66, 51, 78, 101, 58, 37, 39, 10, 35, 55, 57, 
    95, 111, 99, 108, 172, 93, 87, 98, 75, 49, 31, 42, 46, 60, 51, 
    54, 102, 118, 143, 110, 48, 37, 36, 40, 43, 48, 53, 62, 64, 61, 
    67, 47, 102, 129, 85, 54, 50, 47, 48, 50, 61, 65, 64, 64, 84, 
    68, 54, 49, 115, 60, 60, 59, 47, 49, 56, 60, 57, 62, 65, 64, 
    73, 57, 46, 53, 42, 35, 47, 58, 62, 71, 60, 60, 83, 97, 67, 
    
    -- channel=12
    61, 56, 61, 65, 66, 60, 61, 64, 65, 56, 42, 39, 49, 54, 52, 
    66, 59, 63, 65, 67, 97, 78, 47, 34, 48, 70, 50, 33, 38, 51, 
    34, 35, 61, 65, 66, 76, 53, 44, 31, 75, 82, 72, 67, 29, 39, 
    79, 60, 67, 67, 60, 67, 83, 58, 57, 58, 86, 55, 47, 30, 31, 
    118, 118, 82, 81, 134, 120, 92, 57, 43, 56, 106, 75, 56, 51, 24, 
    107, 112, 81, 53, 62, 82, 112, 86, 68, 65, 113, 64, 55, 63, 48, 
    112, 124, 54, 51, 71, 92, 115, 99, 73, 91, 108, 70, 62, 67, 66, 
    118, 126, 100, 76, 84, 90, 103, 69, 57, 83, 96, 69, 50, 58, 60, 
    139, 127, 97, 76, 74, 69, 74, 73, 72, 103, 37, 37, 28, 54, 64, 
    125, 132, 109, 103, 73, 53, 84, 120, 79, 29, 43, 21, 48, 72, 72, 
    108, 126, 115, 115, 190, 116, 93, 92, 74, 66, 52, 60, 71, 72, 64, 
    76, 98, 124, 174, 143, 61, 63, 56, 56, 59, 68, 74, 80, 91, 82, 
    99, 70, 103, 154, 83, 70, 70, 67, 72, 74, 86, 89, 89, 86, 104, 
    94, 80, 66, 113, 74, 82, 83, 68, 67, 75, 85, 80, 87, 87, 89, 
    95, 78, 79, 73, 68, 56, 62, 71, 83, 96, 87, 84, 106, 128, 94, 
    
    -- channel=13
    92, 92, 97, 100, 98, 90, 98, 102, 102, 89, 73, 70, 78, 87, 91, 
    95, 95, 99, 102, 97, 106, 103, 93, 65, 48, 54, 47, 43, 64, 89, 
    86, 53, 100, 102, 102, 52, 67, 39, 46, 23, 43, 32, 44, 34, 61, 
    79, 41, 92, 97, 103, 62, 73, 55, 36, 3, 49, 32, 33, 39, 22, 
    57, 46, 93, 62, 99, 72, 53, 53, 32, 0, 47, 61, 37, 46, 27, 
    38, 25, 90, 83, 0, 31, 65, 50, 56, 6, 58, 42, 24, 37, 42, 
    39, 34, 45, 100, 15, 46, 47, 53, 51, 0, 45, 46, 25, 31, 50, 
    44, 25, 45, 73, 43, 37, 47, 20, 45, 16, 42, 40, 17, 31, 46, 
    41, 14, 59, 19, 74, 0, 32, 49, 25, 41, 34, 28, 14, 36, 82, 
    27, 16, 53, 0, 51, 39, 16, 56, 43, 39, 27, 15, 24, 60, 81, 
    0, 23, 40, 3, 88, 72, 28, 14, 38, 24, 18, 21, 6, 7, 26, 
    0, 0, 31, 19, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 40, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=14
    100, 109, 109, 104, 105, 105, 110, 115, 104, 83, 78, 89, 92, 93, 88, 
    106, 112, 113, 108, 106, 120, 80, 97, 73, 57, 31, 39, 65, 80, 87, 
    79, 102, 109, 112, 112, 110, 61, 38, 26, 57, 11, 17, 18, 49, 92, 
    0, 98, 92, 110, 97, 71, 40, 15, 26, 55, 26, 31, 14, 22, 87, 
    0, 62, 65, 84, 54, 49, 27, 18, 26, 67, 23, 5, 28, 8, 59, 
    0, 51, 57, 104, 98, 37, 35, 11, 11, 99, 13, 0, 28, 10, 16, 
    0, 39, 54, 62, 102, 72, 30, 23, 0, 101, 0, 5, 30, 23, 15, 
    0, 6, 12, 39, 58, 63, 16, 35, 15, 96, 24, 4, 30, 40, 54, 
    0, 16, 0, 50, 34, 48, 25, 32, 35, 60, 34, 15, 47, 65, 87, 
    26, 20, 0, 53, 0, 38, 47, 16, 27, 27, 15, 8, 47, 90, 76, 
    50, 18, 0, 69, 0, 0, 35, 2, 0, 0, 0, 0, 0, 3, 0, 
    0, 19, 0, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 31, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 16, 0, 12, 3, 0, 0, 0, 
    13, 0, 0, 0, 0, 24, 25, 6, 0, 0, 39, 14, 22, 0, 0, 
    60, 0, 0, 0, 0, 0, 23, 5, 0, 0, 50, 17, 16, 0, 0, 
    80, 12, 9, 0, 59, 23, 70, 24, 10, 0, 45, 35, 0, 8, 0, 
    66, 62, 23, 0, 67, 59, 77, 35, 29, 0, 80, 46, 2, 8, 0, 
    52, 103, 23, 15, 0, 5, 104, 44, 61, 0, 92, 30, 0, 0, 8, 
    65, 101, 25, 26, 0, 48, 84, 43, 31, 0, 62, 41, 0, 10, 0, 
    95, 84, 70, 32, 0, 36, 42, 20, 0, 19, 35, 33, 0, 0, 0, 
    83, 76, 107, 9, 81, 0, 0, 68, 11, 35, 33, 0, 0, 0, 0, 
    59, 75, 108, 0, 111, 48, 32, 104, 81, 13, 0, 0, 14, 32, 43, 
    53, 64, 81, 37, 195, 91, 50, 47, 46, 22, 25, 26, 29, 34, 39, 
    41, 27, 12, 137, 120, 29, 33, 23, 22, 17, 21, 27, 44, 41, 33, 
    57, 33, 0, 167, 45, 23, 32, 27, 24, 27, 32, 44, 40, 26, 72, 
    57, 37, 30, 77, 27, 20, 32, 26, 21, 30, 40, 23, 13, 67, 68, 
    
    
    others => 0);
end ifmap_package;
