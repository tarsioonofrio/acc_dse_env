library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    158, 159, 165, 166, 160, 156, 162, 159, 158, 159, 161, 160, 161, 166, 169, 170, 167, 162, 160, 160, 156, 149, 150, 148, 149, 143, 140, 141, 143, 137, 126, 116, 
    152, 151, 159, 166, 162, 160, 164, 162, 163, 156, 155, 159, 163, 170, 171, 171, 169, 160, 154, 151, 145, 139, 140, 141, 149, 147, 145, 142, 143, 136, 125, 119, 
    151, 151, 158, 167, 160, 163, 165, 165, 163, 162, 158, 157, 161, 166, 167, 169, 170, 159, 145, 121, 110, 98, 101, 114, 120, 134, 143, 140, 142, 139, 130, 120, 
    155, 155, 160, 174, 167, 167, 169, 169, 165, 165, 167, 191, 177, 157, 162, 164, 158, 149, 104, 103, 98, 92, 80, 74, 86, 83, 113, 132, 140, 140, 136, 127, 
    155, 156, 161, 170, 169, 163, 169, 166, 164, 164, 173, 246, 195, 151, 146, 142, 111, 78, 85, 113, 112, 106, 97, 93, 74, 84, 85, 105, 128, 138, 133, 129, 
    148, 133, 130, 147, 161, 165, 167, 167, 163, 165, 163, 180, 157, 128, 97, 66, 69, 66, 89, 118, 122, 119, 114, 94, 99, 91, 58, 67, 108, 140, 138, 134, 
    127, 109, 47, 88, 153, 170, 168, 170, 169, 166, 164, 147, 129, 127, 100, 68, 78, 72, 83, 132, 146, 124, 105, 107, 115, 85, 63, 46, 79, 132, 141, 134, 
    131, 99, 42, 70, 143, 167, 165, 168, 171, 161, 140, 120, 130, 144, 116, 88, 91, 85, 77, 124, 163, 136, 102, 106, 100, 85, 54, 49, 57, 107, 138, 136, 
    170, 103, 54, 124, 153, 161, 163, 166, 165, 174, 113, 125, 157, 156, 121, 86, 82, 84, 80, 81, 138, 146, 113, 87, 83, 86, 71, 56, 40, 74, 133, 137, 
    180, 134, 94, 154, 174, 158, 156, 153, 207, 237, 207, 156, 174, 148, 125, 93, 86, 74, 59, 76, 137, 143, 133, 106, 86, 87, 84, 75, 50, 40, 95, 132, 
    183, 108, 142, 165, 177, 155, 159, 122, 213, 237, 220, 164, 183, 156, 125, 120, 78, 80, 45, 91, 175, 157, 155, 107, 87, 103, 88, 78, 59, 41, 59, 104, 
    188, 100, 135, 170, 187, 166, 173, 134, 117, 194, 199, 170, 185, 189, 134, 117, 102, 84, 38, 125, 210, 160, 146, 93, 83, 94, 104, 85, 73, 55, 62, 76, 
    189, 90, 127, 175, 174, 166, 178, 159, 97, 168, 168, 137, 186, 216, 160, 123, 120, 115, 50, 150, 194, 155, 123, 91, 84, 84, 95, 86, 84, 73, 79, 73, 
    189, 93, 152, 185, 119, 136, 173, 167, 103, 147, 145, 167, 189, 226, 180, 141, 126, 117, 71, 154, 186, 149, 114, 87, 80, 72, 80, 99, 100, 90, 97, 94, 
    194, 108, 168, 186, 105, 99, 156, 167, 100, 115, 138, 198, 190, 172, 145, 154, 146, 103, 71, 152, 179, 137, 130, 110, 85, 91, 95, 109, 115, 100, 97, 117, 
    197, 132, 172, 184, 130, 78, 140, 155, 115, 130, 143, 230, 242, 145, 135, 131, 121, 108, 95, 144, 168, 152, 112, 87, 71, 87, 105, 112, 120, 103, 121, 136, 
    203, 146, 168, 191, 168, 78, 126, 138, 138, 96, 154, 173, 162, 140, 113, 113, 101, 105, 112, 171, 156, 148, 135, 109, 78, 79, 94, 101, 107, 125, 151, 144, 
    214, 163, 164, 183, 176, 94, 96, 156, 148, 106, 129, 118, 114, 116, 102, 115, 86, 101, 144, 118, 68, 128, 133, 75, 60, 58, 71, 102, 116, 143, 150, 140, 
    212, 178, 167, 173, 176, 124, 86, 141, 153, 135, 104, 77, 134, 124, 129, 147, 85, 92, 150, 132, 117, 107, 75, 64, 44, 65, 86, 133, 155, 160, 154, 151, 
    199, 187, 171, 174, 177, 144, 86, 119, 122, 137, 144, 70, 129, 108, 145, 184, 116, 73, 131, 137, 134, 89, 51, 52, 47, 90, 121, 163, 171, 164, 158, 149, 
    165, 195, 179, 177, 181, 152, 99, 131, 171, 103, 93, 80, 93, 122, 178, 191, 150, 100, 89, 87, 60, 46, 38, 24, 46, 60, 108, 144, 144, 128, 127, 120, 
    117, 195, 177, 178, 181, 138, 83, 150, 245, 219, 133, 134, 149, 176, 190, 194, 168, 125, 110, 61, 35, 34, 49, 58, 61, 58, 69, 72, 78, 69, 59, 55, 
    79, 175, 174, 176, 177, 140, 109, 211, 253, 252, 208, 124, 114, 124, 116, 122, 104, 68, 68, 60, 52, 50, 51, 56, 56, 51, 43, 51, 59, 48, 43, 42, 
    41, 96, 144, 168, 178, 165, 165, 246, 253, 227, 110, 60, 53, 49, 49, 48, 45, 42, 46, 42, 38, 46, 46, 43, 42, 46, 46, 50, 55, 53, 51, 45, 
    29, 29, 59, 131, 166, 132, 194, 254, 241, 141, 61, 50, 50, 51, 49, 50, 47, 42, 39, 34, 35, 39, 38, 42, 45, 56, 62, 59, 56, 50, 46, 51, 
    48, 30, 34, 73, 128, 128, 215, 256, 187, 66, 54, 50, 52, 52, 46, 45, 43, 41, 36, 39, 40, 40, 43, 46, 59, 62, 64, 59, 54, 50, 70, 83, 
    52, 35, 31, 41, 66, 128, 224, 240, 124, 58, 49, 56, 54, 44, 44, 47, 46, 43, 43, 44, 44, 45, 54, 58, 54, 46, 43, 36, 51, 73, 85, 76, 
    50, 35, 29, 35, 44, 78, 202, 211, 97, 65, 54, 48, 58, 48, 40, 45, 47, 48, 47, 46, 51, 39, 39, 48, 47, 39, 28, 40, 67, 67, 46, 51, 
    50, 35, 32, 33, 41, 46, 104, 170, 64, 54, 52, 53, 61, 58, 54, 45, 42, 41, 46, 49, 46, 42, 40, 39, 37, 40, 44, 63, 47, 31, 15, 51, 
    68, 42, 31, 38, 37, 43, 42, 71, 49, 31, 27, 38, 49, 56, 58, 53, 56, 60, 57, 53, 50, 45, 39, 33, 42, 62, 79, 73, 56, 38, 13, 40, 
    61, 49, 35, 43, 39, 42, 44, 40, 42, 27, 23, 30, 27, 29, 36, 47, 56, 62, 66, 75, 69, 49, 43, 43, 60, 85, 109, 93, 60, 26, 29, 20, 
    54, 56, 45, 43, 40, 40, 40, 38, 36, 26, 22, 29, 25, 29, 19, 18, 32, 47, 61, 74, 66, 53, 52, 45, 67, 89, 105, 89, 48, 24, 34, 21, 
    
    -- channel=1
    112, 111, 116, 118, 112, 109, 115, 113, 111, 113, 116, 111, 111, 117, 117, 119, 117, 113, 111, 112, 109, 107, 107, 106, 107, 101, 98, 97, 97, 95, 91, 85, 
    112, 110, 114, 116, 112, 113, 117, 114, 116, 110, 111, 110, 113, 119, 117, 115, 115, 111, 112, 115, 110, 104, 102, 100, 105, 102, 102, 97, 98, 95, 91, 88, 
    110, 109, 111, 111, 106, 115, 117, 117, 115, 115, 114, 109, 111, 115, 114, 113, 116, 114, 111, 96, 90, 78, 77, 85, 86, 96, 103, 99, 99, 98, 95, 89, 
    107, 110, 109, 112, 110, 117, 120, 119, 115, 117, 123, 146, 130, 111, 115, 114, 112, 111, 80, 87, 90, 90, 75, 63, 70, 62, 85, 98, 102, 101, 99, 94, 
    107, 114, 115, 114, 114, 113, 120, 116, 113, 116, 128, 214, 156, 114, 111, 108, 80, 53, 69, 103, 110, 114, 102, 94, 72, 78, 73, 83, 96, 101, 94, 93, 
    109, 104, 100, 112, 115, 113, 116, 115, 111, 116, 118, 138, 122, 102, 75, 50, 58, 56, 83, 113, 121, 122, 116, 96, 100, 91, 58, 58, 84, 105, 98, 95, 
    100, 95, 37, 74, 117, 118, 115, 118, 117, 116, 120, 107, 98, 108, 87, 67, 83, 75, 84, 130, 142, 118, 99, 102, 111, 83, 71, 47, 61, 98, 99, 93, 
    115, 96, 43, 64, 111, 117, 114, 116, 119, 113, 109, 94, 110, 131, 106, 87, 95, 88, 77, 118, 153, 124, 93, 98, 93, 81, 60, 53, 47, 83, 103, 97, 
    161, 105, 58, 121, 124, 113, 117, 122, 121, 135, 89, 105, 141, 143, 111, 80, 81, 85, 78, 71, 125, 135, 103, 79, 77, 82, 73, 57, 35, 59, 106, 103, 
    176, 139, 100, 154, 149, 116, 116, 118, 180, 214, 180, 131, 153, 131, 110, 85, 84, 74, 57, 68, 125, 133, 124, 98, 81, 85, 85, 76, 49, 30, 75, 103, 
    183, 116, 151, 169, 156, 112, 118, 89, 197, 224, 191, 135, 159, 137, 108, 111, 76, 80, 44, 85, 165, 147, 147, 100, 83, 102, 88, 79, 59, 36, 46, 81, 
    191, 108, 144, 175, 167, 120, 123, 93, 95, 182, 171, 142, 161, 171, 119, 107, 98, 84, 38, 121, 201, 152, 139, 89, 80, 93, 104, 87, 75, 53, 55, 56, 
    194, 96, 134, 180, 156, 123, 123, 109, 68, 154, 144, 114, 166, 202, 149, 113, 114, 114, 50, 147, 187, 149, 118, 88, 83, 84, 95, 87, 87, 73, 74, 55, 
    192, 95, 154, 188, 110, 106, 124, 116, 72, 132, 125, 149, 174, 216, 172, 131, 117, 114, 71, 152, 181, 144, 110, 85, 80, 73, 80, 100, 101, 88, 89, 73, 
    196, 107, 167, 186, 109, 89, 119, 122, 74, 106, 123, 185, 180, 165, 140, 143, 136, 100, 71, 152, 175, 133, 128, 109, 86, 93, 96, 110, 116, 96, 85, 95, 
    197, 129, 167, 178, 137, 83, 120, 125, 94, 120, 131, 221, 236, 138, 130, 121, 112, 104, 88, 134, 159, 147, 108, 85, 72, 88, 104, 109, 110, 86, 96, 104, 
    203, 146, 164, 182, 170, 86, 125, 126, 121, 80, 143, 163, 152, 132, 106, 106, 101, 101, 90, 143, 138, 141, 130, 105, 76, 79, 93, 91, 83, 88, 108, 104, 
    215, 166, 167, 184, 182, 102, 96, 149, 137, 93, 116, 105, 102, 105, 91, 110, 91, 103, 128, 96, 56, 120, 126, 69, 56, 56, 70, 93, 94, 112, 116, 110, 
    211, 184, 175, 181, 184, 131, 88, 139, 148, 128, 90, 64, 121, 111, 117, 143, 92, 96, 139, 117, 109, 99, 68, 59, 41, 62, 69, 105, 119, 120, 115, 111, 
    192, 189, 176, 179, 182, 149, 90, 121, 124, 136, 134, 59, 118, 97, 134, 176, 118, 75, 119, 124, 129, 86, 49, 51, 49, 90, 91, 118, 121, 113, 111, 107, 
    156, 193, 178, 173, 181, 157, 103, 135, 175, 105, 90, 77, 90, 118, 173, 182, 148, 100, 78, 77, 61, 52, 46, 33, 57, 71, 100, 125, 123, 109, 113, 105, 
    120, 200, 178, 169, 179, 144, 87, 153, 247, 222, 140, 141, 156, 182, 196, 192, 172, 133, 109, 62, 49, 54, 70, 81, 85, 84, 99, 101, 104, 96, 92, 90, 
    105, 197, 183, 172, 177, 146, 112, 211, 252, 253, 224, 143, 132, 141, 133, 133, 124, 93, 87, 82, 84, 84, 85, 93, 94, 91, 96, 104, 108, 97, 97, 95, 
    89, 137, 168, 174, 182, 170, 166, 245, 251, 231, 136, 88, 80, 76, 75, 72, 79, 81, 81, 82, 86, 90, 89, 87, 89, 93, 94, 96, 96, 94, 95, 90, 
    91, 87, 102, 153, 179, 136, 189, 250, 245, 159, 94, 84, 84, 85, 83, 84, 86, 84, 82, 79, 83, 86, 85, 89, 92, 103, 103, 101, 102, 99, 94, 103, 
    111, 94, 85, 106, 148, 136, 213, 253, 198, 93, 91, 88, 90, 90, 83, 82, 82, 81, 80, 83, 86, 89, 92, 95, 108, 110, 109, 108, 108, 105, 123, 137, 
    114, 99, 86, 83, 95, 145, 229, 245, 143, 92, 87, 94, 92, 82, 82, 83, 84, 83, 86, 88, 90, 97, 106, 110, 105, 97, 95, 91, 108, 130, 138, 125, 
    110, 98, 89, 86, 83, 106, 219, 228, 126, 104, 94, 87, 97, 87, 80, 82, 84, 87, 89, 89, 97, 92, 93, 102, 101, 93, 85, 101, 129, 126, 98, 96, 
    108, 97, 92, 88, 88, 84, 133, 197, 100, 97, 94, 95, 103, 100, 96, 83, 79, 80, 88, 92, 92, 95, 93, 92, 90, 93, 102, 125, 110, 90, 60, 93, 
    124, 100, 88, 91, 87, 89, 79, 107, 89, 77, 71, 82, 93, 100, 102, 92, 94, 99, 99, 97, 95, 94, 88, 83, 91, 112, 132, 131, 116, 97, 64, 85, 
    116, 102, 85, 91, 90, 92, 88, 81, 85, 72, 67, 74, 71, 73, 80, 86, 95, 101, 109, 119, 113, 95, 88, 88, 105, 130, 156, 145, 115, 82, 82, 64, 
    107, 105, 89, 86, 89, 92, 87, 81, 79, 69, 66, 73, 69, 73, 63, 58, 70, 87, 104, 119, 111, 96, 95, 87, 109, 131, 146, 135, 99, 77, 84, 67, 
    
    -- channel=2
    49, 47, 51, 53, 46, 41, 47, 45, 44, 41, 41, 52, 49, 41, 45, 44, 40, 38, 39, 43, 44, 45, 45, 43, 44, 39, 43, 41, 38, 36, 36, 33, 
    51, 40, 45, 56, 49, 43, 47, 45, 46, 38, 41, 54, 52, 41, 40, 33, 30, 33, 41, 50, 53, 55, 52, 48, 50, 46, 45, 38, 34, 31, 32, 34, 
    47, 33, 36, 48, 42, 44, 45, 45, 43, 43, 48, 57, 51, 38, 37, 35, 39, 47, 54, 49, 52, 50, 47, 50, 48, 55, 51, 39, 35, 34, 34, 33, 
    40, 32, 31, 44, 43, 46, 48, 48, 44, 45, 57, 95, 75, 41, 47, 54, 58, 67, 47, 65, 76, 84, 66, 50, 52, 39, 45, 46, 43, 39, 39, 36, 
    41, 48, 49, 47, 43, 40, 47, 44, 41, 42, 59, 164, 107, 56, 60, 71, 50, 31, 56, 98, 111, 118, 105, 93, 67, 70, 47, 45, 48, 46, 36, 36, 
    54, 64, 57, 53, 44, 39, 41, 41, 37, 39, 42, 85, 78, 58, 43, 31, 43, 45, 76, 110, 120, 122, 116, 96, 97, 86, 47, 37, 49, 58, 44, 40, 
    57, 80, 17, 28, 48, 43, 40, 43, 42, 37, 39, 52, 59, 75, 70, 57, 72, 64, 74, 121, 132, 108, 90, 94, 103, 77, 69, 39, 36, 58, 48, 39, 
    90, 92, 38, 41, 56, 42, 36, 39, 49, 51, 51, 49, 77, 107, 93, 79, 88, 82, 69, 107, 140, 112, 81, 88, 84, 74, 58, 49, 32, 50, 51, 39, 
    144, 105, 59, 113, 82, 43, 41, 50, 66, 95, 59, 78, 121, 128, 101, 74, 77, 82, 73, 61, 112, 123, 93, 70, 69, 76, 67, 53, 27, 35, 59, 45, 
    163, 143, 105, 149, 112, 51, 47, 60, 146, 198, 166, 119, 145, 125, 107, 79, 79, 71, 53, 58, 112, 122, 114, 89, 74, 78, 78, 71, 43, 15, 44, 57, 
    175, 122, 158, 168, 122, 50, 51, 47, 179, 226, 188, 131, 155, 132, 104, 104, 69, 77, 40, 77, 154, 137, 138, 92, 77, 96, 79, 73, 59, 33, 31, 46, 
    189, 116, 153, 178, 136, 59, 55, 44, 80, 188, 164, 133, 151, 159, 106, 95, 89, 79, 34, 113, 192, 142, 130, 82, 75, 88, 94, 81, 78, 55, 48, 26, 
    194, 105, 144, 185, 133, 68, 53, 47, 44, 152, 126, 94, 148, 183, 129, 98, 105, 109, 47, 140, 178, 140, 111, 83, 79, 80, 85, 81, 89, 73, 64, 24, 
    193, 103, 163, 192, 98, 66, 58, 50, 39, 120, 103, 127, 155, 200, 157, 117, 107, 109, 68, 147, 174, 136, 104, 80, 76, 70, 72, 94, 99, 81, 69, 34, 
    196, 112, 172, 188, 109, 67, 62, 55, 34, 88, 103, 169, 169, 159, 140, 134, 125, 95, 70, 149, 170, 127, 122, 105, 83, 91, 90, 104, 111, 80, 53, 47, 
    197, 136, 174, 181, 142, 77, 88, 77, 52, 93, 116, 211, 230, 137, 130, 112, 101, 95, 75, 118, 146, 138, 101, 80, 68, 87, 99, 99, 93, 54, 48, 48, 
    204, 160, 178, 188, 172, 90, 126, 113, 82, 37, 133, 155, 141, 117, 88, 90, 92, 87, 58, 104, 109, 126, 118, 97, 72, 77, 94, 82, 55, 45, 55, 46, 
    215, 180, 184, 194, 186, 105, 102, 145, 111, 61, 105, 95, 89, 89, 73, 98, 88, 95, 102, 64, 32, 105, 115, 61, 51, 53, 65, 78, 64, 68, 64, 54, 
    205, 192, 189, 193, 188, 133, 96, 143, 141, 111, 80, 55, 108, 96, 100, 133, 93, 93, 120, 93, 92, 86, 58, 52, 39, 60, 40, 59, 62, 54, 45, 46, 
    180, 187, 181, 185, 184, 152, 99, 132, 130, 135, 126, 51, 108, 86, 123, 168, 118, 73, 103, 105, 118, 78, 44, 50, 52, 93, 60, 68, 64, 52, 50, 46, 
    146, 187, 175, 172, 180, 160, 111, 146, 185, 111, 87, 73, 86, 116, 173, 177, 148, 101, 66, 63, 57, 54, 51, 41, 69, 83, 75, 82, 76, 61, 69, 63, 
    124, 200, 176, 168, 179, 147, 91, 159, 250, 225, 144, 147, 164, 192, 208, 197, 181, 143, 109, 62, 58, 68, 87, 102, 110, 111, 122, 119, 120, 112, 112, 115, 
    133, 213, 192, 177, 182, 150, 113, 209, 247, 252, 232, 157, 149, 162, 156, 152, 148, 119, 104, 101, 111, 110, 115, 125, 131, 130, 135, 141, 142, 132, 137, 132, 
    135, 168, 188, 188, 192, 174, 164, 237, 241, 228, 153, 111, 105, 105, 107, 101, 115, 120, 113, 116, 125, 125, 126, 128, 132, 139, 137, 137, 135, 134, 139, 133, 
    141, 130, 134, 176, 191, 137, 181, 242, 245, 175, 127, 118, 119, 121, 120, 116, 117, 117, 115, 113, 120, 125, 125, 130, 134, 145, 142, 142, 146, 144, 140, 149, 
    162, 140, 124, 136, 167, 143, 209, 249, 205, 118, 128, 125, 127, 127, 121, 115, 113, 112, 113, 117, 123, 131, 134, 138, 150, 152, 147, 149, 154, 152, 167, 182, 
    165, 147, 130, 122, 126, 164, 234, 247, 153, 114, 123, 131, 129, 119, 119, 119, 119, 119, 123, 127, 131, 141, 150, 154, 150, 141, 140, 138, 158, 178, 182, 169, 
    162, 149, 138, 133, 126, 138, 233, 234, 140, 126, 129, 124, 133, 123, 116, 119, 122, 126, 130, 132, 140, 138, 139, 148, 147, 139, 133, 153, 182, 176, 142, 139, 
    161, 147, 143, 141, 138, 125, 159, 211, 119, 121, 128, 130, 139, 135, 131, 120, 118, 120, 130, 135, 136, 139, 138, 136, 135, 138, 151, 178, 164, 140, 103, 136, 
    177, 148, 137, 146, 139, 132, 113, 133, 114, 105, 105, 117, 128, 135, 137, 128, 131, 137, 139, 138, 137, 136, 131, 125, 133, 154, 179, 181, 168, 146, 108, 127, 
    168, 148, 132, 143, 139, 134, 125, 112, 115, 104, 102, 109, 106, 108, 115, 120, 128, 135, 144, 156, 152, 134, 127, 127, 144, 170, 197, 190, 164, 130, 126, 107, 
    160, 149, 132, 134, 134, 132, 123, 115, 114, 105, 101, 108, 104, 108, 98, 89, 100, 118, 137, 152, 145, 131, 130, 123, 145, 167, 182, 175, 145, 124, 129, 110, 
    
    -- channel=3
    235, 231, 232, 232, 232, 232, 232, 232, 232, 232, 233, 233, 233, 233, 233, 233, 233, 232, 231, 230, 232, 232, 232, 233, 232, 233, 232, 232, 232, 233, 233, 232, 
    238, 235, 235, 235, 235, 235, 235, 235, 235, 235, 236, 236, 236, 236, 236, 236, 237, 236, 236, 234, 234, 234, 235, 236, 236, 236, 235, 235, 235, 236, 236, 235, 
    237, 234, 234, 234, 234, 234, 234, 234, 234, 234, 234, 234, 234, 234, 235, 235, 236, 236, 235, 234, 227, 231, 231, 234, 234, 234, 234, 234, 234, 235, 235, 234, 
    238, 235, 235, 235, 235, 235, 235, 235, 234, 234, 234, 234, 234, 234, 235, 235, 233, 232, 228, 223, 186, 209, 207, 228, 236, 234, 234, 234, 234, 235, 235, 235, 
    237, 234, 235, 235, 235, 235, 235, 235, 234, 234, 235, 235, 234, 234, 235, 235, 236, 233, 219, 203, 163, 195, 214, 230, 237, 235, 235, 235, 235, 236, 236, 236, 
    239, 236, 236, 236, 236, 236, 235, 235, 234, 235, 237, 237, 234, 232, 235, 229, 208, 194, 185, 174, 165, 184, 207, 226, 236, 236, 236, 236, 236, 237, 237, 237, 
    228, 228, 232, 231, 234, 237, 237, 236, 237, 237, 239, 239, 225, 224, 233, 221, 183, 161, 159, 154, 144, 143, 156, 198, 233, 236, 235, 235, 235, 236, 237, 239, 
    212, 224, 230, 227, 229, 234, 237, 238, 239, 239, 239, 240, 201, 219, 233, 214, 193, 185, 184, 173, 165, 159, 162, 186, 229, 234, 233, 233, 234, 236, 237, 238, 
    216, 221, 225, 225, 227, 231, 236, 238, 238, 238, 237, 239, 197, 220, 233, 230, 209, 209, 219, 208, 209, 210, 217, 218, 225, 228, 228, 230, 230, 235, 237, 238, 
    118, 119, 124, 136, 172, 225, 235, 237, 236, 235, 235, 233, 214, 226, 232, 236, 228, 227, 231, 225, 225, 217, 201, 185, 172, 167, 167, 186, 223, 235, 236, 238, 
    109, 103, 108, 111, 146, 222, 227, 229, 236, 234, 231, 230, 229, 231, 232, 230, 231, 231, 229, 223, 191, 164, 146, 137, 134, 128, 121, 149, 216, 234, 235, 237, 
    195, 188, 199, 200, 209, 223, 213, 211, 216, 220, 219, 210, 209, 211, 216, 220, 225, 226, 225, 218, 183, 175, 181, 178, 186, 170, 142, 185, 219, 231, 234, 236, 
    193, 191, 202, 214, 223, 214, 203, 171, 177, 207, 174, 98, 93, 101, 111, 122, 137, 153, 202, 223, 218, 220, 223, 217, 221, 212, 196, 222, 219, 221, 232, 235, 
    113, 111, 113, 125, 138, 170, 191, 190, 208, 216, 158, 54, 45, 49, 53, 66, 102, 159, 221, 234, 233, 227, 223, 207, 202, 211, 212, 199, 179, 188, 211, 221, 
    61, 69, 63, 68, 123, 139, 151, 195, 214, 206, 163, 103, 95, 101, 138, 181, 207, 221, 219, 205, 183, 158, 147, 131, 125, 130, 136, 133, 128, 138, 182, 197, 
    40, 58, 85, 127, 132, 96, 119, 163, 173, 184, 182, 181, 183, 198, 218, 200, 174, 159, 145, 132, 116, 98, 94, 99, 105, 107, 122, 138, 150, 157, 188, 185, 
    13, 26, 134, 206, 138, 118, 141, 172, 181, 207, 220, 228, 224, 230, 226, 176, 144, 138, 142, 145, 154, 149, 149, 154, 157, 160, 173, 187, 190, 178, 165, 157, 
    5, 58, 200, 225, 197, 199, 212, 226, 229, 233, 232, 230, 209, 223, 221, 210, 198, 180, 193, 188, 189, 194, 192, 184, 172, 171, 161, 144, 136, 131, 128, 138, 
    39, 145, 190, 186, 184, 192, 194, 194, 194, 191, 192, 190, 177, 180, 154, 147, 145, 156, 146, 113, 114, 132, 126, 111, 92, 91, 93, 94, 105, 121, 129, 129, 
    122, 162, 143, 137, 131, 128, 127, 130, 131, 128, 127, 129, 129, 124, 104, 100, 102, 118, 112, 94, 94, 94, 87, 83, 80, 83, 93, 101, 108, 115, 121, 130, 
    73, 76, 77, 80, 84, 87, 87, 90, 94, 102, 107, 113, 115, 118, 118, 120, 115, 110, 106, 100, 95, 85, 79, 80, 80, 77, 80, 82, 92, 113, 125, 136, 
    13, 3, 9, 18, 18, 21, 20, 22, 26, 34, 42, 48, 52, 60, 66, 70, 71, 72, 67, 60, 55, 53, 53, 57, 57, 57, 72, 87, 104, 120, 130, 137, 
    36, 11, 8, 32, 36, 22, 8, 3, 1, 0, 0, 0, 6, 5, 1, 3, 13, 24, 21, 21, 21, 22, 30, 39, 57, 85, 113, 123, 116, 122, 134, 153, 
    35, 26, 13, 27, 71, 70, 49, 27, 15, 5, 2, 0, 17, 57, 31, 10, 4, 4, 7, 14, 25, 41, 62, 86, 122, 144, 132, 114, 117, 132, 146, 172, 
    16, 13, 4, 3, 45, 65, 54, 36, 18, 4, 2, 0, 7, 118, 161, 131, 112, 105, 105, 109, 118, 138, 154, 151, 127, 105, 106, 120, 129, 142, 164, 184, 
    40, 12, 0, 0, 12, 30, 32, 21, 7, 2, 2, 3, 0, 68, 182, 205, 196, 194, 195, 187, 172, 150, 123, 103, 95, 104, 122, 129, 132, 152, 171, 185, 
    69, 26, 1, 1, 4, 12, 18, 12, 4, 2, 2, 4, 1, 32, 153, 203, 195, 191, 179, 155, 119, 91, 81, 94, 117, 125, 125, 129, 144, 162, 173, 184, 
    83, 47, 1, 2, 2, 5, 7, 4, 1, 1, 1, 3, 1, 27, 142, 205, 198, 169, 121, 85, 74, 85, 102, 121, 128, 122, 121, 132, 147, 165, 176, 186, 
    92, 54, 6, 3, 2, 1, 1, 1, 1, 1, 1, 1, 0, 15, 102, 157, 117, 74, 56, 74, 99, 115, 122, 124, 123, 125, 128, 136, 148, 162, 177, 188, 
    87, 43, 19, 11, 8, 5, 2, 2, 3, 3, 3, 2, 0, 4, 42, 71, 53, 57, 80, 113, 132, 134, 123, 116, 120, 131, 139, 143, 156, 169, 182, 188, 
    82, 46, 36, 31, 27, 22, 17, 16, 18, 19, 20, 19, 19, 23, 37, 64, 87, 104, 116, 128, 139, 131, 117, 115, 123, 131, 139, 148, 159, 174, 185, 187, 
    85, 62, 58, 55, 51, 47, 46, 48, 49, 51, 53, 55, 59, 68, 81, 104, 116, 127, 133, 127, 127, 118, 114, 122, 129, 136, 141, 149, 158, 168, 180, 186, 
    
    -- channel=4
    235, 231, 232, 232, 232, 232, 232, 232, 232, 232, 233, 233, 233, 233, 233, 232, 231, 231, 233, 233, 232, 231, 232, 233, 233, 233, 232, 232, 232, 233, 233, 232, 
    238, 235, 235, 235, 235, 235, 235, 235, 235, 235, 236, 236, 236, 236, 236, 236, 234, 234, 236, 236, 235, 234, 236, 236, 236, 236, 235, 235, 235, 236, 236, 235, 
    237, 234, 234, 234, 234, 234, 234, 234, 234, 234, 234, 234, 234, 234, 235, 234, 233, 234, 235, 235, 230, 235, 233, 234, 234, 234, 234, 234, 234, 235, 235, 234, 
    238, 235, 235, 235, 235, 235, 235, 235, 234, 234, 234, 234, 234, 234, 235, 235, 233, 232, 230, 226, 192, 216, 210, 228, 235, 234, 234, 234, 234, 235, 235, 235, 
    237, 234, 235, 235, 235, 235, 235, 235, 234, 234, 235, 235, 234, 234, 235, 235, 238, 237, 225, 210, 172, 205, 218, 229, 235, 235, 235, 235, 236, 236, 236, 236, 
    239, 235, 235, 235, 235, 235, 236, 235, 234, 235, 236, 236, 235, 233, 237, 231, 216, 205, 198, 188, 179, 196, 215, 228, 235, 236, 236, 236, 236, 237, 237, 237, 
    229, 227, 230, 228, 232, 236, 237, 237, 235, 235, 236, 237, 229, 228, 237, 226, 197, 180, 180, 176, 163, 159, 169, 206, 238, 237, 236, 235, 236, 238, 237, 237, 
    220, 230, 234, 232, 234, 237, 238, 237, 237, 237, 236, 238, 204, 222, 236, 218, 204, 201, 201, 191, 182, 174, 176, 199, 239, 239, 238, 238, 239, 239, 239, 238, 
    234, 236, 238, 239, 240, 238, 237, 236, 236, 236, 237, 239, 198, 221, 234, 231, 213, 216, 228, 218, 221, 224, 233, 235, 240, 238, 239, 240, 240, 240, 240, 238, 
    140, 138, 142, 155, 188, 234, 236, 234, 233, 235, 237, 237, 216, 228, 234, 237, 230, 230, 236, 232, 237, 233, 219, 204, 189, 179, 180, 199, 235, 241, 240, 240, 
    130, 121, 125, 127, 159, 229, 228, 226, 232, 234, 236, 237, 234, 235, 237, 235, 236, 237, 237, 232, 206, 184, 165, 156, 149, 140, 133, 162, 228, 241, 240, 240, 
    212, 202, 211, 211, 217, 227, 213, 209, 213, 222, 226, 221, 219, 221, 225, 229, 234, 236, 237, 231, 204, 198, 200, 194, 197, 178, 151, 195, 230, 240, 241, 240, 
    207, 202, 211, 217, 225, 219, 208, 174, 180, 213, 184, 112, 114, 121, 129, 138, 152, 167, 216, 236, 232, 233, 234, 226, 228, 219, 203, 230, 227, 230, 239, 241, 
    130, 125, 125, 131, 145, 182, 201, 199, 219, 230, 172, 71, 70, 73, 73, 84, 114, 168, 227, 239, 237, 231, 228, 211, 208, 218, 219, 206, 186, 197, 221, 231, 
    81, 86, 79, 85, 141, 155, 157, 200, 228, 223, 180, 121, 112, 117, 151, 192, 212, 222, 219, 203, 186, 166, 154, 138, 133, 139, 146, 142, 137, 153, 197, 212, 
    53, 70, 98, 144, 151, 107, 115, 158, 180, 194, 194, 193, 194, 209, 228, 210, 181, 165, 150, 136, 125, 111, 106, 111, 118, 121, 135, 151, 164, 174, 206, 203, 
    15, 29, 140, 216, 150, 123, 133, 162, 181, 209, 224, 234, 234, 241, 238, 189, 159, 154, 158, 163, 171, 165, 165, 171, 174, 177, 190, 204, 207, 196, 183, 175, 
    5, 62, 207, 232, 205, 207, 212, 224, 230, 236, 238, 238, 221, 238, 238, 228, 217, 200, 216, 213, 212, 214, 212, 204, 193, 191, 181, 165, 156, 146, 143, 154, 
    45, 155, 204, 196, 197, 211, 211, 208, 206, 203, 207, 207, 193, 198, 176, 169, 161, 171, 163, 133, 137, 157, 150, 135, 115, 112, 114, 116, 125, 133, 141, 142, 
    135, 179, 160, 154, 152, 152, 150, 150, 150, 147, 147, 149, 149, 145, 126, 122, 120, 134, 128, 109, 112, 117, 112, 103, 97, 103, 111, 117, 121, 125, 133, 144, 
    87, 90, 90, 93, 98, 102, 102, 105, 111, 119, 124, 131, 137, 136, 132, 133, 136, 133, 127, 119, 109, 101, 97, 92, 94, 100, 100, 98, 104, 119, 135, 149, 
    25, 11, 16, 26, 26, 25, 25, 30, 36, 43, 51, 59, 69, 75, 77, 79, 87, 88, 81, 72, 67, 68, 69, 69, 71, 78, 89, 100, 113, 124, 136, 146, 
    46, 16, 13, 44, 45, 25, 11, 8, 4, 2, 2, 4, 13, 18, 19, 23, 29, 38, 33, 31, 38, 44, 50, 58, 70, 90, 115, 123, 115, 123, 139, 160, 
    41, 27, 19, 41, 81, 70, 50, 31, 15, 5, 2, 0, 17, 64, 50, 36, 30, 30, 30, 35, 43, 55, 71, 97, 124, 131, 120, 105, 111, 134, 152, 179, 
    15, 10, 10, 12, 44, 52, 43, 33, 18, 4, 2, 1, 8, 117, 158, 128, 112, 105, 103, 105, 107, 115, 126, 126, 106, 86, 94, 116, 130, 147, 172, 194, 
    40, 10, 3, 4, 6, 12, 12, 10, 6, 1, 1, 2, 0, 58, 128, 130, 127, 123, 119, 113, 110, 96, 75, 66, 71, 93, 118, 132, 141, 162, 182, 197, 
    77, 29, 1, 1, 1, 2, 3, 2, 1, 0, 0, 0, 1, 12, 45, 47, 46, 48, 50, 49, 42, 38, 48, 77, 110, 126, 128, 135, 153, 176, 187, 198, 
    94, 52, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 2, 3, 25, 32, 25, 25, 25, 29, 41, 66, 92, 113, 124, 126, 127, 139, 157, 179, 191, 201, 
    102, 60, 7, 2, 2, 3, 3, 2, 1, 0, 0, 1, 3, 1, 19, 31, 17, 13, 27, 58, 90, 115, 126, 124, 123, 130, 135, 145, 159, 176, 192, 202, 
    99, 51, 23, 12, 10, 11, 10, 7, 4, 4, 4, 3, 6, 5, 13, 21, 27, 50, 77, 98, 113, 126, 126, 125, 128, 138, 148, 154, 168, 184, 197, 202, 
    96, 57, 44, 35, 30, 28, 26, 23, 21, 21, 22, 23, 27, 31, 40, 55, 70, 88, 102, 112, 121, 122, 122, 127, 133, 139, 149, 160, 172, 189, 200, 202, 
    101, 75, 67, 61, 56, 53, 53, 55, 55, 56, 58, 62, 67, 71, 84, 96, 103, 109, 116, 121, 127, 124, 125, 131, 136, 145, 152, 162, 171, 183, 195, 200, 
    
    -- channel=5
    235, 231, 232, 232, 232, 232, 232, 232, 232, 232, 233, 233, 233, 233, 233, 233, 233, 233, 233, 232, 234, 234, 232, 230, 231, 233, 232, 232, 232, 233, 233, 232, 
    238, 235, 235, 235, 235, 235, 235, 235, 235, 235, 236, 236, 236, 236, 236, 236, 233, 233, 234, 234, 237, 238, 237, 235, 234, 236, 235, 235, 235, 236, 236, 235, 
    237, 234, 234, 234, 234, 234, 234, 234, 234, 234, 234, 234, 234, 234, 235, 234, 231, 231, 234, 236, 233, 238, 235, 234, 234, 234, 234, 234, 234, 235, 235, 234, 
    238, 235, 235, 235, 235, 235, 235, 235, 234, 234, 234, 234, 234, 234, 235, 234, 230, 231, 232, 231, 197, 219, 213, 230, 235, 234, 234, 234, 234, 235, 235, 235, 
    237, 234, 235, 235, 235, 235, 235, 235, 234, 234, 235, 235, 234, 234, 235, 235, 236, 237, 230, 219, 179, 208, 221, 232, 237, 235, 235, 235, 236, 236, 236, 236, 
    238, 235, 235, 235, 235, 235, 235, 235, 234, 235, 236, 236, 236, 234, 237, 232, 218, 210, 207, 200, 189, 202, 220, 232, 237, 235, 235, 235, 236, 237, 237, 237, 
    229, 228, 231, 230, 233, 236, 235, 235, 236, 236, 237, 238, 230, 229, 238, 228, 204, 190, 191, 190, 177, 171, 177, 211, 239, 234, 233, 235, 236, 237, 237, 238, 
    222, 233, 238, 234, 234, 236, 235, 236, 238, 238, 237, 239, 203, 221, 235, 218, 210, 210, 211, 203, 196, 187, 185, 204, 240, 238, 237, 238, 238, 238, 238, 238, 
    241, 243, 246, 243, 240, 237, 235, 235, 237, 237, 237, 239, 196, 218, 231, 229, 217, 222, 235, 227, 234, 235, 240, 241, 243, 240, 240, 240, 239, 239, 239, 238, 
    149, 148, 153, 161, 191, 233, 233, 232, 234, 235, 236, 235, 214, 226, 232, 236, 232, 235, 241, 239, 247, 243, 226, 211, 195, 186, 185, 201, 235, 239, 239, 239, 
    141, 133, 137, 137, 165, 231, 225, 224, 233, 234, 234, 235, 235, 236, 238, 236, 238, 240, 241, 238, 213, 191, 172, 163, 159, 153, 143, 166, 229, 239, 238, 239, 
    224, 215, 224, 223, 227, 231, 211, 206, 214, 222, 225, 219, 223, 225, 230, 233, 237, 239, 241, 237, 208, 203, 207, 202, 211, 196, 164, 202, 233, 238, 239, 239, 
    222, 217, 224, 234, 241, 227, 208, 174, 183, 214, 188, 121, 126, 132, 139, 147, 161, 174, 220, 237, 235, 238, 240, 233, 237, 229, 212, 237, 234, 233, 242, 242, 
    152, 147, 141, 151, 165, 193, 205, 204, 226, 234, 183, 92, 91, 91, 90, 98, 129, 179, 233, 241, 241, 237, 233, 217, 212, 220, 223, 214, 196, 205, 227, 234, 
    108, 114, 100, 102, 155, 164, 164, 207, 234, 228, 190, 138, 131, 135, 168, 207, 223, 232, 227, 212, 195, 174, 163, 147, 140, 144, 152, 151, 147, 160, 203, 216, 
    77, 94, 116, 153, 156, 110, 118, 161, 182, 197, 198, 200, 202, 217, 236, 217, 186, 172, 159, 149, 138, 123, 118, 123, 128, 130, 145, 161, 174, 184, 213, 208, 
    35, 47, 151, 220, 150, 123, 134, 162, 180, 211, 225, 233, 232, 240, 238, 190, 163, 162, 170, 177, 187, 182, 182, 187, 189, 191, 204, 217, 218, 208, 193, 183, 
    24, 79, 217, 239, 212, 211, 218, 229, 237, 246, 245, 239, 220, 239, 241, 234, 228, 214, 230, 229, 231, 234, 232, 224, 212, 209, 197, 179, 169, 161, 158, 165, 
    71, 179, 222, 216, 217, 229, 230, 227, 227, 228, 228, 221, 207, 215, 193, 188, 184, 195, 186, 156, 161, 180, 173, 158, 138, 135, 133, 131, 140, 151, 158, 156, 
    161, 207, 194, 189, 187, 190, 192, 193, 192, 190, 189, 189, 188, 186, 163, 154, 154, 170, 163, 145, 148, 153, 144, 136, 130, 134, 139, 141, 144, 146, 148, 156, 
    109, 113, 122, 127, 134, 142, 147, 150, 152, 160, 165, 172, 181, 186, 180, 175, 172, 168, 163, 155, 148, 139, 132, 127, 129, 133, 129, 122, 126, 138, 146, 156, 
    41, 25, 35, 48, 52, 56, 58, 61, 62, 70, 77, 87, 106, 121, 126, 126, 127, 126, 120, 112, 106, 104, 103, 102, 105, 110, 115, 119, 128, 136, 141, 149, 
    55, 20, 19, 53, 58, 41, 30, 24, 17, 15, 15, 20, 42, 56, 60, 62, 71, 81, 77, 76, 78, 79, 83, 90, 101, 118, 138, 138, 125, 128, 137, 158, 
    45, 26, 18, 41, 84, 76, 57, 37, 21, 11, 7, 7, 35, 91, 78, 62, 60, 62, 63, 69, 74, 83, 99, 123, 146, 149, 135, 114, 116, 133, 146, 175, 
    17, 9, 8, 11, 46, 57, 47, 35, 20, 7, 4, 3, 15, 134, 179, 148, 131, 125, 124, 127, 126, 133, 144, 141, 116, 91, 97, 116, 129, 144, 165, 190, 
    35, 7, 3, 4, 7, 17, 17, 12, 7, 3, 2, 3, 2, 64, 146, 148, 144, 141, 137, 129, 122, 106, 83, 69, 70, 88, 113, 126, 135, 158, 176, 194, 
    64, 21, 1, 2, 0, 5, 9, 5, 2, 0, 0, 1, 1, 11, 59, 68, 67, 69, 67, 59, 49, 42, 46, 71, 102, 116, 120, 128, 147, 171, 183, 196, 
    82, 43, 1, 2, 0, 2, 5, 2, 0, 0, 0, 0, 0, 2, 38, 54, 46, 43, 36, 34, 39, 56, 82, 105, 115, 115, 118, 131, 150, 174, 187, 199, 
    93, 50, 3, 1, 0, 1, 3, 2, 1, 0, 0, 1, 2, 0, 28, 47, 23, 12, 22, 55, 81, 99, 111, 112, 113, 119, 126, 137, 151, 171, 188, 201, 
    89, 37, 11, 4, 2, 4, 4, 2, 1, 1, 1, 2, 6, 2, 13, 24, 25, 41, 62, 82, 101, 113, 112, 111, 115, 126, 137, 145, 161, 179, 193, 201, 
    82, 36, 22, 17, 15, 15, 13, 12, 12, 13, 14, 15, 20, 21, 27, 45, 67, 81, 85, 88, 105, 110, 107, 112, 119, 127, 138, 151, 164, 183, 196, 200, 
    83, 48, 38, 37, 35, 33, 34, 38, 40, 41, 44, 46, 45, 48, 59, 74, 83, 92, 97, 97, 107, 106, 108, 117, 123, 133, 141, 153, 163, 178, 191, 199, 
    
    -- channel=6
    158, 158, 139, 132, 166, 182, 187, 193, 199, 205, 209, 206, 218, 223, 227, 230, 213, 226, 231, 235, 236, 232, 234, 234, 236, 226, 230, 238, 232, 228, 237, 238, 
    170, 172, 151, 137, 174, 193, 197, 199, 206, 215, 217, 210, 225, 231, 233, 237, 219, 228, 232, 242, 245, 234, 236, 242, 241, 228, 235, 243, 233, 232, 246, 246, 
    174, 176, 157, 142, 181, 201, 206, 199, 209, 223, 218, 212, 224, 230, 230, 239, 221, 228, 233, 239, 232, 213, 236, 243, 245, 231, 238, 248, 237, 230, 250, 245, 
    180, 178, 160, 147, 186, 203, 212, 207, 214, 228, 221, 214, 220, 231, 223, 240, 224, 228, 233, 228, 177, 172, 230, 243, 248, 232, 238, 250, 238, 228, 249, 244, 
    186, 185, 165, 147, 189, 204, 217, 207, 211, 231, 222, 214, 218, 231, 211, 235, 226, 224, 232, 212, 159, 168, 224, 237, 247, 231, 235, 246, 232, 234, 248, 242, 
    193, 190, 170, 142, 191, 203, 219, 211, 215, 234, 221, 214, 214, 228, 199, 205, 207, 206, 235, 193, 112, 158, 222, 230, 245, 229, 226, 241, 228, 231, 243, 235, 
    196, 191, 172, 133, 191, 202, 222, 217, 223, 235, 218, 214, 215, 227, 188, 176, 187, 186, 205, 187, 120, 137, 172, 183, 219, 223, 216, 235, 226, 225, 240, 235, 
    204, 197, 174, 140, 203, 218, 224, 224, 232, 237, 220, 220, 220, 221, 201, 205, 172, 138, 100, 83, 71, 62, 65, 60, 104, 182, 209, 228, 218, 212, 239, 236, 
    175, 170, 157, 137, 176, 186, 175, 197, 209, 212, 206, 210, 212, 201, 193, 193, 142, 105, 89, 91, 84, 83, 94, 69, 78, 121, 162, 183, 174, 163, 207, 195, 
    114, 115, 113, 104, 105, 107, 111, 128, 139, 146, 151, 155, 157, 147, 151, 150, 118, 100, 99, 99, 85, 86, 86, 83, 139, 128, 154, 153, 118, 109, 132, 123, 
    66, 76, 75, 68, 83, 90, 84, 90, 93, 106, 102, 103, 106, 107, 114, 108, 90, 90, 91, 85, 72, 66, 95, 114, 128, 110, 147, 199, 125, 103, 92, 94, 
    53, 65, 75, 77, 111, 106, 85, 70, 93, 113, 95, 93, 108, 115, 107, 97, 98, 95, 98, 97, 90, 85, 149, 187, 179, 146, 112, 204, 154, 95, 87, 85, 
    58, 86, 94, 74, 100, 100, 77, 85, 120, 133, 127, 108, 105, 110, 98, 87, 81, 81, 87, 95, 95, 112, 170, 195, 208, 193, 127, 173, 178, 80, 85, 79, 
    74, 89, 87, 75, 82, 68, 71, 80, 89, 103, 118, 111, 101, 106, 105, 98, 96, 98, 98, 109, 114, 142, 180, 184, 191, 192, 160, 132, 170, 80, 60, 67, 
    77, 79, 82, 78, 79, 72, 70, 86, 109, 121, 129, 133, 137, 136, 135, 131, 146, 148, 146, 150, 148, 163, 179, 181, 185, 176, 170, 101, 90, 73, 55, 59, 
    96, 94, 106, 104, 109, 131, 132, 138, 144, 152, 155, 154, 155, 155, 158, 148, 150, 157, 156, 146, 119, 130, 146, 169, 177, 168, 167, 105, 69, 98, 86, 72, 
    106, 101, 115, 131, 129, 135, 144, 143, 146, 150, 154, 154, 154, 153, 151, 144, 130, 134, 139, 127, 94, 117, 146, 159, 167, 163, 162, 132, 144, 192, 154, 105, 
    95, 108, 118, 109, 95, 93, 129, 145, 149, 151, 150, 144, 134, 126, 122, 123, 122, 133, 155, 148, 131, 147, 162, 156, 157, 151, 153, 149, 159, 164, 157, 148, 
    102, 89, 73, 70, 86, 111, 123, 140, 143, 129, 120, 117, 120, 126, 133, 141, 150, 142, 153, 159, 151, 157, 165, 161, 153, 152, 154, 144, 131, 121, 125, 149, 
    86, 61, 71, 110, 128, 138, 130, 123, 118, 108, 118, 132, 143, 152, 156, 153, 149, 137, 145, 154, 153, 154, 160, 164, 152, 144, 125, 105, 92, 75, 86, 132, 
    104, 103, 107, 114, 115, 116, 123, 118, 116, 134, 141, 144, 143, 141, 133, 117, 98, 89, 130, 150, 151, 154, 152, 145, 117, 96, 90, 80, 65, 71, 73, 65, 
    99, 107, 111, 111, 114, 119, 125, 126, 117, 125, 125, 129, 131, 130, 91, 61, 57, 56, 115, 148, 139, 130, 114, 95, 86, 83, 73, 58, 60, 75, 51, 27, 
    62, 104, 116, 114, 116, 117, 102, 91, 84, 81, 78, 112, 133, 130, 96, 76, 83, 86, 107, 108, 96, 88, 83, 81, 70, 61, 51, 45, 52, 46, 30, 24, 
    57, 96, 106, 105, 107, 104, 65, 53, 59, 64, 68, 110, 135, 133, 115, 98, 88, 79, 78, 80, 81, 80, 70, 55, 44, 49, 45, 41, 34, 30, 27, 24, 
    65, 90, 104, 105, 109, 109, 79, 73, 85, 88, 98, 106, 98, 83, 68, 65, 70, 74, 81, 82, 72, 51, 41, 44, 61, 55, 39, 35, 32, 30, 27, 25, 
    67, 87, 105, 103, 102, 99, 88, 81, 76, 69, 59, 57, 58, 63, 66, 70, 72, 68, 62, 54, 46, 47, 49, 44, 56, 46, 30, 28, 29, 25, 24, 30, 
    54, 58, 65, 58, 55, 50, 45, 44, 46, 51, 55, 58, 62, 64, 62, 58, 51, 38, 37, 48, 49, 48, 42, 38, 41, 32, 27, 28, 27, 25, 28, 31, 
    30, 29, 26, 27, 31, 32, 33, 39, 49, 52, 53, 51, 46, 40, 38, 40, 38, 44, 66, 55, 41, 37, 36, 37, 31, 27, 26, 27, 28, 30, 33, 23, 
    33, 31, 27, 28, 28, 30, 31, 32, 35, 33, 30, 30, 34, 39, 41, 45, 42, 52, 73, 49, 30, 35, 38, 32, 27, 26, 27, 29, 30, 38, 26, 13, 
    31, 30, 26, 26, 25, 25, 26, 27, 29, 32, 37, 40, 42, 41, 40, 42, 39, 46, 64, 38, 28, 36, 30, 29, 26, 25, 27, 28, 33, 37, 9, 4, 
    23, 27, 25, 28, 30, 32, 34, 37, 39, 39, 40, 39, 38, 35, 30, 33, 28, 36, 57, 36, 30, 29, 29, 29, 24, 24, 23, 27, 36, 19, 4, 5, 
    28, 30, 32, 34, 33, 34, 35, 37, 38, 38, 36, 34, 30, 24, 15, 12, 8, 19, 45, 32, 25, 27, 27, 28, 24, 21, 20, 34, 25, 5, 4, 7, 
    
    -- channel=7
    190, 187, 166, 158, 193, 208, 211, 216, 219, 221, 222, 218, 229, 232, 235, 237, 220, 233, 238, 239, 241, 239, 241, 241, 242, 231, 235, 243, 237, 231, 239, 241, 
    200, 199, 176, 160, 199, 217, 218, 218, 223, 229, 229, 219, 233, 238, 239, 243, 225, 234, 238, 245, 247, 237, 239, 245, 245, 233, 239, 248, 236, 232, 246, 247, 
    201, 200, 179, 162, 201, 220, 223, 214, 221, 233, 226, 219, 229, 234, 234, 244, 226, 233, 238, 243, 235, 214, 234, 241, 247, 233, 240, 250, 238, 229, 249, 244, 
    203, 199, 179, 164, 201, 217, 225, 217, 223, 235, 227, 217, 221, 232, 226, 244, 228, 231, 237, 235, 184, 175, 228, 241, 248, 232, 238, 250, 237, 227, 247, 242, 
    207, 204, 181, 161, 201, 214, 225, 213, 215, 237, 226, 215, 217, 229, 212, 236, 227, 225, 236, 225, 170, 174, 224, 236, 247, 231, 235, 246, 231, 231, 245, 239, 
    208, 205, 183, 154, 201, 212, 226, 215, 218, 238, 223, 215, 215, 229, 199, 205, 209, 208, 239, 204, 124, 167, 227, 233, 246, 229, 225, 239, 226, 230, 241, 232, 
    204, 199, 179, 139, 194, 203, 221, 213, 219, 233, 216, 212, 216, 230, 188, 176, 190, 192, 212, 192, 129, 151, 183, 190, 224, 224, 214, 229, 219, 222, 235, 224, 
    205, 198, 175, 138, 192, 203, 206, 204, 212, 223, 208, 210, 213, 216, 199, 206, 178, 149, 113, 93, 85, 80, 80, 69, 108, 183, 206, 222, 208, 197, 221, 212, 
    173, 168, 154, 133, 165, 172, 160, 179, 190, 194, 189, 195, 199, 191, 193, 198, 152, 121, 107, 108, 104, 104, 110, 79, 82, 122, 159, 175, 163, 149, 190, 175, 
    115, 116, 114, 105, 109, 110, 112, 127, 135, 136, 140, 147, 151, 143, 158, 161, 134, 119, 120, 120, 108, 108, 102, 92, 143, 128, 151, 145, 110, 106, 130, 120, 
    78, 87, 86, 82, 99, 105, 97, 100, 101, 109, 106, 111, 114, 118, 132, 127, 109, 109, 110, 107, 96, 87, 108, 119, 132, 111, 144, 191, 120, 111, 102, 104, 
    74, 85, 95, 98, 128, 122, 98, 81, 104, 129, 113, 115, 132, 139, 134, 123, 120, 115, 116, 119, 113, 104, 158, 189, 183, 148, 109, 197, 149, 103, 99, 99, 
    81, 107, 113, 93, 117, 115, 93, 102, 137, 152, 149, 131, 130, 136, 125, 113, 108, 108, 114, 123, 118, 127, 175, 194, 206, 189, 118, 162, 167, 80, 98, 101, 
    97, 110, 106, 93, 98, 84, 89, 100, 110, 123, 138, 134, 126, 131, 130, 124, 123, 127, 126, 135, 134, 153, 181, 180, 184, 183, 151, 122, 160, 77, 72, 89, 
    102, 101, 102, 97, 95, 88, 88, 107, 130, 142, 151, 158, 163, 164, 161, 157, 171, 173, 170, 169, 162, 169, 177, 174, 176, 168, 164, 98, 87, 70, 63, 75, 
    123, 118, 127, 124, 126, 148, 152, 160, 167, 175, 179, 180, 183, 184, 185, 174, 173, 178, 175, 160, 128, 133, 142, 161, 169, 162, 166, 108, 70, 95, 89, 82, 
    133, 125, 138, 152, 148, 154, 166, 167, 170, 174, 179, 182, 185, 185, 181, 171, 152, 152, 154, 139, 102, 120, 144, 155, 165, 162, 163, 136, 145, 187, 153, 108, 
    124, 133, 141, 131, 116, 114, 152, 170, 175, 175, 176, 173, 167, 160, 154, 151, 144, 150, 168, 160, 140, 152, 165, 158, 163, 155, 156, 151, 158, 158, 152, 147, 
    129, 113, 96, 93, 110, 135, 148, 164, 169, 159, 150, 146, 148, 153, 159, 165, 170, 160, 168, 172, 161, 164, 168, 164, 160, 158, 158, 146, 132, 121, 125, 150, 
    112, 85, 96, 135, 155, 165, 156, 147, 142, 141, 151, 160, 167, 173, 174, 171, 167, 155, 162, 168, 163, 161, 163, 166, 158, 151, 130, 111, 98, 82, 92, 138, 
    133, 132, 135, 143, 143, 143, 150, 142, 138, 161, 169, 171, 169, 165, 151, 134, 116, 107, 148, 164, 163, 163, 159, 152, 128, 108, 102, 91, 75, 78, 80, 72, 
    132, 140, 144, 143, 144, 147, 151, 150, 139, 146, 148, 154, 159, 156, 110, 78, 75, 74, 132, 163, 153, 143, 126, 109, 103, 100, 90, 76, 75, 82, 57, 33, 
    94, 137, 148, 146, 146, 145, 129, 115, 106, 102, 99, 135, 157, 154, 114, 93, 101, 104, 125, 124, 113, 106, 102, 101, 88, 79, 69, 63, 67, 53, 37, 31, 
    86, 125, 134, 134, 137, 133, 92, 77, 82, 89, 92, 131, 153, 150, 132, 115, 106, 97, 96, 97, 99, 101, 95, 79, 60, 64, 60, 57, 47, 38, 34, 31, 
    90, 116, 129, 131, 137, 138, 106, 97, 108, 116, 124, 126, 113, 95, 84, 83, 89, 92, 98, 100, 92, 74, 67, 69, 74, 66, 51, 46, 43, 38, 35, 32, 
    92, 112, 130, 127, 124, 120, 110, 102, 97, 90, 80, 76, 75, 80, 84, 91, 95, 89, 81, 73, 65, 65, 67, 61, 69, 58, 42, 40, 42, 40, 35, 37, 
    76, 79, 86, 78, 74, 69, 64, 63, 65, 70, 74, 77, 81, 82, 81, 80, 73, 59, 55, 68, 67, 63, 54, 50, 54, 45, 40, 40, 41, 40, 39, 37, 
    45, 43, 40, 42, 49, 52, 53, 58, 68, 71, 72, 70, 65, 59, 58, 59, 56, 63, 85, 73, 57, 51, 47, 47, 44, 40, 39, 40, 41, 42, 42, 29, 
    43, 40, 36, 38, 44, 48, 49, 50, 53, 52, 49, 49, 53, 59, 62, 61, 55, 69, 94, 66, 44, 46, 47, 40, 39, 39, 40, 42, 41, 46, 32, 18, 
    40, 39, 35, 36, 39, 41, 41, 43, 46, 51, 56, 58, 61, 61, 60, 55, 46, 60, 85, 54, 40, 46, 37, 36, 38, 38, 40, 42, 43, 40, 13, 7, 
    34, 38, 36, 40, 44, 47, 49, 51, 54, 57, 59, 57, 57, 55, 51, 43, 31, 48, 78, 50, 41, 37, 35, 35, 37, 37, 36, 41, 45, 20, 6, 7, 
    41, 43, 45, 47, 48, 48, 48, 49, 50, 51, 49, 45, 40, 34, 26, 17, 8, 27, 63, 44, 33, 34, 34, 35, 35, 34, 34, 44, 31, 6, 5, 8, 
    
    -- channel=8
    222, 218, 194, 186, 222, 236, 238, 241, 243, 245, 244, 235, 240, 241, 242, 245, 227, 240, 245, 248, 249, 243, 243, 243, 245, 235, 239, 247, 241, 234, 243, 246, 
    229, 226, 201, 184, 223, 240, 240, 238, 243, 247, 245, 232, 243, 245, 245, 248, 230, 239, 243, 251, 251, 238, 238, 244, 248, 236, 243, 252, 240, 236, 250, 251, 
    225, 222, 199, 181, 219, 238, 239, 228, 235, 244, 236, 228, 235, 239, 238, 247, 229, 236, 241, 246, 236, 215, 232, 239, 248, 235, 242, 252, 241, 232, 251, 247, 
    222, 216, 194, 179, 214, 228, 235, 225, 229, 239, 230, 221, 225, 236, 230, 247, 230, 234, 240, 238, 186, 176, 229, 241, 248, 233, 239, 251, 238, 228, 248, 243, 
    223, 217, 193, 172, 210, 221, 231, 217, 218, 235, 225, 215, 219, 232, 214, 238, 229, 227, 238, 228, 176, 178, 229, 239, 247, 231, 234, 245, 231, 232, 246, 240, 
    220, 213, 191, 164, 206, 213, 225, 213, 214, 230, 218, 214, 214, 227, 200, 206, 208, 206, 237, 207, 130, 173, 230, 233, 244, 225, 219, 232, 221, 231, 242, 230, 
    212, 202, 185, 150, 196, 201, 217, 208, 211, 219, 208, 211, 212, 221, 185, 175, 187, 189, 210, 197, 137, 157, 184, 187, 221, 220, 206, 218, 209, 219, 231, 216, 
    211, 201, 179, 147, 197, 204, 206, 203, 208, 210, 198, 205, 206, 206, 192, 203, 179, 155, 122, 106, 100, 94, 88, 73, 111, 183, 202, 215, 198, 185, 206, 193, 
    179, 173, 160, 140, 170, 175, 161, 179, 187, 184, 180, 189, 195, 185, 186, 196, 159, 137, 128, 128, 126, 126, 128, 90, 88, 124, 158, 172, 156, 137, 176, 159, 
    123, 126, 123, 112, 114, 114, 114, 128, 134, 134, 137, 144, 152, 146, 160, 167, 147, 139, 144, 140, 130, 131, 120, 104, 149, 131, 150, 141, 106, 105, 128, 117, 
    89, 102, 98, 88, 107, 115, 104, 106, 107, 118, 113, 115, 123, 134, 151, 146, 128, 127, 127, 120, 111, 104, 122, 128, 134, 110, 139, 182, 114, 117, 109, 112, 
    88, 104, 110, 106, 142, 137, 113, 94, 116, 146, 127, 125, 148, 165, 165, 151, 142, 130, 127, 127, 123, 114, 165, 191, 180, 142, 100, 184, 140, 109, 108, 108, 
    100, 130, 132, 104, 129, 130, 109, 118, 154, 171, 168, 151, 155, 165, 154, 139, 130, 125, 129, 140, 134, 137, 179, 193, 203, 185, 112, 152, 160, 84, 105, 109, 
    120, 134, 126, 106, 113, 101, 108, 121, 131, 145, 161, 159, 153, 161, 158, 149, 146, 147, 145, 155, 150, 161, 182, 177, 181, 181, 148, 118, 157, 80, 78, 96, 
    127, 128, 125, 114, 116, 113, 115, 134, 159, 168, 176, 184, 190, 191, 190, 185, 197, 196, 190, 184, 172, 173, 175, 168, 171, 165, 163, 99, 87, 71, 67, 81, 
    151, 149, 154, 145, 153, 179, 184, 193, 201, 205, 207, 208, 209, 210, 212, 200, 198, 201, 195, 171, 134, 135, 139, 155, 165, 161, 168, 113, 73, 92, 90, 86, 
    165, 159, 167, 176, 175, 185, 198, 201, 205, 208, 210, 210, 210, 208, 201, 190, 170, 170, 169, 148, 108, 122, 142, 153, 167, 165, 167, 142, 147, 181, 152, 111, 
    157, 170, 174, 157, 141, 143, 182, 202, 208, 211, 209, 202, 191, 181, 167, 162, 155, 160, 178, 169, 147, 157, 167, 160, 169, 162, 161, 156, 158, 150, 150, 148, 
    162, 148, 128, 121, 138, 164, 177, 194, 199, 188, 178, 171, 170, 172, 172, 176, 180, 168, 176, 181, 170, 173, 175, 172, 168, 165, 163, 150, 133, 118, 125, 153, 
    143, 117, 127, 166, 188, 197, 186, 176, 169, 163, 171, 178, 185, 190, 191, 186, 180, 165, 172, 177, 173, 172, 175, 178, 164, 156, 136, 116, 103, 87, 98, 144, 
    166, 165, 168, 176, 176, 174, 179, 170, 164, 184, 190, 189, 185, 181, 168, 150, 129, 118, 157, 173, 173, 173, 171, 162, 133, 112, 106, 95, 80, 84, 86, 78, 
    165, 172, 177, 175, 174, 176, 179, 176, 164, 171, 171, 173, 175, 171, 126, 94, 88, 85, 142, 172, 162, 152, 136, 117, 108, 104, 94, 80, 79, 88, 63, 39, 
    124, 166, 178, 175, 175, 173, 154, 139, 130, 126, 122, 154, 174, 169, 131, 108, 114, 114, 134, 133, 121, 113, 109, 108, 95, 86, 75, 69, 73, 59, 43, 38, 
    111, 150, 160, 159, 163, 158, 116, 100, 104, 112, 115, 151, 172, 168, 149, 131, 119, 107, 106, 106, 106, 108, 100, 84, 69, 73, 68, 65, 55, 44, 40, 37, 
    113, 138, 151, 154, 161, 162, 128, 119, 129, 136, 144, 146, 132, 114, 101, 98, 101, 103, 109, 108, 99, 80, 72, 75, 85, 77, 61, 58, 52, 45, 41, 39, 
    116, 136, 154, 151, 148, 143, 132, 124, 118, 103, 91, 87, 86, 91, 99, 101, 101, 99, 94, 82, 72, 72, 74, 69, 78, 68, 52, 50, 51, 48, 47, 48, 
    96, 100, 106, 99, 92, 86, 82, 81, 82, 79, 81, 84, 87, 91, 94, 88, 77, 68, 68, 76, 74, 72, 64, 59, 63, 54, 49, 50, 49, 48, 52, 48, 
    59, 57, 54, 55, 60, 61, 62, 68, 78, 79, 79, 77, 72, 68, 69, 66, 61, 71, 97, 82, 65, 60, 56, 57, 53, 49, 48, 49, 50, 50, 50, 35, 
    50, 48, 44, 45, 49, 53, 53, 55, 58, 59, 56, 56, 60, 66, 71, 68, 59, 75, 104, 75, 53, 56, 58, 51, 49, 48, 49, 51, 50, 53, 37, 20, 
    45, 44, 40, 41, 44, 46, 46, 48, 51, 57, 63, 65, 68, 68, 68, 61, 50, 66, 93, 63, 49, 56, 48, 47, 47, 47, 49, 51, 52, 46, 14, 5, 
    39, 43, 41, 45, 50, 54, 56, 59, 62, 64, 66, 64, 64, 61, 58, 49, 36, 53, 85, 59, 50, 48, 47, 47, 46, 46, 45, 50, 54, 24, 3, 3, 
    47, 50, 52, 54, 56, 56, 56, 58, 58, 55, 53, 50, 45, 39, 30, 20, 11, 33, 72, 54, 44, 45, 45, 46, 44, 44, 43, 52, 37, 8, 3, 7, 
    
    -- channel=9
    155, 167, 176, 190, 177, 166, 168, 166, 170, 179, 187, 187, 187, 187, 184, 184, 182, 180, 184, 186, 187, 187, 188, 189, 187, 187, 188, 195, 201, 201, 202, 192, 
    153, 163, 171, 187, 179, 155, 154, 159, 159, 165, 171, 175, 169, 171, 162, 165, 170, 164, 166, 165, 167, 173, 169, 168, 169, 173, 190, 202, 204, 202, 203, 189, 
    155, 160, 168, 184, 187, 174, 176, 188, 182, 179, 177, 190, 192, 194, 188, 185, 193, 194, 193, 194, 195, 197, 193, 191, 191, 197, 206, 207, 208, 206, 204, 189, 
    151, 157, 166, 177, 180, 185, 199, 197, 182, 204, 205, 198, 210, 197, 196, 203, 205, 207, 210, 203, 207, 210, 197, 204, 208, 198, 204, 201, 209, 207, 206, 192, 
    151, 158, 168, 174, 177, 181, 191, 196, 183, 194, 189, 185, 196, 185, 185, 202, 199, 199, 200, 192, 195, 199, 190, 188, 201, 199, 201, 196, 206, 204, 207, 196, 
    148, 156, 167, 174, 171, 174, 196, 195, 192, 190, 189, 184, 187, 189, 189, 191, 190, 195, 187, 198, 192, 188, 192, 193, 205, 206, 203, 209, 212, 208, 209, 196, 
    148, 153, 165, 174, 168, 176, 203, 195, 188, 188, 187, 190, 182, 194, 197, 195, 196, 193, 200, 205, 198, 197, 197, 201, 197, 200, 198, 195, 197, 203, 207, 195, 
    153, 155, 163, 172, 172, 188, 199, 209, 196, 190, 189, 191, 193, 188, 187, 196, 202, 194, 196, 206, 194, 201, 196, 200, 181, 187, 200, 201, 200, 196, 199, 189, 
    160, 159, 163, 172, 174, 176, 176, 190, 180, 175, 176, 176, 181, 170, 172, 182, 187, 178, 181, 187, 177, 188, 180, 187, 199, 196, 188, 188, 197, 192, 194, 184, 
    171, 167, 162, 172, 170, 171, 180, 176, 155, 156, 150, 156, 150, 146, 153, 158, 166, 166, 164, 157, 157, 162, 156, 166, 200, 199, 188, 189, 197, 193, 194, 182, 
    175, 180, 168, 176, 173, 177, 182, 174, 156, 160, 159, 154, 159, 163, 168, 173, 170, 164, 160, 162, 160, 168, 167, 172, 194, 195, 196, 196, 197, 191, 193, 183, 
    181, 187, 178, 187, 183, 170, 174, 182, 179, 179, 180, 181, 184, 187, 193, 193, 193, 192, 188, 185, 184, 186, 192, 192, 187, 188, 192, 189, 190, 191, 196, 186, 
    185, 190, 186, 171, 153, 132, 149, 193, 198, 191, 186, 188, 191, 193, 195, 196, 195, 192, 190, 188, 188, 190, 192, 191, 191, 193, 195, 197, 202, 202, 204, 193, 
    186, 194, 188, 158, 132, 116, 94, 109, 145, 177, 194, 194, 191, 193, 196, 199, 199, 199, 200, 198, 196, 196, 199, 198, 197, 196, 196, 196, 198, 197, 198, 185, 
    186, 197, 196, 198, 194, 184, 141, 92, 84, 104, 142, 179, 195, 201, 204, 204, 204, 204, 204, 199, 194, 194, 194, 191, 189, 190, 190, 190, 191, 190, 192, 181, 
    184, 199, 198, 200, 197, 200, 201, 177, 117, 84, 93, 128, 173, 202, 208, 205, 202, 200, 199, 199, 195, 196, 197, 195, 193, 195, 194, 191, 191, 189, 190, 178, 
    185, 201, 203, 208, 205, 206, 208, 214, 175, 92, 76, 91, 105, 140, 181, 203, 206, 202, 197, 194, 193, 194, 194, 194, 194, 195, 193, 191, 193, 190, 190, 180, 
    187, 204, 207, 214, 212, 212, 211, 208, 203, 124, 71, 87, 84, 84, 99, 132, 167, 190, 203, 203, 195, 192, 197, 196, 194, 194, 192, 191, 193, 191, 192, 183, 
    190, 207, 207, 214, 212, 211, 211, 208, 211, 137, 72, 87, 83, 84, 86, 83, 89, 107, 131, 155, 163, 182, 203, 204, 202, 198, 194, 191, 193, 192, 191, 182, 
    191, 210, 209, 215, 213, 212, 212, 213, 204, 113, 47, 58, 63, 76, 87, 93, 90, 80, 70, 62, 58, 77, 122, 159, 180, 194, 201, 200, 200, 196, 196, 185, 
    191, 208, 207, 211, 209, 210, 209, 212, 157, 101, 65, 37, 51, 68, 74, 88, 91, 86, 85, 73, 55, 46, 62, 72, 78, 107, 133, 158, 184, 195, 196, 186, 
    186, 202, 203, 209, 207, 206, 209, 200, 149, 140, 151, 100, 45, 53, 50, 96, 156, 160, 128, 72, 98, 112, 89, 66, 67, 131, 166, 163, 173, 183, 188, 178, 
    185, 201, 202, 210, 210, 208, 209, 209, 210, 211, 215, 189, 144, 146, 148, 168, 202, 206, 192, 154, 163, 178, 177, 159, 156, 178, 191, 194, 196, 193, 188, 176, 
    176, 188, 192, 196, 192, 188, 185, 183, 182, 178, 179, 173, 170, 170, 171, 173, 169, 160, 161, 167, 165, 161, 165, 170, 170, 160, 152, 150, 157, 163, 164, 156, 
    114, 99, 110, 107, 102, 97, 94, 93, 88, 85, 88, 80, 77, 78, 83, 101, 113, 108, 106, 107, 108, 110, 111, 113, 117, 119, 120, 119, 120, 121, 122, 124, 
    122, 109, 113, 117, 115, 112, 114, 113, 111, 112, 111, 109, 110, 109, 110, 108, 115, 112, 105, 107, 108, 106, 101, 104, 106, 107, 109, 109, 103, 102, 94, 101, 
    120, 97, 107, 112, 109, 104, 98, 94, 94, 93, 88, 86, 82, 79, 80, 78, 80, 79, 72, 69, 67, 66, 65, 65, 64, 65, 66, 64, 67, 63, 53, 77, 
    91, 55, 65, 69, 66, 66, 63, 61, 66, 64, 60, 57, 57, 60, 61, 63, 63, 66, 64, 58, 56, 57, 59, 60, 58, 57, 56, 57, 52, 49, 75, 92, 
    93, 60, 66, 68, 67, 67, 64, 65, 69, 65, 62, 59, 59, 59, 60, 61, 64, 63, 58, 56, 55, 55, 56, 56, 57, 58, 56, 53, 65, 93, 97, 81, 
    89, 57, 61, 57, 57, 59, 57, 59, 60, 58, 56, 54, 60, 61, 59, 61, 65, 61, 58, 57, 60, 60, 61, 61, 66, 62, 57, 70, 97, 89, 59, 67, 
    89, 60, 63, 62, 62, 62, 62, 63, 62, 61, 65, 82, 84, 81, 78, 81, 88, 84, 85, 83, 80, 67, 66, 64, 52, 56, 86, 103, 76, 57, 61, 75, 
    92, 60, 61, 60, 63, 66, 67, 65, 66, 67, 65, 72, 73, 73, 72, 70, 73, 74, 75, 75, 75, 64, 64, 62, 65, 86, 88, 64, 57, 60, 64, 73, 
    
    -- channel=10
    156, 176, 179, 192, 185, 171, 173, 173, 175, 179, 182, 184, 185, 184, 182, 181, 179, 179, 183, 185, 186, 186, 187, 189, 187, 187, 188, 195, 197, 196, 202, 183, 
    155, 179, 184, 195, 190, 162, 159, 164, 163, 165, 169, 176, 171, 174, 164, 167, 172, 166, 168, 166, 169, 175, 171, 169, 170, 174, 191, 204, 206, 208, 215, 190, 
    154, 178, 185, 196, 203, 193, 178, 168, 160, 175, 190, 196, 195, 197, 190, 188, 196, 195, 194, 195, 196, 198, 193, 191, 192, 196, 205, 205, 206, 208, 215, 191, 
    154, 178, 188, 195, 202, 197, 188, 128, 108, 152, 154, 155, 158, 149, 149, 148, 167, 161, 163, 173, 168, 163, 174, 159, 188, 208, 204, 206, 204, 205, 212, 188, 
    154, 177, 187, 191, 198, 196, 189, 126, 128, 139, 106, 107, 115, 120, 118, 113, 119, 114, 114, 126, 118, 112, 136, 112, 160, 203, 201, 206, 206, 205, 214, 190, 
    151, 174, 187, 189, 197, 200, 183, 147, 169, 168, 145, 165, 170, 146, 149, 157, 180, 178, 176, 189, 176, 179, 188, 177, 196, 208, 207, 208, 208, 209, 216, 190, 
    152, 172, 185, 189, 194, 198, 147, 96, 149, 151, 144, 152, 152, 121, 128, 139, 156, 151, 170, 162, 150, 173, 150, 164, 156, 166, 204, 210, 211, 207, 212, 188, 
    155, 172, 182, 187, 194, 181, 119, 101, 123, 131, 131, 120, 146, 135, 135, 127, 123, 123, 131, 123, 109, 132, 123, 159, 123, 132, 191, 199, 201, 201, 208, 186, 
    161, 175, 180, 185, 192, 186, 171, 175, 162, 165, 172, 166, 175, 172, 173, 170, 172, 178, 178, 175, 163, 172, 178, 190, 172, 176, 200, 205, 200, 201, 209, 185, 
    172, 183, 180, 186, 190, 192, 194, 183, 160, 165, 162, 163, 159, 158, 164, 162, 167, 174, 172, 162, 160, 163, 165, 182, 200, 198, 202, 205, 202, 202, 208, 184, 
    177, 196, 186, 190, 192, 193, 193, 183, 163, 167, 165, 159, 164, 166, 170, 172, 168, 166, 166, 171, 168, 173, 171, 178, 199, 198, 199, 199, 200, 200, 208, 184, 
    183, 204, 195, 200, 201, 187, 190, 198, 194, 193, 193, 193, 193, 194, 198, 198, 198, 195, 195, 198, 197, 196, 196, 197, 201, 203, 201, 201, 202, 200, 209, 187, 
    185, 205, 198, 178, 166, 141, 154, 196, 202, 202, 199, 197, 197, 199, 201, 202, 201, 199, 198, 196, 196, 198, 199, 198, 199, 202, 203, 206, 207, 206, 212, 189, 
    186, 208, 200, 165, 144, 124, 95, 107, 143, 179, 199, 199, 197, 198, 201, 204, 204, 205, 206, 204, 201, 201, 205, 205, 204, 203, 203, 203, 202, 202, 207, 183, 
    186, 212, 208, 204, 206, 193, 143, 91, 81, 101, 142, 181, 198, 204, 207, 207, 207, 207, 207, 202, 197, 197, 198, 197, 197, 197, 197, 197, 196, 197, 204, 181, 
    184, 214, 210, 206, 209, 212, 207, 179, 116, 83, 93, 128, 174, 203, 210, 206, 204, 202, 202, 201, 198, 199, 201, 201, 200, 202, 201, 199, 198, 198, 203, 180, 
    186, 215, 214, 213, 214, 214, 212, 217, 175, 91, 73, 86, 101, 138, 181, 204, 208, 203, 199, 198, 199, 201, 201, 200, 200, 202, 201, 201, 202, 200, 204, 182, 
    187, 216, 216, 217, 219, 217, 214, 211, 204, 123, 68, 82, 79, 81, 97, 130, 165, 188, 201, 202, 196, 193, 199, 198, 198, 199, 200, 200, 201, 199, 204, 182, 
    188, 217, 213, 214, 216, 216, 214, 210, 212, 136, 70, 83, 78, 80, 80, 77, 83, 102, 126, 151, 159, 178, 201, 204, 203, 201, 200, 198, 199, 197, 201, 180, 
    187, 218, 214, 213, 215, 216, 215, 216, 204, 112, 45, 55, 58, 69, 77, 81, 80, 77, 70, 62, 59, 79, 124, 160, 181, 196, 205, 205, 203, 200, 202, 180, 
    188, 216, 210, 209, 211, 214, 212, 212, 154, 95, 58, 33, 48, 62, 65, 77, 82, 84, 84, 72, 56, 47, 63, 72, 78, 107, 132, 158, 181, 193, 202, 182, 
    184, 210, 206, 207, 209, 211, 212, 200, 145, 133, 143, 97, 45, 50, 46, 90, 150, 158, 127, 71, 97, 112, 88, 65, 67, 130, 165, 162, 168, 181, 197, 176, 
    183, 210, 205, 208, 211, 212, 213, 210, 209, 209, 212, 191, 148, 147, 147, 166, 200, 208, 195, 157, 166, 181, 180, 162, 159, 180, 193, 197, 195, 193, 199, 177, 
    174, 196, 195, 194, 194, 190, 187, 185, 184, 181, 183, 181, 178, 176, 174, 173, 170, 164, 166, 172, 170, 166, 170, 176, 175, 165, 157, 155, 157, 163, 175, 158, 
    112, 108, 112, 105, 103, 100, 97, 96, 92, 90, 94, 87, 84, 83, 87, 103, 115, 112, 111, 112, 113, 115, 116, 118, 122, 123, 124, 123, 121, 122, 132, 124, 
    117, 115, 113, 112, 113, 111, 113, 113, 111, 112, 111, 110, 110, 109, 110, 107, 115, 115, 108, 110, 111, 109, 104, 107, 109, 110, 112, 112, 100, 95, 98, 101, 
    113, 102, 105, 106, 106, 102, 97, 93, 95, 94, 89, 85, 82, 78, 79, 78, 80, 79, 71, 68, 67, 65, 65, 65, 65, 66, 66, 65, 60, 55, 71, 100, 
    84, 60, 65, 64, 64, 64, 62, 60, 66, 64, 61, 56, 57, 60, 61, 63, 64, 67, 65, 59, 56, 58, 59, 60, 58, 57, 56, 56, 56, 72, 117, 128, 
    83, 59, 63, 62, 63, 65, 61, 63, 67, 62, 60, 57, 58, 58, 60, 61, 65, 68, 64, 62, 61, 60, 62, 61, 58, 58, 61, 65, 91, 136, 137, 99, 
    79, 53, 61, 57, 55, 59, 58, 60, 61, 60, 57, 55, 60, 62, 61, 63, 67, 63, 60, 59, 62, 62, 64, 63, 62, 60, 71, 110, 142, 119, 79, 74, 
    82, 58, 66, 65, 63, 62, 62, 62, 63, 62, 65, 79, 79, 76, 74, 77, 84, 80, 80, 78, 76, 63, 62, 65, 66, 86, 124, 141, 102, 66, 64, 69, 
    78, 52, 58, 58, 58, 58, 59, 57, 58, 59, 58, 69, 71, 71, 70, 69, 72, 72, 73, 74, 73, 63, 63, 68, 90, 128, 128, 88, 66, 63, 65, 68, 
    
    -- channel=11
    149, 187, 193, 205, 202, 183, 181, 180, 182, 189, 193, 192, 192, 192, 189, 189, 186, 185, 189, 192, 193, 193, 192, 190, 187, 187, 188, 195, 202, 209, 212, 171, 
    157, 204, 215, 227, 224, 190, 179, 179, 179, 187, 195, 195, 187, 190, 180, 183, 188, 183, 184, 183, 185, 191, 188, 188, 190, 194, 211, 224, 223, 222, 227, 183, 
    153, 201, 213, 219, 223, 213, 196, 184, 177, 195, 211, 212, 208, 210, 204, 202, 209, 209, 208, 209, 210, 212, 208, 208, 208, 213, 222, 223, 218, 215, 224, 184, 
    166, 207, 211, 222, 226, 220, 201, 131, 119, 158, 166, 177, 178, 167, 166, 171, 183, 178, 178, 186, 185, 186, 180, 165, 207, 228, 220, 221, 224, 223, 230, 186, 
    167, 203, 202, 218, 224, 225, 214, 142, 153, 152, 120, 129, 129, 126, 124, 131, 134, 132, 130, 138, 136, 136, 141, 123, 186, 227, 218, 217, 222, 220, 227, 185, 
    164, 201, 203, 217, 220, 218, 209, 165, 196, 181, 156, 180, 179, 160, 163, 172, 191, 193, 190, 201, 191, 192, 198, 190, 212, 225, 225, 225, 223, 225, 232, 188, 
    164, 198, 200, 217, 217, 214, 172, 104, 158, 165, 166, 175, 165, 144, 151, 160, 178, 173, 189, 182, 170, 183, 173, 185, 166, 178, 220, 226, 221, 224, 231, 188, 
    169, 201, 199, 216, 218, 203, 146, 111, 134, 149, 157, 144, 155, 143, 143, 144, 147, 142, 148, 142, 127, 141, 142, 176, 137, 149, 209, 220, 217, 220, 228, 186, 
    177, 206, 199, 217, 219, 205, 193, 197, 184, 183, 187, 184, 192, 186, 187, 189, 192, 194, 194, 191, 178, 186, 188, 200, 193, 198, 214, 219, 219, 221, 228, 185, 
    186, 212, 197, 214, 215, 214, 220, 210, 185, 187, 182, 186, 182, 180, 185, 186, 193, 198, 195, 184, 181, 182, 182, 198, 222, 222, 221, 223, 223, 222, 227, 183, 
    188, 222, 200, 216, 215, 212, 214, 204, 181, 184, 182, 176, 181, 184, 188, 191, 189, 186, 184, 185, 182, 184, 186, 201, 223, 221, 220, 219, 219, 220, 227, 184, 
    191, 226, 207, 224, 220, 209, 215, 222, 217, 215, 214, 215, 217, 219, 223, 223, 223, 221, 219, 218, 216, 214, 217, 219, 219, 219, 217, 214, 215, 219, 227, 186, 
    188, 220, 212, 206, 181, 153, 172, 217, 226, 225, 221, 220, 222, 223, 225, 226, 225, 221, 220, 218, 217, 219, 220, 218, 217, 220, 222, 224, 224, 224, 230, 187, 
    189, 223, 214, 193, 157, 126, 99, 115, 157, 198, 221, 221, 218, 220, 223, 226, 226, 224, 225, 223, 220, 221, 224, 224, 223, 222, 222, 222, 221, 221, 226, 183, 
    189, 226, 222, 233, 220, 196, 146, 90, 84, 113, 161, 202, 218, 224, 227, 228, 226, 225, 224, 220, 215, 215, 216, 217, 216, 216, 216, 216, 215, 218, 225, 182, 
    187, 229, 224, 234, 225, 225, 218, 179, 115, 88, 106, 145, 192, 221, 228, 225, 223, 219, 218, 217, 214, 214, 217, 219, 219, 221, 220, 218, 217, 220, 226, 183, 
    190, 233, 222, 233, 228, 226, 224, 225, 181, 98, 80, 91, 106, 146, 192, 217, 224, 225, 221, 218, 217, 218, 218, 217, 218, 221, 221, 221, 221, 220, 227, 188, 
    191, 234, 221, 233, 231, 227, 226, 221, 213, 130, 73, 79, 75, 80, 100, 136, 173, 200, 215, 220, 217, 217, 223, 222, 221, 221, 219, 219, 218, 219, 227, 189, 
    189, 232, 217, 228, 227, 225, 226, 220, 221, 144, 74, 80, 74, 76, 78, 76, 83, 100, 129, 161, 176, 201, 225, 226, 223, 220, 217, 215, 215, 217, 225, 187, 
    187, 232, 215, 225, 224, 225, 227, 226, 213, 119, 50, 56, 59, 69, 77, 82, 80, 72, 66, 63, 65, 91, 133, 162, 184, 204, 218, 223, 221, 221, 227, 188, 
    183, 231, 222, 223, 223, 230, 228, 225, 162, 98, 60, 39, 53, 67, 68, 78, 81, 82, 83, 72, 57, 49, 63, 67, 75, 109, 139, 168, 198, 215, 223, 195, 
    176, 226, 226, 222, 222, 226, 226, 212, 155, 139, 150, 106, 53, 57, 51, 94, 154, 161, 130, 73, 99, 114, 90, 67, 69, 134, 171, 169, 183, 197, 208, 190, 
    175, 225, 225, 223, 223, 222, 222, 222, 222, 224, 228, 204, 159, 159, 160, 179, 214, 220, 207, 169, 178, 193, 192, 173, 171, 195, 210, 214, 216, 209, 210, 189, 
    166, 212, 215, 209, 206, 204, 201, 199, 199, 195, 197, 194, 192, 193, 194, 196, 196, 194, 196, 202, 200, 196, 200, 205, 206, 197, 192, 191, 197, 197, 201, 181, 
    101, 120, 130, 120, 118, 112, 107, 106, 101, 98, 102, 99, 98, 101, 108, 128, 144, 146, 146, 147, 148, 150, 152, 158, 164, 166, 168, 168, 168, 165, 167, 146, 
    111, 130, 134, 134, 138, 136, 137, 136, 132, 134, 131, 126, 127, 128, 131, 131, 138, 134, 127, 129, 129, 128, 124, 126, 129, 130, 132, 132, 119, 115, 115, 96, 
    104, 113, 120, 120, 122, 118, 108, 100, 96, 91, 85, 89, 88, 85, 87, 86, 86, 79, 70, 67, 66, 65, 63, 60, 59, 60, 60, 59, 54, 50, 63, 75, 
    61, 55, 61, 57, 58, 63, 59, 54, 56, 51, 47, 47, 48, 50, 49, 50, 51, 55, 53, 47, 45, 46, 50, 55, 54, 52, 52, 52, 48, 58, 104, 104, 
    68, 61, 65, 60, 62, 61, 55, 57, 61, 56, 55, 58, 59, 56, 56, 54, 57, 59, 55, 52, 51, 51, 52, 52, 51, 53, 55, 57, 75, 113, 120, 75, 
    62, 52, 59, 53, 57, 57, 52, 54, 54, 50, 48, 50, 57, 56, 52, 53, 57, 54, 52, 51, 54, 55, 53, 48, 50, 52, 61, 95, 124, 101, 62, 50, 
    62, 53, 58, 55, 59, 61, 60, 60, 57, 55, 58, 75, 76, 72, 68, 69, 75, 74, 75, 73, 70, 58, 55, 53, 51, 69, 107, 127, 91, 58, 54, 51, 
    64, 51, 51, 46, 51, 56, 57, 53, 52, 51, 50, 62, 64, 62, 60, 57, 60, 62, 64, 64, 64, 53, 52, 55, 70, 103, 105, 72, 53, 50, 52, 50, 
    
    -- channel=12
    65, 70, 48, 30, 23, 40, 44, 45, 45, 40, 10, 15, 44, 53, 51, 48, 65, 90, 93, 91, 95, 81, 60, 55, 112, 111, 41, 68, 77, 51, 54, 67, 
    69, 79, 60, 30, 41, 65, 49, 49, 49, 35, 7, 25, 65, 69, 55, 49, 77, 85, 83, 80, 87, 81, 55, 59, 131, 121, 31, 47, 56, 54, 65, 61, 
    73, 84, 72, 41, 64, 74, 50, 54, 54, 32, 11, 36, 60, 67, 47, 39, 75, 77, 59, 62, 83, 85, 48, 63, 139, 128, 23, 41, 70, 78, 73, 48, 
    88, 75, 80, 54, 80, 68, 55, 63, 58, 28, 17, 37, 43, 51, 40, 39, 85, 98, 75, 70, 86, 84, 50, 68, 142, 137, 47, 75, 100, 93, 65, 38, 
    95, 89, 111, 66, 81, 61, 61, 68, 62, 22, 15, 22, 31, 35, 51, 63, 72, 75, 72, 71, 77, 83, 51, 78, 149, 156, 87, 87, 99, 95, 75, 88, 
    82, 83, 82, 77, 71, 58, 64, 57, 59, 20, 17, 28, 50, 61, 71, 71, 69, 67, 68, 56, 41, 83, 70, 78, 156, 172, 98, 89, 94, 111, 112, 99, 
    69, 64, 32, 59, 72, 74, 73, 49, 49, 18, 29, 62, 82, 85, 86, 63, 34, 52, 95, 43, 25, 94, 85, 78, 166, 180, 109, 107, 108, 131, 86, 47, 
    59, 53, 25, 70, 81, 78, 80, 61, 40, 10, 53, 94, 87, 88, 75, 25, 13, 45, 92, 57, 50, 101, 89, 98, 144, 179, 120, 124, 124, 128, 52, 24, 
    68, 47, 49, 102, 119, 89, 63, 79, 66, 34, 81, 96, 89, 90, 41, 14, 52, 92, 67, 71, 111, 113, 110, 115, 136, 156, 121, 127, 124, 115, 31, 22, 
    77, 53, 55, 114, 128, 123, 65, 55, 79, 82, 111, 110, 106, 69, 20, 37, 92, 105, 83, 97, 118, 120, 115, 92, 144, 147, 125, 127, 119, 95, 14, 23, 
    85, 58, 54, 112, 129, 132, 100, 49, 39, 84, 104, 109, 125, 93, 63, 83, 97, 94, 104, 110, 109, 127, 85, 57, 152, 150, 123, 124, 114, 93, 12, 21, 
    108, 53, 50, 107, 126, 131, 128, 75, 51, 91, 85, 107, 138, 110, 129, 147, 132, 120, 113, 119, 117, 115, 90, 93, 160, 141, 113, 125, 121, 101, 14, 9, 
    96, 42, 43, 92, 106, 128, 130, 119, 120, 123, 114, 137, 148, 110, 105, 132, 146, 135, 128, 134, 140, 120, 126, 119, 152, 145, 99, 106, 130, 99, 18, 40, 
    97, 66, 59, 89, 100, 111, 133, 136, 147, 140, 150, 145, 142, 136, 131, 127, 125, 123, 136, 147, 151, 142, 156, 136, 146, 144, 109, 112, 130, 92, 50, 83, 
    105, 72, 75, 95, 104, 94, 133, 133, 143, 135, 128, 133, 147, 150, 160, 152, 145, 144, 132, 135, 138, 138, 162, 165, 163, 127, 126, 119, 118, 95, 59, 77, 
    94, 68, 68, 91, 101, 98, 123, 131, 147, 193, 138, 79, 124, 147, 147, 162, 180, 171, 152, 144, 144, 121, 148, 179, 180, 160, 128, 123, 112, 63, 26, 84, 
    88, 79, 74, 89, 110, 120, 120, 129, 120, 184, 192, 87, 114, 156, 164, 166, 154, 161, 183, 182, 187, 173, 148, 143, 181, 195, 142, 124, 107, 44, 41, 118, 
    91, 89, 103, 96, 116, 100, 111, 106, 114, 128, 187, 168, 140, 153, 172, 172, 167, 164, 157, 163, 161, 165, 171, 156, 161, 145, 167, 114, 106, 74, 42, 94, 
    101, 97, 120, 122, 114, 78, 95, 91, 115, 110, 129, 204, 167, 137, 160, 153, 179, 186, 170, 178, 179, 156, 162, 165, 156, 140, 104, 72, 84, 89, 70, 114, 
    110, 107, 122, 96, 90, 76, 72, 100, 109, 127, 87, 140, 189, 159, 166, 180, 174, 173, 190, 188, 162, 153, 162, 161, 153, 149, 75, 74, 66, 62, 112, 138, 
    119, 106, 89, 78, 89, 71, 60, 103, 75, 95, 114, 66, 127, 181, 174, 190, 186, 171, 184, 193, 164, 160, 171, 165, 146, 139, 104, 92, 77, 94, 112, 115, 
    126, 94, 58, 103, 106, 76, 72, 95, 94, 65, 120, 99, 91, 161, 196, 188, 182, 193, 167, 167, 170, 160, 154, 161, 145, 138, 110, 81, 105, 136, 109, 100, 
    111, 82, 70, 104, 113, 94, 69, 84, 116, 109, 85, 125, 127, 155, 186, 200, 187, 187, 177, 157, 148, 162, 164, 166, 162, 149, 121, 97, 120, 115, 97, 97, 
    101, 92, 140, 180, 151, 123, 85, 76, 103, 124, 90, 84, 146, 175, 173, 200, 188, 173, 173, 159, 159, 172, 163, 173, 164, 139, 131, 131, 112, 95, 100, 96, 
    119, 144, 192, 209, 194, 157, 127, 108, 106, 94, 106, 111, 124, 175, 176, 197, 184, 170, 176, 165, 156, 197, 175, 163, 147, 131, 122, 101, 100, 96, 107, 102, 
    110, 116, 138, 169, 197, 196, 160, 136, 129, 99, 92, 138, 146, 159, 180, 169, 142, 141, 175, 178, 166, 188, 179, 151, 143, 154, 112, 58, 91, 101, 102, 73, 
    91, 87, 74, 107, 165, 185, 191, 163, 134, 128, 106, 102, 118, 132, 146, 116, 77, 99, 161, 182, 183, 159, 173, 167, 156, 135, 94, 43, 91, 92, 68, 77, 
    81, 95, 50, 44, 95, 148, 166, 187, 174, 144, 126, 114, 104, 114, 119, 107, 81, 82, 157, 182, 169, 178, 169, 150, 152, 108, 44, 63, 97, 69, 80, 86, 
    90, 95, 52, 21, 28, 109, 146, 176, 202, 181, 142, 127, 120, 119, 114, 130, 129, 118, 144, 169, 159, 173, 180, 152, 119, 68, 44, 85, 51, 114, 167, 106, 
    95, 91, 57, 52, 24, 49, 119, 156, 187, 203, 186, 155, 141, 133, 116, 117, 109, 119, 139, 153, 159, 167, 156, 125, 101, 65, 68, 64, 55, 144, 170, 122, 
    94, 75, 32, 73, 46, 33, 54, 115, 150, 176, 195, 194, 177, 155, 136, 146, 139, 101, 94, 119, 101, 95, 96, 105, 131, 118, 107, 109, 128, 143, 154, 106, 
    78, 35, 24, 76, 65, 40, 27, 59, 120, 136, 150, 176, 192, 183, 165, 186, 207, 170, 107, 86, 66, 85, 112, 140, 169, 149, 137, 137, 150, 143, 154, 128, 
    
    -- channel=13
    68, 81, 64, 46, 33, 57, 75, 80, 83, 70, 20, 34, 71, 75, 70, 66, 87, 120, 124, 121, 126, 108, 84, 82, 136, 129, 59, 91, 96, 67, 76, 87, 
    80, 102, 74, 47, 56, 92, 84, 84, 88, 62, 18, 48, 93, 92, 77, 73, 107, 117, 111, 106, 117, 108, 77, 83, 151, 139, 45, 65, 71, 66, 90, 81, 
    95, 109, 88, 56, 84, 105, 86, 90, 92, 53, 20, 60, 89, 88, 66, 60, 103, 102, 78, 84, 114, 114, 66, 86, 158, 143, 35, 55, 84, 98, 98, 59, 
    116, 100, 100, 73, 109, 102, 88, 96, 94, 45, 26, 56, 65, 67, 54, 55, 106, 117, 97, 98, 118, 114, 69, 91, 160, 150, 64, 93, 120, 126, 94, 50, 
    120, 104, 128, 93, 114, 94, 90, 94, 93, 39, 26, 36, 47, 55, 73, 86, 105, 113, 107, 101, 103, 109, 74, 103, 162, 172, 112, 116, 129, 132, 103, 108, 
    105, 102, 98, 98, 95, 89, 91, 78, 88, 35, 27, 43, 77, 93, 106, 108, 103, 101, 100, 78, 57, 110, 98, 102, 167, 186, 130, 127, 129, 144, 132, 120, 
    94, 96, 48, 79, 90, 100, 93, 63, 74, 29, 38, 90, 126, 129, 130, 99, 58, 71, 115, 57, 37, 123, 113, 106, 183, 193, 141, 140, 137, 160, 101, 59, 
    86, 84, 47, 105, 103, 97, 94, 71, 56, 20, 73, 139, 138, 140, 114, 41, 26, 65, 115, 79, 59, 125, 120, 140, 176, 195, 150, 148, 144, 155, 63, 24, 
    98, 78, 74, 140, 149, 114, 80, 92, 71, 44, 113, 144, 136, 134, 63, 23, 69, 124, 94, 86, 112, 139, 155, 165, 170, 177, 150, 150, 146, 142, 41, 22, 
    116, 81, 78, 148, 163, 155, 84, 69, 81, 90, 137, 142, 138, 93, 33, 56, 124, 143, 115, 128, 151, 156, 156, 129, 167, 173, 152, 154, 148, 121, 22, 24, 
    120, 79, 73, 145, 165, 166, 127, 65, 54, 114, 142, 127, 126, 93, 71, 108, 135, 133, 146, 161, 156, 165, 117, 87, 169, 175, 151, 156, 145, 116, 19, 23, 
    123, 69, 66, 138, 161, 168, 165, 95, 75, 140, 138, 112, 109, 102, 136, 162, 153, 154, 151, 135, 124, 133, 118, 136, 189, 170, 146, 157, 148, 119, 20, 11, 
    106, 57, 60, 121, 135, 164, 173, 152, 144, 147, 127, 118, 115, 92, 102, 139, 141, 138, 133, 116, 120, 107, 119, 136, 176, 174, 135, 145, 161, 114, 26, 43, 
    116, 85, 78, 116, 127, 140, 172, 171, 153, 124, 130, 120, 119, 118, 113, 110, 105, 108, 119, 125, 131, 122, 129, 117, 144, 162, 141, 154, 166, 112, 65, 95, 
    132, 96, 99, 120, 130, 114, 165, 168, 139, 107, 104, 112, 124, 129, 142, 132, 122, 119, 107, 111, 115, 118, 141, 144, 142, 123, 146, 159, 157, 112, 72, 94, 
    121, 90, 93, 118, 127, 124, 151, 166, 153, 171, 121, 69, 107, 124, 123, 139, 155, 144, 128, 119, 122, 103, 131, 167, 159, 140, 128, 160, 149, 75, 34, 104, 
    112, 100, 100, 126, 141, 152, 149, 163, 138, 163, 166, 71, 100, 133, 139, 141, 129, 136, 160, 158, 163, 151, 125, 126, 169, 177, 122, 143, 143, 61, 51, 139, 
    112, 112, 131, 129, 147, 124, 144, 137, 143, 121, 168, 153, 122, 127, 146, 147, 141, 139, 132, 138, 134, 143, 153, 134, 145, 130, 146, 122, 134, 100, 58, 111, 
    121, 118, 149, 142, 141, 97, 123, 118, 143, 126, 121, 187, 145, 110, 136, 130, 154, 161, 148, 154, 151, 134, 150, 145, 134, 123, 97, 87, 103, 119, 97, 134, 
    136, 135, 151, 111, 122, 101, 93, 125, 134, 153, 96, 125, 169, 136, 146, 160, 150, 148, 166, 167, 141, 128, 144, 145, 132, 130, 75, 94, 83, 87, 149, 169, 
    148, 140, 112, 94, 121, 104, 84, 130, 102, 116, 141, 74, 118, 163, 155, 170, 165, 149, 157, 167, 146, 137, 147, 145, 127, 124, 109, 113, 96, 119, 156, 161, 
    152, 119, 72, 125, 129, 101, 99, 121, 120, 91, 154, 125, 93, 150, 181, 169, 162, 173, 145, 143, 143, 135, 129, 139, 125, 120, 117, 102, 129, 171, 154, 153, 
    136, 104, 82, 123, 136, 118, 98, 115, 150, 141, 117, 148, 129, 149, 173, 179, 165, 168, 159, 143, 126, 139, 140, 141, 136, 133, 122, 109, 152, 164, 150, 149, 
    125, 111, 150, 191, 172, 158, 121, 111, 145, 153, 115, 105, 148, 161, 154, 172, 161, 155, 156, 141, 137, 147, 136, 143, 137, 140, 123, 134, 156, 149, 158, 149, 
    149, 162, 200, 220, 209, 189, 170, 147, 145, 122, 125, 136, 139, 159, 150, 164, 155, 155, 159, 142, 133, 169, 147, 136, 127, 126, 107, 114, 154, 143, 160, 156, 
    139, 137, 157, 190, 213, 215, 191, 176, 169, 132, 117, 163, 173, 151, 154, 143, 124, 129, 153, 152, 145, 163, 149, 124, 119, 131, 96, 74, 145, 149, 151, 120, 
    115, 111, 97, 134, 191, 207, 211, 193, 177, 173, 145, 127, 144, 143, 134, 104, 73, 92, 139, 155, 161, 138, 148, 142, 131, 117, 85, 60, 146, 145, 111, 109, 
    106, 114, 65, 64, 120, 178, 195, 213, 202, 185, 173, 153, 142, 150, 141, 125, 108, 96, 142, 154, 144, 161, 149, 127, 131, 98, 49, 97, 147, 108, 118, 117, 
    116, 112, 62, 38, 41, 135, 180, 199, 212, 204, 183, 178, 171, 164, 158, 161, 157, 139, 135, 141, 135, 153, 156, 126, 103, 66, 59, 124, 84, 136, 197, 131, 
    127, 123, 79, 78, 37, 66, 149, 191, 208, 219, 214, 194, 184, 180, 165, 159, 135, 125, 123, 131, 138, 147, 135, 114, 108, 79, 85, 91, 78, 172, 201, 143, 
    125, 104, 52, 107, 67, 48, 78, 151, 189, 203, 217, 218, 205, 195, 180, 182, 165, 116, 94, 122, 97, 89, 89, 111, 150, 138, 130, 134, 159, 181, 188, 129, 
    102, 51, 40, 115, 96, 58, 41, 78, 160, 181, 185, 207, 218, 210, 196, 206, 214, 180, 124, 113, 86, 102, 132, 160, 186, 167, 167, 167, 180, 179, 185, 156, 
    
    -- channel=14
    50, 64, 46, 30, 22, 36, 55, 57, 59, 54, 12, 18, 43, 44, 49, 50, 58, 77, 81, 77, 83, 78, 56, 57, 97, 93, 31, 58, 65, 41, 53, 66, 
    58, 81, 57, 29, 35, 61, 59, 60, 64, 47, 7, 27, 56, 62, 59, 47, 68, 74, 74, 68, 78, 81, 51, 60, 111, 96, 21, 39, 45, 44, 69, 66, 
    72, 87, 70, 35, 53, 72, 60, 65, 69, 38, 7, 35, 52, 65, 48, 33, 67, 66, 50, 55, 77, 82, 45, 62, 116, 99, 16, 38, 63, 75, 77, 51, 
    94, 76, 80, 47, 71, 72, 65, 74, 72, 30, 12, 34, 40, 52, 35, 30, 75, 87, 68, 69, 81, 77, 46, 67, 119, 107, 42, 73, 95, 96, 68, 34, 
    97, 79, 106, 60, 75, 68, 72, 76, 73, 24, 12, 17, 28, 37, 51, 59, 72, 79, 75, 71, 71, 73, 45, 77, 128, 129, 82, 85, 94, 97, 73, 80, 
    82, 77, 75, 67, 61, 69, 77, 61, 67, 19, 13, 22, 44, 59, 71, 73, 72, 72, 73, 53, 34, 73, 62, 77, 136, 147, 96, 91, 92, 110, 104, 92, 
    72, 70, 25, 51, 62, 79, 79, 50, 56, 15, 24, 54, 73, 75, 77, 62, 34, 51, 96, 42, 22, 88, 72, 74, 149, 161, 104, 108, 107, 131, 81, 43, 
    63, 59, 21, 70, 77, 72, 75, 58, 41, 8, 47, 81, 75, 75, 62, 18, 6, 39, 89, 64, 42, 94, 72, 83, 131, 162, 114, 120, 118, 133, 52, 21, 
    73, 53, 49, 104, 121, 88, 57, 70, 51, 23, 71, 83, 78, 79, 34, 7, 40, 81, 60, 62, 80, 99, 91, 93, 115, 141, 120, 121, 121, 124, 33, 20, 
    86, 58, 56, 118, 131, 127, 64, 51, 59, 64, 97, 99, 94, 58, 13, 28, 83, 93, 73, 80, 98, 105, 95, 74, 116, 132, 119, 126, 127, 101, 13, 23, 
    91, 59, 53, 116, 132, 135, 103, 48, 32, 75, 96, 97, 102, 74, 50, 73, 90, 82, 89, 97, 98, 108, 71, 49, 119, 124, 119, 138, 123, 91, 10, 20, 
    101, 51, 47, 110, 129, 135, 135, 72, 46, 84, 82, 79, 94, 86, 117, 135, 120, 102, 93, 94, 92, 88, 74, 88, 132, 115, 118, 141, 119, 91, 11, 7, 
    88, 40, 40, 96, 107, 131, 139, 119, 107, 102, 87, 89, 95, 74, 81, 108, 118, 110, 100, 93, 102, 85, 87, 95, 124, 120, 101, 113, 123, 89, 15, 32, 
    95, 63, 55, 92, 100, 110, 139, 137, 123, 97, 101, 92, 90, 88, 86, 86, 85, 88, 100, 108, 114, 108, 110, 95, 109, 117, 107, 115, 128, 88, 49, 76, 
    106, 69, 71, 96, 104, 86, 134, 135, 116, 87, 81, 88, 96, 96, 110, 106, 98, 95, 87, 92, 97, 107, 127, 128, 122, 94, 116, 119, 122, 92, 53, 70, 
    96, 64, 64, 92, 103, 95, 121, 133, 129, 150, 100, 51, 88, 101, 98, 113, 131, 119, 101, 95, 96, 83, 113, 152, 148, 120, 98, 124, 118, 57, 13, 72, 
    87, 76, 71, 90, 115, 124, 120, 130, 110, 142, 150, 58, 84, 116, 119, 120, 108, 113, 133, 134, 137, 126, 103, 110, 159, 163, 99, 114, 117, 42, 33, 107, 
    86, 88, 100, 93, 117, 99, 117, 105, 110, 102, 155, 139, 107, 111, 129, 129, 124, 119, 109, 118, 113, 118, 124, 113, 131, 117, 131, 99, 105, 72, 39, 87, 
    95, 96, 120, 115, 109, 71, 99, 86, 108, 99, 106, 176, 130, 94, 123, 117, 137, 141, 129, 136, 131, 111, 120, 121, 117, 107, 80, 67, 72, 81, 67, 110, 
    109, 112, 125, 87, 88, 72, 71, 94, 100, 121, 73, 115, 152, 118, 135, 148, 133, 130, 148, 149, 125, 113, 121, 122, 114, 113, 58, 78, 61, 56, 115, 138, 
    119, 116, 89, 67, 88, 72, 60, 102, 72, 87, 109, 55, 101, 146, 141, 156, 152, 136, 140, 152, 134, 123, 127, 124, 109, 105, 93, 98, 77, 98, 122, 119, 
    126, 97, 50, 93, 96, 70, 75, 96, 90, 59, 118, 97, 73, 131, 162, 151, 150, 163, 132, 127, 125, 118, 110, 117, 105, 102, 94, 79, 107, 142, 112, 106, 
    112, 81, 55, 89, 92, 78, 69, 89, 119, 107, 83, 118, 107, 125, 151, 156, 148, 155, 148, 126, 108, 123, 120, 117, 114, 102, 84, 86, 129, 121, 99, 105, 
    98, 86, 120, 154, 119, 95, 69, 78, 115, 126, 87, 78, 125, 139, 132, 150, 141, 142, 146, 126, 121, 132, 118, 123, 115, 88, 82, 111, 121, 101, 106, 103, 
    116, 136, 167, 182, 159, 119, 96, 92, 102, 90, 102, 111, 112, 136, 131, 143, 134, 142, 150, 128, 117, 156, 132, 119, 102, 89, 78, 83, 106, 96, 113, 108, 
    108, 109, 113, 146, 166, 158, 123, 105, 102, 82, 85, 140, 145, 126, 134, 123, 104, 115, 138, 137, 131, 150, 138, 106, 97, 111, 74, 45, 96, 101, 105, 75, 
    88, 85, 55, 86, 139, 151, 151, 126, 104, 104, 87, 87, 111, 110, 110, 82, 53, 75, 121, 140, 145, 120, 129, 122, 116, 98, 62, 32, 97, 98, 65, 64, 
    82, 92, 34, 32, 75, 117, 134, 156, 141, 109, 98, 87, 82, 90, 91, 95, 82, 70, 121, 139, 129, 143, 128, 107, 113, 78, 29, 63, 99, 71, 71, 66, 
    90, 86, 35, 13, 15, 78, 114, 148, 162, 139, 111, 98, 97, 91, 86, 113, 120, 106, 115, 126, 118, 135, 135, 106, 79, 42, 38, 91, 44, 96, 153, 83, 
    92, 86, 45, 37, 13, 31, 87, 122, 150, 173, 158, 122, 117, 114, 93, 92, 77, 85, 103, 113, 126, 133, 115, 91, 78, 50, 59, 60, 42, 108, 134, 98, 
    82, 71, 24, 56, 36, 23, 35, 84, 118, 146, 165, 165, 150, 130, 111, 121, 108, 66, 63, 98, 78, 69, 70, 86, 117, 108, 96, 98, 120, 116, 123, 89, 
    65, 27, 17, 64, 52, 29, 15, 37, 89, 100, 116, 150, 170, 152, 136, 156, 166, 121, 69, 74, 47, 71, 102, 127, 156, 139, 131, 130, 147, 136, 146, 117, 
    
    -- channel=15
    179, 139, 77, 88, 141, 157, 156, 151, 156, 158, 144, 151, 151, 136, 121, 118, 126, 108, 84, 84, 98, 98, 94, 83, 90, 86, 84, 96, 117, 87, 76, 77, 
    184, 133, 128, 146, 159, 159, 158, 167, 165, 162, 153, 154, 150, 150, 136, 125, 129, 109, 90, 82, 93, 98, 94, 88, 78, 76, 91, 106, 118, 98, 91, 90, 
    180, 152, 176, 170, 164, 152, 155, 164, 162, 170, 162, 159, 156, 151, 146, 140, 146, 124, 88, 71, 85, 98, 103, 107, 101, 109, 111, 111, 111, 101, 93, 95, 
    175, 174, 184, 181, 168, 152, 164, 163, 166, 179, 167, 168, 174, 162, 159, 164, 151, 137, 89, 58, 72, 90, 99, 107, 117, 128, 125, 121, 105, 97, 109, 111, 
    175, 174, 167, 172, 162, 161, 176, 175, 178, 178, 179, 180, 176, 168, 160, 164, 173, 156, 120, 69, 66, 90, 99, 94, 105, 124, 127, 123, 112, 104, 113, 116, 
    181, 174, 144, 170, 169, 166, 176, 179, 180, 180, 180, 181, 176, 174, 159, 150, 181, 175, 155, 116, 96, 125, 131, 112, 117, 120, 122, 121, 121, 120, 118, 124, 
    192, 156, 138, 178, 175, 174, 176, 175, 184, 180, 186, 184, 187, 187, 173, 153, 166, 173, 173, 167, 150, 149, 148, 121, 115, 117, 109, 111, 120, 122, 123, 128, 
    185, 125, 156, 171, 173, 175, 175, 184, 188, 183, 193, 194, 189, 185, 184, 166, 164, 172, 177, 176, 170, 137, 143, 122, 107, 110, 96, 103, 117, 118, 123, 125, 
    155, 149, 159, 160, 172, 173, 178, 180, 187, 186, 186, 191, 187, 175, 172, 160, 154, 151, 166, 176, 183, 155, 166, 133, 104, 104, 112, 119, 118, 122, 122, 125, 
    154, 152, 147, 169, 178, 178, 183, 170, 176, 188, 198, 193, 174, 167, 165, 169, 157, 140, 146, 169, 179, 160, 171, 141, 95, 104, 117, 119, 116, 123, 118, 125, 
    134, 112, 159, 177, 174, 184, 184, 186, 186, 194, 191, 176, 155, 158, 167, 187, 174, 147, 134, 151, 160, 156, 155, 124, 74, 102, 105, 102, 107, 117, 123, 127, 
    65, 91, 174, 157, 147, 177, 191, 190, 188, 176, 172, 176, 184, 174, 148, 163, 176, 154, 133, 149, 152, 149, 131, 80, 66, 97, 103, 102, 103, 113, 120, 125, 
    21, 92, 191, 177, 188, 202, 189, 182, 179, 156, 165, 188, 200, 174, 152, 114, 95, 127, 120, 137, 151, 136, 114, 78, 64, 73, 89, 98, 98, 113, 117, 118, 
    44, 99, 168, 173, 200, 195, 188, 187, 165, 149, 180, 194, 185, 168, 168, 154, 107, 146, 145, 138, 156, 127, 100, 72, 57, 64, 83, 96, 98, 106, 108, 111, 
    105, 118, 117, 159, 196, 190, 180, 187, 173, 173, 198, 193, 171, 165, 180, 188, 174, 187, 173, 179, 160, 128, 105, 72, 67, 69, 87, 108, 99, 100, 97, 102, 
    138, 113, 104, 157, 198, 196, 180, 168, 180, 191, 203, 205, 210, 191, 196, 200, 192, 187, 188, 190, 168, 153, 113, 80, 70, 64, 96, 135, 120, 90, 90, 98, 
    150, 138, 115, 147, 190, 187, 176, 150, 171, 199, 211, 198, 211, 194, 190, 203, 191, 186, 184, 189, 190, 166, 100, 70, 47, 56, 106, 143, 149, 92, 74, 94, 
    155, 155, 146, 165, 189, 192, 191, 145, 156, 210, 169, 149, 192, 194, 178, 168, 169, 181, 170, 167, 154, 117, 67, 43, 34, 49, 104, 143, 156, 106, 63, 80, 
    165, 162, 138, 166, 196, 190, 186, 137, 116, 201, 157, 169, 210, 182, 128, 143, 124, 147, 127, 97, 82, 56, 47, 51, 43, 64, 105, 157, 157, 123, 57, 65, 
    169, 150, 120, 158, 190, 190, 190, 152, 60, 153, 188, 185, 195, 165, 144, 206, 177, 137, 101, 61, 55, 51, 71, 80, 55, 74, 110, 160, 176, 142, 54, 50, 
    170, 160, 150, 166, 186, 188, 186, 154, 32, 49, 126, 146, 155, 140, 140, 192, 204, 156, 97, 62, 73, 73, 82, 87, 58, 62, 107, 166, 188, 167, 72, 51, 
    178, 171, 151, 156, 181, 178, 163, 124, 36, 29, 40, 55, 78, 99, 101, 130, 144, 123, 95, 55, 52, 51, 60, 85, 78, 77, 102, 153, 187, 177, 89, 55, 
    181, 171, 146, 152, 169, 167, 149, 105, 79, 94, 66, 46, 47, 71, 92, 120, 90, 55, 56, 41, 35, 34, 30, 55, 82, 86, 97, 119, 173, 174, 106, 60, 
    177, 156, 158, 163, 156, 160, 148, 137, 143, 118, 102, 107, 110, 109, 125, 103, 47, 17, 16, 19, 24, 28, 14, 19, 43, 65, 96, 99, 140, 173, 133, 67, 
    158, 139, 167, 182, 151, 140, 171, 192, 172, 116, 133, 136, 146, 141, 127, 101, 65, 37, 32, 25, 24, 17, 10, 15, 20, 66, 97, 78, 98, 148, 156, 105, 
    160, 164, 174, 171, 158, 136, 148, 177, 184, 147, 169, 151, 127, 139, 142, 125, 103, 77, 63, 43, 33, 24, 17, 26, 31, 62, 72, 50, 72, 90, 120, 136, 
    160, 163, 167, 167, 177, 168, 140, 120, 171, 143, 118, 130, 123, 156, 166, 145, 124, 105, 91, 78, 76, 66, 56, 67, 70, 65, 65, 73, 100, 123, 81, 106, 
    156, 159, 140, 147, 180, 170, 153, 123, 139, 156, 115, 126, 131, 158, 168, 162, 127, 119, 123, 120, 112, 104, 105, 119, 116, 105, 104, 109, 122, 134, 92, 104, 
    164, 158, 123, 139, 173, 156, 141, 140, 141, 121, 130, 161, 151, 157, 166, 168, 144, 138, 143, 132, 129, 133, 138, 148, 143, 137, 134, 132, 120, 100, 115, 147, 
    142, 149, 144, 168, 167, 161, 158, 158, 165, 144, 151, 169, 161, 160, 158, 162, 153, 145, 137, 127, 141, 149, 150, 158, 159, 150, 148, 143, 123, 119, 139, 159, 
    152, 166, 179, 185, 167, 167, 170, 168, 167, 164, 173, 178, 169, 157, 137, 133, 146, 143, 140, 136, 140, 151, 152, 157, 166, 156, 153, 144, 133, 131, 144, 153, 
    159, 178, 183, 171, 139, 125, 145, 159, 162, 139, 149, 156, 158, 152, 131, 115, 132, 142, 148, 143, 144, 157, 156, 161, 167, 159, 148, 156, 156, 150, 153, 152, 
    
    -- channel=16
    118, 96, 49, 59, 96, 95, 84, 83, 95, 97, 83, 90, 92, 82, 75, 79, 91, 80, 59, 50, 55, 56, 56, 51, 60, 56, 51, 58, 76, 53, 47, 47, 
    130, 88, 89, 105, 108, 96, 93, 104, 101, 98, 90, 91, 84, 87, 79, 72, 82, 72, 61, 50, 55, 56, 55, 51, 43, 40, 53, 65, 75, 61, 58, 57, 
    132, 104, 129, 122, 108, 89, 95, 106, 98, 105, 98, 94, 85, 80, 79, 76, 85, 76, 54, 42, 51, 58, 63, 66, 60, 66, 67, 66, 67, 62, 56, 57, 
    129, 127, 136, 132, 112, 90, 104, 105, 101, 113, 101, 102, 103, 90, 87, 93, 79, 78, 51, 31, 42, 51, 57, 62, 70, 77, 75, 74, 60, 55, 67, 69, 
    128, 127, 121, 127, 109, 99, 114, 114, 111, 111, 112, 113, 108, 99, 89, 92, 94, 89, 78, 44, 39, 52, 56, 46, 53, 67, 71, 73, 66, 59, 69, 71, 
    137, 131, 104, 127, 118, 106, 113, 116, 115, 117, 116, 113, 109, 105, 90, 84, 106, 104, 103, 79, 58, 77, 82, 61, 62, 63, 67, 70, 73, 72, 70, 75, 
    152, 119, 102, 135, 122, 117, 115, 111, 121, 123, 124, 112, 115, 113, 102, 92, 100, 101, 109, 110, 92, 87, 91, 67, 62, 64, 56, 59, 69, 72, 74, 78, 
    147, 89, 120, 126, 120, 118, 114, 121, 128, 122, 124, 115, 115, 109, 108, 100, 101, 104, 109, 106, 102, 75, 87, 72, 59, 60, 46, 53, 66, 68, 73, 75, 
    118, 111, 120, 114, 119, 116, 117, 119, 128, 122, 111, 109, 115, 103, 97, 94, 94, 89, 97, 100, 109, 95, 114, 89, 62, 58, 64, 71, 70, 72, 72, 75, 
    119, 113, 105, 120, 124, 122, 123, 111, 118, 123, 125, 121, 118, 109, 101, 111, 105, 85, 82, 96, 106, 100, 122, 103, 61, 62, 71, 73, 71, 75, 68, 75, 
    100, 72, 114, 126, 120, 127, 124, 126, 127, 129, 128, 123, 121, 119, 120, 144, 131, 99, 79, 88, 95, 97, 108, 91, 46, 62, 61, 59, 64, 70, 73, 76, 
    34, 52, 127, 105, 93, 122, 132, 131, 129, 115, 120, 140, 166, 151, 116, 133, 141, 110, 86, 97, 96, 92, 86, 49, 42, 60, 62, 60, 62, 66, 69, 74, 
    4, 64, 142, 125, 140, 154, 140, 132, 127, 107, 123, 156, 178, 147, 119, 83, 64, 91, 83, 100, 111, 92, 77, 49, 41, 47, 55, 57, 59, 67, 66, 68, 
    24, 72, 122, 123, 156, 150, 143, 141, 119, 106, 143, 160, 151, 129, 128, 119, 77, 116, 115, 109, 123, 90, 68, 45, 35, 43, 51, 55, 59, 62, 58, 62, 
    69, 82, 74, 112, 150, 145, 134, 143, 131, 132, 161, 156, 125, 114, 133, 151, 145, 160, 146, 152, 129, 93, 75, 47, 47, 48, 56, 68, 60, 60, 54, 57, 
    87, 65, 59, 112, 152, 150, 134, 125, 143, 155, 167, 165, 155, 132, 143, 160, 162, 158, 159, 161, 137, 120, 84, 57, 51, 43, 64, 95, 81, 55, 54, 57, 
    88, 78, 64, 102, 144, 141, 129, 108, 139, 165, 175, 157, 158, 134, 134, 159, 154, 148, 147, 152, 154, 135, 73, 49, 30, 35, 75, 103, 111, 61, 44, 57, 
    86, 87, 87, 116, 143, 147, 145, 105, 128, 179, 133, 108, 145, 139, 122, 121, 125, 135, 124, 121, 114, 88, 42, 24, 19, 29, 73, 102, 117, 80, 39, 46, 
    92, 92, 77, 118, 156, 153, 145, 98, 92, 170, 116, 122, 165, 131, 75, 98, 76, 97, 85, 64, 54, 27, 17, 27, 26, 40, 69, 117, 127, 100, 36, 40, 
    94, 84, 60, 110, 156, 163, 155, 115, 39, 124, 148, 137, 149, 113, 87, 156, 120, 80, 61, 39, 39, 24, 34, 46, 31, 45, 69, 120, 153, 123, 34, 32, 
    97, 93, 89, 114, 150, 162, 152, 117, 13, 29, 100, 116, 115, 86, 73, 124, 134, 91, 47, 27, 49, 50, 49, 50, 25, 30, 66, 125, 162, 150, 56, 32, 
    106, 104, 87, 99, 141, 150, 129, 87, 15, 11, 22, 37, 54, 57, 41, 62, 83, 72, 54, 26, 32, 35, 34, 51, 40, 43, 62, 112, 155, 158, 74, 31, 
    112, 104, 79, 90, 123, 137, 115, 66, 47, 66, 40, 23, 27, 38, 44, 69, 54, 31, 38, 29, 25, 22, 15, 31, 49, 51, 58, 78, 134, 148, 87, 31, 
    109, 88, 89, 96, 105, 129, 115, 94, 97, 71, 54, 60, 66, 62, 75, 60, 26, 10, 9, 14, 17, 19, 11, 12, 23, 31, 58, 59, 94, 136, 105, 35, 
    91, 70, 96, 112, 96, 104, 137, 147, 117, 58, 69, 67, 74, 69, 63, 53, 41, 25, 19, 13, 12, 9, 13, 18, 12, 36, 62, 39, 52, 104, 121, 71, 
    91, 92, 98, 98, 97, 86, 105, 134, 142, 107, 124, 97, 68, 73, 78, 73, 62, 43, 38, 28, 22, 14, 11, 20, 20, 42, 48, 20, 37, 56, 88, 100, 
    91, 94, 97, 98, 113, 111, 91, 76, 132, 110, 80, 81, 71, 95, 99, 84, 72, 61, 56, 51, 53, 43, 32, 43, 46, 40, 37, 40, 64, 90, 48, 66, 
    87, 96, 80, 82, 113, 109, 98, 72, 92, 115, 69, 70, 74, 94, 96, 88, 69, 71, 76, 74, 66, 60, 61, 75, 73, 64, 63, 65, 76, 94, 54, 58, 
    96, 97, 67, 76, 105, 90, 78, 80, 87, 72, 76, 98, 87, 92, 93, 90, 79, 84, 85, 70, 66, 72, 77, 87, 83, 82, 80, 79, 67, 53, 70, 94, 
    73, 84, 81, 101, 97, 91, 88, 91, 105, 89, 91, 99, 89, 93, 93, 90, 88, 85, 73, 60, 73, 82, 84, 91, 93, 86, 87, 85, 67, 68, 87, 100, 
    83, 96, 106, 113, 96, 95, 96, 95, 102, 105, 109, 104, 91, 90, 82, 74, 82, 78, 77, 74, 77, 85, 87, 92, 100, 89, 90, 84, 78, 77, 87, 90, 
    92, 107, 113, 104, 82, 66, 77, 92, 95, 81, 91, 90, 88, 91, 77, 61, 70, 77, 86, 82, 83, 92, 91, 96, 101, 92, 87, 91, 92, 90, 91, 87, 
    
    -- channel=17
    83, 61, 26, 36, 65, 67, 58, 54, 63, 65, 52, 59, 62, 53, 46, 52, 71, 65, 43, 39, 47, 47, 45, 38, 47, 45, 42, 50, 69, 46, 41, 41, 
    97, 53, 58, 70, 70, 67, 68, 77, 68, 65, 56, 57, 52, 57, 50, 46, 60, 52, 43, 38, 47, 47, 44, 40, 32, 30, 43, 56, 67, 53, 51, 49, 
    100, 71, 92, 81, 68, 57, 68, 78, 64, 71, 63, 59, 52, 48, 49, 48, 59, 50, 33, 30, 43, 48, 53, 56, 51, 56, 57, 56, 57, 53, 47, 49, 
    96, 95, 97, 89, 73, 55, 73, 72, 65, 78, 66, 66, 67, 55, 54, 63, 47, 46, 26, 18, 34, 41, 47, 53, 61, 68, 64, 62, 48, 45, 58, 60, 
    92, 97, 84, 87, 73, 63, 76, 75, 74, 74, 75, 75, 67, 59, 53, 59, 59, 52, 51, 30, 31, 41, 46, 39, 46, 59, 61, 61, 52, 48, 58, 60, 
    101, 102, 71, 89, 81, 70, 76, 76, 76, 81, 78, 71, 68, 67, 53, 49, 67, 65, 72, 57, 43, 62, 66, 50, 56, 54, 56, 58, 60, 61, 60, 65, 
    120, 89, 73, 99, 83, 80, 81, 75, 81, 87, 85, 66, 76, 79, 67, 53, 60, 64, 74, 77, 65, 64, 65, 47, 53, 54, 45, 48, 58, 61, 63, 66, 
    117, 59, 91, 91, 81, 81, 79, 84, 87, 86, 86, 72, 77, 76, 74, 63, 66, 73, 76, 73, 71, 47, 56, 47, 44, 49, 35, 42, 55, 57, 62, 64, 
    92, 84, 91, 81, 83, 79, 80, 80, 88, 83, 73, 70, 81, 72, 67, 61, 67, 65, 70, 70, 79, 64, 79, 60, 44, 45, 52, 59, 58, 61, 61, 64, 
    97, 88, 76, 90, 91, 86, 83, 71, 79, 82, 84, 83, 88, 83, 77, 85, 81, 62, 57, 70, 80, 72, 89, 75, 43, 49, 58, 60, 58, 63, 57, 64, 
    81, 48, 86, 98, 89, 91, 82, 84, 91, 84, 80, 80, 94, 101, 103, 126, 107, 73, 55, 67, 75, 76, 81, 68, 32, 49, 47, 45, 51, 58, 62, 65, 
    20, 31, 99, 77, 64, 86, 90, 90, 95, 69, 69, 95, 143, 136, 103, 121, 118, 82, 63, 80, 82, 77, 66, 33, 33, 48, 48, 46, 48, 54, 59, 63, 
    0, 50, 112, 92, 110, 122, 105, 98, 96, 72, 84, 119, 157, 125, 95, 73, 52, 71, 65, 84, 96, 79, 65, 42, 37, 37, 41, 41, 45, 56, 57, 58, 
    20, 60, 97, 92, 125, 120, 112, 111, 89, 76, 110, 128, 127, 100, 98, 108, 68, 99, 98, 91, 106, 76, 58, 41, 33, 35, 37, 38, 46, 52, 50, 53, 
    59, 70, 58, 88, 123, 117, 106, 115, 102, 103, 130, 125, 95, 80, 102, 137, 131, 140, 126, 132, 111, 78, 64, 42, 43, 40, 42, 50, 47, 50, 46, 49, 
    73, 53, 50, 94, 126, 124, 108, 98, 114, 125, 138, 136, 123, 98, 113, 140, 143, 137, 138, 140, 117, 105, 73, 51, 47, 35, 50, 77, 67, 45, 45, 50, 
    72, 65, 58, 86, 119, 117, 105, 83, 110, 137, 147, 130, 130, 107, 109, 135, 132, 127, 126, 131, 135, 119, 61, 42, 26, 27, 60, 85, 97, 51, 36, 51, 
    71, 72, 81, 102, 120, 124, 122, 80, 99, 151, 106, 84, 124, 121, 101, 92, 99, 115, 104, 101, 94, 72, 31, 17, 14, 21, 58, 85, 104, 70, 31, 41, 
    79, 78, 68, 100, 134, 136, 125, 75, 71, 147, 91, 97, 142, 113, 55, 72, 53, 79, 69, 50, 42, 20, 13, 22, 20, 35, 55, 96, 111, 91, 30, 35, 
    81, 72, 50, 88, 135, 153, 138, 93, 31, 111, 127, 113, 124, 92, 71, 141, 103, 65, 51, 33, 36, 25, 36, 44, 26, 43, 54, 96, 137, 115, 30, 26, 
    83, 82, 79, 95, 130, 150, 134, 98, 10, 23, 86, 99, 101, 76, 66, 116, 122, 78, 39, 23, 46, 47, 47, 46, 20, 27, 52, 103, 146, 137, 47, 25, 
    92, 92, 78, 83, 123, 135, 110, 70, 12, 8, 16, 29, 47, 52, 37, 56, 70, 57, 43, 18, 25, 28, 29, 44, 33, 38, 49, 94, 140, 141, 61, 24, 
    97, 93, 70, 78, 107, 118, 96, 48, 37, 58, 34, 19, 19, 31, 38, 59, 39, 19, 27, 18, 17, 17, 10, 24, 42, 44, 48, 64, 120, 128, 70, 24, 
    94, 77, 82, 88, 91, 107, 95, 75, 74, 55, 48, 57, 58, 53, 67, 51, 16, 4, 3, 8, 14, 19, 7, 6, 17, 23, 48, 47, 81, 115, 87, 27, 
    75, 59, 87, 105, 83, 82, 117, 126, 85, 34, 57, 62, 66, 61, 57, 46, 36, 23, 18, 13, 15, 14, 12, 14, 7, 28, 54, 30, 40, 85, 104, 62, 
    77, 77, 81, 86, 85, 69, 87, 112, 111, 79, 100, 79, 59, 67, 69, 58, 51, 38, 32, 21, 17, 12, 6, 14, 15, 34, 41, 15, 31, 46, 76, 90, 
    79, 81, 82, 85, 101, 96, 74, 57, 109, 87, 58, 62, 61, 88, 90, 68, 59, 53, 47, 42, 44, 35, 24, 35, 38, 29, 27, 31, 57, 82, 39, 56, 
    76, 87, 74, 74, 102, 95, 83, 57, 77, 99, 55, 58, 63, 84, 87, 77, 57, 60, 67, 68, 59, 49, 49, 63, 60, 49, 48, 51, 63, 84, 45, 47, 
    85, 90, 64, 69, 94, 78, 65, 68, 76, 60, 66, 90, 74, 78, 83, 81, 67, 71, 76, 64, 59, 57, 62, 72, 68, 66, 64, 62, 50, 41, 61, 83, 
    61, 75, 73, 92, 87, 81, 78, 80, 93, 76, 80, 89, 74, 76, 78, 80, 74, 69, 62, 53, 64, 66, 68, 75, 77, 72, 72, 68, 50, 56, 78, 89, 
    70, 81, 90, 100, 86, 85, 87, 85, 86, 87, 93, 90, 74, 70, 63, 60, 66, 60, 62, 62, 65, 70, 71, 76, 85, 77, 78, 71, 62, 65, 77, 79, 
    79, 93, 95, 89, 70, 57, 70, 81, 83, 64, 71, 71, 74, 76, 61, 47, 56, 63, 72, 70, 69, 76, 75, 80, 86, 79, 73, 78, 79, 76, 79, 73, 
    
    -- channel=18
    160, 185, 209, 217, 230, 246, 249, 246, 248, 243, 230, 221, 218, 221, 216, 199, 188, 187, 184, 180, 166, 144, 121, 139, 106, 102, 102, 79, 94, 101, 91, 94, 
    225, 239, 242, 230, 232, 245, 243, 235, 237, 230, 216, 205, 201, 203, 200, 186, 175, 171, 161, 127, 142, 141, 122, 135, 118, 82, 37, 52, 95, 107, 97, 100, 
    252, 249, 241, 220, 217, 226, 223, 214, 213, 207, 195, 184, 179, 182, 179, 167, 159, 152, 148, 129, 128, 140, 128, 114, 87, 40, 4, 38, 99, 115, 105, 105, 
    233, 225, 222, 211, 211, 203, 200, 192, 187, 183, 174, 164, 160, 165, 160, 153, 145, 141, 140, 138, 125, 125, 127, 105, 59, 37, 26, 55, 112, 120, 112, 109, 
    207, 195, 207, 201, 190, 180, 179, 171, 163, 159, 153, 146, 145, 151, 147, 141, 135, 136, 131, 135, 129, 122, 132, 90, 58, 61, 48, 86, 117, 120, 114, 109, 
    182, 171, 170, 162, 153, 156, 159, 151, 144, 141, 140, 138, 139, 141, 138, 138, 135, 140, 134, 138, 140, 137, 102, 69, 75, 62, 67, 116, 129, 128, 112, 110, 
    141, 136, 136, 134, 136, 134, 140, 133, 135, 137, 139, 141, 143, 146, 142, 145, 145, 145, 138, 143, 142, 107, 47, 33, 72, 75, 108, 127, 132, 132, 111, 112, 
    118, 125, 128, 129, 136, 131, 138, 132, 136, 140, 144, 147, 150, 158, 154, 153, 146, 149, 147, 148, 128, 66, 13, 17, 80, 117, 128, 122, 123, 128, 114, 112, 
    115, 126, 132, 133, 139, 135, 143, 137, 139, 145, 149, 152, 148, 154, 163, 170, 158, 162, 157, 148, 115, 44, 14, 30, 105, 139, 136, 126, 119, 122, 116, 111, 
    118, 128, 136, 136, 141, 136, 145, 141, 141, 147, 154, 165, 157, 154, 162, 167, 155, 147, 145, 138, 99, 56, 46, 55, 109, 124, 122, 126, 115, 116, 117, 110, 
    125, 132, 139, 137, 142, 136, 144, 140, 139, 144, 150, 153, 131, 139, 144, 152, 166, 186, 211, 214, 128, 92, 69, 42, 85, 95, 99, 115, 112, 111, 113, 107, 
    133, 137, 142, 138, 141, 136, 142, 138, 137, 143, 136, 132, 142, 182, 201, 203, 210, 206, 207, 192, 162, 189, 146, 42, 27, 40, 103, 114, 109, 106, 108, 104, 
    140, 139, 143, 139, 143, 140, 138, 137, 135, 133, 144, 164, 171, 160, 137, 115, 106, 93, 75, 59, 111, 220, 201, 95, 13, 7, 62, 116, 99, 101, 105, 100, 
    144, 138, 143, 140, 146, 146, 130, 135, 130, 145, 140, 110, 94, 92, 49, 19, 29, 50, 25, 18, 120, 209, 210, 157, 38, 6, 19, 68, 69, 82, 99, 95, 
    145, 139, 146, 142, 144, 142, 121, 128, 133, 127, 84, 68, 86, 82, 46, 22, 19, 50, 30, 65, 175, 201, 205, 203, 102, 16, 18, 22, 35, 56, 79, 88, 
    143, 139, 148, 144, 138, 132, 139, 131, 117, 66, 72, 86, 106, 78, 40, 34, 36, 70, 115, 182, 203, 197, 205, 195, 108, 61, 37, 18, 24, 79, 100, 83, 
    142, 139, 147, 144, 133, 114, 132, 121, 81, 89, 60, 69, 85, 68, 83, 155, 192, 219, 237, 235, 215, 215, 211, 114, 48, 93, 53, 20, 65, 139, 143, 84, 
    143, 141, 142, 137, 116, 69, 58, 67, 81, 75, 29, 28, 36, 25, 140, 242, 236, 235, 227, 220, 219, 223, 149, 58, 57, 84, 78, 78, 133, 161, 167, 91, 
    143, 140, 136, 134, 141, 71, 45, 52, 67, 33, 23, 22, 47, 41, 155, 217, 199, 190, 191, 208, 220, 223, 173, 103, 93, 115, 135, 149, 152, 148, 165, 89, 
    143, 140, 126, 181, 189, 76, 33, 43, 57, 21, 16, 23, 57, 66, 158, 194, 182, 179, 196, 201, 194, 206, 222, 179, 151, 156, 149, 151, 150, 146, 136, 66, 
    140, 133, 154, 234, 181, 90, 38, 42, 52, 11, 11, 11, 20, 49, 160, 186, 176, 185, 185, 115, 69, 90, 161, 196, 183, 170, 160, 153, 147, 136, 77, 38, 
    130, 128, 163, 163, 139, 106, 45, 46, 28, 3, 9, 15, 30, 54, 162, 180, 172, 190, 113, 21, 20, 21, 48, 149, 187, 171, 142, 133, 128, 67, 21, 39, 
    124, 132, 103, 26, 72, 108, 52, 48, 18, 7, 11, 59, 90, 99, 165, 176, 177, 169, 42, 29, 47, 38, 14, 70, 149, 136, 117, 117, 60, 14, 21, 48, 
    121, 124, 73, 30, 59, 114, 68, 31, 13, 14, 24, 72, 79, 108, 187, 187, 191, 139, 27, 43, 30, 27, 28, 27, 108, 132, 123, 89, 22, 21, 42, 59, 
    109, 102, 71, 63, 60, 113, 77, 28, 16, 31, 48, 71, 70, 136, 189, 179, 180, 116, 31, 54, 53, 41, 27, 14, 72, 133, 124, 60, 18, 34, 50, 59, 
    87, 81, 61, 60, 58, 105, 75, 21, 20, 46, 76, 96, 97, 145, 164, 163, 170, 113, 32, 57, 71, 49, 37, 17, 41, 108, 96, 33, 12, 29, 40, 50, 
    73, 73, 64, 60, 57, 95, 87, 47, 61, 98, 137, 165, 169, 176, 183, 182, 182, 124, 34, 54, 96, 92, 51, 27, 17, 70, 59, 12, 6, 18, 29, 40, 
    73, 73, 69, 78, 65, 89, 69, 47, 52, 60, 74, 86, 91, 96, 98, 96, 98, 83, 32, 60, 59, 62, 29, 20, 4, 17, 10, 3, 7, 10, 17, 33, 
    75, 83, 72, 54, 45, 39, 15, 4, 3, 2, 5, 7, 7, 8, 10, 11, 11, 13, 8, 66, 67, 47, 56, 15, 2, 2, 1, 3, 6, 10, 15, 32, 
    80, 89, 81, 47, 21, 10, 16, 25, 14, 10, 14, 14, 14, 14, 14, 12, 10, 9, 6, 23, 62, 72, 42, 7, 3, 4, 5, 5, 7, 11, 21, 33, 
    73, 79, 73, 55, 46, 47, 59, 58, 26, 17, 25, 28, 31, 32, 29, 28, 24, 21, 16, 12, 20, 22, 8, 6, 8, 7, 8, 8, 11, 15, 27, 31, 
    69, 72, 76, 78, 88, 83, 72, 56, 32, 38, 43, 42, 47, 51, 50, 49, 44, 38, 30, 28, 34, 34, 19, 12, 14, 16, 15, 13, 18, 26, 30, 29, 
    
    -- channel=19
    37, 49, 57, 58, 66, 78, 80, 81, 86, 82, 73, 66, 65, 67, 67, 56, 50, 50, 64, 115, 52, 56, 50, 39, 22, 34, 46, 36, 29, 18, 21, 19, 
    67, 72, 77, 68, 67, 74, 72, 66, 68, 64, 57, 52, 50, 54, 55, 46, 41, 42, 39, 41, 40, 35, 30, 33, 34, 46, 30, 27, 28, 21, 22, 18, 
    72, 68, 72, 62, 58, 61, 56, 49, 48, 45, 43, 40, 38, 42, 43, 38, 34, 35, 30, 28, 35, 33, 31, 34, 48, 34, 13, 14, 21, 20, 19, 17, 
    56, 54, 61, 60, 62, 48, 43, 36, 35, 35, 34, 32, 31, 33, 34, 32, 29, 30, 27, 29, 32, 28, 29, 37, 42, 18, 11, 15, 22, 19, 16, 17, 
    57, 57, 66, 59, 52, 36, 32, 27, 28, 29, 28, 26, 26, 26, 28, 30, 28, 28, 28, 28, 28, 48, 67, 42, 25, 18, 13, 25, 27, 31, 19, 17, 
    59, 58, 47, 33, 26, 26, 25, 22, 23, 25, 26, 25, 24, 24, 27, 31, 29, 30, 33, 30, 33, 93, 94, 60, 41, 27, 30, 44, 43, 45, 24, 19, 
    34, 28, 23, 20, 22, 23, 22, 21, 22, 22, 25, 26, 24, 25, 29, 35, 32, 31, 35, 30, 51, 89, 55, 37, 56, 40, 43, 45, 36, 30, 23, 21, 
    17, 17, 16, 18, 22, 23, 22, 22, 24, 23, 26, 27, 25, 27, 29, 39, 40, 45, 51, 48, 65, 64, 18, 11, 34, 37, 31, 32, 25, 22, 22, 21, 
    17, 18, 18, 18, 21, 22, 23, 23, 25, 24, 28, 30, 37, 56, 51, 59, 59, 58, 55, 54, 61, 40, 17, 16, 26, 25, 24, 27, 26, 23, 21, 20, 
    19, 18, 18, 18, 21, 20, 22, 24, 24, 25, 32, 49, 62, 76, 57, 52, 49, 46, 50, 58, 56, 49, 48, 44, 41, 35, 25, 25, 25, 24, 20, 20, 
    20, 18, 19, 18, 21, 21, 21, 23, 25, 25, 36, 53, 49, 66, 62, 74, 104, 137, 166, 184, 124, 104, 75, 33, 56, 61, 38, 25, 24, 25, 18, 19, 
    21, 18, 20, 19, 24, 24, 22, 24, 25, 29, 31, 48, 85, 151, 178, 190, 205, 205, 202, 197, 178, 208, 152, 22, 24, 37, 70, 40, 21, 22, 17, 17, 
    20, 20, 22, 21, 24, 24, 25, 26, 25, 32, 66, 112, 144, 155, 140, 117, 100, 88, 71, 61, 117, 232, 213, 78, 15, 10, 50, 70, 26, 21, 17, 16, 
    20, 22, 25, 22, 23, 23, 25, 26, 26, 72, 103, 91, 80, 86, 52, 18, 17, 34, 15, 16, 124, 221, 224, 155, 36, 7, 22, 59, 33, 19, 18, 16, 
    24, 23, 27, 22, 24, 25, 19, 21, 55, 85, 58, 41, 61, 78, 50, 24, 11, 43, 30, 73, 191, 216, 209, 205, 103, 14, 16, 23, 27, 22, 20, 18, 
    26, 22, 26, 23, 25, 37, 60, 52, 76, 52, 56, 59, 80, 77, 46, 38, 35, 73, 124, 196, 223, 216, 217, 210, 118, 57, 21, 14, 31, 71, 62, 17, 
    25, 20, 25, 23, 33, 53, 96, 92, 73, 93, 62, 66, 81, 71, 90, 162, 196, 223, 245, 245, 227, 228, 222, 121, 37, 59, 17, 9, 72, 140, 117, 19, 
    25, 21, 24, 26, 40, 44, 53, 69, 88, 82, 37, 41, 49, 32, 148, 251, 246, 242, 233, 226, 225, 226, 139, 31, 11, 25, 40, 67, 133, 162, 151, 34, 
    22, 19, 22, 38, 93, 70, 46, 54, 75, 38, 24, 27, 56, 49, 163, 227, 214, 205, 203, 218, 229, 228, 163, 74, 57, 90, 128, 149, 151, 150, 160, 51, 
    19, 15, 38, 124, 175, 90, 36, 42, 63, 23, 11, 21, 64, 79, 170, 208, 199, 197, 211, 214, 206, 217, 227, 177, 152, 168, 167, 162, 154, 151, 136, 42, 
    18, 10, 101, 220, 190, 111, 47, 46, 57, 10, 9, 14, 31, 66, 177, 204, 194, 202, 198, 124, 79, 102, 172, 211, 200, 184, 177, 169, 156, 140, 74, 17, 
    14, 20, 132, 165, 150, 128, 55, 52, 30, 3, 10, 22, 45, 72, 180, 198, 190, 205, 123, 25, 26, 30, 56, 163, 202, 184, 158, 147, 136, 68, 13, 17, 
    10, 35, 83, 33, 83, 130, 62, 53, 19, 7, 16, 72, 108, 117, 183, 194, 195, 183, 47, 30, 49, 43, 20, 79, 161, 148, 132, 129, 64, 10, 9, 24, 
    10, 33, 55, 35, 70, 136, 78, 36, 15, 17, 34, 88, 97, 126, 205, 205, 208, 152, 32, 43, 32, 31, 32, 31, 117, 145, 138, 99, 23, 12, 25, 33, 
    10, 21, 54, 65, 71, 136, 87, 33, 21, 39, 63, 87, 86, 154, 207, 197, 198, 129, 37, 56, 55, 44, 28, 15, 77, 147, 139, 67, 14, 20, 28, 31, 
    7, 14, 47, 62, 69, 128, 86, 28, 30, 60, 94, 111, 111, 162, 182, 180, 188, 127, 41, 60, 75, 53, 35, 15, 44, 122, 111, 38, 7, 13, 16, 22, 
    11, 17, 39, 59, 70, 117, 104, 61, 81, 121, 159, 183, 185, 195, 201, 199, 198, 136, 42, 60, 102, 98, 52, 28, 21, 79, 69, 16, 3, 7, 12, 22, 
    19, 20, 29, 67, 73, 103, 85, 60, 69, 80, 91, 100, 104, 113, 113, 109, 109, 89, 37, 65, 64, 66, 31, 23, 8, 20, 14, 5, 6, 6, 11, 24, 
    23, 28, 29, 37, 44, 44, 22, 7, 10, 10, 12, 12, 13, 16, 17, 16, 15, 15, 9, 67, 68, 48, 56, 16, 4, 3, 3, 4, 6, 9, 14, 25, 
    33, 37, 39, 32, 23, 18, 25, 32, 23, 21, 23, 23, 23, 21, 19, 15, 11, 10, 7, 24, 62, 71, 41, 8, 4, 5, 5, 6, 9, 14, 24, 29, 
    35, 37, 41, 50, 60, 67, 81, 77, 44, 36, 45, 48, 49, 44, 39, 35, 29, 27, 21, 16, 23, 25, 10, 9, 11, 9, 10, 11, 14, 20, 31, 30, 
    42, 42, 59, 87, 109, 111, 102, 82, 55, 62, 69, 71, 74, 72, 70, 67, 59, 51, 43, 41, 47, 44, 24, 18, 20, 22, 21, 19, 22, 28, 32, 30, 
    
    -- channel=20
    13, 11, 14, 10, 9, 10, 5, 2, 3, 3, 1, 2, 4, 6, 5, 0, 1, 0, 35, 86, 22, 23, 29, 8, 13, 27, 39, 29, 19, 8, 6, 5, 
    13, 12, 10, 4, 7, 8, 3, 0, 4, 2, 1, 1, 2, 4, 4, 1, 1, 1, 16, 19, 7, 6, 6, 7, 33, 46, 23, 22, 19, 8, 4, 6, 
    7, 4, 3, 0, 4, 4, 1, 0, 4, 4, 4, 4, 4, 6, 5, 3, 4, 3, 12, 9, 4, 7, 6, 10, 40, 35, 13, 12, 15, 6, 3, 6, 
    1, 3, 8, 11, 18, 4, 3, 3, 5, 6, 8, 7, 8, 9, 6, 6, 7, 5, 10, 9, 4, 10, 16, 23, 30, 22, 17, 14, 15, 6, 5, 8, 
    12, 19, 29, 26, 23, 6, 7, 8, 7, 8, 9, 8, 9, 10, 7, 8, 9, 7, 8, 7, 8, 37, 64, 39, 16, 16, 14, 21, 14, 15, 13, 9, 
    24, 30, 22, 12, 9, 6, 9, 8, 5, 5, 9, 10, 11, 10, 7, 9, 10, 11, 11, 7, 20, 85, 93, 59, 34, 14, 19, 32, 23, 27, 16, 9, 
    12, 11, 10, 7, 8, 8, 10, 7, 6, 5, 10, 14, 13, 12, 10, 12, 9, 14, 14, 7, 37, 86, 60, 40, 53, 28, 28, 28, 20, 16, 6, 7, 
    3, 6, 6, 7, 11, 10, 12, 9, 9, 8, 12, 14, 14, 18, 16, 19, 16, 21, 26, 22, 49, 62, 20, 10, 30, 26, 16, 13, 9, 8, 4, 7, 
    7, 10, 9, 8, 11, 10, 14, 11, 13, 12, 14, 15, 19, 36, 34, 40, 36, 32, 34, 34, 51, 43, 15, 9, 20, 12, 9, 10, 8, 8, 8, 8, 
    12, 12, 11, 8, 12, 10, 14, 13, 14, 14, 20, 34, 39, 49, 40, 38, 32, 27, 39, 50, 54, 59, 52, 38, 35, 21, 11, 12, 6, 9, 11, 10, 
    12, 11, 11, 9, 12, 10, 13, 13, 13, 16, 27, 40, 32, 50, 50, 63, 88, 119, 161, 180, 121, 113, 84, 34, 50, 49, 29, 17, 9, 10, 12, 10, 
    9, 10, 14, 11, 14, 12, 13, 12, 12, 18, 24, 39, 77, 147, 175, 186, 200, 200, 210, 202, 177, 213, 158, 28, 19, 34, 70, 37, 10, 9, 11, 9, 
    8, 10, 15, 13, 16, 14, 13, 14, 12, 24, 62, 108, 142, 162, 147, 125, 110, 94, 84, 74, 126, 241, 215, 84, 12, 9, 52, 73, 25, 13, 9, 8, 
    11, 11, 15, 14, 17, 16, 12, 14, 20, 68, 103, 93, 86, 95, 61, 25, 22, 35, 17, 23, 137, 235, 235, 167, 42, 7, 23, 66, 40, 17, 9, 7, 
    15, 13, 18, 14, 16, 18, 11, 18, 54, 83, 59, 46, 68, 83, 55, 27, 12, 39, 28, 76, 200, 232, 231, 224, 115, 22, 19, 26, 31, 22, 13, 8, 
    16, 13, 19, 14, 14, 30, 57, 55, 79, 53, 57, 60, 82, 78, 50, 41, 35, 71, 124, 200, 231, 230, 236, 221, 126, 68, 26, 14, 32, 73, 63, 9, 
    17, 14, 19, 17, 24, 47, 93, 92, 79, 98, 60, 61, 76, 71, 94, 166, 198, 226, 250, 252, 237, 240, 231, 124, 42, 74, 28, 12, 76, 149, 126, 17, 
    18, 16, 18, 21, 36, 42, 56, 72, 96, 88, 36, 36, 45, 34, 154, 256, 250, 249, 244, 237, 237, 238, 150, 39, 21, 46, 59, 77, 142, 174, 163, 38, 
    17, 16, 16, 34, 92, 73, 60, 66, 84, 44, 28, 33, 62, 55, 174, 240, 225, 217, 217, 231, 239, 238, 177, 86, 69, 106, 146, 164, 164, 161, 169, 55, 
    13, 10, 32, 125, 180, 98, 53, 56, 72, 28, 14, 27, 73, 89, 185, 224, 213, 213, 228, 227, 215, 225, 242, 192, 165, 180, 181, 176, 166, 159, 141, 42, 
    12, 7, 101, 229, 201, 123, 62, 57, 65, 15, 9, 15, 38, 79, 191, 218, 208, 219, 216, 138, 88, 109, 184, 228, 218, 201, 191, 181, 166, 147, 77, 14, 
    13, 24, 139, 179, 162, 141, 69, 61, 35, 4, 11, 27, 54, 86, 194, 212, 204, 219, 136, 36, 32, 34, 64, 177, 221, 204, 173, 159, 144, 73, 15, 13, 
    9, 39, 91, 49, 96, 143, 76, 62, 21, 7, 21, 81, 121, 131, 197, 208, 209, 193, 56, 38, 55, 46, 25, 89, 178, 169, 149, 141, 72, 14, 8, 20, 
    5, 34, 59, 48, 83, 149, 92, 45, 15, 19, 42, 100, 111, 140, 219, 219, 222, 160, 38, 51, 37, 35, 36, 39, 130, 164, 155, 110, 29, 12, 22, 30, 
    7, 23, 58, 77, 84, 148, 101, 42, 22, 43, 74, 101, 100, 168, 221, 211, 212, 137, 43, 64, 63, 52, 35, 21, 86, 162, 154, 78, 19, 18, 24, 28, 
    9, 21, 55, 76, 82, 140, 101, 37, 33, 67, 108, 127, 126, 176, 195, 194, 201, 135, 48, 70, 86, 65, 46, 21, 50, 131, 123, 49, 11, 10, 11, 20, 
    11, 23, 49, 73, 87, 132, 120, 75, 93, 134, 177, 200, 200, 207, 212, 213, 214, 148, 53, 72, 113, 110, 64, 34, 24, 85, 76, 22, 7, 9, 13, 22, 
    15, 22, 37, 78, 87, 115, 96, 72, 82, 93, 105, 114, 119, 125, 126, 123, 124, 102, 48, 76, 75, 78, 41, 27, 9, 24, 16, 6, 8, 10, 15, 25, 
    21, 31, 35, 43, 50, 48, 25, 12, 14, 14, 17, 17, 20, 24, 26, 25, 24, 20, 13, 74, 78, 59, 65, 18, 3, 5, 4, 3, 5, 9, 13, 26, 
    33, 40, 44, 37, 30, 23, 30, 37, 28, 25, 28, 28, 27, 24, 23, 19, 15, 9, 6, 28, 71, 83, 47, 8, 2, 5, 5, 4, 6, 11, 21, 28, 
    37, 41, 48, 59, 73, 79, 92, 89, 56, 47, 56, 59, 57, 48, 43, 40, 35, 27, 21, 21, 33, 37, 16, 8, 8, 9, 10, 10, 13, 18, 29, 28, 
    44, 49, 70, 101, 128, 128, 118, 99, 71, 78, 84, 85, 87, 83, 81, 79, 71, 60, 49, 49, 58, 56, 32, 19, 19, 24, 24, 21, 25, 31, 34, 28, 
    
    -- channel=21
    83, 82, 81, 77, 81, 85, 91, 92, 92, 95, 101, 92, 87, 82, 80, 76, 68, 65, 63, 62, 60, 56, 52, 47, 42, 37, 35, 34, 36, 29, 25, 21, 
    84, 83, 83, 77, 80, 84, 90, 93, 90, 88, 95, 97, 88, 82, 78, 76, 71, 68, 64, 66, 61, 54, 52, 46, 42, 38, 36, 35, 36, 30, 29, 31, 
    82, 81, 80, 75, 75, 84, 88, 76, 82, 86, 87, 99, 101, 88, 77, 76, 73, 68, 64, 64, 58, 55, 52, 45, 43, 40, 41, 44, 49, 48, 49, 53, 
    83, 81, 80, 78, 74, 87, 80, 50, 85, 97, 87, 91, 104, 102, 88, 80, 73, 64, 63, 63, 59, 56, 57, 58, 61, 63, 68, 71, 73, 71, 69, 69, 
    79, 79, 79, 79, 74, 83, 76, 55, 83, 84, 75, 75, 78, 89, 90, 87, 83, 66, 67, 70, 78, 80, 84, 87, 87, 86, 89, 89, 88, 84, 79, 73, 
    76, 74, 75, 77, 73, 73, 70, 70, 70, 69, 71, 73, 75, 78, 78, 81, 90, 89, 96, 98, 100, 104, 102, 104, 99, 95, 97, 94, 87, 80, 73, 66, 
    74, 72, 71, 73, 74, 62, 43, 51, 68, 64, 68, 71, 75, 74, 81, 94, 96, 98, 110, 114, 102, 100, 104, 109, 99, 91, 85, 80, 76, 73, 70, 67, 
    71, 72, 71, 72, 71, 58, 42, 41, 57, 54, 58, 63, 65, 71, 82, 96, 105, 94, 93, 103, 103, 106, 108, 97, 93, 91, 84, 80, 80, 80, 79, 77, 
    73, 73, 75, 82, 88, 103, 87, 46, 56, 56, 69, 82, 81, 87, 90, 87, 98, 99, 94, 91, 97, 102, 106, 102, 94, 99, 97, 92, 89, 89, 91, 95, 
    86, 95, 109, 123, 136, 153, 104, 51, 60, 59, 73, 97, 101, 108, 102, 90, 95, 97, 97, 93, 93, 99, 105, 110, 103, 105, 108, 108, 109, 110, 110, 110, 
    127, 139, 150, 157, 160, 162, 87, 50, 67, 56, 53, 88, 101, 112, 107, 90, 94, 96, 94, 96, 96, 95, 96, 101, 104, 113, 125, 126, 123, 119, 116, 112, 
    152, 157, 159, 162, 160, 159, 90, 44, 72, 69, 58, 86, 103, 90, 97, 92, 90, 96, 95, 94, 99, 98, 87, 92, 97, 112, 131, 131, 127, 121, 116, 108, 
    155, 158, 160, 157, 152, 148, 114, 48, 68, 88, 94, 103, 115, 96, 88, 93, 89, 101, 98, 94, 99, 101, 84, 85, 105, 110, 125, 132, 127, 118, 107, 95, 
    148, 148, 149, 146, 144, 142, 136, 80, 47, 72, 94, 104, 114, 113, 92, 94, 93, 103, 97, 93, 96, 97, 85, 82, 107, 107, 111, 121, 112, 100, 87, 77, 
    134, 135, 138, 140, 142, 147, 151, 137, 93, 73, 50, 62, 89, 94, 90, 98, 102, 105, 103, 97, 94, 94, 86, 83, 95, 101, 92, 102, 95, 82, 74, 75, 
    131, 134, 139, 144, 152, 159, 154, 152, 158, 118, 53, 57, 103, 100, 95, 102, 110, 116, 111, 106, 97, 91, 87, 85, 84, 98, 85, 83, 83, 85, 90, 95, 
    135, 144, 152, 160, 164, 161, 137, 115, 157, 145, 128, 110, 123, 122, 104, 103, 105, 109, 108, 104, 97, 90, 88, 87, 79, 92, 87, 85, 101, 105, 105, 94, 
    148, 154, 159, 164, 170, 179, 176, 127, 176, 197, 157, 152, 113, 145, 128, 103, 103, 101, 104, 102, 97, 95, 91, 89, 79, 86, 91, 91, 109, 104, 86, 70, 
    155, 164, 178, 197, 221, 238, 248, 196, 156, 200, 176, 184, 108, 142, 137, 106, 100, 99, 100, 101, 101, 99, 95, 89, 80, 81, 92, 83, 88, 82, 73, 71, 
    191, 214, 235, 249, 253, 246, 251, 244, 160, 158, 172, 195, 113, 114, 139, 110, 98, 98, 97, 99, 103, 104, 102, 92, 83, 78, 85, 73, 75, 80, 74, 72, 
    245, 252, 253, 254, 243, 187, 186, 201, 145, 128, 151, 156, 116, 106, 128, 114, 104, 103, 101, 103, 108, 110, 105, 92, 82, 76, 84, 85, 78, 83, 77, 73, 
    251, 252, 252, 256, 233, 126, 107, 114, 105, 115, 120, 110, 99, 99, 104, 103, 109, 110, 107, 107, 112, 110, 96, 86, 78, 76, 90, 104, 91, 82, 82, 79, 
    248, 248, 246, 235, 200, 124, 114, 118, 93, 87, 83, 79, 80, 86, 75, 68, 95, 100, 98, 97, 98, 97, 97, 97, 91, 87, 91, 111, 110, 85, 82, 82, 
    235, 214, 181, 150, 138, 136, 133, 132, 100, 61, 57, 60, 67, 89, 96, 58, 51, 69, 71, 80, 94, 101, 104, 101, 93, 87, 94, 109, 119, 98, 81, 81, 
    153, 130, 122, 120, 124, 122, 111, 103, 106, 90, 57, 52, 69, 102, 106, 83, 64, 71, 77, 85, 100, 103, 102, 109, 106, 87, 93, 99, 113, 115, 92, 80, 
    109, 111, 114, 109, 101, 97, 102, 109, 117, 120, 103, 85, 93, 101, 95, 89, 74, 75, 82, 90, 114, 119, 105, 102, 111, 107, 94, 98, 101, 117, 107, 79, 
    105, 98, 93, 91, 99, 106, 111, 113, 112, 104, 97, 95, 80, 76, 84, 92, 81, 72, 79, 89, 117, 123, 105, 94, 96, 103, 103, 101, 96, 105, 111, 90, 
    87, 87, 94, 101, 108, 110, 107, 100, 91, 81, 86, 104, 93, 73, 76, 92, 88, 77, 79, 79, 91, 100, 93, 86, 87, 92, 97, 96, 96, 96, 102, 101, 
    90, 96, 103, 105, 101, 95, 86, 80, 81, 85, 96, 106, 98, 85, 96, 93, 88, 81, 79, 76, 71, 76, 84, 91, 92, 86, 83, 90, 98, 96, 91, 96, 
    100, 99, 95, 86, 80, 79, 79, 79, 82, 83, 98, 108, 99, 96, 97, 89, 92, 84, 79, 81, 76, 74, 82, 89, 90, 85, 82, 86, 93, 92, 83, 83, 
    87, 78, 73, 71, 77, 87, 89, 83, 81, 79, 97, 106, 100, 103, 89, 92, 96, 87, 88, 89, 82, 79, 84, 83, 86, 90, 86, 83, 86, 86, 79, 73, 
    62, 63, 70, 73, 84, 86, 83, 81, 78, 74, 94, 107, 95, 104, 91, 88, 91, 88, 88, 89, 85, 80, 85, 83, 84, 89, 86, 80, 76, 77, 76, 72, 
    
    -- channel=22
    94, 94, 93, 89, 90, 90, 96, 96, 97, 102, 110, 101, 94, 88, 85, 82, 78, 75, 73, 72, 69, 65, 61, 56, 51, 46, 41, 39, 40, 34, 29, 25, 
    96, 95, 95, 89, 89, 89, 95, 98, 97, 96, 106, 107, 96, 89, 85, 82, 79, 75, 71, 73, 68, 61, 59, 53, 49, 44, 39, 37, 38, 32, 31, 31, 
    94, 92, 92, 87, 84, 90, 93, 81, 89, 96, 99, 110, 112, 98, 86, 84, 79, 73, 68, 70, 63, 58, 54, 48, 46, 43, 41, 43, 47, 46, 48, 49, 
    95, 93, 92, 90, 83, 93, 86, 57, 93, 107, 99, 104, 116, 114, 101, 90, 78, 67, 66, 66, 62, 56, 56, 57, 60, 62, 65, 66, 67, 65, 63, 61, 
    92, 91, 91, 91, 83, 89, 82, 62, 92, 95, 88, 88, 92, 104, 105, 100, 91, 70, 69, 72, 80, 77, 80, 83, 83, 81, 81, 80, 79, 75, 70, 63, 
    88, 86, 87, 89, 82, 79, 76, 77, 80, 82, 85, 87, 90, 94, 94, 95, 99, 94, 98, 99, 100, 100, 96, 98, 93, 88, 88, 83, 76, 69, 62, 55, 
    85, 84, 82, 84, 81, 61, 42, 55, 83, 87, 88, 89, 91, 87, 93, 101, 98, 100, 112, 115, 105, 103, 103, 103, 91, 80, 78, 74, 68, 63, 57, 54, 
    82, 83, 82, 84, 76, 55, 38, 44, 76, 85, 82, 81, 80, 83, 91, 99, 103, 96, 97, 108, 109, 114, 113, 94, 82, 77, 77, 75, 71, 68, 64, 59, 
    81, 82, 84, 91, 94, 104, 85, 49, 73, 84, 91, 99, 97, 100, 101, 94, 101, 104, 101, 98, 106, 111, 114, 103, 87, 85, 82, 78, 74, 70, 71, 72, 
    92, 101, 115, 128, 142, 157, 104, 54, 75, 84, 93, 113, 117, 124, 117, 101, 103, 106, 107, 103, 104, 110, 116, 118, 100, 90, 85, 84, 85, 85, 85, 82, 
    130, 142, 153, 160, 166, 170, 89, 53, 80, 77, 70, 104, 119, 130, 127, 107, 106, 108, 105, 106, 106, 105, 110, 114, 105, 98, 98, 96, 94, 91, 89, 85, 
    154, 159, 162, 164, 167, 169, 93, 46, 81, 86, 74, 103, 123, 112, 122, 114, 106, 109, 106, 103, 107, 105, 103, 110, 102, 97, 101, 99, 96, 94, 90, 85, 
    157, 159, 161, 158, 158, 159, 117, 48, 73, 101, 108, 120, 135, 120, 116, 117, 107, 115, 108, 102, 105, 106, 100, 105, 112, 96, 96, 101, 98, 93, 85, 76, 
    153, 152, 151, 147, 147, 147, 135, 76, 44, 73, 103, 117, 131, 133, 115, 113, 108, 119, 113, 107, 106, 106, 101, 100, 117, 105, 93, 98, 93, 85, 74, 64, 
    143, 142, 142, 142, 143, 148, 149, 131, 84, 65, 53, 70, 99, 107, 104, 109, 114, 124, 125, 117, 110, 108, 101, 98, 108, 111, 88, 90, 85, 72, 65, 63, 
    140, 141, 142, 145, 153, 160, 153, 147, 151, 111, 52, 58, 106, 104, 101, 110, 123, 137, 135, 128, 115, 108, 104, 101, 99, 111, 89, 78, 74, 72, 74, 77, 
    143, 149, 155, 159, 164, 160, 136, 114, 155, 143, 122, 104, 118, 119, 102, 108, 120, 132, 133, 128, 117, 109, 107, 106, 97, 108, 98, 86, 90, 84, 79, 68, 
    154, 157, 159, 161, 167, 177, 176, 129, 179, 199, 151, 142, 104, 137, 123, 108, 121, 126, 131, 128, 119, 115, 112, 110, 99, 105, 106, 94, 92, 74, 52, 39, 
    157, 164, 176, 193, 218, 236, 247, 199, 163, 206, 173, 177, 101, 136, 134, 113, 119, 126, 130, 129, 125, 122, 118, 113, 104, 103, 106, 80, 62, 44, 37, 39, 
    192, 212, 232, 246, 250, 242, 250, 247, 169, 170, 174, 193, 110, 112, 139, 120, 118, 126, 128, 128, 128, 127, 126, 116, 108, 102, 96, 62, 42, 37, 39, 43, 
    245, 251, 250, 251, 241, 186, 190, 210, 161, 146, 156, 160, 125, 115, 135, 122, 120, 127, 129, 128, 127, 127, 125, 116, 106, 98, 87, 66, 45, 42, 41, 41, 
    251, 251, 251, 254, 234, 131, 116, 130, 127, 138, 130, 124, 122, 119, 114, 107, 118, 128, 130, 127, 125, 119, 111, 108, 99, 90, 82, 80, 61, 47, 44, 41, 
    252, 252, 249, 239, 203, 128, 123, 131, 111, 108, 102, 103, 106, 105, 81, 68, 102, 117, 120, 116, 110, 107, 112, 115, 104, 89, 75, 84, 81, 52, 45, 45, 
    245, 223, 191, 160, 144, 137, 137, 138, 109, 75, 81, 87, 90, 102, 99, 58, 58, 86, 95, 101, 109, 116, 122, 116, 97, 77, 70, 80, 89, 66, 47, 47, 
    165, 141, 134, 132, 130, 123, 112, 105, 107, 94, 74, 71, 83, 110, 111, 86, 72, 90, 102, 108, 118, 123, 123, 124, 108, 73, 66, 68, 82, 84, 61, 48, 
    117, 120, 122, 117, 106, 97, 101, 106, 112, 115, 106, 87, 92, 104, 104, 97, 84, 95, 108, 114, 134, 142, 130, 122, 119, 100, 69, 64, 69, 87, 79, 50, 
    108, 102, 96, 94, 101, 107, 110, 107, 103, 93, 86, 81, 66, 72, 93, 104, 94, 95, 107, 113, 137, 148, 133, 122, 114, 107, 81, 66, 64, 75, 85, 63, 
    88, 87, 93, 99, 107, 108, 101, 87, 73, 60, 65, 83, 74, 63, 78, 94, 89, 87, 95, 93, 105, 123, 122, 114, 109, 104, 78, 59, 60, 63, 74, 75, 
    93, 95, 97, 95, 91, 84, 69, 56, 50, 49, 66, 85, 83, 73, 85, 72, 62, 62, 67, 68, 69, 88, 100, 104, 101, 90, 64, 51, 53, 54, 58, 69, 
    96, 91, 81, 68, 59, 55, 52, 48, 47, 46, 64, 82, 82, 79, 77, 57, 53, 50, 52, 58, 58, 63, 71, 74, 72, 65, 52, 46, 48, 49, 48, 54, 
    73, 60, 49, 43, 44, 48, 52, 48, 48, 44, 58, 73, 75, 79, 62, 53, 50, 46, 52, 57, 52, 47, 51, 47, 47, 49, 46, 42, 43, 45, 43, 42, 
    41, 37, 39, 37, 42, 41, 41, 45, 47, 43, 54, 71, 67, 76, 59, 46, 43, 42, 45, 48, 47, 45, 49, 45, 43, 45, 42, 39, 37, 40, 40, 38, 
    
    -- channel=23
    85, 84, 83, 79, 80, 82, 93, 95, 90, 85, 79, 72, 75, 78, 84, 79, 68, 62, 60, 61, 60, 59, 56, 51, 46, 41, 37, 35, 36, 30, 25, 21, 
    86, 85, 85, 79, 78, 80, 90, 93, 84, 73, 70, 71, 68, 69, 71, 72, 70, 67, 62, 62, 56, 53, 52, 46, 41, 37, 34, 32, 33, 27, 26, 27, 
    84, 83, 82, 78, 73, 80, 86, 72, 70, 65, 56, 67, 72, 63, 54, 60, 66, 65, 61, 58, 48, 47, 45, 38, 36, 33, 34, 37, 42, 41, 42, 44, 
    85, 83, 82, 80, 72, 82, 77, 43, 67, 69, 50, 52, 65, 63, 50, 47, 50, 52, 57, 54, 45, 43, 43, 44, 47, 50, 56, 59, 60, 59, 56, 55, 
    82, 81, 81, 81, 72, 76, 70, 44, 61, 51, 34, 29, 31, 39, 38, 35, 41, 43, 57, 59, 61, 61, 65, 68, 68, 66, 71, 72, 71, 67, 62, 56, 
    77, 76, 76, 79, 71, 66, 62, 56, 44, 33, 26, 23, 22, 20, 15, 14, 31, 53, 79, 84, 83, 82, 78, 80, 76, 72, 77, 75, 68, 60, 53, 46, 
    73, 71, 70, 72, 71, 55, 32, 32, 38, 24, 20, 19, 18, 11, 14, 21, 24, 41, 70, 89, 86, 80, 79, 82, 75, 72, 72, 67, 59, 52, 45, 42, 
    68, 69, 68, 69, 67, 51, 28, 17, 23, 12, 10, 11, 9, 11, 17, 24, 28, 22, 33, 63, 77, 79, 77, 64, 65, 73, 72, 66, 60, 54, 47, 43, 
    68, 69, 71, 78, 82, 93, 70, 19, 18, 12, 25, 37, 32, 33, 33, 20, 22, 24, 25, 33, 49, 56, 60, 59, 59, 75, 73, 63, 57, 52, 52, 53, 
    80, 89, 103, 117, 128, 141, 85, 22, 21, 15, 33, 56, 57, 61, 53, 28, 21, 22, 22, 20, 24, 35, 45, 58, 61, 72, 70, 65, 65, 64, 63, 61, 
    119, 131, 142, 149, 152, 152, 71, 24, 30, 17, 21, 49, 60, 68, 63, 33, 25, 27, 21, 17, 15, 20, 28, 43, 55, 70, 77, 74, 73, 71, 68, 65, 
    143, 148, 150, 153, 153, 153, 79, 23, 40, 34, 25, 46, 61, 48, 55, 39, 29, 36, 31, 21, 19, 21, 18, 31, 42, 59, 76, 77, 77, 76, 74, 69, 
    146, 149, 151, 148, 146, 146, 107, 32, 43, 55, 52, 59, 71, 52, 44, 41, 34, 50, 44, 30, 26, 28, 18, 25, 46, 50, 69, 81, 81, 79, 73, 66, 
    144, 143, 143, 139, 138, 137, 126, 64, 26, 46, 61, 65, 70, 64, 40, 36, 36, 54, 51, 40, 33, 29, 18, 19, 47, 51, 60, 78, 79, 74, 64, 55, 
    133, 132, 134, 134, 134, 136, 137, 119, 71, 49, 27, 33, 46, 42, 32, 34, 40, 57, 61, 50, 39, 28, 17, 17, 36, 51, 48, 65, 70, 62, 54, 50, 
    125, 127, 129, 133, 140, 145, 136, 129, 132, 90, 30, 30, 64, 51, 39, 39, 49, 69, 69, 61, 44, 28, 20, 19, 25, 48, 41, 45, 53, 57, 60, 61, 
    125, 132, 139, 145, 149, 145, 117, 90, 128, 114, 98, 80, 87, 77, 49, 40, 46, 63, 68, 60, 45, 31, 25, 23, 21, 42, 43, 45, 64, 66, 62, 50, 
    136, 140, 144, 147, 154, 164, 158, 104, 149, 166, 122, 119, 80, 103, 75, 41, 45, 56, 65, 60, 48, 40, 31, 27, 21, 35, 47, 50, 65, 57, 35, 20, 
    144, 151, 164, 182, 210, 230, 235, 178, 133, 171, 138, 149, 77, 103, 85, 45, 43, 56, 63, 60, 53, 48, 39, 29, 23, 29, 47, 39, 39, 31, 22, 21, 
    183, 205, 225, 240, 248, 242, 242, 230, 141, 132, 132, 159, 83, 77, 86, 49, 42, 55, 60, 58, 57, 55, 47, 33, 25, 26, 39, 28, 25, 29, 28, 27, 
    241, 248, 247, 249, 236, 176, 171, 181, 120, 98, 114, 118, 77, 60, 71, 52, 46, 54, 57, 58, 59, 57, 48, 32, 24, 23, 37, 37, 28, 32, 31, 26, 
    248, 249, 249, 253, 224, 106, 83, 85, 71, 78, 81, 65, 48, 46, 52, 49, 51, 55, 54, 57, 61, 51, 36, 27, 21, 22, 39, 54, 40, 31, 31, 28, 
    247, 248, 245, 235, 194, 109, 96, 94, 65, 53, 35, 25, 28, 43, 45, 32, 46, 51, 47, 47, 48, 45, 43, 41, 34, 30, 36, 58, 57, 33, 29, 30, 
    236, 215, 182, 152, 136, 129, 122, 116, 81, 35, 13, 9, 20, 52, 73, 34, 17, 28, 26, 32, 47, 59, 59, 49, 35, 26, 34, 52, 63, 44, 28, 29, 
    154, 130, 122, 120, 123, 118, 104, 92, 90, 70, 31, 18, 29, 61, 69, 52, 34, 36, 36, 40, 58, 71, 65, 61, 48, 23, 31, 40, 56, 60, 39, 28, 
    105, 107, 109, 104, 95, 88, 91, 93, 96, 98, 86, 62, 56, 56, 47, 49, 40, 37, 42, 48, 76, 91, 72, 57, 54, 44, 29, 35, 42, 61, 55, 29, 
    95, 89, 83, 81, 86, 88, 91, 88, 83, 73, 68, 62, 40, 35, 44, 52, 40, 30, 39, 49, 81, 95, 71, 50, 41, 42, 37, 35, 34, 48, 58, 40, 
    75, 73, 79, 85, 87, 83, 76, 64, 51, 39, 42, 59, 50, 34, 41, 49, 38, 30, 36, 39, 55, 69, 60, 45, 38, 38, 34, 29, 32, 36, 48, 51, 
    76, 78, 79, 77, 68, 57, 44, 33, 29, 30, 46, 61, 55, 41, 50, 38, 29, 26, 29, 30, 29, 37, 46, 48, 46, 37, 25, 24, 30, 32, 36, 47, 
    80, 74, 64, 50, 38, 32, 30, 27, 27, 27, 45, 60, 53, 47, 44, 29, 28, 23, 23, 28, 25, 24, 32, 37, 35, 29, 21, 21, 26, 30, 28, 34, 
    58, 45, 33, 26, 26, 29, 33, 28, 27, 24, 39, 51, 49, 50, 33, 28, 27, 21, 25, 29, 24, 21, 25, 23, 23, 26, 22, 18, 21, 26, 25, 23, 
    27, 23, 24, 21, 26, 25, 24, 25, 26, 22, 33, 48, 42, 51, 35, 24, 21, 20, 21, 24, 23, 23, 29, 25, 24, 27, 22, 18, 17, 22, 24, 22, 
    
    -- channel=24
    23, 19, 21, 65, 164, 188, 183, 178, 170, 172, 186, 186, 184, 183, 182, 183, 180, 164, 127, 92, 107, 110, 153, 194, 195, 201, 197, 198, 201, 200, 199, 197, 
    23, 19, 21, 46, 153, 202, 191, 178, 164, 158, 169, 183, 186, 184, 180, 178, 180, 173, 138, 86, 74, 106, 180, 206, 207, 213, 208, 206, 207, 205, 204, 202, 
    23, 20, 23, 31, 127, 200, 185, 168, 159, 158, 154, 162, 178, 178, 179, 178, 181, 190, 182, 125, 71, 114, 197, 209, 213, 216, 213, 211, 212, 211, 208, 206, 
    23, 21, 24, 23, 99, 189, 175, 160, 168, 168, 166, 149, 170, 186, 191, 195, 195, 200, 188, 141, 99, 146, 210, 214, 213, 212, 212, 213, 217, 217, 215, 214, 
    25, 23, 23, 21, 72, 170, 165, 151, 175, 183, 185, 155, 146, 157, 169, 188, 197, 196, 178, 141, 121, 172, 211, 219, 221, 217, 217, 217, 214, 212, 209, 206, 
    26, 27, 26, 23, 49, 143, 164, 154, 169, 194, 200, 166, 130, 125, 128, 151, 165, 165, 148, 143, 147, 182, 188, 201, 212, 217, 213, 219, 220, 215, 215, 211, 
    30, 26, 27, 25, 37, 125, 180, 171, 169, 197, 202, 179, 139, 113, 122, 130, 119, 133, 122, 140, 185, 203, 191, 201, 215, 218, 215, 219, 220, 218, 220, 224, 
    94, 48, 31, 36, 100, 175, 193, 168, 163, 192, 198, 195, 174, 145, 142, 132, 106, 121, 122, 139, 192, 209, 189, 213, 242, 237, 239, 232, 208, 213, 222, 229, 
    180, 158, 114, 122, 177, 190, 190, 160, 133, 173, 197, 200, 194, 185, 167, 146, 129, 129, 133, 141, 177, 201, 189, 220, 241, 235, 232, 213, 189, 199, 225, 234, 
    197, 192, 178, 186, 193, 195, 197, 157, 128, 163, 185, 191, 193, 195, 178, 151, 114, 129, 131, 134, 170, 194, 208, 234, 236, 240, 235, 201, 185, 187, 208, 235, 
    202, 196, 187, 192, 200, 205, 197, 151, 149, 175, 184, 189, 193, 187, 168, 136, 117, 128, 128, 129, 167, 181, 205, 240, 243, 243, 238, 206, 186, 187, 193, 221, 
    205, 205, 197, 192, 203, 208, 194, 160, 168, 191, 193, 191, 193, 172, 146, 119, 124, 142, 133, 135, 167, 176, 191, 234, 243, 241, 236, 215, 186, 184, 185, 196, 
    206, 204, 200, 193, 197, 199, 191, 180, 172, 179, 183, 173, 174, 174, 152, 131, 141, 166, 142, 154, 169, 172, 191, 230, 240, 241, 239, 228, 200, 186, 184, 192, 
    210, 202, 198, 191, 201, 180, 177, 202, 171, 154, 142, 142, 168, 168, 147, 156, 175, 169, 150, 164, 158, 160, 197, 230, 241, 241, 244, 242, 226, 191, 195, 215, 
    211, 201, 199, 192, 207, 170, 161, 215, 189, 186, 173, 172, 190, 177, 137, 127, 180, 174, 150, 160, 175, 176, 193, 236, 245, 242, 243, 251, 239, 201, 212, 225, 
    211, 196, 197, 193, 209, 181, 154, 217, 206, 197, 195, 185, 170, 173, 166, 152, 163, 184, 166, 152, 192, 181, 175, 204, 238, 243, 244, 247, 223, 213, 226, 226, 
    214, 194, 180, 181, 197, 196, 155, 198, 214, 192, 174, 183, 173, 161, 174, 178, 128, 164, 189, 147, 167, 180, 156, 118, 157, 215, 239, 235, 206, 214, 234, 228, 
    215, 198, 166, 163, 180, 202, 190, 185, 207, 210, 205, 214, 193, 174, 176, 173, 129, 137, 191, 153, 163, 200, 171, 135, 116, 144, 184, 193, 187, 210, 239, 235, 
    216, 205, 174, 164, 185, 203, 210, 194, 191, 211, 218, 226, 225, 203, 190, 179, 151, 121, 168, 158, 167, 194, 170, 172, 154, 131, 153, 169, 162, 184, 222, 236, 
    216, 208, 192, 180, 197, 202, 209, 210, 186, 189, 197, 204, 209, 213, 207, 181, 178, 149, 146, 175, 183, 174, 156, 171, 163, 148, 169, 180, 166, 160, 172, 204, 
    218, 213, 202, 182, 191, 203, 201, 202, 202, 195, 193, 192, 178, 198, 207, 199, 211, 203, 166, 187, 177, 155, 147, 166, 167, 171, 182, 175, 156, 156, 159, 167, 
    217, 215, 209, 186, 179, 200, 208, 200, 209, 215, 210, 186, 161, 182, 196, 194, 203, 207, 190, 185, 155, 142, 155, 166, 172, 179, 173, 159, 150, 158, 158, 143, 
    214, 213, 214, 192, 169, 197, 218, 217, 215, 217, 212, 195, 170, 179, 195, 191, 190, 192, 192, 170, 132, 142, 167, 170, 170, 179, 173, 157, 157, 147, 134, 125, 
    213, 209, 211, 202, 168, 193, 216, 222, 223, 222, 211, 205, 194, 194, 201, 198, 198, 196, 188, 153, 134, 155, 171, 167, 166, 189, 178, 165, 163, 142, 133, 137, 
    211, 206, 206, 202, 175, 191, 211, 213, 214, 216, 198, 171, 194, 206, 201, 201, 200, 197, 177, 150, 144, 158, 167, 157, 159, 181, 176, 168, 152, 150, 149, 144, 
    210, 204, 201, 193, 181, 188, 208, 210, 205, 206, 160, 122, 177, 208, 198, 194, 193, 184, 166, 150, 139, 156, 160, 153, 155, 160, 159, 155, 152, 152, 140, 131, 
    210, 202, 198, 187, 174, 178, 205, 214, 209, 203, 164, 131, 180, 202, 187, 182, 182, 169, 157, 139, 134, 153, 154, 144, 151, 141, 131, 141, 157, 155, 150, 147, 
    210, 200, 194, 181, 168, 168, 196, 215, 212, 199, 189, 184, 203, 185, 173, 172, 163, 155, 147, 118, 131, 148, 145, 141, 144, 132, 127, 133, 149, 163, 162, 156, 
    208, 194, 189, 180, 162, 158, 189, 211, 211, 197, 194, 199, 191, 172, 163, 164, 158, 147, 130, 109, 137, 144, 144, 145, 144, 132, 124, 134, 151, 162, 159, 147, 
    194, 177, 176, 181, 159, 143, 179, 205, 208, 199, 194, 190, 181, 165, 156, 161, 149, 136, 112, 114, 137, 133, 138, 146, 146, 131, 131, 144, 150, 149, 148, 141, 
    172, 157, 165, 178, 167, 133, 156, 199, 206, 199, 199, 194, 160, 133, 132, 139, 140, 126, 107, 126, 130, 129, 138, 149, 141, 140, 145, 142, 136, 140, 149, 152, 
    151, 134, 144, 155, 158, 125, 130, 183, 197, 191, 183, 165, 128, 103, 94, 105, 119, 112, 117, 124, 121, 125, 139, 143, 139, 140, 129, 125, 132, 149, 155, 150, 
    
    -- channel=25
    19, 21, 16, 47, 131, 147, 147, 142, 135, 137, 144, 142, 141, 140, 140, 143, 140, 126, 96, 73, 95, 93, 130, 164, 155, 156, 155, 157, 158, 155, 152, 151, 
    20, 20, 17, 31, 122, 161, 155, 146, 138, 136, 139, 149, 152, 150, 146, 151, 159, 150, 117, 73, 65, 88, 156, 175, 168, 169, 171, 173, 172, 168, 164, 163, 
    20, 20, 20, 21, 102, 162, 151, 140, 141, 149, 136, 139, 154, 153, 152, 159, 166, 171, 161, 109, 58, 97, 177, 183, 179, 178, 177, 178, 177, 173, 169, 166, 
    20, 20, 21, 17, 79, 153, 140, 130, 151, 164, 157, 135, 153, 166, 169, 176, 176, 175, 161, 118, 82, 133, 196, 195, 189, 183, 180, 179, 179, 177, 173, 171, 
    21, 20, 21, 19, 56, 137, 130, 119, 156, 178, 179, 146, 132, 139, 148, 167, 175, 169, 152, 120, 109, 167, 206, 210, 209, 201, 195, 191, 186, 182, 177, 172, 
    22, 22, 23, 22, 38, 115, 130, 120, 146, 185, 195, 158, 118, 108, 107, 132, 146, 143, 129, 132, 143, 183, 190, 199, 207, 209, 204, 209, 209, 202, 199, 194, 
    24, 19, 21, 20, 30, 113, 161, 148, 151, 186, 194, 170, 128, 98, 105, 113, 104, 116, 107, 128, 178, 202, 192, 197, 206, 207, 209, 215, 216, 214, 215, 218, 
    88, 41, 24, 29, 96, 174, 186, 156, 149, 181, 189, 186, 164, 132, 129, 118, 92, 107, 108, 124, 180, 204, 187, 206, 230, 224, 231, 228, 205, 211, 220, 226, 
    177, 153, 109, 117, 175, 189, 183, 147, 120, 161, 188, 192, 184, 173, 154, 131, 115, 115, 119, 127, 166, 197, 188, 216, 233, 226, 227, 211, 188, 198, 224, 232, 
    194, 188, 175, 182, 191, 194, 190, 144, 115, 152, 177, 182, 183, 182, 164, 138, 102, 118, 119, 123, 160, 189, 208, 233, 232, 235, 234, 203, 187, 189, 209, 235, 
    199, 192, 183, 187, 198, 205, 191, 138, 136, 165, 176, 181, 184, 175, 154, 124, 107, 118, 119, 120, 158, 176, 205, 240, 243, 244, 242, 212, 192, 192, 198, 224, 
    201, 201, 193, 187, 201, 209, 188, 146, 155, 182, 185, 183, 183, 159, 132, 107, 115, 133, 124, 126, 158, 170, 189, 235, 246, 246, 242, 222, 194, 192, 192, 202, 
    203, 201, 197, 189, 196, 198, 183, 165, 159, 170, 176, 165, 164, 162, 138, 120, 133, 159, 135, 146, 161, 165, 189, 231, 244, 248, 247, 234, 208, 195, 193, 199, 
    208, 202, 196, 185, 193, 167, 156, 185, 161, 145, 135, 135, 161, 158, 137, 143, 164, 164, 149, 162, 153, 157, 195, 228, 242, 247, 249, 245, 232, 199, 204, 222, 
    210, 204, 197, 182, 191, 142, 125, 193, 181, 177, 166, 167, 184, 170, 130, 114, 165, 170, 152, 158, 171, 174, 189, 231, 242, 244, 245, 251, 242, 207, 221, 233, 
    212, 200, 197, 185, 189, 145, 112, 192, 199, 190, 189, 180, 164, 167, 160, 137, 146, 176, 162, 145, 184, 177, 168, 195, 232, 241, 245, 249, 228, 221, 236, 235, 
    216, 199, 182, 174, 176, 155, 110, 173, 208, 186, 168, 178, 168, 155, 167, 164, 110, 150, 177, 134, 154, 171, 144, 104, 145, 209, 238, 237, 210, 221, 243, 237, 
    219, 206, 169, 158, 163, 167, 149, 162, 202, 205, 200, 209, 188, 168, 170, 161, 112, 120, 173, 135, 147, 186, 155, 115, 98, 132, 178, 188, 185, 212, 243, 239, 
    221, 214, 179, 161, 175, 181, 179, 177, 189, 207, 212, 221, 220, 197, 184, 171, 139, 103, 149, 140, 151, 177, 148, 147, 131, 112, 138, 156, 151, 177, 217, 234, 
    223, 218, 198, 178, 194, 194, 190, 200, 186, 184, 191, 199, 203, 208, 200, 177, 171, 135, 127, 158, 168, 155, 131, 143, 137, 126, 148, 159, 147, 144, 158, 197, 
    225, 221, 208, 183, 191, 199, 190, 194, 198, 188, 190, 186, 171, 193, 198, 191, 207, 191, 148, 169, 160, 135, 123, 141, 142, 149, 159, 152, 135, 136, 140, 154, 
    222, 221, 214, 190, 179, 195, 200, 190, 198, 205, 209, 178, 151, 179, 182, 181, 197, 196, 174, 165, 134, 124, 137, 147, 153, 161, 153, 139, 131, 139, 139, 125, 
    219, 218, 219, 198, 170, 191, 210, 207, 203, 206, 207, 180, 156, 174, 180, 176, 182, 181, 176, 150, 111, 125, 150, 152, 152, 161, 154, 138, 138, 128, 115, 106, 
    218, 214, 217, 207, 170, 188, 210, 213, 212, 211, 199, 182, 174, 186, 186, 181, 186, 182, 171, 133, 114, 137, 154, 149, 148, 171, 159, 146, 144, 123, 115, 118, 
    216, 212, 212, 209, 179, 189, 207, 205, 205, 205, 177, 138, 167, 195, 187, 182, 185, 181, 158, 130, 125, 141, 150, 140, 141, 163, 157, 149, 133, 131, 130, 124, 
    215, 210, 208, 200, 187, 190, 206, 204, 198, 196, 131, 80, 145, 194, 184, 174, 174, 165, 147, 131, 120, 139, 143, 136, 137, 142, 140, 136, 133, 133, 121, 112, 
    215, 208, 205, 194, 181, 183, 205, 209, 204, 194, 129, 81, 142, 186, 171, 161, 161, 149, 137, 120, 115, 135, 137, 126, 133, 123, 112, 122, 138, 136, 131, 128, 
    214, 205, 200, 188, 176, 175, 198, 212, 208, 192, 160, 142, 170, 168, 155, 149, 141, 133, 127, 100, 113, 131, 128, 123, 126, 114, 108, 114, 130, 144, 144, 137, 
    210, 196, 192, 183, 169, 166, 192, 210, 209, 192, 182, 180, 171, 153, 141, 140, 134, 125, 111, 92, 120, 126, 126, 127, 126, 114, 105, 116, 133, 144, 141, 129, 
    196, 179, 179, 185, 166, 151, 181, 204, 205, 194, 186, 179, 166, 146, 133, 136, 126, 114, 93, 97, 120, 115, 120, 128, 128, 113, 113, 126, 132, 131, 130, 123, 
    177, 161, 170, 184, 174, 140, 156, 195, 201, 193, 191, 182, 145, 113, 108, 115, 118, 106, 89, 110, 114, 112, 120, 131, 123, 122, 127, 124, 117, 122, 130, 134, 
    157, 140, 151, 161, 166, 130, 128, 177, 191, 183, 175, 154, 112, 83, 71, 83, 99, 94, 101, 110, 108, 108, 121, 126, 121, 122, 111, 107, 115, 132, 137, 132, 
    
    -- channel=26
    23, 28, 19, 40, 113, 115, 109, 116, 113, 103, 106, 105, 105, 105, 105, 107, 106, 99, 76, 58, 84, 86, 114, 137, 124, 125, 124, 125, 127, 125, 122, 120, 
    24, 27, 20, 26, 106, 130, 118, 124, 125, 114, 109, 117, 120, 118, 114, 121, 133, 131, 106, 68, 62, 81, 140, 150, 138, 140, 137, 136, 136, 133, 129, 128, 
    24, 26, 23, 18, 88, 131, 116, 123, 139, 141, 116, 116, 129, 127, 125, 132, 142, 154, 152, 105, 55, 89, 159, 158, 151, 151, 146, 142, 142, 139, 136, 132, 
    24, 25, 25, 18, 69, 124, 106, 115, 156, 166, 146, 120, 137, 148, 149, 151, 150, 156, 148, 109, 74, 122, 177, 169, 161, 157, 152, 149, 150, 148, 145, 142, 
    25, 24, 25, 23, 51, 109, 96, 104, 161, 184, 178, 141, 124, 128, 134, 147, 151, 150, 137, 108, 96, 152, 183, 181, 179, 174, 168, 164, 160, 156, 152, 147, 
    26, 26, 27, 28, 35, 89, 95, 102, 150, 193, 199, 159, 116, 102, 98, 118, 130, 131, 119, 122, 132, 167, 166, 170, 178, 183, 179, 183, 183, 177, 175, 169, 
    26, 22, 25, 26, 29, 92, 128, 123, 147, 195, 199, 171, 126, 94, 99, 106, 96, 109, 101, 122, 172, 192, 170, 176, 195, 196, 197, 202, 197, 191, 191, 194, 
    77, 33, 17, 25, 88, 154, 155, 126, 140, 190, 193, 185, 163, 129, 123, 113, 88, 103, 104, 121, 177, 198, 165, 189, 228, 219, 224, 218, 186, 187, 196, 205, 
    149, 128, 86, 96, 155, 167, 153, 119, 111, 168, 191, 191, 183, 170, 148, 127, 112, 112, 116, 124, 163, 187, 162, 193, 223, 213, 207, 187, 157, 166, 196, 210, 
    161, 158, 146, 155, 167, 169, 159, 117, 104, 155, 179, 181, 182, 180, 159, 135, 100, 116, 117, 121, 158, 178, 178, 204, 216, 214, 203, 167, 147, 150, 176, 207, 
    170, 165, 158, 165, 175, 176, 160, 112, 123, 164, 177, 180, 182, 172, 149, 121, 106, 116, 117, 118, 156, 166, 175, 209, 222, 216, 205, 169, 145, 147, 159, 186, 
    172, 174, 169, 166, 176, 176, 157, 122, 141, 177, 185, 182, 182, 157, 127, 104, 115, 132, 123, 125, 159, 164, 163, 206, 224, 217, 205, 181, 146, 142, 147, 156, 
    167, 167, 165, 160, 165, 164, 153, 143, 145, 163, 174, 164, 163, 159, 133, 118, 134, 159, 135, 146, 163, 163, 168, 205, 223, 220, 214, 199, 163, 144, 144, 152, 
    169, 162, 160, 155, 163, 136, 131, 164, 146, 136, 132, 133, 159, 158, 135, 146, 167, 162, 144, 158, 152, 152, 176, 203, 215, 216, 221, 218, 197, 159, 162, 182, 
    174, 164, 162, 157, 168, 120, 109, 178, 166, 167, 161, 163, 182, 171, 132, 120, 169, 163, 140, 149, 166, 164, 170, 204, 211, 213, 218, 228, 214, 176, 187, 199, 
    175, 160, 161, 159, 170, 132, 104, 183, 188, 182, 184, 176, 162, 168, 163, 141, 145, 165, 146, 133, 175, 165, 150, 169, 202, 212, 217, 221, 196, 186, 199, 199, 
    179, 159, 146, 148, 161, 151, 109, 168, 199, 181, 164, 174, 165, 156, 170, 166, 105, 136, 159, 119, 143, 158, 126, 80, 118, 183, 209, 205, 175, 183, 201, 197, 
    181, 164, 133, 131, 149, 165, 151, 159, 194, 199, 196, 205, 185, 168, 172, 162, 104, 105, 155, 119, 134, 173, 136, 92, 75, 111, 152, 158, 152, 176, 203, 200, 
    183, 172, 142, 133, 159, 176, 177, 170, 177, 197, 207, 217, 217, 198, 187, 170, 131, 90, 133, 126, 139, 162, 130, 126, 111, 96, 118, 132, 124, 146, 184, 199, 
    185, 176, 161, 149, 175, 183, 182, 188, 170, 170, 185, 194, 201, 208, 202, 175, 164, 123, 113, 145, 157, 140, 113, 123, 119, 112, 134, 142, 127, 121, 132, 166, 
    189, 183, 173, 155, 171, 186, 177, 178, 180, 172, 178, 177, 164, 188, 195, 189, 201, 182, 136, 157, 147, 120, 106, 124, 128, 138, 148, 138, 120, 119, 122, 130, 
    189, 188, 183, 161, 158, 183, 187, 176, 184, 191, 192, 164, 139, 166, 173, 177, 192, 188, 162, 150, 118, 107, 121, 133, 142, 150, 141, 125, 117, 124, 125, 108, 
    186, 186, 187, 166, 148, 180, 199, 197, 193, 195, 192, 168, 145, 159, 169, 170, 175, 172, 163, 134, 93, 108, 134, 139, 141, 151, 142, 124, 124, 114, 101, 91, 
    186, 181, 183, 172, 143, 176, 201, 207, 206, 203, 189, 175, 165, 171, 174, 172, 178, 171, 158, 117, 97, 120, 138, 136, 138, 161, 146, 132, 130, 109, 100, 104, 
    184, 178, 175, 169, 146, 170, 198, 202, 200, 197, 171, 136, 161, 180, 171, 170, 173, 168, 144, 115, 108, 124, 134, 126, 130, 153, 145, 135, 119, 117, 116, 111, 
    184, 176, 168, 157, 147, 162, 192, 200, 191, 185, 129, 82, 141, 179, 166, 159, 159, 150, 132, 116, 105, 122, 127, 122, 127, 132, 128, 122, 119, 119, 107, 98, 
    184, 172, 163, 148, 134, 146, 186, 202, 192, 178, 130, 88, 140, 172, 152, 144, 145, 132, 122, 105, 100, 119, 121, 112, 122, 113, 100, 108, 124, 122, 117, 114, 
    183, 169, 158, 142, 126, 132, 178, 204, 195, 175, 157, 144, 164, 152, 135, 131, 124, 116, 111, 84, 97, 115, 113, 109, 114, 102, 95, 100, 116, 130, 130, 123, 
    177, 161, 153, 142, 119, 122, 178, 204, 197, 180, 170, 168, 157, 135, 122, 123, 119, 109, 94, 75, 104, 111, 112, 113, 112, 100, 92, 102, 119, 130, 126, 115, 
    163, 144, 141, 145, 116, 107, 169, 200, 194, 183, 172, 163, 150, 129, 115, 121, 112, 100, 78, 81, 104, 101, 106, 114, 114, 99, 99, 112, 118, 117, 116, 110, 
    142, 126, 131, 143, 124, 95, 145, 192, 190, 183, 178, 168, 130, 98, 92, 101, 104, 92, 75, 95, 99, 97, 106, 116, 109, 108, 113, 110, 103, 108, 116, 119, 
    123, 104, 112, 120, 116, 87, 118, 174, 181, 174, 164, 141, 99, 69, 57, 70, 87, 81, 88, 96, 93, 94, 107, 112, 107, 108, 97, 93, 101, 118, 123, 118, 
    
    -- channel=27
    217, 210, 205, 199, 218, 214, 207, 189, 187, 174, 166, 169, 150, 154, 140, 143, 167, 191, 219, 223, 219, 215, 226, 225, 219, 190, 175, 187, 200, 170, 161, 162, 
    222, 221, 220, 215, 216, 225, 211, 179, 180, 192, 190, 188, 199, 206, 209, 219, 229, 235, 236, 236, 233, 226, 225, 229, 231, 212, 208, 205, 216, 183, 186, 200, 
    234, 233, 231, 232, 233, 239, 217, 173, 164, 180, 173, 183, 190, 188, 212, 224, 218, 235, 227, 225, 229, 223, 214, 225, 234, 232, 230, 216, 209, 202, 208, 211, 
    245, 244, 244, 242, 244, 243, 228, 158, 146, 157, 131, 159, 145, 136, 162, 159, 169, 203, 195, 211, 209, 203, 208, 226, 230, 233, 228, 213, 199, 219, 224, 212, 
    245, 243, 244, 244, 245, 241, 207, 117, 99, 108, 89, 107, 100, 91, 100, 92, 102, 124, 124, 149, 182, 185, 202, 233, 225, 226, 227, 205, 194, 213, 226, 222, 
    245, 244, 244, 243, 245, 237, 216, 126, 72, 90, 91, 102, 101, 103, 107, 99, 89, 89, 91, 93, 126, 190, 216, 235, 231, 223, 216, 196, 174, 189, 217, 236, 
    245, 243, 243, 244, 241, 219, 217, 158, 80, 114, 132, 151, 140, 132, 143, 138, 130, 122, 114, 120, 110, 155, 221, 233, 235, 224, 198, 192, 167, 171, 204, 235, 
    244, 243, 243, 246, 227, 199, 215, 153, 81, 146, 187, 202, 207, 158, 131, 131, 129, 141, 131, 132, 159, 132, 159, 215, 229, 215, 212, 209, 197, 171, 178, 221, 
    244, 243, 244, 245, 227, 206, 218, 130, 81, 130, 128, 129, 184, 145, 116, 125, 124, 137, 142, 125, 153, 147, 144, 198, 214, 219, 233, 220, 184, 164, 169, 201, 
    243, 243, 244, 242, 228, 190, 168, 110, 83, 134, 119, 110, 143, 128, 115, 120, 125, 131, 146, 125, 149, 155, 140, 196, 233, 240, 240, 233, 200, 200, 215, 220, 
    239, 241, 244, 245, 220, 133, 130, 95, 78, 116, 116, 108, 109, 107, 109, 108, 115, 120, 120, 115, 136, 150, 143, 167, 208, 228, 245, 243, 244, 245, 245, 244, 
    222, 233, 242, 244, 216, 169, 165, 89, 61, 67, 91, 100, 95, 95, 98, 96, 96, 95, 90, 97, 105, 121, 129, 126, 155, 216, 248, 243, 244, 244, 244, 244, 
    208, 223, 236, 227, 191, 183, 181, 100, 55, 56, 88, 101, 111, 99, 86, 84, 82, 84, 93, 113, 109, 98, 112, 129, 174, 226, 245, 244, 244, 244, 244, 244, 
    200, 204, 219, 195, 170, 154, 156, 102, 104, 99, 108, 102, 115, 117, 94, 85, 90, 106, 122, 140, 128, 104, 108, 124, 150, 179, 195, 212, 239, 245, 244, 244, 
    200, 210, 207, 169, 164, 148, 147, 138, 129, 92, 106, 93, 89, 93, 84, 77, 76, 81, 81, 81, 79, 74, 75, 82, 101, 123, 140, 143, 191, 244, 244, 244, 
    210, 226, 196, 119, 112, 150, 186, 192, 108, 77, 77, 55, 45, 47, 60, 63, 59, 63, 59, 54, 49, 50, 61, 64, 71, 75, 91, 103, 135, 225, 246, 244, 
    199, 193, 180, 96, 93, 145, 192, 161, 86, 73, 92, 98, 104, 79, 79, 71, 37, 28, 30, 27, 52, 50, 22, 28, 24, 53, 91, 104, 128, 206, 247, 243, 
    211, 199, 194, 113, 120, 157, 159, 71, 68, 90, 116, 124, 149, 121, 128, 102, 78, 98, 112, 100, 148, 147, 92, 99, 94, 108, 135, 142, 156, 183, 242, 245, 
    220, 202, 183, 102, 110, 165, 132, 30, 57, 98, 107, 83, 82, 101, 129, 100, 153, 174, 158, 159, 172, 168, 162, 163, 160, 175, 156, 119, 114, 135, 228, 247, 
    219, 207, 188, 98, 83, 141, 111, 42, 58, 72, 76, 62, 53, 56, 64, 93, 160, 124, 91, 101, 116, 107, 103, 103, 99, 155, 126, 67, 81, 118, 217, 248, 
    217, 210, 199, 101, 56, 88, 93, 60, 56, 46, 63, 70, 60, 54, 64, 65, 99, 114, 105, 103, 100, 96, 93, 97, 102, 111, 100, 73, 82, 114, 212, 249, 
    209, 205, 202, 117, 83, 70, 81, 68, 50, 35, 43, 51, 68, 77, 87, 63, 52, 71, 82, 72, 64, 67, 62, 93, 88, 60, 83, 108, 112, 108, 204, 250, 
    205, 202, 197, 104, 93, 111, 71, 73, 63, 41, 38, 34, 75, 99, 142, 79, 30, 86, 147, 118, 99, 114, 102, 153, 178, 63, 74, 141, 119, 90, 195, 246, 
    198, 194, 185, 87, 49, 108, 97, 99, 95, 51, 39, 36, 40, 50, 87, 55, 32, 79, 151, 127, 122, 136, 116, 156, 159, 55, 53, 74, 62, 78, 194, 240, 
    182, 180, 169, 77, 37, 59, 108, 144, 106, 60, 43, 32, 29, 28, 30, 33, 39, 42, 58, 88, 106, 121, 122, 117, 67, 47, 51, 50, 51, 80, 186, 225, 
    168, 165, 164, 125, 91, 96, 111, 141, 96, 74, 55, 36, 30, 30, 29, 31, 35, 24, 64, 174, 205, 203, 179, 181, 87, 38, 43, 48, 66, 91, 174, 211, 
    162, 163, 175, 180, 152, 118, 108, 141, 91, 83, 78, 48, 25, 24, 25, 29, 39, 38, 71, 164, 184, 177, 169, 166, 81, 30, 30, 49, 78, 95, 169, 206, 
    154, 172, 179, 166, 146, 117, 103, 146, 87, 85, 82, 54, 32, 30, 33, 37, 54, 77, 86, 101, 107, 121, 142, 137, 60, 30, 33, 54, 78, 91, 165, 199, 
    166, 169, 158, 148, 143, 133, 103, 113, 79, 81, 75, 60, 42, 39, 42, 44, 48, 54, 65, 77, 90, 110, 131, 139, 53, 29, 38, 54, 70, 91, 169, 196, 
    162, 151, 147, 141, 137, 133, 107, 78, 72, 78, 70, 60, 50, 42, 46, 48, 49, 51, 59, 66, 76, 89, 101, 113, 69, 29, 35, 52, 63, 98, 174, 186, 
    148, 141, 142, 140, 143, 140, 106, 60, 66, 74, 66, 55, 57, 52, 54, 58, 58, 58, 65, 70, 73, 80, 87, 93, 77, 37, 38, 55, 74, 131, 179, 180, 
    144, 149, 160, 162, 158, 146, 126, 61, 57, 57, 58, 67, 70, 69, 73, 72, 68, 73, 89, 98, 94, 97, 99, 97, 82, 69, 64, 71, 119, 164, 182, 186, 
    
    -- channel=28
    215, 208, 208, 202, 215, 209, 202, 185, 184, 168, 152, 160, 157, 167, 154, 157, 181, 203, 225, 225, 222, 219, 229, 228, 221, 197, 184, 196, 208, 184, 176, 165, 
    226, 224, 225, 217, 213, 221, 204, 171, 180, 189, 178, 177, 196, 205, 208, 224, 236, 240, 242, 243, 238, 229, 228, 231, 231, 214, 212, 210, 222, 190, 191, 197, 
    235, 234, 234, 235, 234, 239, 214, 166, 166, 177, 168, 177, 184, 183, 206, 223, 220, 236, 227, 232, 235, 228, 217, 224, 233, 233, 230, 221, 217, 206, 209, 210, 
    245, 244, 244, 243, 244, 244, 227, 153, 146, 155, 130, 159, 144, 138, 162, 160, 172, 205, 194, 220, 222, 211, 211, 224, 230, 233, 229, 219, 207, 223, 226, 212, 
    245, 244, 244, 244, 245, 240, 205, 112, 98, 109, 91, 109, 101, 92, 100, 92, 104, 125, 124, 154, 194, 194, 201, 227, 220, 222, 227, 211, 203, 220, 232, 225, 
    245, 244, 244, 243, 246, 235, 212, 123, 71, 93, 95, 105, 103, 106, 110, 102, 91, 89, 91, 93, 129, 197, 217, 230, 221, 218, 214, 198, 180, 197, 226, 237, 
    245, 243, 243, 244, 240, 214, 213, 156, 79, 119, 137, 154, 144, 139, 155, 150, 142, 128, 121, 126, 114, 160, 225, 233, 233, 218, 192, 186, 165, 176, 212, 236, 
    244, 243, 243, 247, 226, 193, 211, 150, 81, 152, 188, 200, 205, 165, 141, 144, 142, 150, 141, 143, 167, 140, 163, 214, 224, 209, 211, 210, 199, 174, 175, 220, 
    244, 243, 244, 245, 225, 202, 216, 127, 81, 134, 132, 135, 185, 151, 124, 135, 134, 145, 150, 136, 164, 158, 142, 192, 207, 216, 231, 215, 177, 158, 156, 196, 
    242, 242, 244, 242, 227, 189, 168, 110, 83, 140, 128, 118, 147, 135, 124, 129, 133, 139, 151, 134, 158, 164, 145, 193, 229, 239, 239, 230, 193, 190, 204, 215, 
    232, 239, 243, 244, 218, 129, 128, 94, 79, 122, 122, 112, 113, 112, 115, 115, 124, 128, 127, 126, 144, 158, 153, 170, 206, 227, 246, 244, 243, 243, 245, 244, 
    205, 227, 242, 242, 211, 161, 159, 88, 60, 69, 94, 102, 98, 97, 103, 102, 104, 100, 95, 103, 113, 127, 137, 128, 153, 215, 248, 243, 244, 244, 244, 244, 
    188, 213, 228, 220, 180, 170, 173, 99, 55, 57, 90, 102, 114, 103, 88, 85, 85, 85, 93, 115, 112, 101, 118, 134, 176, 225, 245, 244, 244, 244, 244, 244, 
    184, 188, 202, 181, 152, 134, 141, 99, 103, 102, 111, 103, 118, 120, 96, 86, 92, 107, 125, 146, 132, 106, 110, 127, 152, 179, 195, 210, 238, 245, 244, 244, 
    182, 194, 189, 152, 146, 123, 127, 126, 124, 93, 105, 94, 90, 93, 85, 79, 78, 83, 84, 85, 81, 75, 76, 83, 101, 122, 138, 138, 188, 244, 244, 244, 
    189, 204, 167, 101, 101, 125, 169, 174, 103, 77, 79, 54, 43, 47, 59, 62, 59, 62, 57, 52, 47, 48, 61, 64, 70, 74, 90, 97, 128, 223, 246, 244, 
    174, 164, 151, 84, 82, 124, 172, 146, 83, 73, 87, 90, 100, 75, 76, 68, 33, 23, 26, 23, 48, 47, 20, 25, 21, 50, 86, 100, 120, 202, 247, 243, 
    192, 180, 179, 104, 104, 135, 142, 64, 65, 87, 108, 120, 149, 118, 125, 98, 70, 89, 106, 96, 144, 144, 89, 96, 90, 103, 130, 139, 151, 178, 241, 244, 
    209, 189, 171, 94, 98, 146, 118, 28, 54, 95, 103, 79, 83, 100, 128, 95, 146, 170, 155, 158, 171, 168, 160, 161, 158, 172, 155, 119, 111, 128, 226, 247, 
    208, 193, 176, 91, 76, 127, 100, 40, 53, 68, 73, 57, 50, 53, 61, 89, 156, 119, 87, 98, 113, 104, 99, 100, 96, 152, 122, 63, 77, 112, 214, 248, 
    202, 195, 190, 95, 51, 78, 83, 56, 51, 39, 60, 68, 57, 51, 59, 61, 95, 110, 102, 101, 99, 95, 92, 96, 100, 108, 96, 70, 79, 108, 208, 249, 
    194, 192, 192, 110, 76, 62, 73, 63, 46, 29, 40, 48, 65, 72, 83, 59, 48, 67, 77, 67, 60, 64, 59, 88, 82, 54, 78, 105, 107, 101, 201, 249, 
    195, 190, 187, 97, 85, 99, 65, 67, 58, 38, 35, 32, 72, 96, 141, 76, 25, 79, 140, 113, 94, 109, 97, 146, 171, 58, 69, 138, 116, 83, 192, 244, 
    189, 183, 176, 82, 44, 99, 89, 94, 90, 48, 36, 33, 38, 47, 85, 52, 28, 74, 145, 123, 119, 134, 113, 151, 156, 51, 50, 71, 59, 71, 192, 238, 
    174, 173, 163, 72, 34, 54, 101, 139, 102, 58, 40, 30, 26, 25, 26, 30, 37, 38, 53, 86, 104, 117, 118, 114, 62, 43, 48, 46, 47, 75, 184, 223, 
    162, 160, 158, 120, 87, 89, 103, 136, 92, 72, 52, 34, 28, 27, 27, 29, 32, 21, 61, 175, 207, 202, 177, 180, 84, 34, 40, 44, 62, 87, 171, 209, 
    156, 156, 168, 176, 147, 112, 102, 136, 86, 81, 75, 45, 22, 22, 23, 26, 35, 34, 69, 164, 185, 177, 169, 165, 78, 25, 26, 45, 75, 92, 167, 204, 
    149, 167, 173, 161, 141, 113, 99, 142, 83, 83, 79, 51, 29, 28, 31, 34, 50, 72, 81, 97, 102, 116, 138, 133, 55, 27, 29, 50, 76, 89, 164, 198, 
    164, 166, 155, 144, 139, 130, 99, 108, 76, 80, 72, 56, 38, 36, 39, 41, 45, 51, 61, 72, 84, 103, 124, 131, 49, 26, 33, 50, 69, 89, 169, 195, 
    160, 148, 146, 141, 135, 130, 102, 73, 69, 77, 66, 56, 47, 40, 43, 45, 46, 48, 54, 61, 70, 84, 94, 106, 64, 26, 31, 48, 61, 98, 175, 186, 
    147, 141, 142, 140, 143, 139, 104, 57, 64, 74, 63, 52, 55, 49, 51, 54, 54, 54, 61, 66, 68, 74, 81, 87, 72, 33, 35, 52, 72, 132, 182, 181, 
    146, 150, 161, 163, 157, 145, 124, 58, 55, 56, 57, 65, 67, 66, 70, 69, 67, 72, 87, 95, 92, 95, 96, 94, 81, 68, 62, 70, 118, 163, 182, 185, 
    
    -- channel=29
    209, 202, 191, 182, 209, 209, 198, 175, 171, 165, 157, 160, 149, 154, 141, 143, 164, 188, 214, 219, 209, 202, 217, 214, 208, 177, 161, 173, 183, 157, 149, 149, 
    212, 212, 210, 205, 207, 219, 200, 163, 165, 182, 184, 182, 194, 201, 205, 215, 223, 227, 227, 228, 221, 212, 211, 215, 223, 205, 195, 187, 198, 170, 173, 186, 
    230, 229, 227, 226, 227, 236, 211, 164, 159, 173, 183, 184, 188, 191, 207, 224, 219, 229, 224, 214, 214, 208, 200, 211, 222, 224, 219, 197, 185, 188, 197, 198, 
    245, 244, 244, 241, 242, 241, 227, 175, 168, 176, 161, 187, 174, 160, 184, 182, 185, 213, 208, 202, 185, 186, 196, 212, 215, 220, 213, 187, 169, 197, 212, 200, 
    245, 243, 244, 244, 245, 241, 205, 132, 139, 161, 138, 167, 159, 139, 155, 141, 142, 166, 153, 164, 169, 169, 196, 224, 209, 209, 212, 177, 160, 184, 204, 210, 
    245, 244, 244, 243, 246, 238, 215, 129, 113, 156, 160, 170, 170, 170, 177, 167, 157, 157, 152, 143, 148, 179, 205, 228, 218, 206, 193, 170, 147, 160, 192, 223, 
    245, 243, 243, 244, 241, 221, 221, 180, 131, 180, 196, 207, 200, 203, 217, 211, 204, 195, 192, 191, 163, 166, 205, 225, 227, 213, 177, 169, 145, 146, 178, 218, 
    244, 242, 242, 247, 230, 202, 217, 192, 134, 194, 224, 232, 234, 215, 206, 209, 207, 208, 202, 207, 224, 180, 154, 204, 220, 201, 196, 188, 171, 146, 154, 199, 
    245, 243, 243, 245, 227, 209, 223, 174, 135, 186, 193, 193, 221, 204, 193, 201, 202, 205, 205, 198, 220, 208, 163, 188, 203, 209, 223, 203, 161, 139, 148, 178, 
    242, 241, 243, 242, 229, 205, 194, 164, 140, 193, 189, 184, 202, 196, 192, 196, 199, 202, 208, 198, 215, 224, 188, 200, 230, 238, 237, 227, 188, 186, 202, 211, 
    234, 238, 243, 244, 223, 160, 169, 156, 134, 177, 179, 172, 174, 174, 180, 183, 187, 190, 188, 190, 205, 220, 208, 196, 217, 230, 246, 244, 244, 244, 244, 244, 
    211, 230, 242, 242, 216, 182, 190, 151, 106, 110, 147, 160, 158, 159, 166, 170, 169, 163, 158, 166, 173, 189, 198, 175, 183, 224, 248, 243, 244, 244, 244, 244, 
    196, 218, 233, 225, 189, 180, 195, 159, 93, 92, 141, 160, 186, 168, 143, 140, 139, 137, 146, 167, 152, 131, 143, 150, 188, 227, 243, 244, 244, 244, 244, 244, 
    195, 199, 211, 193, 164, 149, 162, 137, 150, 170, 178, 166, 189, 205, 166, 146, 153, 172, 192, 211, 175, 128, 128, 138, 160, 177, 191, 211, 239, 245, 243, 243, 
    194, 207, 200, 162, 156, 136, 142, 137, 162, 178, 177, 159, 150, 163, 149, 139, 141, 146, 146, 147, 134, 124, 127, 133, 149, 163, 173, 166, 204, 245, 243, 244, 
    195, 208, 173, 110, 113, 139, 180, 185, 133, 154, 127, 87, 73, 76, 89, 95, 92, 96, 94, 88, 86, 86, 99, 103, 109, 116, 143, 155, 175, 232, 245, 245, 
    183, 170, 161, 101, 96, 136, 181, 161, 128, 132, 129, 135, 140, 125, 125, 106, 53, 43, 44, 39, 77, 71, 35, 40, 32, 80, 145, 151, 167, 219, 246, 243, 
    202, 193, 194, 124, 120, 146, 153, 73, 105, 135, 131, 148, 184, 159, 169, 131, 102, 118, 132, 122, 175, 170, 111, 115, 111, 145, 178, 181, 187, 197, 242, 244, 
    216, 200, 184, 114, 115, 157, 130, 36, 79, 149, 129, 99, 111, 129, 157, 132, 177, 193, 183, 185, 200, 193, 186, 189, 181, 199, 182, 151, 148, 162, 232, 246, 
    217, 204, 187, 113, 96, 139, 113, 61, 78, 112, 115, 93, 85, 83, 94, 125, 191, 159, 127, 138, 160, 149, 140, 143, 138, 189, 159, 99, 115, 154, 226, 247, 
    213, 208, 199, 117, 73, 92, 99, 84, 75, 65, 97, 105, 95, 87, 103, 95, 134, 162, 153, 151, 150, 144, 137, 143, 147, 153, 143, 111, 115, 146, 222, 247, 
    204, 206, 204, 131, 101, 81, 92, 90, 70, 45, 57, 69, 98, 111, 125, 87, 74, 102, 112, 103, 98, 101, 94, 125, 115, 82, 113, 149, 154, 137, 212, 248, 
    209, 208, 206, 117, 105, 122, 86, 94, 86, 54, 51, 47, 102, 131, 173, 99, 45, 100, 158, 130, 121, 138, 124, 171, 187, 75, 95, 171, 152, 117, 207, 250, 
    221, 214, 204, 104, 59, 116, 114, 128, 124, 65, 52, 48, 56, 70, 108, 75, 48, 95, 166, 143, 145, 167, 143, 175, 175, 74, 72, 98, 84, 104, 214, 251, 
    215, 212, 201, 99, 47, 68, 128, 176, 135, 80, 56, 45, 40, 39, 43, 47, 55, 60, 80, 110, 125, 147, 144, 139, 92, 67, 70, 67, 69, 109, 217, 251, 
    207, 207, 203, 157, 115, 117, 133, 170, 126, 101, 72, 48, 40, 41, 41, 45, 50, 39, 83, 192, 218, 220, 199, 201, 107, 52, 56, 63, 90, 126, 210, 247, 
    188, 192, 206, 216, 191, 154, 134, 161, 121, 115, 104, 62, 33, 34, 35, 41, 51, 49, 85, 179, 199, 192, 190, 187, 96, 39, 38, 66, 111, 133, 209, 245, 
    191, 198, 205, 198, 181, 158, 132, 160, 114, 118, 111, 70, 39, 38, 44, 49, 68, 93, 105, 126, 135, 150, 173, 166, 72, 40, 42, 71, 113, 130, 207, 242, 
    206, 209, 198, 184, 171, 163, 130, 133, 107, 111, 104, 77, 50, 47, 53, 57, 63, 72, 87, 104, 120, 145, 168, 176, 69, 40, 48, 71, 102, 126, 212, 238, 
    199, 194, 194, 189, 178, 166, 134, 101, 99, 105, 96, 79, 62, 54, 59, 62, 65, 69, 78, 87, 100, 116, 129, 143, 87, 39, 44, 71, 89, 133, 223, 232, 
    193, 188, 190, 188, 189, 188, 144, 80, 90, 99, 88, 70, 73, 69, 74, 78, 78, 78, 86, 93, 97, 102, 109, 114, 94, 48, 48, 74, 100, 173, 232, 231, 
    196, 199, 208, 205, 200, 187, 165, 85, 76, 76, 78, 84, 84, 89, 98, 99, 94, 99, 114, 124, 125, 129, 128, 127, 112, 91, 84, 96, 148, 204, 225, 223, 
    
    
    others => 0);
end ifmap_package;
