-gN_BRAM_IWGHT=15 -gN_BRAM_IFMAP=3