library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -- layer=3
    -6197, -1875, 218, 1837, 8123, -5510, 6866, -6140, 4071, -1814,

    -- weights
    -- layer=3 filter=0 channel=0
    -10, 3, 15, 4, -18, -23, -30, 2, -18, -6, -68, 4, 21, -27, -23, 30, 42, 12, 41, 29, -37, -20, -8, -26, 0, -30, 0, -27, -23, 4, -19, -17, 14, 18, -8, -2, -13, 20, 5, 39, -5, 12, -8, -41, -18, 0, 16, -10, -17, -26, 9, -32, -17, -15, 9, -5, 2, -4, 23, -2, 22, 12, -1, 17, 13, -6, -7, 9, -17, -8, -7, 5, 39, 12, -9, 35, -7, -9, -24, -21, 24, -2, -24, 7, -9, 40, 11, 11, 10, -11, 23, -12, -23, 19, -7, 20, -21, -6, 63, -5, 20, 9, -24, 42, 38, 27, -17, 12, 15, 13, 38, 22, -19, -29, 23, -29, 9, -6, -21, 14, -4, 0, 5, 1, 18, -22, 0, 5, -16, 42, 8, 10, 1, -27, -14, -21, 25, -10, -26, -3, -31, 15, -36, -12, -22, -6, -53, 20, -13, -2, 0, 5, 19, -22, 6, -13, -31, -30, 1, -2, -19, 4, -31, 30, -35, 17, -4, -3, 5, 23, -49, -1, 3, 4, -3, 20, 10, -10, 12, -53, -32, 20, 7, 1, -11, -18, 12, -37, -10, 13, 32, 5, -27, 29, 1, -30, 0, 37, -28, -19, -31, -16, -48, -24, 15, -9, 32, 9, -27, -1, 57, 15, -46, -10, 9, -32, -8, -4, 9, -35, 30, -17, 42, 0, 10, -10, 25, -28, 2, 14, -6, -15, 17, 9, 29, -3, 1, 16, -10, 30, 29, -8, 17, 4, 1, -35, -16, -16, 15, -7, -4, -14, -67, 15, 3, -30, 3, 18, 2, -27, -2, 0, 17, -4, -36, -15, -9, -9, 3, 8, -2, 12, 2, 33, 1, -15, 17, 12, -21, -16, -22, -33, -14, -14, 25, 11, -6, -4, 2, 15, 39, 10, -31, 21, 1, -27, 0, -10, 28, -6, -39, 19, -23, 7, -37, -19, 28, 18, -8, -13, -11, -4, -13, -5, 22, -40, -36, 2, 24, 15, -4, -11, 24, -14, 52, 11, 20, 4, -4, 4, -21, 8, -11, -36, 0, 2, -44, 0, 49, 16, -6, -10, 21, -35, 20, 6, 12, -41, -33, -43, -3, 6, 22, -9, -18, 2, -22, -13, 10, -12, -3, -11, -2, 30, -12, 21, -27, 31, 25, 18, -5, -22, -23, -46, -9, 7, 1, -6, 19, -30, -13, -8, 25, -28, 4, 24, 11, -14, -34, 24, 12, 19, 31, 41, -45, 18, -12, 22, 37, -3, 18, 13, -22, -3, 22, 9, 39, -22, 34, 10, 10, 26, -18, -56, -16, 20, 8, 14, -61, 11, 36, 3, -29, 16, 26, 13, -29, -25, 34, -16, 10, 28, -50, -23, -22, -34, 1, 0, -11, -16, -8, 8, -4, 53, 10, 8, 19, 0, -4, 9, -7, -40, 4, 31, 26, 16, -10, 21, 4, 3, 20, -19, 31, 0, 24, 30, -40, -10, -7, 34, -17, -14, 0, 7, -21, 19, 28, 20, -12, -8, 25, -10, -35, 20, 3, -19, 12, 4, -16, -19, -16, -4, -17, -10, -17, 1, -13, -12, -18, -13, 17, 32, -20, 4, -3, 36, 14, 30, -23, 17, -11, 33, 4, -52, 1, -39, 11, 12, -4, -21, -10, -10, -76, 9, -14, 13, -8, 37, -16, -8, 34, -6, 12, 38, -6, -45, -26, 0, 17, 24, -19, 15, -39, 4, -2, -25, 22, 19, 2, -5, -24, 22, 33, 44, 7, -19, -56, -2, 1, 42, 3, 12, -7, -45, -11, -9, 4, 50, -31, 24, -19, -10, -1, -28, -22, -2,
    -- layer=3 filter=0 channel=1
    -23, -4, -30, 18, -9, 26, -10, 9, 14, -9, -8, 3, 2, 13, 20, 0, -1, -22, 2, -4, 3, -27, -8, -18, 3, -12, -4, 15, -5, 0, 18, -8, 12, 0, -16, -3, 28, 5, -34, -12, 12, -20, -17, 18, 33, -11, 0, 9, 31, -10, -32, -15, -6, -3, 21, 4, 7, -21, -17, -1, -9, 11, 9, -11, -62, -10, -47, -41, 11, 41, -6, 15, -13, -27, 5, -1, 0, -13, 15, 28, 0, -34, -19, -1, 48, -21, 8, 4, -13, 36, 10, 20, -18, -3, -4, -7, -5, -2, 31, -30, -11, 24, -16, -8, -12, 32, -3, -5, -13, -21, 18, 23, 7, -24, 11, -6, -8, -14, -15, -34, 6, 16, 24, 2, -30, -2, -20, 26, -3, -19, 5, 21, 19, 33, -4, -20, -15, -26, -2, -32, -24, -30, 8, 27, -8, 12, 9, 2, 5, 6, 3, 4, 0, 38, 0, -7, -16, 32, -14, -6, -22, 16, 25, -14, -18, -40, -9, -2, -37, 15, 0, 39, 11, 12, -2, -2, 15, -22, 26, 32, -5, -31, 17, 8, -10, -29, -5, 1, -15, 22, -52, -14, -2, -45, -10, -12, 8, -1, -3, -9, -5, -11, 31, -5, 34, -11, 21, -20, 9, -13, -27, 40, -30, -25, 1, -46, -35, -29, 20, 32, 15, -27, 16, 19, 3, 14, -29, 22, 7, 32, 14, -28, 37, -12, -3, -52, -26, 13, -18, 11, -21, -7, 27, 42, 41, -13, -6, -59, -16, 21, 35, 19, 7, -18, -43, 46, -21, 54, 35, -33, 34, 13, 37, 4, -16, 23, 10, 19, 9, 16, -24, 23, -17, -9, -24, -8, -40, -35, -22, -23, 18, -47, 13, 9, 29, -33, -24, -21, 19, -10, -22, 14, 15, 2, 12, -19, 8, 28, -24, -57, -3, 20, -43, 19, 12, 7, 14, 6, 29, -70, -2, 10, 5, 29, 48, -57, -32, 23, -42, 10, -16, 25, 7, -42, 0, 4, 29, 0, -12, 10, -11, -12, -30, 18, -16, 8, -12, 18, -39, 16, -35, -42, 26, -26, 14, 0, 6, 23, -16, -4, -15, -4, 23, 21, -37, -15, -25, 3, 19, -18, -4, -31, -8, -25, -25, -15, -23, 13, -27, 18, 19, -2, -4, -49, 23, 24, -25, 6, 23, -34, -30, 0, -6, 71, 35, -23, -1, -55, -13, 13, -64, 18, -24, -44, -35, 10, 12, -43, -26, 16, -37, -17, 23, 1, -7, -10, 0, -20, -53, -43, -51, 28, 34, -27, -1, 13, -24, 34, 75, -10, -23, 15, -8, 3, -2, 7, 48, -29, -87, 19, -55, -5, -23, -3, 15, -4, 17, 9, 20, 14, -20, 31, 13, 23, 3, 15, -16, -47, -4, 18, -12, 7, 3, 38, 25, 12, 18, -20, -27, 7, 14, 13, 19, 39, -46, 46, -26, 18, 32, -15, 8, -11, 10, 6, 3, -9, 20, 25, 13, -18, -11, 38, -1, 28, -40, 45, 14, -12, 2, 23, 22, 22, -32, -15, 2, -5, -36, -17, 26, 22, -1, -29, 8, -15, 1, 14, -6, -16, 9, -13, -41, -41, -18, 39, -8, -31, 18, 21, -20, 10, 40, 8, 10, 14, -65, -25, 49, -40, -7, 40, -31, 22, -7, -42, 55, -16, -5, 17, -23, -21, 24, -23, -26, 24, -20, 51, -46, 20, -17, 35, 0, -21, 1, -43, -30, 28, -40, -11, -17, 8, -53, 25, 26, -36, -12, -33, 13, -52, -9, 37, 4, 8, 31, 21, -25, -5,
    -- layer=3 filter=0 channel=2
    -11, -4, -16, -11, 0, -7, -12, -17, 1, 12, -32, -9, -20, -7, -11, 12, 7, 27, 0, -13, 0, 25, -23, 4, 5, 37, 0, -8, -20, 1, -15, -11, 11, 5, 8, -35, -2, 18, 21, 9, 13, 23, 31, -37, -3, 6, 1, -12, 0, 50, -18, -12, -14, 25, 25, 26, 15, -17, 21, -14, 0, 17, 5, 2, -23, -22, -14, 7, -30, -5, -1, 13, 21, -10, 5, 9, -9, 11, -30, 5, 0, -13, 54, 29, -35, -38, 24, 0, 19, -5, -5, -16, 1, 2, -32, 2, 11, -5, 0, 21, 7, -21, 14, 23, -27, 12, 21, -9, 9, 24, -8, -7, 42, -11, 19, 0, -13, -25, 21, -6, 10, -6, 1, -6, 8, 13, -9, -5, -10, 9, -13, 4, -45, -34, -5, 13, 21, -10, 1, -17, 5, 0, 11, -7, 3, -28, 30, -17, 1, -10, 2, 16, 17, 6, -11, 1, 4, 9, 6, -7, 25, -4, 5, -24, -17, -7, -4, 12, 15, -21, 16, -8, -20, -23, -7, 1, 0, 0, -18, -7, 16, 22, -19, 21, -28, 8, -17, -23, 54, -9, 2, 4, -20, -7, -8, 15, -24, -19, 35, -24, 41, 17, -18, 37, 1, -27, 10, 38, 23, 21, 14, -20, 16, 17, 12, 16, -26, -29, 18, 18, -19, -19, 33, -15, -19, -16, 38, -48, 40, -5, -10, 8, 36, 36, 6, -12, -3, -21, 16, 11, 9, 2, 1, 10, -44, 19, -6, 11, -23, 25, -23, 7, 10, -7, -9, -46, -27, 5, 35, 8, 5, 21, -4, -4, 0, -13, 31, 22, -30, -22, -12, 6, 35, 11, 37, -27, -19, -13, 0, -18, -3, 4, -93, -26, 1, -27, 13, 8, -25, 28, 11, 18, 8, 0, -3, 6, -40, 0, 6, 6, -9, 18, 16, -26, 52, -19, -18, -9, -3, -23, 8, 1, 16, -7, -15, 4, 10, 23, 26, 16, -51, 30, -11, -20, 12, -37, -29, -18, -13, 12, -19, 48, 16, -8, 28, -23, 35, 19, 56, -11, -12, -10, 7, 13, 36, 0, 32, -7, -18, 8, -21, 2, 6, -31, 48, 19, -1, 17, 4, 30, -6, 17, -16, 44, -8, 14, 19, 34, 28, 10, 6, -29, -3, -9, 0, 7, 2, -10, -3, -19, 37, 18, 17, -16, -43, 23, 5, -3, -22, -4, 35, 20, 25, 13, 16, 23, 20, 30, 1, 0, 19, 6, 22, 0, 14, 10, 27, -12, -14, -19, 45, 0, -42, -33, 12, -9, 22, -27, -25, -27, -8, 16, 30, 29, -5, 29, -39, -5, 30, 20, -12, 30, 3, -2, 0, 15, 0, 9, -2, -7, 10, -8, 4, 18, -6, -18, 48, 19, 9, 3, 42, -17, 17, -23, -28, 22, -26, -15, 18, 20, -4, 53, -21, -29, 5, -23, -2, -33, -18, 5, -8, -7, -49, -10, -31, -16, -23, 4, 30, 23, -7, 10, -32, 2, 6, -9, -7, 15, 18, -28, -33, -50, 3, 8, -16, -18, 48, 18, 3, -24, -8, 6, -16, -26, -17, -17, -4, -18, 31, -22, 24, 25, -12, -32, -22, 8, -21, -45, -11, 13, -27, 0, 35, 5, 12, 15, -25, 8, -7, -28, 4, -16, -12, -13, 4, 16, -27, -10, -4, -30, -23, -1, 0, 11, 15, -33, 37, 2, -16, 12, -3, 37, 18, 29, -11, -30, 28, 2, 22, 38, -5, 6, -34, 27, -22, 27, 5, 6, 19, 20, -1, -37, 12, -2, -5, 2,
    -- layer=3 filter=0 channel=3
    -9, 17, 28, 4, 9, -9, 20, -18, -31, 2, -29, 0, -2, -9, -13, -27, -15, 10, 14, -6, 1, -31, -13, 11, 40, -7, -21, -7, 24, 37, 8, 4, -23, 12, 16, -12, 9, 13, 28, 13, 10, -38, 37, -6, 30, 3, 26, 10, 14, -23, -10, -2, 12, -5, -1, 13, 8, 1, -33, 5, 25, 17, 3, -26, 22, -23, 15, -11, 8, -7, -10, 0, -19, -22, 17, 10, 13, -15, 35, -20, 6, -14, -7, -11, 3, 2, 0, 18, -13, 8, -22, 7, -4, -16, 11, -5, -16, 18, -9, -5, 9, -1, 16, -16, -9, 1, 16, 18, 0, -14, 11, 9, 6, 11, 6, -9, 21, 17, -5, -34, -4, -12, -32, -24, 17, 0, 29, -17, 36, -7, 23, 6, -13, 4, -19, -7, -17, 6, -10, 0, 3, -11, -22, -11, 0, 12, -34, -9, 11, -39, -29, -4, -3, 4, -7, -1, -17, 17, 20, 27, -23, 11, 3, -24, -20, 14, 26, -18, -17, -16, 12, 14, -6, 23, 1, -30, -15, 11, -31, -25, -17, 13, -18, -43, -7, -16, 6, 14, 28, -17, -3, -12, 10, -4, 8, 5, -13, -17, 11, 1, 1, -22, -17, -12, -45, 14, -18, -20, -3, 21, -6, 4, 11, -2, 17, -22, -26, 22, 5, 18, -13, 3, -20, -22, 12, 12, -15, 13, 15, -36, -8, 8, 21, -9, -21, -9, -4, -11, 34, -20, 8, -22, 2, 8, 4, -4, 16, -8, 25, -13, 0, 15, 16, 7, 33, -3, -19, -43, -5, 38, -24, -15, -11, -19, 15, 3, -14, -19, -31, 15, 20, -26, 25, -37, 14, 0, 24, -11, 17, 21, 11, -9, 4, -5, -27, -2, -9, 0, -16, -26, 24, -15, -22, -31, 0, 20, 15, 13, -19, 18, -16, -10, 17, -2, 3, 23, -70, 36, -1, 12, 5, -9, -23, -6, -38, -17, 0, 14, 62, 28, 24, -44, 13, 26, -42, 1, 3, 14, -12, -3, -32, -17, -16, 16, -16, -16, 5, -17, 0, -23, 19, 3, 5, -3, 10, 27, -12, -8, -19, -25, 14, -18, -16, -37, 9, -3, -8, -1, 8, 25, -12, -17, 2, 27, 20, -12, 3, 11, -7, 35, -14, 14, 11, 26, 23, 2, 7, 4, 1, 30, 29, 16, 14, -2, -7, 6, 18, -16, -40, 6, 9, 13, -16, 0, 16, 43, -20, 14, -24, -17, 2, 12, -3, -24, -6, -11, 13, -4, 11, 27, 3, -28, 0, 27, 3, 14, -1, -36, -3, 9, -4, 19, -23, 5, 27, 25, -17, 27, -4, -9, -4, -2, 16, -15, -6, -6, -6, 20, 5, -16, -10, 15, -3, -43, 53, -25, 11, 35, -8, -26, -25, -23, 9, -16, -3, 11, 15, -1, 17, -4, -13, -16, -29, 28, 2, 0, 37, 7, -9, -39, 12, 11, -11, 12, 17, 15, 5, -7, 7, -4, -23, -39, -2, -24, -15, -15, -25, -6, 7, 22, -16, 7, 10, 12, 3, 15, 16, -23, -9, 12, 5, 1, -26, 2, -14, 2, -11, 0, 0, -23, -2, 13, -34, -25, 6, 16, -45, -41, 15, -31, 1, 4, 14, -1, -17, 33, -43, 5, 5, 3, 26, 8, 8, 14, 11, -37, -16, 0, 30, -30, 18, 15, 27, -7, 12, 6, 8, -7, 14, 25, -6, -22, -11, 31, 10, -3, 23, 3, 11, -20, 17, -21, -38, 11, -12, -5, -2, 13, -8, -5, 16, -7, -14, -23, 0, 18,
    -- layer=3 filter=0 channel=4
    8, -17, -37, 1, 16, -10, -1, 12, -37, -40, -6, -8, 15, -25, 0, 5, 13, 40, -23, -28, 37, 0, 0, 33, 6, 12, -24, -20, 39, 15, -31, 15, 2, -54, -45, -3, 14, -12, -8, -24, -18, -35, 8, -9, -5, -18, 8, -3, -48, 10, 26, 6, 15, 25, 11, -10, -18, 6, -1, -30, 0, 10, -4, -20, -4, -1, -12, -7, -18, -56, 4, -1, 24, 22, -27, -11, 0, -5, 20, -2, 24, 22, -49, -11, -13, 42, -11, 46, -6, -16, -8, -3, -26, 37, 12, -22, 10, -18, -2, -26, -33, 11, -18, 14, -20, 13, -9, -15, 8, -3, -1, -16, -78, 14, 11, -2, -1, 28, 23, 27, -14, -9, 25, 15, -5, 7, -10, -100, -13, -2, 0, -7, 2, -22, 14, -6, -2, 0, -2, 43, -21, -14, 36, 10, 8, 0, -106, -3, 23, 52, 23, 25, -19, 16, -15, 17, 28, 6, -20, -17, 7, -20, 16, -23, -17, -21, 1, -28, 10, 20, -11, -4, 30, -13, -34, 14, -85, 32, 2, 6, -15, -19, -19, -12, 3, -30, -24, -18, -19, -22, 20, -40, -16, 34, -7, -19, 13, -4, 12, 17, 15, 8, 22, 31, -18, 23, -30, -9, -27, 40, -18, 1, 33, 0, 26, -9, -23, 22, 12, 11, 28, 6, 5, -23, -8, -18, -61, -8, 6, 5, -5, -13, 0, 30, -14, 6, -13, 20, -9, 13, -25, 10, -11, -30, 8, -27, -5, 12, -3, 14, 12, 7, -54, -4, -11, 1, -2, 13, -21, 20, -6, 24, 10, 24, -1, -8, -15, -9, 16, -9, -9, -26, 7, -37, -40, 25, -5, -78, 36, -7, -16, 31, -9, -19, 12, 19, 5, 14, 18, 27, -35, 54, 1, -17, -21, -4, -15, -1, 26, -4, -23, 0, -9, -21, 17, -11, -67, -32, -4, -34, -14, -15, 14, -25, 11, -13, -24, 7, 15, -5, -29, -3, 9, 16, 0, 0, 11, 0, 5, 20, 23, 1, -1, 0, -33, -29, 24, -9, -38, 25, -12, -4, -44, 11, -3, -11, -8, -13, 8, -25, -17, -27, 16, 2, -3, 43, 11, 12, -17, -24, 16, 13, -36, -27, 19, 1, 30, -3, 11, -16, -35, 24, 18, 14, 3, -20, -15, 2, 21, 16, -11, -12, 12, -33, -2, 43, 43, 20, 11, -35, 4, -17, 36, 19, 4, -20, 14, -2, 4, 21, 28, -15, -36, -14, 39, -13, -9, 24, 18, 0, -7, -27, -5, -18, 31, -12, 21, 15, -25, 5, 13, -33, -33, 30, -14, 0, -31, 29, -16, 25, 6, 32, -50, 2, 6, -4, 15, -21, 13, 15, -29, -31, 15, -5, -26, 18, -8, 14, -7, 11, 37, 11, 5, -24, 7, 24, 42, -1, -18, -40, -29, -14, 22, -34, 30, 14, -18, -10, 18, -14, -34, 0, -12, 4, 8, -27, -11, 16, 8, 8, -17, -20, -26, -44, 44, -32, 2, 24, -8, -28, 23, -5, 23, -15, 0, -52, -1, 17, -20, 9, -25, 32, -4, 8, 11, -76, -33, -1, 0, -14, -5, 0, 9, 15, -11, 6, -8, -8, 21, 6, 24, 19, 9, -21, 26, 12, -8, 0, 10, -23, -7, 6, -18, -25, -29, 31, 18, -18, -25, -3, 18, 17, -20, -26, 11, -42, -1, -11, 30, -52, 12, 13, 10, -4, -5, 0, -29, -12, 26, 0, -37, 19, -37, 34, -12, 18, -25, 4, 3, 28, -21, 16, -13, -1, -26, 15,
    -- layer=3 filter=0 channel=5
    -5, 16, 39, 34, 28, -19, 29, 3, 7, -18, -3, 0, 1, -18, -25, -41, -19, -3, 25, 23, -12, 0, 11, -1, -5, -11, 1, 33, -11, 5, -31, -21, -1, 21, 25, -31, -46, 32, 19, -10, 5, -30, 18, 5, -19, 11, 0, -29, 23, 22, -33, 17, -12, -27, -6, 0, 22, -2, -17, -25, 6, 10, -28, 0, 40, 22, 13, 34, 40, 20, 11, 4, -43, -25, 31, 10, 17, 4, -12, -13, 12, 10, 22, 34, 10, -91, 24, -23, -8, -32, 2, 13, 14, -9, -22, -23, -21, 15, -4, -2, 31, 0, 25, -12, 27, 25, 0, 3, 17, 8, 21, 4, 21, -13, -18, 28, 29, -1, 6, -38, 9, 2, -60, -19, -35, -13, -3, -21, -9, 21, 19, 20, -28, 8, 2, -16, 0, 16, -6, 0, 12, -7, 16, -5, 36, 13, 18, 8, 0, -40, -46, -37, -23, 6, -40, 2, 31, -2, 25, 13, -9, 0, -14, -19, 43, -18, -16, -11, -3, 11, 30, -33, 19, -12, -22, -52, 16, 6, -38, -4, 49, 17, 9, 1, 8, 19, -43, -3, 30, -26, -7, 17, -16, 13, 1, 9, -18, -27, 0, -12, 28, 13, -22, -2, -29, 4, -16, -50, -3, 28, -15, -19, -3, -15, 19, -1, 28, 4, -9, 5, 4, -7, -23, -3, 21, -19, 2, 14, -30, -17, -1, 26, 17, 15, 5, 9, 13, -4, 11, -48, -22, 16, -34, 41, -5, 7, -14, -6, 2, -36, -10, 17, 30, -21, -30, 3, 13, -15, -15, 1, 17, 12, 1, 25, -2, -33, -38, -13, -26, 13, 1, -10, -14, 1, 23, 12, 21, -14, 12, -5, -13, 33, 15, -15, 15, -5, -9, 15, -5, 15, 1, 15, -21, -27, -15, -11, -19, -29, 42, 36, -13, -12, -13, -24, -40, -13, -34, 33, -13, 4, 0, -34, -10, -30, -10, 30, -6, 5, 3, -43, -22, -14, 17, 12, -34, -38, -23, 11, 8, 31, -5, -26, -26, 21, -12, 10, 45, -37, -47, -1, -13, 13, -35, -8, -21, 16, -9, 2, -21, 15, 0, 12, 21, -27, 0, -17, 2, 14, 0, 8, -7, -9, 13, 24, 0, 5, 0, -32, 6, -18, -39, 2, 18, 22, 9, 9, 21, -22, 2, 3, 32, 10, 8, 3, -59, -11, 29, 2, -33, -16, -16, 10, 2, 14, -19, 2, -30, -5, -22, 9, -18, 46, 18, -15, 7, -6, -9, 0, 46, 10, 3, -12, -18, 25, -29, -26, 7, -5, -4, -9, -6, 4, -16, 5, 7, -1, -36, 31, -6, -12, 36, -39, 29, -7, 4, -9, -37, -4, -13, -5, -14, -14, 19, -5, -6, 1, -19, 43, -12, -49, 2, -19, -4, -13, 26, 7, 0, 8, 0, -16, -1, 6, 7, -27, -25, -15, 11, 3, 13, -50, -22, 14, 19, -12, 21, -11, 52, 3, 4, -26, -6, -23, 9, 1, 13, -1, 6, 2, 1, 1, -17, -11, 7, -16, 13, 5, 8, -43, -58, 0, -2, 9, 21, -14, -25, -26, 3, 17, 20, 8, -42, 13, -14, -20, 2, -9, -46, -28, 24, -11, -23, -15, 14, -64, -21, 34, -12, -10, 13, -14, 5, 23, -12, -24, -36, 0, -1, -8, 3, 17, -3, 22, 5, 0, -2, -39, -35, 10, 24, -6, 15, 0, 17, 17, 6, 10, 31, -22, 8, -62, 3, -42, -27, -13, -17, 13, 2, 27, 21, -28, 5, -19, -10, -28, 3, 20,
    -- layer=3 filter=0 channel=6
    6, -31, -22, 2, 5, 8, -38, -14, 25, -28, -7, 0, -13, 9, 42, -19, -31, -11, -8, -14, -11, 24, 16, 48, -20, -7, 25, -15, -21, 28, -11, 19, 6, 29, -52, -33, 31, -4, 3, -10, -16, 0, 11, -42, 40, 15, -20, -50, 16, -4, -15, 31, -22, -21, -4, 11, -24, -31, -12, -4, 32, 10, 22, 18, 23, -49, 10, -28, -42, 11, 23, -28, 26, -10, 37, 19, 31, -57, 40, -16, 16, -25, 20, -57, -11, -17, -14, -4, 4, 21, 4, 3, 14, 12, 10, 5, -24, -5, -69, -2, -13, -50, -22, -3, -43, 1, -21, -22, -12, 14, -40, 21, -21, 36, 17, -4, -1, -21, 6, 32, 10, 17, 10, 24, -7, 16, -24, 18, 10, -65, -53, 26, -30, 2, -49, 4, -3, -39, 19, 17, 0, -10, -20, -49, 13, -20, -28, -16, -35, 29, -14, 16, 13, -4, -18, -13, -1, 3, 27, -22, 0, 41, -12, 5, 12, -23, -3, 1, -30, -24, 12, -24, 7, -6, -20, 9, -1, 29, -14, 18, -2, -5, 19, -29, -6, -30, -21, -3, -66, 22, -12, -24, -4, -47, -26, 17, -57, 26, -36, 14, -19, -6, 1, 12, 13, 14, 0, 8, 14, 1, 13, -54, -31, -1, 9, 16, -38, 51, -33, -32, -22, 36, -5, -25, -16, -7, 37, -30, 14, -27, 10, -20, -17, 32, -6, -29, 0, 10, -31, -62, 4, -9, 18, -5, 4, 26, 17, 0, 1, 28, -13, 6, 58, -2, 5, -42, 9, -70, 8, -1, -82, -12, -22, 17, 2, 43, 9, -40, 32, 0, -15, -18, 17, 17, 30, -15, -26, -17, 20, 2, -18, -37, 9, -17, -101, 10, 11, 9, 23, -5, -2, -39, 27, -11, -25, 8, 30, 32, -46, -60, 11, 20, 19, -18, 21, 41, 19, 13, -38, 40, -2, 60, -20, -18, -15, 35, 85, -5, -4, -1, -11, -29, 3, 8, -65, -7, -21, -12, 7, -25, -7, -29, 2, 25, 45, -37, 16, -3, 52, -2, -2, -21, -12, 24, 2, -2, -18, -4, -46, -41, 46, 3, 8, -14, -21, 40, -6, 26, -14, -21, -3, -10, 65, 5, -13, 19, -15, -51, 49, 42, 10, 7, 0, -3, -24, -2, -22, -15, -15, 28, -27, 12, -63, -36, 13, -54, -4, 22, -62, -25, 22, 19, -25, -8, -26, -14, 19, -14, -17, 10, -13, 10, -5, -22, 16, -29, 29, -2, -37, 32, 14, 16, 12, 51, 12, 27, 15, -23, 8, -73, 31, -27, -5, -13, 37, 38, 25, -8, -21, 21, -7, -58, -2, -25, 9, -11, 7, 17, 22, 18, 9, 1, -9, 1, -21, 18, -4, -54, 3, -1, -35, 1, 1, 5, 2, 23, -14, -23, -1, -45, 41, 27, 25, -10, -4, 5, 8, -15, -3, -21, 40, -8, 2, 40, 14, 7, -44, -4, -22, 16, 16, -30, 24, 27, 11, 2, 2, -37, 60, 2, 37, 23, 28, 19, -13, -30, -13, 0, 0, 20, 39, -12, 0, 9, -4, -25, -7, -13, -4, -12, -14, 7, 2, -39, -26, -5, 9, -48, -8, -7, -7, -21, -24, -11, 37, 36, 10, -36, -15, 17, -21, 7, 35, -5, -21, 11, 22, 55, 68, 5, -8, 18, -5, 16, 16, 14, -20, -7, 11, -3, -33, -13, 41, 11, -15, 23, 51, -26, -16, -50, -11, -2, 0, -10, 48, -22, -15, -30, -15, -26, 5, -1, 0, 0, 14, -50,
    -- layer=3 filter=0 channel=7
    -25, 2, 13, -34, -16, 31, -16, 18, -12, -27, 32, -35, -19, -10, -12, -23, 21, -12, -17, 34, 23, 16, 38, -28, 2, 8, 10, -24, 22, -11, -13, 0, 16, -17, -18, 49, 5, -6, -15, -52, -30, 12, 14, 33, -6, 4, -49, 12, -33, 1, -1, 30, -6, -30, -6, 13, -1, 19, -7, -21, -33, 13, -44, 19, 15, 56, 10, 10, -42, -23, 19, -14, 18, -11, -12, 19, -26, 47, -64, 24, -11, -3, 11, 6, -9, 1, 37, -18, -30, 9, 1, -43, 28, -1, -33, 7, -22, -13, 8, 5, -2, 41, 9, -37, 68, -42, 34, 26, 6, -1, -2, -44, -14, -58, -8, 1, 39, -28, -22, -41, -5, 17, 11, -4, 22, 1, -16, 8, -41, -5, 0, 3, -17, 1, 23, 16, 14, -20, 22, 1, 16, -9, -8, 42, -60, 14, 2, 27, -6, 31, 28, -8, -24, -43, -16, -9, 4, -11, -29, -13, 19, -24, -29, 42, 0, 9, -16, -50, 3, 11, -2, -18, -7, -20, -16, 2, -22, -61, -12, -16, 30, 0, 18, -27, -14, 19, 34, 28, -27, 3, -3, 38, -10, 44, 1, 46, 37, -40, 6, -23, -18, -26, 10, -35, -16, 33, 14, -20, -14, 8, -9, 2, 50, 17, -24, -23, 48, -16, -22, 12, 5, -12, -7, 7, -19, 9, -23, 12, -31, -33, -27, -2, -31, -50, 34, 1, 35, -13, 16, -19, 26, 26, -24, -35, -30, 14, -15, 8, 0, 0, -6, 6, -82, -2, 11, 36, 2, 21, -15, 23, -51, -3, 8, -19, -23, 34, 43, -19, 3, -36, 20, 20, -19, -55, -53, 6, 0, -69, -51, -31, 1, -13, 60, 7, 2, -6, -1, -11, -14, 9, -11, 2, 14, 22, 12, -11, -6, 3, -7, 30, -41, -14, 43, 13, -29, -7, -13, -18, 47, -19, 10, -12, -24, -47, -43, -24, -52, 19, -74, -41, -23, 30, 21, 33, -41, -2, 37, 20, 0, -17, -7, 24, -18, -28, 27, 1, 10, -43, -6, 21, 18, -3, -4, 16, -42, 12, -16, 6, 32, 37, -39, 12, 21, -30, 31, -6, 27, -37, 10, 33, 1, 28, -62, -17, -14, -10, 13, -43, 7, -36, -36, -10, 20, 26, -7, -42, 0, -14, 10, 21, -16, 11, -68, 32, 21, 29, 24, 32, 37, -24, 14, -27, 6, -21, -28, -31, 12, 31, 40, 38, 42, -4, -79, 19, 38, -43, 1, 1, 43, -3, 23, -12, -10, 25, 42, -10, -18, 2, -52, 32, 12, -21, -9, 14, -10, -55, -19, -6, 16, -4, 1, 7, -63, 1, 4, -37, -28, 26, 8, 9, 0, -27, -22, 4, -39, -15, 5, 15, -14, -5, 35, 23, 14, -23, -59, -16, 29, 31, -42, 41, 18, -25, 24, 16, 33, 30, -61, 5, 23, -1, -15, 34, 16, -28, -11, 0, 0, 8, 16, -7, -8, -35, -33, -33, -16, -50, -13, 31, -44, 2, -21, -18, 19, -15, -3, 0, -2, 32, -31, -49, -50, 31, -3, 35, -19, 21, -13, 28, 6, 20, -50, 45, -19, 0, 26, 31, -15, -7, -17, -23, -18, 0, -17, 11, 37, -28, 14, -13, -8, 29, 2, 2, -8, -1, -12, 32, -9, -33, -32, -42, -31, 6, 18, 1, -15, -71, -33, 22, 8, -18, -16, 46, -28, -16, 5, -4, -34, -8, 6, 5, -37, 23, -6, 40, -28, 2, 2, -27, -1, -22, -21, -2, 22, 10, -65, 26,
    -- layer=3 filter=0 channel=8
    0, 17, -2, -34, 0, 33, -15, 3, 10, 27, -40, -17, -18, -12, -32, 13, -12, 21, -32, 18, 32, -14, -3, -6, 9, -5, 48, -8, -15, -20, -20, -16, 0, -24, -6, 19, 41, -14, -33, 31, 1, 15, -64, -9, 0, 17, 11, 26, -59, -25, 3, -5, -34, -18, 5, 9, 17, -6, -9, 3, -69, 1, 32, 28, -22, 21, -6, 7, 26, 5, 9, -1, 3, -11, 0, -14, -24, 17, -41, 4, 29, 17, -12, -22, 5, -5, 14, 9, -13, -19, 29, -57, -34, -9, 3, 6, -9, -2, -5, 18, -12, -34, -11, 46, 3, 11, -31, -2, -21, 21, 1, -6, -35, -24, 32, -18, -11, 30, -5, 29, 0, -28, -1, -31, -43, 4, -29, 16, -3, -12, -29, -18, 46, 6, -6, -16, 18, 25, -5, -11, 9, -5, -20, 2, 6, -2, -6, 9, -2, 5, 20, 9, -1, -3, -1, 6, -15, -58, 1, 9, -10, 8, 8, 26, -12, -1, -11, 4, 36, 28, -27, 12, 0, -10, 31, 40, -20, -35, -5, 14, -21, -1, 3, 2, -13, -6, 14, 15, -21, -14, 3, 6, 25, 15, 3, -3, 26, 16, 12, 7, 8, -16, -1, -4, -34, -22, -26, -15, 5, 7, -18, 24, 4, -25, 0, 31, -6, -28, 8, 2, 32, -11, -15, 16, 3, 11, -41, -15, -22, -3, -13, 21, -34, 2, -19, 34, -15, -5, -10, 3, -62, -42, 14, -17, -20, 4, 8, -2, -15, 8, 6, -33, -61, -15, 35, 44, 17, -26, -12, -4, -22, 23, -8, -22, 0, 6, -47, -12, -10, -6, -56, 20, 24, 16, -16, -1, 0, 18, 2, -7, 13, 24, -46, -27, 16, 3, 25, -13, 23, 24, -15, -5, -10, 2, -16, 33, 1, -11, 14, 0, -8, -6, -1, 32, -50, -61, 10, -21, -14, -10, -4, 27, -3, 14, 31, 9, -27, 9, 10, 3, -29, -8, -43, -3, -20, 36, -16, 6, -14, 24, -13, 8, -14, 8, -54, 0, 8, -35, 5, 1, -16, -2, 17, -16, 2, -39, 3, -32, 59, -5, -24, -5, 12, 16, -21, 32, 10, 0, 3, 12, 19, 24, 19, -13, 12, 19, 1, 20, -19, -74, -4, 11, -6, 23, -7, 6, 4, -26, -17, -7, -35, 17, 42, 4, -14, -11, 27, -40, 29, 14, 29, -12, -51, -17, -8, -19, -28, -8, -62, 13, -37, 17, 72, 5, -62, -43, 21, -16, -18, 31, -39, 4, -19, 32, -74, -7, -20, 10, -33, -52, -20, -27, 1, -29, -40, 34, 3, 15, -2, -12, -21, 6, 99, -54, 13, -8, -6, 18, 7, 55, -10, 16, 37, -69, 38, 9, 8, 23, 27, -22, -4, -60, 1, 22, 28, 14, -2, 13, 53, 3, 32, -16, -38, -11, 0, -9, 22, -4, -77, -20, 27, 6, 50, 22, 35, 5, -21, -55, 29, -20, -5, -12, 21, -15, -19, 12, -5, 1, -11, 48, -37, -56, 28, 8, 22, 47, 29, 13, 36, 33, 25, -19, -23, 2, -14, 20, 29, -11, 7, 18, 46, -53, -12, -6, -14, -40, -23, 21, 26, -19, 4, 9, 17, 33, -50, 53, -69, -25, -2, 4, 20, 12, -43, -26, -14, -35, 22, 10, -4, -33, 25, -34, 43, 2, -17, 12, -6, -21, 3, 48, -5, -35, -22, 4, 4, -30, 64, 26, 0, -1, 29, -43, 6, 23, -13, -20, 0, -23, -4, -7, 23, 7, -45, -2, 91, 29,
    -- layer=3 filter=0 channel=9
    -44, -4, 58, -16, -24, 24, 44, 0, 34, 17, 38, -6, -20, 31, 14, 23, 0, -12, 13, -5, -1, -40, 1, -3, 24, 31, -25, -51, -18, -20, 10, 18, 4, 24, 11, 45, 27, 7, -13, 18, 8, 8, 3, 14, 7, -5, 10, 15, 7, -47, 3, 16, 13, 16, -11, -20, 12, 2, -7, -14, -59, 18, -55, 9, -40, -3, 14, -20, -16, 19, 21, 21, -7, 25, 7, -13, -10, 4, -20, 16, -7, 24, 32, 17, 0, -40, 17, 15, -10, -1, -26, -58, -6, 15, 21, -25, 19, 7, -7, -10, 13, -22, -14, -36, -44, 21, 12, 12, -10, 18, 15, -7, 27, -12, 20, -19, 1, 12, 9, 9, -15, 12, 16, 21, -15, 11, -15, -22, -37, 21, -4, -29, -36, 6, -9, 16, -25, -5, 26, -11, 12, 42, -7, 30, -13, 39, 42, -11, -6, -41, -8, -21, 38, -22, 10, -31, -5, -18, 16, -14, -11, -2, -1, 19, -3, 31, -33, -19, -7, 26, -12, 29, 12, 10, 27, -17, 26, -43, 16, 16, -13, 24, 14, -9, -26, 24, 37, -10, -11, -14, -19, -26, 5, 10, -21, -18, 19, -14, 16, -22, -61, -17, -19, 2, 13, -21, -16, -6, 28, -15, -26, 25, 11, -52, -31, -43, 26, 7, 15, -12, 6, -35, -5, 21, -20, 18, 27, 28, -40, 22, -23, 22, -6, -16, 0, 2, 2, -26, 21, -20, -38, -37, 17, -25, 17, -29, -1, 21, -2, 18, 11, 6, -17, 13, -15, -25, 7, 5, 14, 26, -10, -39, -16, 9, 11, -2, -74, -6, 31, 7, 45, -2, 45, 69, -35, 37, -35, 43, -4, 26, 20, -23, 50, 1, -37, 31, -7, 16, 7, -19, -38, 16, -21, 40, -3, 0, 19, 25, -6, 16, -9, -8, 0, 11, 7, 0, 26, -6, 11, 13, 7, 16, 4, 12, 1, 25, -25, -17, -48, -53, 19, 14, 7, 21, 43, 11, 32, 2, 9, 0, -41, -34, -1, 1, 19, -3, -42, 43, -1, -7, -25, 9, 30, 14, 14, 11, 2, 23, 24, 3, -25, 6, 8, -4, -10, -26, -10, 7, -29, -14, 12, 3, -5, -30, -38, -10, 0, -1, -38, -27, 15, 13, -20, 13, -16, 24, -16, -6, -1, 13, -10, 12, -56, -6, 18, -25, -69, 0, 29, 17, -44, -12, -29, -43, -31, -18, -9, -44, 1, -7, 6, -53, -27, -8, 10, -47, -35, -59, -38, -45, -37, 10, 13, -36, -24, -13, 13, 37, 37, 49, -16, 21, -12, -80, 18, -46, 37, 2, -22, 20, -83, 0, -17, -4, 21, 43, 6, -8, 11, -73, 12, -12, 0, -6, -6, -2, 35, -25, 12, 3, -34, -16, 38, 33, -44, -24, -3, -5, -53, -12, -18, -15, 26, -8, 15, -24, -8, 16, -18, -36, 22, -39, -3, -16, -31, 5, -13, -9, -32, 9, -12, 20, 14, -2, 0, 32, -7, 1, -31, -5, -3, 14, -43, -16, -58, 5, -14, -21, 10, 2, 5, -14, -2, -4, -2, -24, -1, 24, -9, 9, 37, -24, 52, 32, -42, 12, 24, 14, -25, 26, 37, -19, -7, -23, -33, -37, 50, 3, -78, -33, -52, -5, -14, -16, 34, -32, -51, 0, -53, 10, 20, 11, -27, 16, 21, 34, 0, 0, -52, 4, -18, -4, -34, -25, 21, -7, -37, -14, -82, 20, -61, -2, 1, 10, 6, -28, -9, -35, 7, -35, -47, 16, 22, -7, 32, -2,

    others => 0);
end iwght_package;
