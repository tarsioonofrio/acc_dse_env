library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package inmem_package is
  type mem is array(0 to 4000000) of integer;

  constant input_mem : mem := (
    -- bias
    28383, 475, 834, -13, -9146, 1779, -21610, -12738, 17147, -7762,

    -- weights
    -- filter=0 channel=0
    21, 22, 10, 3, -1, 6, 9, -1, 2, 2, -3, 4, -5, -5, 1, 7, 7, -2, -1, 0, 6, 0, -1, -1, 4, 7, 10, 17, 24, 29, 3, 7, -6, 2, 4, -6, 2, -11, -11, -10, 0, -8, -3, 1, 3, 0, 2, -4, 0, -5, -1, -11, -8, 1, 5, -7, 0, 4, 13, 21, 4, 4, 4, -9, -11, -5, -7, -10, -1, -9, -8, -4, -1, 1, -10, -3, 2, -9, -13, -6, -12, -6, -16, -15, -4, -6, -1, 6, 1, 24, 6, -10, -11, 0, -6, -4, -2, -8, -11, 6, -7, 0, -6, 5, -6, 0, 4, -14, -4, -17, -8, -12, -10, -11, -1, -5, -2, 0, -4, 19, -5, -4, -4, -8, -4, -4, 0, 1, 0, 5, 5, 7, 0, 9, -4, -1, -5, -7, 0, -6, -20, -20, -16, -13, -16, -2, 2, -4, 3, 7, -4, 1, -2, -8, -3, -3, -12, -1, -8, -5, -5, 0, -3, 4, 5, -2, 7, -4, -1, -17, -18, -15, -10, -12, -10, -10, -9, -5, -3, 5, -3, -6, -12, -2, -6, -12, -15, -7, -7, -7, -5, -3, 12, 13, 7, 12, 4, 3, -3, -8, -17, -16, -14, -9, -9, -12, 0, -3, 2, 11, -5, -4, -3, -8, -12, -4, -14, -17, -9, -13, -10, -2, -2, 13, 14, 4, 2, 1, -8, -10, -2, -6, -10, -5, -18, -4, -11, -9, -10, 1, -4, -1, -3, -16, -11, -8, -15, -16, -13, -12, -2, -1, 7, 8, 20, 19, 14, 8, 2, -3, 2, -11, -16, -13, -15, -18, -16, -5, -8, 0, -4, -8, -4, -9, -10, -8, -9, -16, -11, -5, -10, 8, 3, 10, 7, 8, 20, 15, 4, 3, -3, -11, -5, -13, -9, -9, -17, -14, -10, 10, 0, 0, -4, -13, -8, -12, -9, -4, -6, -1, 1, 8, 15, 14, 18, 22, 8, 6, 4, 3, -2, 0, -7, -7, -12, -13, -15, -13, -12, 12, 3, 0, -9, -16, -6, -17, -19, -10, -16, -8, 0, 5, 1, 22, 11, 28, 17, 20, 16, 7, -3, -13, -1, -5, -10, -5, -16, -16, -1, -3, 9, -9, -5, -1, -2, -2, -11, -7, -14, -15, 3, 1, 8, 21, 16, 29, 27, 27, 18, 7, -1, -10, -10, -18, -7, -14, -5, -15, -10, 6, -6, 0, -15, -8, -18, -18, -12, -11, -14, -8, -6, 0, 14, 22, 20, 32, 30, 24, 29, 19, 0, 1, -6, -7, -12, -21, -16, -5, -9, 3, 4, 4, -2, -2, -16, -9, -5, -4, -4, -2, -9, 4, 1, 13, 26, 31, 28, 21, 29, 13, 6, -2, -11, -20, -6, -9, -19, -4, -4, 6, 0, 3, -2, -16, -7, -3, -13, -18, -12, -3, -3, -3, 3, 25, 23, 29, 28, 24, 20, 19, 2, 0, -13, -7, -10, -19, -19, -18, -12, -1, 9, -9, -2, -2, -14, -16, -6, -15, -1, -11, 1, -5, 6, 11, 28, 24, 29, 32, 25, 4, 4, -4, -1, -19, -17, -19, -10, -9, -10, 5, 9, -6, -12, -8, -11, -17, -9, -11, -4, -4, 1, 6, 5, 13, 18, 18, 16, 14, 12, 11, 5, 4, -5, -9, -11, -13, -18, -2, -11, -2, 5, -7, -13, -1, -2, -8, -16, -4, -3, 0, -3, -4, 0, 7, 19, 25, 15, 17, 3, 0, 2, -3, -12, -8, -7, -4, -7, -7, -7, 1, -2, 2, -13, -10, -11, -17, -9, -9, -6, -6, -10, 3, 12, 14, 16, 23, 13, 5, 12, 0, -5, -7, -13, -6, -9, -12, -17, -9, -1, 1, 3, -6, -10, -15, -3, -14, -19, -16, -16, -12, -10, 8, 0, 11, 9, 19, 19, 7, 0, 0, -1, -7, -5, -11, -12, -4, -17, -5, 0, 9, -2, 0, -2, -12, -10, -9, -3, -18, -7, 1, 1, -7, 2, 7, 4, 8, 12, 0, -2, 4, -6, -6, -4, -14, -13, -6, -8, -13, -8, 13, -2, -7, -14, -12, -2, -6, -6, -5, -6, 0, -5, 1, -1, 1, 12, 9, 11, 9, 6, -7, -5, -13, -4, -18, -11, -18, -10, -2, -8, 15, -4, -5, 0, -4, -14, -15, -10, 0, -5, 2, 6, -7, 10, 7, -1, -2, 0, 6, -11, -8, -16, -20, -9, -5, -4, -16, -7, -4, -7, 14, 8, -3, -4, -15, -1, -4, -5, -12, -3, -7, 4, 0, 1, 8, 11, 3, 8, 1, -7, -8, -12, -6, -21, -7, -5, -2, -6, -1, -7, 17, 9, -2, -7, 0, -3, -10, -7, 0, 0, -8, -4, 2, 4, 2, 1, -2, 3, -4, -8, -8, -16, -5, -9, -12, -6, -9, -6, -6, -8, 12, -4, 7, -10, -10, -13, -6, -4, 2, -4, -4, 3, 1, -8, 5, 5, 0, -5, -11, -7, -2, -5, -20, -4, -8, -15, -2, -10, -11, -6, 20, 3, 1, -6, -3, -7, -4, -5, -4, -2, 0, 0, -2, 5, -1, 1, 4, -11, -1, -11, -13, -10, -4, -2, -14, -10, -9, 1, -5, 5, 14, 14, 8, 7, 0, -8, -7, -8, -8, 3, -4, 1, -8, 1, -1, 5, -2, -9, -1, 0, 0, -10, -8, 1, -11, -7, 3, 4, 0, 18, 31, 23, 23, 18, 12, 4, 10, 5, 1, 6, 3, 5, 3, -4, 10, 4, 0, 4, 6, -2, 6, 8, -3, 9, 5, 6, 1, 21, 18, 24, 33,
    -- filter=0 channel=1
    0, 9, 9, 3, 10, 15, 5, 14, 7, 9, 0, -2, 0, -6, -9, -7, -14, -5, -5, -8, 0, -7, -2, -7, -10, 1, 0, -10, -8, -10, -1, 0, 15, 14, 17, 12, 14, 11, 8, 0, 0, 1, -11, -6, -7, -1, -13, -6, -8, 1, -10, 0, 0, 1, 0, -4, -9, -13, -9, -8, 5, 3, -1, 11, 0, 3, 6, 0, -4, 1, 2, -12, -7, -7, -15, -16, -8, 2, -5, -4, 0, 5, 1, -3, -3, 2, -3, -15, -9, -9, 10, 1, 9, 10, 4, 16, 1, 12, 5, 2, 0, -2, -15, -19, -12, -14, 1, -8, 1, 5, 2, -2, 6, -1, -3, -8, 0, -5, -9, -1, -1, -3, 10, 4, 4, 16, 4, 13, -2, 4, -3, -2, -6, -22, -9, -9, -2, 1, 2, -2, 0, 11, 6, -1, -1, 3, -11, -6, 1, -11, -7, 0, -1, 8, 1, 11, 15, 4, -1, -3, -7, -8, -20, -24, -22, -4, -6, 0, 6, 0, 12, 3, 11, 6, 12, 7, 0, -3, 1, 4, 2, -5, 0, 14, 13, 6, 8, 15, 2, -4, -4, -15, -19, -20, -10, -4, -8, 6, -1, 8, 4, 1, 12, 8, 9, 7, -7, -8, -9, -1, -4, 5, 3, 13, 0, 10, 11, 13, 4, 5, 0, -9, -12, -24, -22, -21, -10, 1, -2, 13, 14, 8, 11, 22, 9, 3, 2, -3, -5, 3, -6, 0, 11, 10, 0, 13, 18, 6, -1, -5, 0, -19, -12, -16, -12, -12, -11, 2, -4, 3, 11, 20, 14, 20, 6, 8, 11, -6, -8, -7, 0, 8, 4, 5, 2, 3, 5, 11, 8, 5, -10, -12, -20, -25, -21, -10, -8, 1, -1, 4, 3, 9, 8, 22, 24, 15, 15, 3, -4, -7, -6, 11, 10, 8, 8, 17, 2, 0, 9, 0, -6, -21, -21, -32, -30, -15, -5, 3, -5, -2, 15, 7, 23, 17, 13, 14, 0, 2, -5, -3, 4, 5, 0, 14, 12, 3, 17, 10, 7, 3, -16, -19, -20, -19, -31, -17, -15, -6, 4, 0, 2, 14, 12, 11, 14, 8, 2, 7, 0, 4, 0, 12, 14, 9, 6, 10, 8, 8, 2, -7, -4, -25, -19, -20, -23, -20, -4, -5, -4, 10, 10, 17, 5, 23, 20, 12, 8, 1, -3, -1, 5, 0, 10, 17, 5, 11, 6, 0, 6, 0, -18, -15, -33, -33, -22, -19, -15, -6, -1, 7, 14, 1, 18, 17, 19, 21, 9, 10, 1, 6, -5, 11, 15, 12, 13, 4, 16, 6, 6, -10, -8, -27, -29, -31, -38, -23, -10, -10, 5, 13, 1, 7, 11, 22, 23, 8, 15, 12, 8, -2, 2, 8, 12, 11, 17, 14, 13, 15, 0, 0, -20, -22, -27, -38, -24, -18, -11, -4, 1, 7, 9, 12, 14, 19, 9, 17, 5, 8, 3, 2, 1, -2, 8, 8, 11, 16, 8, 7, 0, -6, -13, -21, -24, -25, -21, -17, -13, -12, 3, 9, 13, 2, 12, 14, 19, 13, 16, 7, 6, 0, 5, 11, 8, 4, 13, 13, 7, 8, 6, 0, -11, -14, -19, -29, -29, -27, -11, -6, 2, 8, 7, 16, 9, 23, 23, 18, 17, 12, 6, -4, 2, -3, 14, 3, 10, 11, 10, 10, 8, -2, -3, -15, -32, -27, -32, -21, -13, -4, -7, -1, 14, 11, 13, 13, 14, 11, 13, 2, -4, 1, 5, 9, 10, 10, 3, 8, 16, 7, -3, -5, -7, -18, -21, -18, -22, -8, -7, -3, 6, 10, 12, 7, 11, 9, 11, 6, 2, 4, 5, 1, 9, 4, 0, 9, 7, 11, 19, 9, 7, 0, 0, -8, -13, -22, -24, -12, -14, 5, 2, 12, 12, 19, 15, 18, 10, 19, 10, 0, 6, 2, 0, 12, 7, 7, 12, 8, 14, 5, 7, 0, -12, -16, -21, -15, -13, -20, 0, 2, 8, 9, 7, 4, 15, 8, 9, 5, -1, 0, -3, -10, -1, 3, 2, 17, 13, 6, 20, 18, 5, -5, -5, -13, -19, -15, -24, -11, -10, -6, 3, 12, 8, 3, 21, 14, 14, 12, -3, -4, 2, -3, -2, 1, 0, 6, 16, 20, 15, 7, 10, 3, -4, -18, -14, -11, -9, -19, -9, 1, 8, 0, 17, 5, 11, 11, 11, 1, -4, 5, -2, -8, 6, 10, -2, 16, 3, 6, 13, 4, 2, 0, -9, -16, -24, -23, -19, -10, 1, 7, 0, 9, 0, 11, 4, 10, 0, 0, 3, -10, 1, -9, -3, 9, 2, 12, 14, 17, 3, 6, 5, 4, -4, -1, -5, -9, -18, -17, -4, 4, 4, 7, 0, 4, 6, 0, -2, -3, -8, -9, -11, -6, -1, 7, 2, 4, 9, 6, 1, 4, 0, -1, -2, -14, -17, -12, -17, -17, 0, 4, 5, 1, 4, 10, 0, 3, 1, 2, -9, -6, -1, -4, 4, -1, 0, 12, 10, 8, -1, 9, 3, 7, 0, -12, -7, -8, -16, -10, -6, -7, -6, -9, -4, -7, 4, -2, -9, 0, -10, -17, -1, 0, 12, 10, -2, 13, 8, 12, -3, 9, 2, -8, -9, 2, -2, -11, -5, 0, -11, -4, 2, 0, -6, -3, 3, -10, -2, -8, -13, -3, -11, 1, 9, 0, 8, -1, 10, 2, 3, 2, 5, -2, -1, -5, -1, -6, -4, 0, -3, 0, 0, -7, 1, -10, 3, -2, -8, 3, -7, -9, -6, -8,
    -- filter=0 channel=2
    -2, 0, -6, 6, 5, 6, 0, 0, -6, 3, 3, -8, -4, -11, 0, -6, -10, 1, 0, 1, -5, 4, 4, -3, -7, 0, 3, 1, -7, 6, 2, -4, 3, 8, 4, 6, -9, -1, 4, 0, -9, -4, -7, -12, -3, 3, -6, -1, -8, -11, -5, -12, -2, -2, 3, 5, 7, -3, 2, 4, 8, -3, -7, 3, 0, 0, -7, 4, 2, -5, 2, -5, -3, -4, -10, -7, -6, -7, -13, -14, 2, 2, 2, -1, -5, 5, -6, 6, -2, 3, -7, 4, -1, 0, 4, 5, -6, 0, 1, -10, 0, -9, -5, -3, -8, -15, 0, -13, -5, -11, -3, -9, -4, -2, 2, -1, 5, 4, -3, 4, -6, 3, 7, 3, 2, 5, -1, -1, 0, -2, -7, -2, -3, 0, -15, -7, -14, -8, -9, -5, -10, -2, -12, -13, 3, -3, 0, 6, 1, -2, -4, -2, -4, -4, -5, 0, -8, 0, -9, -11, -6, -8, -5, -1, -9, -3, -18, -7, -10, -14, -2, -12, -2, -1, -3, 5, 1, 0, 5, 4, 4, -5, -2, 7, -3, 6, -2, -8, 1, 0, -14, -11, -15, -10, -16, -11, -3, -17, -14, -6, -10, -8, -9, 0, -6, 3, 2, -7, -7, 0, -2, 1, -5, -1, 3, -6, 0, -7, -5, 3, -13, -3, -12, -14, -4, 0, -7, 0, -5, 0, -3, -11, -13, -1, -3, -3, 3, 0, -1, -4, 6, 3, 2, 8, 6, -5, 7, -6, 2, 5, -3, 1, 0, -5, 4, 0, -4, -5, -10, 0, 0, -4, -3, -3, 1, -2, -5, 8, -4, 3, 0, -3, 9, 7, -3, 5, 6, 0, 4, 0, -4, 4, -6, 4, -3, 1, 6, -5, -3, -4, -7, -1, -3, 0, 2, 0, 0, 7, 5, 8, 7, 1, 2, -6, -4, 4, -4, 3, -4, 8, -3, -2, 5, -3, 10, 3, -5, 4, -6, 0, 4, 4, -6, 0, -9, -4, -3, -2, -3, 0, 0, -1, -1, 6, 6, 6, 2, -3, 12, 14, 12, 4, 2, 1, 15, 11, 12, 2, 11, -4, 0, -3, 3, 6, -4, -1, 4, 0, 6, 0, -5, -4, 7, 4, 8, 6, 2, 0, 12, 6, 19, 4, 7, 4, 17, 0, 3, 11, 2, 7, -3, -3, 4, 7, 9, -3, 2, -2, 11, 11, 1, 2, 5, 9, -1, 7, 12, 12, 13, 18, 7, 14, 24, 20, 5, 8, 2, 8, 14, 14, 0, 2, 2, 0, -1, 11, 10, -2, 7, -1, -4, -2, 2, 3, -2, -5, 3, 2, 13, 11, 13, 21, 17, 9, 11, 9, 17, 18, 8, 15, 14, 11, 6, 8, 4, -3, -1, 4, -2, -1, -3, 0, -1, -2, 8, -3, 11, 13, 13, 15, 14, 25, 21, 10, 11, 17, 13, 6, 12, 15, 3, -2, 5, 9, -1, 5, 1, -2, -2, 10, 9, 9, 0, 9, -1, 10, 0, 0, 15, 16, 21, 20, 18, 16, 16, 19, 12, 9, 11, 7, 9, 11, -3, 2, -4, 11, 1, 2, 1, 11, 6, 6, 3, 7, 4, -3, 6, 14, 5, 13, 13, 13, 8, 13, 13, 11, 6, 9, 15, 12, -2, -2, 7, -5, 0, 5, 0, 13, 11, 0, 6, 0, 1, -5, -4, 1, -3, 8, 9, 3, 7, 11, 15, 11, 9, 13, 6, 8, 10, -2, 7, -5, 0, 0, -5, 3, 7, -2, 4, 4, 0, 5, -1, 11, -4, -2, -3, 2, -2, 9, 8, 11, -3, -1, 7, -1, -2, 12, 8, -4, 7, -6, -3, 0, -8, 0, 6, -3, 6, -1, 9, 9, 0, 1, 6, 10, -2, 0, 0, -4, 7, -1, 2, 6, 6, 1, 6, 3, -4, 3, 2, 0, -4, -8, -10, 7, 2, 6, -2, 12, -1, -5, 8, 2, -3, -2, 5, -8, 5, -5, -8, 0, -3, -1, -1, 0, -9, -1, -10, 0, 0, 0, -1, 2, 5, -3, -1, 6, -4, 9, 1, -2, 12, 10, 5, -2, -3, 0, 2, 1, -9, -11, -4, 0, -5, -9, -6, 0, -7, -10, -3, -4, -10, -6, -6, 3, 8, 5, 4, 5, 2, -2, 2, -2, 3, 5, 4, 7, 6, 0, -3, 3, -11, -5, -16, -1, -4, -4, -5, -1, -4, -1, -6, 1, 3, 1, 7, -3, 0, 0, 4, 1, 1, 3, 10, 2, 0, 7, 1, 2, -6, -1, -10, -7, -8, -12, -16, -11, -1, -7, -12, -1, -10, -10, -9, -3, 6, -5, -2, 6, -2, 10, 9, 4, 6, -2, 0, -8, 2, -8, 3, -2, -6, -4, -8, -10, -1, -14, -11, -14, -4, -2, -1, 0, 2, 6, 8, -3, 0, -6, -1, 4, 2, 8, -2, -2, -4, 2, 3, 1, -8, -2, -4, -12, -4, 0, -11, -12, -9, 2, -6, -4, -9, -9, -3, -2, -1, 0, -2, 6, 7, 9, -6, 7, 5, -5, -1, 5, -6, -1, -4, -5, -7, -5, -9, -7, -12, -8, -2, -11, -11, 3, 1, -5, -3, -1, 5, 2, -6, -5, -1, 3, 0, -6, -1, 6, 3, 5, -8, 2, 5, 1, 3, -8, 2, 0, 0, 3, 1, -12, 0, -1, -8, 1, -8, -2, -3, 4, -2, 8, 5, 3, -5, -5, -1, 5, -1, -9, -2, -6, 5, -9, 0, -5, -8, -4, -3, -2, -1, -11, -4, -4, -4, 1, 0, -7, 8, -2, 2, 6,
    -- filter=0 channel=3
    7, -5, 7, 4, 3, -5, 6, -2, -3, -4, 3, -5, 1, -4, 9, 11, 9, 7, 11, 5, 0, 0, 4, -2, -1, 0, 7, 5, 4, 0, 0, 9, 0, -4, -4, 9, 0, 8, 7, 5, 6, 11, 1, 0, 5, -3, 10, 11, 11, 8, 4, 1, 4, 13, -3, -2, 5, -1, -1, -1, -5, 2, 1, 1, 1, -2, 1, 7, -4, -6, 3, 0, 11, 11, 4, 7, 12, 2, 0, 10, 5, 2, 1, 10, 9, 10, 8, 4, 6, 2, 0, 2, 0, -2, 8, -3, 6, -1, 4, 0, -6, 0, 10, 3, 12, 11, 13, 0, 13, 6, 8, 1, -1, -1, 11, 0, 2, 2, -4, 7, 9, 4, 4, 4, -3, 9, 1, 5, 2, 7, -1, 6, 5, 7, 6, 5, 8, -2, -3, 0, -3, 1, 6, 3, 0, -3, -5, 7, 2, -1, 9, 0, 10, 0, -2, -3, -4, 6, 6, -2, 7, 2, 2, 3, 1, 4, 10, 2, 9, 5, 8, -4, 0, 3, 5, -3, -5, 0, 0, -3, 10, 11, 7, -3, 7, -2, -4, -1, -3, 12, 9, 14, 1, 1, 10, 3, 10, 0, -5, 7, -1, 0, 7, -4, 0, 2, 2, -8, 0, -9, 9, 9, 11, 11, 3, 10, 11, 5, 13, 1, 3, 6, 9, 4, 4, 0, 9, 1, -3, 0, 1, -5, 3, -1, -3, -3, -6, -3, -1, 1, 1, 15, 14, 8, 15, 8, 4, 6, 3, 7, 12, 7, 0, 5, 1, 9, 1, 0, 4, 0, -6, -8, 6, -8, -4, 4, 1, 1, -11, -4, 0, 3, 2, 4, 14, 8, 5, 11, 4, 11, 9, 1, 6, 8, 2, -5, 6, 0, 1, -2, 6, 0, 4, -1, 3, -8, -7, -4, -12, -11, 9, 6, 6, 10, 10, 18, 11, 16, 4, 15, 5, 15, 13, 0, -4, -4, 6, 2, 4, -4, 4, 2, -12, 1, -9, -13, -8, 0, -5, -7, 13, 8, 19, 21, 17, 16, 19, 7, 16, 13, 13, 0, 9, 5, -4, 0, -9, 3, -11, 0, -8, 2, -9, -6, -10, -7, -7, -4, -1, -3, 2, 14, 11, 13, 9, 17, 9, 13, 13, 15, 2, 12, -1, 4, 4, -6, -10, 0, -7, 1, -9, -5, -7, -2, -11, -2, -5, 0, -14, -7, 8, 18, 8, 22, 14, 13, 17, 14, 8, 16, 5, 4, -4, 2, -2, 0, -8, -13, -10, -14, -12, -11, -17, -15, -15, -10, -14, -12, -9, -16, 9, 5, 10, 8, 24, 17, 8, 20, 5, 8, 11, 9, 9, 5, -5, 2, -8, -13, -7, -4, -12, -12, -7, -19, -17, -16, -5, -18, -7, -11, 12, 16, 20, 10, 20, 13, 9, 13, 14, 14, 1, -2, 2, 2, -8, -12, -11, -6, -4, -7, -10, -15, -15, -19, -5, -19, -12, -10, -16, -3, 8, 13, 16, 12, 11, 10, 7, 9, 11, 1, 13, 0, -4, 4, -6, -10, 0, 1, -8, -13, -13, -17, -16, -4, -20, -21, -8, -11, -16, -8, 11, 14, 18, 7, 9, 16, 17, 12, 7, 12, 3, 6, 2, -8, -5, -4, -4, -5, -13, -12, 0, -10, -12, -16, -13, -19, -5, -4, -16, -10, 14, 7, 6, 15, 17, 21, 20, 5, 3, 10, 10, 0, 8, -6, -8, -8, -6, -2, 1, -13, -7, -9, -16, -9, -9, -16, -19, -15, -18, -4, 13, 3, 16, 10, 12, 10, 6, 16, 7, 3, 6, -3, 6, 0, -9, 4, -3, -7, -9, -1, -2, -15, -12, -8, -18, -7, -18, -9, -11, -8, 12, 1, 6, 1, 12, 9, 11, 14, 4, 3, -3, 8, 2, 0, -4, 4, 4, 2, -8, -2, -11, -8, -11, -16, -9, -15, -9, -13, -7, -3, 0, 1, 1, 12, 9, 0, 0, 5, 1, 9, -1, 0, 7, 0, 0, -6, 4, 0, -9, -1, -3, -10, -8, -7, -4, -11, -3, 0, -2, -10, 3, 3, 5, -1, 7, 0, -2, 6, 2, 4, 9, 8, -2, 0, -5, 0, -7, -4, -11, -10, -14, -11, -2, -8, -6, -3, -13, -9, -3, 0, -1, 0, 6, 3, 4, -8, -9, -2, -7, -6, 4, 8, 6, 6, 4, -2, -10, -6, 1, -4, -9, -7, -3, 1, -6, -4, -9, 0, 0, 0, 4, 2, 3, -7, -2, -9, -5, -3, 5, -8, -5, -6, 6, -1, 8, 1, -1, -3, -9, -11, -3, -2, 2, -5, 0, 0, -1, 2, -10, -8, -6, 6, 4, 2, -3, -1, -1, -6, -10, -4, -1, -5, -3, -1, 4, -6, -5, -2, -1, -1, -10, 5, -3, 4, 1, -3, -6, -6, -7, -11, -1, -7, -10, -1, -2, -1, -11, -6, -12, -5, 1, -3, -6, -8, 6, 6, -8, 6, 4, -5, -9, 0, 0, 4, -7, -8, 5, 1, -8, -11, 0, 6, 1, -10, -3, -5, -9, 1, -2, -3, -2, 4, 0, 3, -1, 0, -6, 0, 3, 7, 3, 5, -6, 4, 3, 4, 0, -2, 2, 2, 3, 4, 5, -5, -10, -10, -7, -8, -6, -4, 4, -6, -5, -3, 7, 0, -1, 1, 5, 0, -1, -1, 6, -5, 7, -3, 0, 2, 0, -5, -5, 5, 0, -2, 0, 3, 5, 2, 0, 0, -6, 1, 3, 2, 6, 4, -7, 6, -3, 9, 5, 0, -4, 7, 0, 5, -1, 0, 0, 1,
    -- filter=0 channel=4
    0, 4, 7, 11, 0, 10, 0, 4, 1, 2, -6, -1, 4, 2, -7, -5, -13, -12, -3, -4, -7, -5, -3, -8, 2, -9, -7, 2, -8, -9, 14, 2, 6, 14, 12, -1, 3, 10, 1, 11, 1, 2, -2, -1, 3, -4, 0, -10, -2, -12, 2, -10, 1, -4, -3, 4, 0, -5, 2, -7, 4, 2, 1, 12, 3, 11, 0, 1, -3, -2, -4, -1, 0, -2, 4, 0, -5, -8, -3, -13, 2, -1, -8, -11, -5, 0, 5, -5, -9, -6, 13, 13, 1, 2, 12, 1, 13, 0, 10, 12, -3, 2, 2, -3, -2, 2, 2, 1, -2, -12, -7, -11, -10, -10, -8, -7, 2, 1, 3, -12, 13, 9, 8, 14, 6, 11, 1, 9, -2, 9, 7, 7, -4, 4, 0, -3, -4, 1, 0, 0, -7, -7, -2, 0, 0, 2, -4, 0, 1, -10, 14, 11, 9, -1, -2, 10, 6, -2, 7, -2, 2, 3, 3, -8, 3, 4, 3, -11, -8, -9, -10, -2, -2, -7, -3, 3, -1, 0, 0, -3, 12, 6, 5, 11, 11, 11, 10, -2, 4, -3, 5, 0, 6, 3, 0, 6, -8, -9, -7, 4, -1, 3, -7, -4, 0, 4, -1, 2, 5, 3, 0, 12, 7, 9, 4, -3, -3, 0, 7, -6, 7, 6, 0, 7, -2, -1, 0, 6, -6, -8, 0, -2, 3, 2, -5, 0, -7, -2, -6, 0, 6, 8, 12, 5, -3, -5, 7, 7, 0, -7, 5, -7, -2, 2, -5, 3, -2, -8, -9, 3, -8, -4, -8, -9, -8, 2, -9, 0, 1, -6, 2, 11, 0, 7, 7, 6, 5, -1, -6, 5, -5, 0, -5, -6, 6, 7, 6, 7, -7, -3, -10, 2, -2, 2, -2, -10, -10, 3, -9, -8, 10, 8, 10, 6, 6, 1, 7, 1, -2, 5, -5, 2, -4, 3, 9, -4, 0, -2, -2, -5, 3, 1, -3, -7, -4, -6, -2, -6, -4, 1, 1, 11, 10, 3, 0, 8, 3, 6, -6, -2, 1, 4, 0, 7, 1, 6, -4, 10, 10, 0, 2, -8, 3, -4, 0, -2, -10, 2, -5, -7, 0, 7, 1, 13, 10, 6, 7, 2, 5, -3, 2, -1, 4, 2, 6, 2, 6, 5, 7, 1, 6, 1, -2, -10, -9, -2, 5, 4, -1, 1, 11, 14, 9, 14, -1, 8, 4, -5, 6, 1, 7, 5, 0, -2, 3, 3, 2, 9, 6, 0, 13, 1, 0, 0, -1, -3, 2, 0, 4, -3, 3, 3, 14, 4, 5, -3, 1, 0, 6, -2, 6, 4, 2, 13, 6, 9, 6, 16, 19, 8, 10, 5, 0, 3, -9, -5, 3, -9, -7, -8, 9, 7, 1, 9, 0, 10, -3, 5, -3, 2, -2, 10, 0, 12, 8, 4, 8, 8, 17, 10, 15, 1, 8, 0, -10, 3, 0, 1, -1, -10, 12, 14, 0, 0, 10, 10, -1, 0, 0, 4, 7, -3, 7, 7, 3, 6, 8, 3, 5, 10, 15, 8, 3, -2, -10, -10, 6, 3, -4, 3, 6, 10, 13, 5, 11, 4, 0, 9, -4, 0, 8, 5, -4, 7, 12, 6, 12, 9, 2, -1, 0, 4, -4, 4, 2, 1, 0, 3, 5, -9, 7, 12, 9, 7, 6, 10, -3, 1, 6, -1, 4, 0, 10, 7, 0, 4, 11, 1, 9, 4, -6, 2, -7, -6, 3, -4, -4, -7, -3, -6, 0, 8, 8, 5, -1, -3, -4, 3, 5, 2, -6, 8, -2, -3, 1, 7, -1, 8, -5, -2, -3, -11, -5, -1, -1, -6, -9, -4, 0, -1, 5, 14, 0, 5, 7, 2, 4, -5, 6, -3, -2, 4, 9, 3, 4, -6, 6, -5, -5, 3, 4, 1, 0, 1, 0, -8, -1, -6, 0, -4, 0, 1, 4, 10, 9, -4, 3, 3, 1, 0, 2, 7, -2, 3, -5, -2, 1, 0, -4, -3, 3, -2, -5, -9, -9, 2, 0, 6, 8, -2, 5, 14, 12, 7, 11, 9, 9, 4, 2, 2, -3, -5, -6, 2, -5, -2, -8, 1, 1, -7, 0, -4, -2, -10, 0, -8, 4, 2, -3, -3, 3, 1, 15, 0, 11, 5, 5, 2, 4, 0, 4, 1, -6, 3, -6, -4, -2, -8, 3, 5, -8, 2, 0, -3, 2, -4, -3, 0, 0, -7, 0, 10, 15, 13, 3, -1, -1, 2, 2, 1, 6, 1, 5, 4, 1, 3, -2, -4, -10, -5, -1, -6, -1, 1, 2, -3, 5, 7, -4, -9, 14, 3, 5, 10, 11, 8, 0, 4, -3, -1, -2, 9, 0, 8, -4, 0, 4, -5, 1, -10, -5, 1, -6, -2, 6, -1, 1, -5, -3, 1, 14, 8, 11, 13, 15, 0, 15, 13, 2, 0, 0, 4, -2, -3, 6, 5, 6, -6, 0, 3, -2, 0, 1, -3, -1, -4, 1, -6, 6, -6, 6, 12, 3, 16, 0, 2, 6, 10, 3, 11, 7, 5, 0, 7, -8, -2, -4, 1, 3, -3, -10, -3, -5, 3, -1, 3, 8, 8, 4, -9, 2, 12, 0, 7, 4, 5, 6, 3, 7, 3, -6, 6, 5, -3, -9, -5, -9, -7, -10, -5, -2, -9, 4, 2, 1, 0, -3, 0, -7, -5, 3, -1, 5, 10, 1, 5, 6, -8, 1, -3, -10, 5, -10, -8, -12, -12, -1, -3, -11, -12, -11, -8, -2, -5, -11, -13, -9, -2, -12, -2,
    -- filter=0 channel=5
    12, 5, 6, 7, 7, 3, 4, -2, 1, 3, 7, 2, 9, 8, 8, -5, 6, -5, 2, -4, 1, 5, 0, 3, 6, 5, -6, 5, 8, 2, 14, 0, 11, 10, 14, 1, 7, 16, 4, 0, 13, 1, 1, 14, 13, 4, 4, 14, -1, 7, 3, 11, 8, -3, 4, 5, 9, 1, 8, -8, 0, 10, 9, 6, 5, 5, 20, 8, 12, 7, 6, 8, 15, 7, 8, 7, 7, 16, 5, 14, 12, 4, 0, -1, 7, 1, 8, -5, -1, -9, 1, 17, 16, 17, 20, 13, 12, 13, 8, 21, 18, 9, 19, 13, 6, 13, 3, 5, 17, 4, 7, 7, 10, 7, 3, 5, 8, 9, -8, -10, 7, 9, 22, 15, 8, 11, 20, 16, 18, 9, 21, 18, 13, 6, 13, 9, 5, 13, 4, 6, 13, 2, 2, -3, 3, 8, 7, 5, -4, -5, 0, 6, 7, 23, 21, 14, 14, 12, 17, 12, 11, 12, 4, 3, 0, 2, 1, 7, 7, 5, -7, -2, 7, 7, 9, -5, 4, 8, 4, -12, -4, 3, 21, 7, 16, 3, 11, 4, 6, 10, 4, 0, 0, -2, 5, 4, 0, -4, -1, 0, 3, 0, 3, -2, -3, 7, 0, 0, -8, -13, -2, 5, 13, 5, 8, 3, 0, 7, 5, 1, -2, 1, 13, -3, 3, 0, -2, -1, 0, -5, -7, -4, -3, -3, -8, 0, -5, 2, -7, -14, 0, 12, 12, -1, -3, -2, 0, -4, 8, 1, 5, 9, 0, -5, -9, -4, -1, -16, -16, -16, -13, -17, -6, -16, -5, 2, -6, 0, -14, -13, -7, 7, 6, -4, 0, -8, 0, -1, 4, -2, -4, 1, -4, 8, 6, 1, -4, -7, -10, -20, -10, -21, -18, -6, -11, -5, -6, -10, -2, -8, -1, 1, 9, 0, -11, 1, -13, -4, -6, -2, -2, -3, 0, -3, -2, -3, -2, -11, -10, -18, -10, -17, -13, -13, -14, 0, -6, -1, -10, -8, -7, 6, 6, -1, -10, -12, -6, 0, -7, 4, 3, 2, 0, -3, 1, -12, -10, -11, -14, -18, -24, -19, -22, -11, -10, -15, 0, -14, -17, -9, -9, 6, 5, 0, -14, -5, -6, -14, -6, -1, 0, -5, 1, 0, 2, -12, -12, -14, -18, -15, -15, -21, -21, -13, -14, -11, 3, -6, -9, -12, -1, -8, -6, -14, -18, -6, -11, -5, -13, -12, -10, 2, 5, -5, -12, -14, -15, -18, -12, -17, -10, -12, -20, -18, -18, -11, 2, -8, -15, -19, -6, 1, -11, -7, -3, -10, -15, -13, -13, 1, -2, 0, 2, -8, -5, -8, -8, -21, -23, -15, -19, -23, -23, -6, -8, -3, -3, -11, -16, -13, -12, 3, 5, -14, -8, -18, -5, -13, -3, -11, -5, -3, -1, -4, 1, -7, -8, -16, -17, -24, -22, -8, -11, -8, -9, -12, 0, 0, -1, -10, -3, -1, 2, -1, -5, -8, -11, -7, -11, -5, 4, 5, 8, -4, -12, -10, -13, -21, -8, -9, -21, -17, -14, -7, -16, -6, -8, -9, -13, -17, 2, 4, -3, -3, -13, -4, -8, 0, 3, 0, 7, 0, 0, -5, -7, -7, -12, -12, -8, -15, -11, -16, -20, -20, -3, -11, -5, -10, -2, -3, -12, 2, 4, -5, 0, -13, -11, -11, 4, 2, 0, 3, -4, -5, -7, -8, -12, -7, -11, -8, -11, -18, -19, -17, -4, -2, -8, 0, -18, -14, -10, 2, -6, 6, -4, -2, 1, 0, -9, -4, 1, 10, 6, -2, -4, -4, -10, -5, -10, -9, -13, -10, -21, -14, -14, -12, 1, 0, -17, -9, 1, -1, 0, 6, 0, -1, -7, 0, -4, -3, 3, -1, 12, -4, -1, 0, -10, -9, -11, -9, -3, -5, -11, -16, -1, -5, -8, -4, -1, -2, 7, 8, 1, 2, 8, 7, 8, 9, 8, 2, 7, 7, 11, 0, 4, -7, 1, -15, -13, -8, -5, -11, -3, -13, -8, -7, 0, 0, -2, -14, 4, 4, 11, 7, 8, 4, 10, 12, 6, 2, 7, 14, 6, -3, 2, -6, 3, 2, -5, -11, 1, 0, 0, 5, 1, -2, -2, -10, -15, -12, 1, 2, 20, 22, 7, 5, 3, 11, 1, 14, 9, 5, 6, 2, 13, 8, -6, 5, 6, -3, 4, -1, 6, -4, -2, 3, 6, -4, -9, 0, 8, 17, 23, 19, 20, 20, 15, 11, 16, 6, 8, 9, 10, 12, 4, 12, 10, 7, 0, -1, 3, -4, 5, 9, 3, 12, 0, -2, -11, -12, 8, 7, 9, 27, 10, 16, 18, 20, 12, 17, 17, 8, 18, 5, 13, 12, 14, 8, 12, 13, 15, 11, 12, 6, 13, 4, 6, -2, -1, -10, 3, 10, 10, 21, 9, 24, 7, 10, 7, 8, 20, 16, 12, 13, 12, 16, 5, 4, 10, 5, 13, 9, 14, 4, 15, 9, 10, -5, -5, 0, 14, 4, 8, 9, 14, 10, 9, 5, 13, 8, 3, 8, 21, 11, 19, 12, 12, 19, 6, 3, 7, 1, 2, 1, -1, 7, 4, 4, -5, 7, 4, 0, 4, 17, 4, 17, 3, 0, 5, 14, 3, 7, 4, 8, 4, 2, 10, 4, 12, 6, 2, -4, -2, 11, 8, 7, 0, 0, -7, -1, 9, 12, 14, 0, 6, 5, 8, 6, 10, 0, 1, 5, 3, -2, 9, -3, -2, -1, 3, -4, -3, -5, 6, 8, 4, 4, -6, -7, -5, 8,
    -- filter=0 channel=6
    -8, 0, -7, -10, -2, -6, -10, 0, 1, -1, 1, -12, 1, 0, -11, -10, 4, -9, -11, -11, 0, -12, -11, -12, -11, -14, -17, -9, -10, -17, -7, 6, 6, 1, 3, 3, -9, -8, 2, 0, -4, -1, -7, 4, 3, 0, 0, -2, 6, 1, -4, -7, 2, -3, -8, -9, -3, -10, 0, -11, -5, -4, 4, -5, -6, -2, 0, -5, -7, -2, -5, 2, 8, 2, 8, 11, 2, 0, 4, 2, 6, -8, 1, -6, 3, 0, -3, -4, -7, -5, 5, 3, 6, 10, 9, 7, 8, 4, 6, -2, 5, 12, 8, 6, 9, 3, 5, 5, 5, -4, -1, -8, 7, -5, 2, -10, 0, -4, -8, -5, 5, 11, 7, 1, -1, 4, -5, 0, -4, 2, 0, 10, 2, 3, 2, 8, 8, 0, 10, 1, 6, -4, -7, -6, 5, -3, 4, 0, -5, -1, 1, 11, 0, -2, 2, -5, -4, -2, 2, 0, 8, 11, 17, 10, 5, 11, 8, 1, 6, -5, -4, 1, -7, -6, -7, -4, -8, 4, -9, -8, 7, 10, 2, 1, 11, 11, -4, -3, 5, 1, 0, 11, 9, 3, 11, 18, 10, 10, 0, 0, 4, 7, -5, -6, -2, -4, -3, 5, 2, -10, 11, 1, 5, 2, 2, 4, 6, 8, 3, -1, 11, 10, 9, 2, 9, 6, 0, 1, -1, 0, 8, 1, 0, -8, 6, -7, 6, 0, 1, -3, -1, 4, 1, 14, 11, 4, -3, 8, 3, 0, 7, 10, 7, -2, 13, 9, 5, 13, 4, 2, 8, 2, -1, 6, 6, 4, 6, 5, -3, -5, 0, 8, 16, 2, -2, 0, 11, -1, 5, -3, 5, 8, 3, -3, -4, 7, 4, -5, 0, 3, 8, 9, 4, 0, -2, -5, -6, 5, -2, -3, 3, 8, 12, 0, 0, 10, 9, 1, -2, 3, 8, -1, -6, 3, -2, 1, 0, -1, 0, 0, 9, 3, -1, 2, 7, 7, -1, 1, -1, 2, 0, 3, 4, 3, 1, 4, 2, 1, 13, 1, -4, -1, 1, -9, -8, -17, -8, -3, 0, -6, 8, 5, 9, -2, 11, 7, 0, 6, -6, -2, 2, 8, 11, 15, 6, 3, 7, 7, 7, -2, 6, -2, -4, 0, -17, -18, -14, -17, -6, 2, 0, 3, 6, 13, 8, 3, 10, -2, 1, 4, 0, 7, 9, 12, 5, 15, 10, 8, 9, 9, -1, -1, -7, -4, -3, -11, -13, -12, -6, 2, 3, 2, 12, 3, -1, 1, 0, 3, -4, 4, 11, 9, 12, 12, 12, 13, 19, 17, 11, 3, 1, -3, -8, -12, -16, -20, -19, -20, -12, -7, 0, 0, 3, 11, 10, 6, 0, 7, -3, -3, -1, 9, 4, 0, 13, 5, 16, 12, 14, 0, 0, 0, -6, -8, -4, -9, -20, -14, -5, -1, -4, 7, 8, 2, 14, 3, 2, -4, 5, 6, 5, 10, 6, 11, 15, 15, 12, 13, 14, 2, 1, 3, -9, -1, -12, -12, -12, -11, -4, -13, 6, 2, 4, 11, 14, 5, 0, -3, 0, -2, 1, 0, 15, 1, 16, 4, 4, 9, 1, 13, 2, 0, 5, -13, -7, -23, -17, -13, -3, 3, -5, 12, 7, 12, 4, 9, -3, -4, -2, 1, -1, 3, 11, 0, 7, 4, 5, 7, 2, 5, -3, -8, -6, -11, -5, -6, -8, -6, 0, -5, -4, 3, 8, 7, 3, 8, 7, 8, 3, -1, 9, 2, 14, 13, 0, 4, 12, 11, 13, -3, -1, -2, 5, 3, -3, -1, 2, 1, -6, -4, 8, 11, 3, 8, 7, 0, -4, 0, 1, 0, 1, 1, 1, 6, 7, 7, 3, 8, 0, 7, 2, -2, 8, 0, 0, -3, -4, 0, 6, 10, 1, 5, 1, 3, 3, 10, 0, 3, 2, -9, 2, 7, 0, 12, 9, 9, 4, 9, 7, 0, 0, -1, 8, 11, 4, 2, 3, -2, 0, 6, 15, 1, 0, -3, 0, 0, 8, 3, 6, 3, 10, 5, 7, 13, 0, 5, 1, 5, 1, 0, 11, 7, 14, 16, 9, 15, 7, 9, 12, -1, 4, 4, -5, -1, 1, -7, 8, 7, 7, 0, -1, 5, 6, 10, 4, -3, -1, -4, 2, 1, 9, 15, 1, 8, 8, 5, 3, 7, -3, 0, 7, -5, 1, 1, -10, -9, 0, -7, -5, -12, 10, 0, 7, 4, 12, -5, 7, 0, -4, 11, 4, 5, 16, 13, 8, 17, 10, 3, 8, 7, -2, -2, 3, -10, 4, 3, -6, -2, -9, -6, 6, 5, 0, 2, 0, 6, 6, 4, 7, -1, 7, 7, 5, 6, 15, 1, 8, -2, -4, 5, -5, 4, 2, 3, 3, 3, -5, -2, -10, -2, 0, 10, -2, 6, 5, 8, -7, -5, 0, -4, 8, -1, 13, 0, 12, 13, 7, 10, 1, -3, -7, 3, 6, -3, -1, -12, 3, 2, 0, -9, -2, 0, 2, -5, 4, -1, 1, 1, -1, 5, -4, 4, -4, 0, 10, 0, 3, 0, 3, -5, 4, 1, -2, -1, -6, -6, -10, 2, -11, -11, -5, -6, 5, -8, 4, 2, 7, -3, 1, -6, -6, -6, 7, -3, 2, 3, 7, 4, 0, 3, -1, -3, -10, -3, -11, 0, -9, -8, -16, -18, -5, -9, -4, -1, -10, -6, 2, -12, -13, -12, -10, -5, 1, -7, -7, -1, -9, -6, 0, -8, -1, -12, -1, -5, -5, -6, -13, -10, -15, -25,
    -- filter=0 channel=7
    -15, -16, -3, -3, 0, 0, 5, -2, -6, -3, -2, 0, -1, 1, 5, -9, 6, 1, -3, 7, -2, -2, 10, 3, 7, 6, -5, -4, 7, 0, -12, -2, -10, -9, 1, -2, 0, -4, 8, -5, -1, -1, 3, -7, -7, -2, 0, 2, -1, -6, 1, -5, 5, 8, 3, 8, 7, 3, 8, -7, 0, -5, -7, -6, 4, 0, 6, 10, 1, 0, -1, 0, -2, 1, -2, -8, -10, 0, 6, 6, 5, 2, 1, 0, 7, -1, -2, 5, 1, 0, -7, -12, -1, 0, 1, 3, -4, 11, -1, 0, 1, 4, 1, -7, -8, 7, -3, 2, -5, -1, 2, -2, -6, -2, 5, 4, 2, -1, 14, -3, -13, -6, 1, 0, 10, 8, 7, 4, 7, 2, -2, 4, 1, 1, -6, -6, -6, -5, -5, -4, 6, -3, -7, -4, 7, -7, 6, 4, 12, 8, -4, 1, 3, 0, 8, 2, 11, 1, 2, 14, 1, 5, -3, 5, 0, 7, -5, 1, 1, -10, 0, -11, -5, -8, -7, 1, -6, 10, 6, 6, -14, -3, -2, 6, 0, 13, 8, 11, 9, 2, 11, 3, 3, 12, -3, -3, 6, -6, 1, -7, -3, -4, -4, 1, -6, -5, -8, 11, 12, -5, -10, -15, -5, 5, 7, 14, 1, 14, 8, 6, 16, 7, 8, 0, 10, 4, 7, -4, -8, -8, -9, -10, -9, -1, -9, -5, -6, 2, -1, -4, -6, -15, 0, -2, 1, 11, 14, 15, 13, 14, 8, 10, 10, 4, 7, -1, 2, 0, -3, -16, -11, -5, -7, 2, -2, 0, 7, 6, 12, 0, -5, -15, -8, -4, 4, 9, 10, 6, 11, 7, 11, 9, 4, 11, 16, 17, -1, 2, -2, -3, -14, -5, 0, -8, -6, 3, 3, 1, 6, -7, -15, -6, -3, -8, -9, 6, 3, -2, 0, 3, 4, 6, 4, 15, 7, 12, 2, 10, -3, 0, -4, -7, -6, -1, -4, 2, -7, -1, 0, -3, -4, -14, -13, -3, -12, -4, -2, 5, 11, 13, 2, 14, 8, 8, 21, 14, 21, -2, 0, -6, -12, -5, -15, -5, -9, -8, -7, -5, -1, 8, -9, -5, -2, -3, -6, -1, -11, -1, 0, 1, 11, 3, 18, 18, 9, 24, 12, -2, 2, -9, -4, -18, -14, -6, 4, -8, -3, -4, -2, 6, -3, -7, -11, -7, -14, -8, -11, 3, 5, 11, 13, 10, 6, 9, 21, 11, 16, -1, -10, -11, -9, -17, -5, -3, -11, 3, 7, -1, 6, 4, -9, -3, -15, -16, -11, -11, -4, -10, -4, 6, 6, 0, 16, 9, 24, 11, 17, -3, -1, -14, -11, -9, -5, -11, -12, -9, -6, 8, -1, -1, -3, -11, -12, -3, -15, -4, -17, 1, 5, -2, 3, 0, 13, 17, 22, 24, 14, -6, -14, -15, -13, -9, -4, -5, -12, 3, -9, 7, -3, 3, -5, -16, -17, -13, -9, -11, -10, -5, 6, 4, 9, 6, 12, 8, 11, 16, 15, 12, 1, -16, -13, -20, -11, -4, -10, -6, -7, -3, -1, 0, -12, -5, -2, -5, 0, -1, -3, -4, 0, 11, 10, 11, 4, 16, 9, 16, 23, 6, -9, -13, -15, -17, -5, 0, 2, 3, 1, -6, 4, 2, -4, -14, -1, -13, -5, 1, -1, -5, 0, 6, 16, 12, 16, 11, 10, 21, 17, 4, -7, -8, -8, -9, 0, 2, -1, -7, 3, 5, 7, 7, -3, -10, -13, -4, 0, -4, -5, 10, 11, 14, 12, 6, 17, 16, 21, 19, 14, 10, -9, -10, -2, -8, -6, 0, 4, -9, -9, 6, 8, 0, -16, -10, -8, -5, 0, 8, 4, 14, 7, 19, 6, 15, 18, 17, 5, 16, 4, 0, 2, -9, -7, -3, -2, -9, -11, -1, 0, -2, 4, 0, -10, -8, -3, -5, 5, 1, 2, 8, 7, 7, 16, 22, 13, 18, 6, 3, 11, -6, -6, -5, -1, -6, -7, -11, 2, -6, 0, 7, 0, -4, -3, -2, 0, -4, 2, 10, 17, 10, 6, 9, 6, 8, 4, 2, 15, -2, -4, 2, -8, -12, -9, -10, -5, -13, -9, -6, 0, -1, -3, 4, 0, -1, -9, -3, 12, 9, 6, 16, 16, 13, 15, 16, 7, 9, 4, 8, 6, 2, -1, -9, -5, -8, -1, -10, 0, -4, 2, 0, 5, 7, -5, -4, 5, -5, 7, 8, 15, 9, 10, 9, 10, -1, -2, -4, -5, 0, 1, -4, -4, 1, -1, 0, 2, -4, -5, 2, 6, -2, -1, -6, -4, -2, 4, 5, 0, -1, 0, 1, 8, 0, -3, -6, -3, 0, 2, 0, 5, 2, -1, -4, -6, 5, 3, 6, 0, 4, 2, 5, 11, 8, -15, -13, -1, 0, 8, 7, 14, 7, 6, 3, 6, -7, -8, -2, -2, -4, -5, -3, -8, -2, 0, 7, 10, -3, 10, 10, 6, 5, 3, 5, -14, -11, -5, -8, 1, 0, 0, 1, -2, 4, 0, 5, -4, 1, -7, 1, 3, 5, 7, -2, 0, -1, 3, 3, -2, 4, 2, 5, 7, -3, -16, -8, -9, -8, 2, 9, -3, 3, 5, -3, -3, 5, -7, 7, -2, 0, -8, 4, 1, 0, 8, 8, -2, 9, 6, 9, 6, 4, 7, 3, -23, -12, -8, -2, -5, 1, -3, 6, 4, 6, 0, 0, 0, -7, -7, -1, -2, 0, 2, 0, -4, -3, -3, 6, -4, -3, 6, 2, 4, -9,
    -- filter=0 channel=8
    3, 0, -1, -17, -16, -3, -7, -6, -15, -3, -4, 0, -2, -10, -6, -6, 1, -2, -5, 3, 0, 0, 3, 4, -1, 12, 7, 6, 12, 28, -9, 0, -10, -10, -21, -6, -6, -18, -4, -2, -14, -11, -14, -8, -9, -3, 0, 0, 0, 7, -3, 0, 1, 6, -8, -2, 6, 2, 16, 17, 1, -14, -8, -6, -21, -12, -9, -21, -5, -9, -15, -3, 0, -9, -1, 1, -12, -10, -3, -1, 1, 5, 4, -3, -1, -2, 8, 9, 1, 12, -2, -4, -2, -20, -12, -19, -21, -5, -15, -17, -9, -5, -3, -9, -4, 2, -10, -7, 0, 8, -7, -4, -3, -4, -5, 1, 3, 12, 6, 5, -7, -8, -8, -12, -23, -16, -8, -17, -14, -18, -15, -3, -16, -14, 0, -4, -5, 5, 6, -1, -4, -3, 0, 4, 7, 1, 8, 6, -1, 4, -2, -12, -8, -12, -11, -7, -19, -11, -19, -5, -17, -6, -10, -13, -2, -5, -6, 4, -1, 1, 5, 5, -2, -1, 3, -2, 0, 1, 7, 17, -6, -1, -16, -17, -13, -10, -13, -10, -16, -11, -16, -5, -7, -13, -10, 2, -2, 7, 11, 0, 10, 4, 11, 0, 0, 0, 5, 9, 15, 7, -13, 0, -3, -5, -9, -21, -15, -10, -17, -18, -11, -13, -7, -9, -10, 3, 4, 6, 10, 3, 12, 8, 12, 10, 12, 4, 0, 13, 4, 14, -10, -14, -9, -6, -13, -8, -19, -23, -16, -9, -11, -9, -11, -17, 0, -2, -3, 0, 0, 16, 5, 19, 5, 12, 0, 12, 3, 10, 2, 20, -11, -2, -18, -12, -9, -11, -9, -13, -16, -11, -12, -21, -6, -15, -6, 7, -1, 10, 7, 8, 12, 13, 15, 17, 2, 7, 11, 3, 4, 11, -7, -7, -4, -15, -6, -11, -18, -21, -23, -24, -12, -12, -10, -11, 3, -2, 1, 4, 4, 7, 15, 7, 12, 16, 4, 8, 14, 16, 13, 10, -4, -10, -10, -10, -10, -22, -13, -23, -18, -23, -13, -15, -12, -7, -1, 3, -6, 9, 5, 8, 12, 7, 11, 15, 3, 11, 12, 16, 11, 7, -12, -1, -10, -16, -22, -18, -19, -12, -22, -24, -14, -6, -8, -7, -1, -7, -5, 3, -2, 12, 6, 8, 13, 9, 16, 10, 5, 11, 9, 22, -3, -14, -7, -16, -6, -22, -17, -13, -12, -24, -16, -21, -16, 1, 4, 0, 0, 0, 2, 2, 9, 14, 4, 9, 8, 5, 7, 4, 18, 18, -11, -6, -9, -15, -8, -10, -20, -22, -23, -10, -15, -8, 0, -1, -2, 4, -2, -6, -3, 11, 4, 13, 13, 6, 9, 0, 3, 16, 12, 13, 2, -7, -5, -9, -6, -19, -21, -14, -11, -20, -19, -17, -14, -8, 6, 2, 3, 1, 3, 12, 13, 8, 19, 2, 17, 15, 9, 11, 18, 23, -5, -12, -7, -8, -22, -12, -16, -15, -27, -24, -22, -6, -9, 2, -7, -8, 8, -5, 7, -2, 8, 9, 14, 5, 10, 7, 12, 18, 8, 7, -12, -9, -19, -11, -19, -10, -20, -23, -12, -21, -19, -7, -12, -8, -6, 5, 6, 8, -4, 2, 15, 10, 18, 12, 2, 5, 2, 10, 16, 14, -3, -2, -10, -9, -9, -16, -25, -20, -20, -19, -24, -14, -14, -2, -3, -2, 0, 3, 2, 12, 3, 7, 17, 11, 11, 8, 7, 16, 13, 11, 2, -13, -6, -8, -17, -6, -23, -14, -17, -22, -13, -10, -13, -11, -7, -5, 2, 4, 0, 14, 6, 7, 16, 18, 4, 6, 5, 12, 8, 11, -6, -12, -3, -15, -8, -18, -20, -12, -22, -11, -18, -20, -5, -3, 2, 2, -2, 0, 11, 17, 8, 15, 21, 14, 3, 16, 3, 16, 19, 15, -2, -14, -7, -17, -6, -14, -20, -10, -13, -23, -18, -19, -18, -1, 2, 5, 4, 6, -1, 12, 9, 4, 11, 7, 4, 0, 15, 5, 13, 17, -14, -9, -15, -9, -18, -21, -6, -17, -6, -17, -9, -10, -12, -3, -5, 0, -8, -4, 10, 15, 2, 7, 11, 7, 8, 4, 12, 9, 15, 12, -1, -13, -21, -20, -20, -18, -8, -9, -18, -10, -4, -8, -9, -1, 1, -5, 6, 3, 3, 6, -1, 3, 2, 8, 9, 9, 12, 12, 3, 15, -4, -4, -12, -22, -12, -18, -17, -17, -12, -19, -9, -14, -8, -12, -8, -3, -4, 2, 5, 0, 2, -2, -3, 9, 0, 4, 0, 2, 1, 14, -3, -11, -19, -20, -20, -6, -13, -7, -18, -16, -2, -8, -16, -8, -1, -4, -1, 2, 0, -2, 6, -3, -5, -4, 1, 5, 0, -1, 1, 17, -9, -14, -15, -16, -5, -12, -11, -14, -6, -11, -13, -17, -7, -13, -5, -6, -2, -4, -4, -5, 5, -1, 6, 3, -4, -1, -2, 6, 11, 13, 0, 0, -9, -16, -13, -8, -9, -9, -7, -10, -2, -8, -8, -2, -2, -3, 1, -10, -7, 2, 0, 0, 0, 1, -3, 0, -2, 10, 4, 16, -2, -11, -9, -15, -11, -12, -4, -13, -3, -6, 0, -8, -9, -1, -1, 0, -10, -1, -6, 3, -7, 0, 6, -4, -6, 5, 4, 0, 15, 21, 9, -1, -6, -6, -12, -8, -10, -8, 0, -11, -8, -7, -4, 0, -4, 3, -8, 2, 6, 0, -7, 0, 6, 8, 11, 1, 17, 5, 7, 26,
    -- filter=0 channel=9
    -20, -6, -13, -5, -2, 0, 6, 0, -6, 4, 14, 12, 12, 23, 14, 18, 14, 13, 11, 5, 14, 13, 4, 6, 0, -2, 2, 0, -6, -17, -4, -11, -5, -5, -9, -1, -4, 3, 6, 7, 4, -3, 6, 16, 9, 8, 14, 4, 16, 17, 17, 12, 10, 11, 6, 1, 0, -11, -10, -12, -3, -10, -18, -11, -18, -2, -8, -4, -5, -2, -8, 8, 10, 1, 4, 9, 5, 15, 9, 9, 12, 0, 11, 8, 5, 0, 5, 4, -6, -5, -10, -13, -15, -19, -12, -8, -11, -18, -5, -5, 2, 0, -5, -3, -3, 6, 5, -1, 4, 1, 12, 10, 8, 0, 0, -2, -4, 3, -4, -4, -11, -20, -19, -13, -12, -9, -11, -6, -6, -1, -11, -9, 2, 3, 6, -2, 2, -2, 4, 15, 5, 14, 14, 14, 1, 0, 1, -5, -4, -2, -6, -10, -25, -17, -20, -9, -16, -4, -10, -4, -4, 3, 6, 0, -1, 7, 9, 6, 1, 16, 5, 17, 10, 13, 12, -3, -6, -4, -5, -9, -6, -17, -12, -8, -10, -10, -13, -1, -4, -6, -1, 2, 6, 7, -2, -1, -2, 8, 2, 11, 9, 9, 16, 9, 4, -2, -6, -5, -4, 0, 0, -10, -21, -11, -19, -12, -1, -3, -2, 3, 6, 0, -3, 5, 1, 1, -5, 6, 9, 0, 4, 14, 9, 4, 12, 10, -1, 0, 9, 4, -15, -13, -13, -13, -8, -8, -1, 0, 0, -2, -4, -1, -1, 2, -5, -9, -4, 2, -1, 2, 10, 7, 13, 15, 14, 9, 6, 2, 2, 7, -6, -18, -16, -17, -7, 2, -6, 4, -10, -4, 8, -3, 7, 2, -8, -9, -8, -4, 0, 7, 6, 16, 11, 14, 6, 12, -2, -2, -3, 6, -13, -13, -10, 0, 2, 6, 0, -4, -7, 6, -2, -3, 9, -9, -8, -8, 2, -7, 9, 2, 9, 11, 2, 18, 12, 4, 1, 3, -2, 5, 2, -4, -12, 1, 0, 1, 3, -1, -3, -2, 1, 8, 6, -10, -6, -13, -12, 4, 6, -1, 9, 15, 0, 16, 3, 10, 13, 10, 3, 5, -7, -9, -6, -1, 4, 9, 1, -5, 0, -4, 3, 0, 0, -10, -5, -11, -3, -1, 2, -4, 2, 4, 12, 1, 9, 1, 8, -2, -1, -8, -2, -16, 0, -5, 5, 5, -1, 9, -6, 8, 1, 2, -5, -4, -7, -17, -7, -14, -8, -5, 5, 12, 14, 10, 8, -1, 5, -1, 4, -7, -7, -17, -13, 1, -3, 4, 11, 10, 6, 5, 3, -6, 2, -12, -7, -23, -23, -4, 0, 5, 11, 12, 9, 6, 5, 0, 4, 7, 1, -9, -11, -16, -9, 4, 0, 2, 2, -1, 0, -4, 2, 7, -10, -8, -6, -25, -15, -6, 3, 4, 10, 0, 7, 13, 13, 10, 2, 4, 0, -6, -8, -18, -2, -2, 6, 11, 9, -1, 1, 10, 5, -4, 5, -5, -3, -20, -12, -7, -3, -2, 4, 0, 15, 3, 0, 6, 7, 1, -5, -4, 0, -15, -6, -5, 8, 9, 5, 8, -1, -4, -2, 4, 0, 0, -11, -12, -16, -3, 1, -3, 13, 9, 13, 1, 16, 3, 0, 3, 2, 5, 2, -17, -2, -8, -6, 2, 5, -2, 4, 4, -1, 1, -5, -1, -2, -14, -10, -6, 0, -3, 14, 13, 13, 11, 8, 6, 4, -4, -2, -1, -1, -12, -16, 0, -1, -6, -5, 6, -3, 5, 5, 5, -2, 3, 3, 0, -2, -5, -1, 2, 6, 7, 1, 17, 13, 0, 5, 8, 11, -3, -12, -10, -16, -3, -11, -5, 1, -7, 0, -1, -2, 1, 0, -7, -3, 4, 0, -7, 6, 11, 6, 12, 3, 8, 6, 5, 5, 2, 10, 0, -7, -10, -21, -10, 0, -9, -9, 0, 4, -7, -3, 3, -5, 5, 3, 2, -1, 4, 12, 2, 4, 18, 7, 12, 15, 3, 9, 2, 10, 0, -10, -20, -16, -21, -12, -7, -1, -1, -13, 4, -3, 5, 1, 4, 0, -4, 8, 10, 8, 3, 3, 10, 14, 12, 8, 14, 11, 9, 1, 2, -15, -15, -19, -14, -10, -10, -12, -4, -13, -2, -7, 4, 8, 9, 6, 0, -1, 14, 3, 16, 12, 11, 10, 3, 8, -1, 7, -1, 0, -1, -9, -17, -12, -14, -7, -11, -18, -6, -7, -1, -6, 7, -3, 3, -3, 2, 5, 8, 14, 13, 7, 7, 8, 0, 11, 3, -7, 1, 6, -8, -2, -9, -23, -15, -11, -19, -10, -16, -4, -10, -8, 6, 5, 2, 11, 5, 2, 8, 6, 10, 3, 16, 7, 8, 4, -5, -3, -6, 4, -12, -10, -14, -10, -23, -21, -15, -15, -14, -2, -5, 0, 2, -1, 0, -3, 0, 5, 12, 14, 14, 11, 4, 8, -2, -1, -2, 5, 2, -6, 2, -12, -12, -8, -8, -18, -7, -10, -8, 2, 2, -5, 10, 11, 5, 7, 8, 16, 16, 8, 9, 16, 3, 7, 3, -1, 5, 2, 5, -1, -3, -6, -7, -8, -11, -6, -4, -3, -9, 0, 9, 11, 9, 16, 7, 5, 8, 13, 11, 21, 21, 9, 4, 0, 8, 9, 2, -4, 3, -2, -2, -12, -6, -11, 0, -13, -9, -1, -5, 5, 6, 10, 9, 16, 11, 16, 11, 23, 12, 13, 17, 10, 12, 10, 0, 7, 0, -11, -4, -15, -10,

    -- ifmap
    -- channel=0
    517, 513, 519, 522, 520, 524, 525, 532, 531, 513, 504, 510, 529, 552, 559, 562, 548, 524, 502, 487, 478, 476, 480, 489, 494, 512, 529, 546, 553, 550, 537, 530, 535, 530, 523, 523, 526, 532, 523, 479, 469, 496, 522, 541, 540, 529, 521, 489, 453, 428, 425, 434, 446, 461, 468, 485, 510, 534, 545, 545, 534, 530, 540, 537, 528, 525, 530, 532, 513, 404, 393, 448, 489, 499, 500, 500, 485, 430, 377, 340, 336, 352, 389, 411, 432, 455, 478, 502, 525, 537, 504, 493, 510, 528, 531, 532, 539, 540, 521, 394, 373, 413, 462, 482, 475, 470, 449, 362, 294, 248, 248, 279, 316, 350, 397, 430, 446, 460, 494, 521, 483, 470, 473, 504, 530, 541, 544, 548, 536, 434, 423, 417, 435, 456, 445, 443, 398, 298, 226, 206, 225, 251, 274, 304, 364, 411, 430, 430, 467, 505, 453, 444, 438, 473, 524, 546, 543, 540, 535, 500, 461, 403, 395, 414, 386, 374, 350, 270, 196, 198, 248, 278, 278, 307, 362, 405, 422, 417, 445, 488, 412, 374, 367, 429, 506, 536, 522, 493, 496, 473, 403, 328, 319, 348, 336, 330, 330, 290, 219, 210, 265, 305, 315, 332, 359, 397, 432, 428, 430, 468, 305, 257, 266, 369, 479, 515, 442, 344, 334, 346, 293, 245, 258, 309, 322, 328, 346, 334, 253, 226, 253, 296, 334, 343, 355, 373, 425, 449, 435, 446, 195, 123, 171, 318, 448, 502, 351, 170, 140, 190, 181, 190, 231, 285, 325, 336, 372, 366, 249, 206, 210, 273, 324, 324, 333, 350, 401, 448, 442, 441, 124, 54, 98, 279, 423, 505, 351, 116, 28, 107, 130, 155, 213, 271, 313, 333, 399, 343, 184, 158, 164, 251, 310, 310, 306, 321, 363, 420, 430, 441, 97, 32, 69, 251, 401, 508, 428, 202, 96, 145, 144, 120, 181, 244, 297, 299, 391, 287, 118, 114, 146, 255, 307, 307, 301, 310, 329, 369, 392, 438, 95, 22, 86, 246, 379, 486, 520, 312, 209, 190, 161, 81, 127, 205, 258, 270, 358, 225, 83, 102, 165, 271, 313, 323, 311, 304, 297, 325, 349, 429, 83, 14, 108, 251, 358, 449, 536, 387, 289, 197, 137, 65, 100, 157, 204, 246, 333, 189, 83, 107, 175, 255, 302, 316, 310, 290, 269, 295, 337, 418, 54, 10, 111, 241, 311, 385, 491, 404, 314, 137, 47, 46, 105, 154, 199, 249, 318, 206, 116, 126, 188, 260, 307, 310, 295, 265, 257, 305, 361, 426, 26, 0, 66, 211, 244, 294, 390, 402, 310, 126, 42, 85, 159, 206, 233, 274, 325, 243, 194, 184, 200, 252, 314, 313, 286, 266, 282, 349, 404, 452, 0, 0, 5, 166, 201, 212, 269, 351, 306, 187, 120, 180, 236, 266, 286, 284, 296, 288, 317, 260, 235, 284, 345, 349, 321, 297, 321, 382, 422, 463, 0, 0, 0, 111, 176, 166, 179, 283, 285, 296, 247, 258, 293, 272, 294, 281, 258, 281, 351, 316, 297, 328, 381, 385, 371, 351, 378, 414, 449, 481, 0, 0, 0, 66, 175, 151, 152, 193, 227, 331, 299, 297, 277, 209, 245, 269, 232, 270, 319, 315, 345, 388, 415, 381, 375, 362, 402, 433, 467, 493, 0, 0, 0, 43, 162, 141, 105, 141, 210, 319, 290, 283, 198, 120, 165, 233, 250, 289, 307, 336, 379, 408, 408, 344, 340, 334, 392, 438, 461, 473, 3, 0, 0, 50, 168, 128, 26, 26, 121, 237, 211, 183, 83, 18, 61, 163, 221, 300, 342, 362, 360, 351, 326, 271, 251, 246, 286, 325, 340, 345, 0, 0, 0, 55, 160, 77, 0, 0, 0, 99, 125, 75, 7, 0, 18, 109, 184, 263, 314, 312, 280, 256, 213, 188, 165, 149, 156, 186, 193, 197, 0, 0, 0, 29, 111, 0, 0, 0, 0, 36, 73, 65, 47, 48, 62, 106, 141, 199, 217, 200, 169, 147, 123, 104, 86, 73, 66, 84, 89, 89, 0, 0, 0, 10, 43, 0, 0, 0, 0, 71, 106, 118, 121, 124, 128, 140, 141, 151, 143, 123, 107, 98, 82, 63, 51, 42, 40, 50, 50, 47, 0, 0, 0, 4, 0, 0, 0, 0, 66, 116, 127, 132, 135, 144, 143, 141, 138, 134, 120, 99, 85, 74, 56, 34, 30, 31, 32, 30, 15, 0, 24, 19, 3, 25, 0, 0, 0, 46, 112, 117, 103, 108, 115, 123, 129, 134, 131, 123, 107, 85, 62, 41, 28, 19, 21, 27, 12, 0, 0, 0, 15, 38, 42, 37, 0, 0, 0, 93, 122, 115, 91, 100, 115, 122, 124, 124, 116, 103, 84, 66, 44, 18, 6, 14, 27, 21, 0, 0, 0, 0, 5, 29, 48, 38, 0, 0, 0, 96, 118, 104, 81, 90, 101, 114, 120, 117, 101, 84, 67, 54, 36, 20, 19, 27, 28, 0, 0, 0, 0, 0, 4, 17, 32, 44, 0, 0, 49, 107, 131, 114, 84, 79, 81, 96, 104, 101, 87, 73, 59, 54, 50, 46, 43, 30, 5, 0, 0, 0, 36, 53, 7, 20, 28, 43, 51, 34, 110, 135, 151, 134, 112, 100, 90, 96, 96, 91, 72, 51, 43, 52, 61, 69, 57, 18, 0, 0, 0, 0, 61, 78, 17, 35, 45, 46, 74, 94, 126, 154, 165, 152, 143, 131, 128, 134, 123, 103, 73, 40, 31, 50, 69, 86, 60, 3, 0, 0, 0, 12, 59, 92, 
    
    
    others => 0);
end inmem_package;
