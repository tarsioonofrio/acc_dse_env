library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 2**16) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 21, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 31, 22, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 20, 25, 15, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 38, 10, 0, 0, 0, 0, 0, 20, 30, 9, 0, 0, 0, 0, 0, 5, 22, 0, 0, 0, 0, 0, 0, 0, 23, 57, 61, 36, 0, 0, 0, 0, 0, 33, 47, 9, 0, 0, 8, 0, 0, 35, 54, 0, 0, 0, 0, 0, 0, 0, 29, 66, 79, 50, 0, 0, 0, 0, 0, 64, 70, 15, 0, 0, 11, 7, 0, 52, 73, 18, 0, 0, 0, 0, 0, 0, 14, 64, 88, 60, 0, 0, 0, 0, 16, 105, 87, 15, 0, 0, 0, 9, 4, 67, 83, 36, 0, 0, 0, 0, 0, 0, 0, 66, 86, 56, 0, 0, 0, 0, 44, 116, 82, 5, 0, 0, 0, 0, 25, 76, 77, 26, 0, 0, 0, 0, 0, 0, 4, 76, 79, 43, 0, 0, 0, 0, 42, 101, 66, 0, 0, 0, 0, 0, 45, 88, 72, 14, 0, 0, 0, 0, 0, 0, 32, 72, 55, 21, 0, 0, 0, 0, 18, 74, 60, 0, 0, 0, 0, 0, 49, 95, 84, 23, 0, 0, 0, 0, 0, 0, 39, 39, 12, 0, 0, 0, 0, 0, 0, 45, 49, 0, 0, 0, 0, 0, 40, 101, 100, 42, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 34, 35, 0, 0, 0, 0, 0, 31, 99, 111, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 13, 0, 0, 0, 0, 0, 20, 88, 103, 56, 0, 0, 24, 16, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 70, 87, 39, 0, 0, 49, 72, 0, 0, 0, 0, 0, 32, 63, 57, 37, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 65, 12, 0, 0, 54, 104, 31, 0, 0, 0, 0, 60, 99, 86, 41, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 27, 0, 0, 0, 71, 146, 82, 0, 0, 0, 6, 68, 99, 78, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 116, 190, 138, 38, 0, 0, 14, 46, 67, 60, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 187, 214, 143, 49, 0, 0, 0, 4, 20, 29, 19, 4, 0, 0, 0, 0, 2, 8, 11, 13, 0, 0, 0, 0, 0, 112, 209, 176, 90, 30, 6, 0, 0, 0, 2, 10, 8, 3, 1, 2, 2, 4, 13, 17, 15, 12, 0, 0, 0, 0, 0, 164, 201, 119, 41, 23, 26, 29, 26, 20, 17, 15, 9, 2, 0, 2, 6, 13, 19, 15, 4, 0, 0, 0, 0, 0, 16, 157, 159, 81, 26, 27, 40, 44, 40, 30, 20, 13, 8, 3, 2, 6, 14, 22, 24, 12, 0, 1, 12, 0, 0, 0, 24, 117, 111, 52, 13, 17, 33, 42, 39, 27, 16, 10, 9, 10, 15, 21, 25, 26, 17, 0, 0, 28, 44, 0, 0, 0, 30, 79, 79, 37, 9, 12, 23, 31, 29, 19, 8, 6, 12, 22, 32, 36, 28, 11, 0, 0, 12, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 16, 67, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 3, 16, 1, 0, 1, 3, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 31, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 43, 72, 75, 36, 10, 0, 23, 50, 37, 10, 0, 2, 4, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 91, 107, 100, 83, 41, 9, 0, 16, 55, 59, 43, 35, 37, 36, 29, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 69, 123, 120, 73, 32, 8, 0, 0, 0, 14, 50, 69, 66, 54, 37, 16, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 28, 78, 63, 12, 0, 0, 0, 0, 0, 0, 39, 74, 70, 52, 25, 0, 0, 0, 0, 25, 17, 10, 16, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 6, 34, 48, 51, 26, 5, 0, 0, 0, 0, 32, 27, 20, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 28, 33, 29, 17, 0, 0, 0, 0, 0, 0, 24, 18, 16, 26, 1, 0, 0, 0, 0, 0, 23, 24, 23, 13, 14, 33, 33, 21, 12, 1, 0, 0, 0, 0, 0, 0, 28, 15, 16, 38, 12, 0, 0, 7, 43, 99, 135, 144, 134, 94, 42, 19, 12, 0, 0, 0, 0, 1, 1, 0, 0, 0, 74, 40, 32, 44, 45, 68, 100, 123, 130, 166, 195, 201, 182, 137, 82, 40, 21, 10, 16, 19, 23, 25, 27, 30, 26, 17, 148, 94, 60, 57, 87, 141, 176, 166, 146, 146, 155, 150, 136, 109, 78, 56, 43, 36, 36, 40, 44, 48, 52, 51, 50, 47, 192, 139, 99, 82, 122, 157, 164, 127, 98, 91, 88, 85, 81, 77, 69, 62, 55, 52, 52, 55, 58, 63, 66, 65, 62, 58, 175, 163, 146, 124, 139, 141, 120, 92, 78, 69, 65, 66, 67, 65, 61, 58, 57, 58, 60, 63, 68, 71, 71, 69, 69, 74, 136, 171, 198, 195, 174, 139, 96, 84, 73, 63, 58, 57, 58, 57, 56, 56, 58, 62, 68, 73, 77, 77, 76, 74, 79, 96, 109, 163, 227, 256, 216, 156, 105, 90, 81, 71, 64, 60, 58, 57, 58, 59, 61, 66, 75, 82, 85, 83, 78, 73, 77, 97, 88, 140, 205, 244, 213, 157, 119, 102, 96, 91, 85, 77, 69, 67, 65, 63, 63, 67, 76, 84, 88, 85, 77, 70, 71, 88, 146, 144, 140, 135, 130, 126, 125, 122, 105, 86, 73, 65, 63, 62, 73, 88, 101, 100, 97, 104, 119, 130, 135, 140, 148, 150, 144, 156, 152, 141, 133, 128, 120, 106, 77, 52, 44, 51, 62, 75, 92, 116, 123, 98, 70, 67, 81, 99, 116, 133, 156, 167, 162, 180, 169, 146, 133, 126, 118, 102, 79, 70, 64, 65, 70, 90, 114, 136, 134, 94, 54, 44, 53, 63, 79, 114, 158, 184, 199, 211, 179, 141, 123, 120, 116, 111, 102, 98, 84, 70, 70, 89, 114, 140, 142, 108, 68, 54, 56, 55, 67, 101, 149, 183, 219, 216, 170, 126, 109, 111, 110, 114, 115, 105, 68, 36, 38, 70, 107, 146, 162, 141, 99, 79, 73, 67, 72, 99, 132, 168, 191, 186, 142, 109, 108, 110, 98, 93, 95, 80, 42, 18, 27, 63, 109, 158, 191, 176, 119, 77, 69, 76, 77, 85, 109, 140, 142, 149, 115, 93, 101, 111, 94, 77, 72, 62, 30, 16, 28, 65, 108, 160, 206, 185, 104, 42, 41, 69, 77, 65, 81, 115, 115, 123, 107, 93, 102, 112, 101, 72, 71, 61, 34, 13, 21, 51, 101, 155, 204, 157, 59, 0, 13, 66, 84, 65, 64, 99, 102, 108, 107, 114, 125, 140, 148, 115, 106, 84, 36, 5, 3, 37, 83, 144, 180, 113, 15, 0, 12, 76, 99, 83, 72, 97, 81, 88, 106, 125, 140, 162, 185, 170, 153, 105, 27, 0, 0, 29, 65, 130, 158, 89, 0, 0, 36, 94, 116, 110, 100, 111, 39, 59, 108, 130, 127, 144, 176, 192, 169, 99, 12, 0, 3, 38, 72, 134, 155, 91, 6, 0, 37, 90, 122, 131, 129, 125, 0, 12, 85, 133, 120, 120, 147, 167, 140, 76, 7, 6, 35, 66, 97, 151, 161, 99, 27, 0, 32, 79, 128, 145, 145, 142, 0, 0, 28, 105, 113, 112, 133, 144, 117, 72, 43, 67, 87, 108, 142, 170, 156, 96, 42, 18, 37, 85, 143, 166, 165, 163, 0, 0, 0, 57, 102, 109, 125, 139, 126, 116, 117, 133, 132, 135, 159, 176, 155, 107, 65, 41, 62, 119, 178, 196, 197, 191, 0, 0, 0, 21, 78, 98, 128, 148, 163, 175, 169, 152, 132, 125, 140, 148, 135, 114, 89, 73, 102, 162, 203, 222, 219, 194, 0, 0, 0, 0, 64, 74, 89, 117, 161, 192, 182, 131, 84, 71, 90, 102, 90, 90, 79, 78, 113, 164, 197, 213, 197, 158, 0, 0, 0, 0, 59, 53, 31, 53, 114, 163, 150, 84, 5, 0, 22, 49, 51, 57, 60, 67, 86, 130, 161, 162, 141, 103, 0, 0, 0, 0, 62, 14, 0, 0, 27, 87, 88, 12, 0, 0, 0, 0, 27, 35, 35, 33, 33, 55, 74, 77, 66, 48, 0, 0, 0, 26, 57, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 32, 46, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 59, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 29, 40, 41, 33, 22, 15, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 28, 33, 42, 39, 31, 19, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 23, 36, 34, 29, 22, 6, 0, 0, 0, 0, 0, 0, 0, 0, 22, 2, 0, 0, 0, 0, 0, 3, 23, 34, 40, 38, 33, 24, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 21, 0, 0, 0, 21, 36, 58, 65, 58, 38, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 11, 0, 0, 20, 53, 83, 90, 80, 56, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 5, 34, 60, 59, 50, 35, 11, 0, 0, 0, 0, 0, 14, 30, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 18, 43, 40, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 22, 30, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 20, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 16, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 32, 38, 38, 41, 23, 0, 0, 0, 0, 0, 0, 6, 19, 13, 0, 0, 0, 0, 0, 0, 0, 0, 10, 18, 27, 34, 46, 57, 55, 42, 17, 0, 0, 0, 0, 0, 27, 45, 41, 20, 0, 0, 0, 0, 0, 0, 0, 22, 55, 54, 62, 73, 66, 50, 27, 0, 0, 0, 0, 0, 18, 53, 67, 62, 51, 29, 9, 0, 2, 0, 0, 0, 0, 46, 58, 48, 34, 18, 0, 0, 0, 0, 0, 0, 0, 45, 88, 89, 80, 65, 53, 39, 26, 30, 42, 0, 0, 0, 11, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 47, 71, 70, 59, 48, 38, 30, 29, 34, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 30, 48, 53, 44, 32, 32, 31, 31, 31, 30, 27, 21, 18, 21, 28, 0, 0, 0, 0, 0, 0, 0, 0, 40, 75, 88, 95, 92, 78, 56, 33, 22, 19, 20, 21, 22, 20, 14, 10, 12, 20, 0, 0, 0, 0, 0, 0, 0, 48, 63, 46, 35, 31, 28, 22, 17, 15, 16, 19, 20, 19, 16, 10, 3, 2, 10, 19, 0, 0, 0, 0, 0, 0, 0, 27, 21, 5, 0, 0, 2, 5, 10, 14, 18, 19, 16, 10, 1, 0, 0, 5, 15, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 11, 16, 17, 14, 6, 0, 0, 0, 4, 20, 24, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 13, 13, 9, 1, 0, 0, 2, 19, 31, 25, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 95, 151, 175, 149, 80, 16, 0, 0, 0, 0, 4, 31, 47, 38, 10, 36, 0, 0, 0, 0, 0, 0, 45, 95, 117, 126, 143, 163, 152, 96, 24, 0, 0, 0, 0, 0, 0, 4, 34, 46, 24, 57, 7, 0, 0, 0, 0, 15, 82, 136, 140, 109, 85, 72, 53, 17, 0, 0, 0, 0, 2, 8, 18, 30, 42, 45, 29, 0, 0, 0, 0, 0, 0, 0, 26, 48, 40, 11, 0, 0, 0, 0, 11, 20, 30, 32, 40, 51, 59, 55, 46, 36, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 56, 60, 51, 31, 26, 40, 45, 39, 21, 18, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 50, 61, 39, 24, 0, 0, 0, 1, 0, 0, 0, 9, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 22, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 85, 156, 182, 132, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 40, 32, 11, 0, 0, 0, 0, 0, 8, 42, 130, 215, 269, 220, 96, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 75, 78, 61, 30, 13, 0, 0, 0, 51, 49, 44, 93, 148, 178, 142, 61, 0, 0, 0, 0, 0, 0, 0, 0, 25, 78, 88, 70, 44, 20, 5, 0, 0, 0, 38, 31, 9, 21, 43, 47, 23, 0, 4, 56, 85, 60, 35, 18, 0, 19, 60, 93, 77, 48, 22, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 71, 155, 223, 236, 183, 118, 62, 40, 73, 114, 130, 97, 66, 43, 27, 17, 11, 0, 0, 0, 0, 0, 0, 0, 10, 122, 252, 348, 351, 298, 212, 128, 63, 59, 123, 185, 207, 179, 146, 116, 86, 61, 34, 0, 0, 0, 0, 0, 0, 0, 32, 181, 329, 387, 328, 212, 116, 53, 9, 28, 113, 206, 261, 262, 222, 164, 104, 54, 15, 0, 0, 0, 0, 0, 0, 0, 24, 138, 230, 235, 155, 64, 0, 0, 0, 10, 86, 183, 265, 285, 234, 142, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 58, 46, 0, 0, 0, 0, 0, 54, 135, 210, 252, 245, 174, 68, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 92, 193, 236, 211, 151, 68, 1, 0, 0, 0, 17, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 78, 79, 84, 114, 155, 165, 107, 40, 0, 0, 0, 0, 6, 43, 46, 0, 0, 0, 0, 0, 0, 0, 43, 122, 216, 294, 320, 278, 199, 118, 64, 28, 0, 0, 0, 0, 0, 0, 0, 1, 131, 39, 0, 0, 0, 21, 145, 223, 266, 299, 357, 414, 417, 343, 221, 92, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 225, 127, 13, 0, 24, 214, 374, 424, 357, 279, 251, 260, 247, 197, 119, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 241, 185, 73, 31, 141, 335, 426, 366, 222, 106, 68, 65, 60, 45, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 169, 165, 120, 128, 244, 344, 328, 206, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 71, 124, 173, 260, 359, 356, 256, 112, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 89, 218, 363, 453, 389, 247, 99, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 61, 187, 334, 416, 355, 223, 105, 53, 38, 28, 14, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 391, 403, 410, 411, 409, 397, 385, 368, 354, 339, 326, 315, 289, 246, 198, 159, 133, 102, 80, 70, 81, 109, 140, 179, 227, 279, 343, 381, 405, 414, 414, 404, 382, 348, 319, 281, 255, 231, 193, 146, 112, 86, 62, 36, 11, 0, 15, 45, 72, 104, 152, 218, 267, 338, 388, 410, 416, 409, 375, 318, 262, 224, 189, 153, 115, 83, 57, 28, 3, 0, 0, 0, 0, 0, 13, 33, 82, 153, 201, 295, 363, 399, 411, 399, 354, 290, 234, 190, 148, 109, 76, 45, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 96, 133, 241, 325, 367, 378, 354, 308, 251, 203, 162, 117, 68, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 70, 191, 275, 316, 310, 274, 225, 174, 138, 104, 64, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 5, 134, 231, 272, 241, 188, 133, 89, 57, 41, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 86, 199, 242, 182, 92, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 159, 224, 172, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 104, 205, 189, 80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 172, 209, 132, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 109, 182, 144, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 17, 113, 121, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 60, 0, 0, 0, 0, 18, 64, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 114, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 100, 174, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 133, 198, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 84, 135, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 134, 127, 125, 125, 124, 123, 131, 144, 130, 105, 104, 118, 119, 107, 102, 108, 106, 88, 60, 50, 62, 88, 120, 154, 170, 164, 177, 160, 140, 128, 123, 121, 133, 159, 169, 143, 110, 94, 87, 69, 67, 77, 89, 68, 34, 21, 35, 53, 77, 111, 150, 174, 207, 196, 159, 131, 123, 117, 116, 130, 148, 132, 85, 47, 32, 24, 35, 67, 93, 69, 28, 17, 32, 43, 50, 73, 113, 157, 164, 189, 164, 139, 128, 115, 90, 71, 78, 68, 32, 0, 0, 13, 43, 84, 111, 86, 30, 1, 11, 22, 22, 34, 68, 124, 101, 143, 142, 141, 140, 112, 54, 12, 21, 33, 15, 0, 0, 24, 49, 78, 115, 112, 52, 0, 0, 0, 0, 0, 29, 81, 82, 114, 117, 132, 157, 129, 36, 0, 0, 3, 2, 0, 0, 2, 23, 48, 88, 104, 51, 0, 0, 0, 0, 0, 0, 42, 98, 111, 90, 104, 165, 182, 105, 1, 0, 0, 0, 0, 0, 0, 0, 20, 62, 78, 25, 0, 0, 0, 9, 1, 0, 11, 118, 119, 66, 61, 119, 195, 201, 111, 38, 15, 0, 0, 0, 0, 0, 14, 66, 71, 8, 0, 0, 11, 39, 26, 1, 0, 121, 130, 72, 26, 23, 87, 151, 138, 92, 53, 0, 0, 0, 0, 0, 17, 81, 78, 0, 0, 0, 10, 46, 40, 17, 2, 82, 125, 97, 48, 0, 9, 68, 106, 99, 78, 14, 0, 0, 0, 0, 28, 86, 71, 0, 0, 0, 0, 37, 45, 34, 22, 3, 69, 94, 91, 38, 18, 67, 112, 107, 64, 28, 0, 0, 0, 1, 49, 87, 65, 0, 0, 0, 0, 33, 52, 51, 47, 0, 0, 52, 105, 84, 51, 88, 144, 131, 62, 22, 3, 17, 28, 30, 62, 85, 71, 0, 0, 0, 0, 45, 78, 89, 87, 0, 0, 0, 99, 111, 70, 88, 147, 147, 79, 20, 3, 27, 50, 55, 70, 83, 76, 20, 0, 0, 0, 45, 91, 113, 112, 0, 0, 0, 60, 124, 88, 62, 87, 106, 77, 29, 8, 16, 47, 71, 73, 70, 67, 35, 0, 0, 0, 24, 73, 105, 106, 0, 0, 0, 0, 110, 95, 24, 0, 17, 27, 8, 0, 0, 23, 72, 78, 51, 14, 0, 0, 0, 0, 17, 65, 98, 103, 0, 0, 0, 0, 42, 73, 0, 0, 0, 9, 32, 9, 0, 0, 35, 82, 57, 0, 0, 0, 0, 0, 41, 98, 127, 136, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 63, 22, 0, 0, 0, 26, 36, 0, 0, 0, 0, 0, 79, 152, 186, 189, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 106, 151, 150, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 100, 71, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 130, 102, 64, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 136, 107, 73, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 114, 93, 69, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 89, 79, 62, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 99, 85, 54, 39, 18, 25, 42, 40, 15, 0, 0, 29, 64, 71, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 127, 114, 75, 51, 57, 86, 132, 144, 120, 70, 31, 18, 17, 21, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 132, 141, 116, 81, 76, 115, 154, 146, 89, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 7, 3, 82, 110, 123, 106, 107, 115, 105, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 17, 26, 29, 33, 34, 49, 87, 106, 113, 99, 58, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 22, 34, 41, 43, 49, 39, 29, 59, 103, 114, 84, 37, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 26, 36, 43, 44, 46, 58, 58, 39, 46, 72, 83, 60, 30, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 23, 34, 38, 36, 32, 40, 65, 62, 55, 37, 15, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 23, 28, 27, 24, 28, 45, 75, 54, 54, 53, 55, 57, 61, 66, 67, 71, 67, 72, 72, 74, 77, 64, 41, 16, 3, 6, 3, 2, 3, 12, 24, 37, 40, 69, 58, 51, 52, 54, 57, 62, 78, 87, 76, 68, 61, 54, 43, 26, 13, 5, 15, 20, 14, 5, 1, 5, 14, 28, 34, 53, 41, 40, 46, 49, 48, 47, 55, 57, 45, 30, 16, 12, 4, 0, 1, 9, 18, 25, 19, 19, 15, 9, 11, 17, 26, 21, 17, 29, 41, 42, 42, 42, 39, 32, 13, 2, 5, 6, 4, 5, 19, 28, 21, 10, 7, 12, 13, 11, 0, 4, 14, 13, 15, 30, 41, 36, 32, 31, 28, 27, 15, 18, 24, 20, 17, 15, 25, 24, 17, 0, 0, 0, 0, 0, 0, 0, 5, 28, 31, 40, 47, 45, 35, 32, 36, 39, 40, 34, 26, 13, 9, 4, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 30, 44, 54, 68, 82, 78, 64, 51, 38, 31, 19, 4, 0, 0, 0, 0, 0, 4, 17, 11, 5, 0, 0, 0, 0, 19, 27, 41, 49, 71, 95, 96, 71, 57, 37, 23, 16, 1, 0, 0, 0, 1, 12, 28, 40, 27, 20, 12, 3, 0, 0, 7, 32, 48, 47, 48, 54, 57, 33, 19, 15, 14, 17, 9, 5, 0, 5, 17, 25, 33, 42, 21, 10, 8, 10, 4, 0, 0, 28, 46, 42, 32, 23, 13, 0, 0, 3, 33, 35, 26, 16, 6, 15, 17, 23, 28, 24, 0, 0, 0, 0, 2, 2, 0, 10, 19, 23, 19, 15, 2, 0, 0, 24, 60, 58, 48, 35, 19, 21, 16, 25, 24, 10, 0, 0, 0, 0, 7, 11, 0, 3, 2, 11, 19, 14, 19, 29, 46, 61, 78, 67, 47, 38, 20, 17, 18, 34, 27, 13, 0, 6, 13, 21, 23, 21, 12, 8, 5, 10, 23, 22, 35, 67, 89, 89, 74, 39, 19, 13, 3, 5, 24, 50, 40, 23, 11, 13, 23, 26, 23, 17, 23, 11, 12, 15, 19, 15, 22, 50, 65, 58, 17, 0, 0, 0, 0, 0, 18, 34, 38, 31, 22, 14, 14, 10, 7, 5, 25, 14, 3, 15, 16, 12, 12, 18, 8, 0, 0, 0, 0, 0, 4, 7, 8, 11, 16, 16, 10, 0, 0, 0, 0, 11, 21, 15, 0, 0, 12, 16, 9, 4, 0, 0, 0, 0, 13, 21, 23, 27, 36, 32, 20, 5, 0, 0, 0, 0, 7, 20, 13, 20, 0, 0, 0, 10, 14, 10, 0, 0, 3, 29, 38, 20, 16, 17, 36, 37, 20, 0, 0, 0, 0, 0, 10, 20, 8, 20, 3, 0, 0, 9, 18, 24, 24, 39, 62, 93, 97, 68, 34, 12, 1, 0, 0, 0, 0, 1, 13, 20, 25, 36, 21, 15, 0, 0, 15, 57, 76, 85, 91, 107, 117, 129, 127, 94, 61, 29, 9, 0, 0, 5, 17, 24, 33, 40, 49, 55, 46, 23, 0, 0, 51, 98, 130, 125, 103, 81, 69, 74, 69, 48, 28, 17, 10, 14, 16, 21, 22, 20, 19, 24, 31, 34, 48, 34, 16, 19, 61, 119, 146, 112, 50, 1, 0, 0, 0, 0, 0, 0, 0, 5, 8, 8, 8, 6, 3, 3, 7, 10, 17, 19, 13, 29, 71, 122, 110, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 49, 90, 100, 64, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 0, 2, 31, 80, 108, 84, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 9, 0, 0, 33, 80, 104, 69, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 0, 0, 7, 39, 55, 32, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 23, 60, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 84, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 97, 114, 88, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 91, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 11, 6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 26, 22, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 23, 25, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 26, 19, 27, 0, 0, 0, 0, 8, 51, 100, 138, 164, 132, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 144, 88, 48, 32, 11, 12, 85, 154, 173, 158, 147, 156, 162, 125, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 231, 187, 124, 65, 46, 97, 199, 228, 166, 84, 31, 11, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 217, 233, 182, 97, 64, 120, 187, 160, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 126, 191, 193, 119, 77, 105, 118, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 133, 190, 174, 141, 133, 97, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 15, 90, 170, 208, 214, 177, 109, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 3, 0, 39, 91, 130, 157, 134, 83, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 35, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 83, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 78, 88, 46, 0, 0, 0, 0, 0, 0, 0, 0, 18, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 32, 0, 0, 0, 0, 0, 0, 0, 0, 8, 40, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 37, 55, 55, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 29, 41, 56, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 31, 6, 0, 0, 0, 0, 0, 0, 0, 7, 36, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 73, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 107, 133, 121, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 137, 188, 179, 118, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 86, 162, 199, 170, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 108, 164, 183, 176, 141, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 83, 156, 187, 180, 147, 112, 66, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 45, 73, 102, 122, 128, 117, 98, 79, 58, 37, 19, 15, 26, 0, 0, 0, 0, 0, 0, 0, 0, 78, 136, 164, 187, 197, 185, 155, 126, 106, 94, 84, 73, 58, 42, 31, 25, 23, 27, 0, 0, 0, 0, 0, 0, 0, 116, 175, 180, 181, 184, 181, 163, 140, 117, 98, 84, 71, 56, 40, 27, 19, 16, 12, 6, 0, 0, 0, 0, 0, 0, 59, 142, 135, 111, 100, 103, 105, 103, 99, 94, 85, 73, 57, 41, 27, 20, 19, 12, 0, 0, 31, 0, 0, 0, 0, 0, 76, 107, 81, 63, 67, 77, 85, 87, 85, 81, 73, 62, 47, 33, 25, 24, 23, 13, 0, 0, 43, 0, 0, 0, 0, 0, 86, 92, 63, 51, 58, 70, 77, 77, 72, 65, 58, 52, 46, 40, 35, 30, 24, 5, 0, 0, 46, 30, 16, 14, 48, 96, 124, 105, 70, 56, 57, 65, 67, 61, 51, 43, 41, 44, 50, 53, 43, 24, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 38, 48, 41, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 39, 57, 75, 73, 56, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 24, 29, 36, 55, 65, 61, 48, 28, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 42, 44, 37, 20, 8, 6, 30, 46, 39, 23, 20, 15, 0, 0, 39, 4, 0, 0, 0, 0, 0, 0, 0, 0, 16, 39, 53, 45, 23, 0, 0, 0, 11, 42, 49, 43, 39, 37, 20, 0, 85, 44, 2, 0, 0, 0, 0, 14, 24, 16, 23, 43, 59, 50, 22, 4, 0, 0, 17, 50, 74, 75, 62, 54, 37, 7, 102, 70, 18, 0, 0, 0, 0, 0, 33, 29, 39, 56, 68, 59, 41, 37, 10, 5, 23, 55, 76, 79, 70, 60, 51, 30, 82, 75, 30, 0, 0, 0, 0, 0, 0, 14, 45, 71, 79, 71, 60, 52, 15, 2, 24, 45, 56, 56, 55, 54, 57, 52, 57, 46, 14, 0, 0, 0, 0, 0, 0, 0, 41, 82, 98, 81, 73, 57, 13, 0, 16, 41, 51, 46, 41, 47, 57, 65, 48, 26, 1, 0, 0, 0, 0, 0, 0, 0, 22, 62, 88, 89, 85, 57, 11, 0, 23, 55, 74, 67, 60, 59, 62, 73, 61, 58, 35, 0, 0, 0, 0, 0, 0, 0, 8, 25, 41, 52, 62, 41, 1, 0, 30, 62, 77, 74, 68, 64, 67, 73, 85, 105, 88, 46, 27, 14, 0, 0, 0, 0, 0, 0, 0, 5, 31, 24, 0, 0, 0, 36, 61, 60, 43, 38, 38, 40, 100, 123, 126, 86, 56, 42, 1, 0, 0, 0, 0, 0, 0, 0, 34, 23, 0, 0, 0, 0, 20, 19, 1, 0, 0, 13, 110, 121, 141, 110, 75, 62, 26, 0, 0, 0, 0, 0, 13, 29, 49, 30, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 111, 116, 136, 120, 81, 57, 43, 6, 0, 0, 0, 29, 38, 53, 52, 33, 15, 0, 0, 0, 0, 0, 6, 19, 8, 0, 101, 106, 124, 127, 84, 53, 42, 43, 24, 7, 22, 35, 46, 67, 56, 20, 0, 0, 0, 0, 0, 0, 15, 20, 6, 0, 92, 91, 105, 129, 92, 53, 63, 82, 58, 33, 21, 24, 51, 82, 80, 30, 0, 0, 0, 0, 0, 18, 22, 9, 0, 0, 89, 91, 108, 125, 90, 54, 79, 113, 109, 46, 0, 0, 0, 4, 43, 37, 9, 0, 4, 25, 44, 54, 50, 39, 18, 2, 64, 104, 135, 128, 61, 28, 63, 78, 50, 0, 0, 0, 0, 0, 0, 26, 54, 55, 52, 51, 50, 53, 63, 64, 59, 52, 0, 70, 131, 115, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 41, 51, 52, 49, 48, 49, 54, 61, 63, 63, 0, 9, 77, 77, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 28, 42, 45, 46, 48, 50, 50, 53, 58, 59, 60, 0, 0, 25, 27, 0, 0, 0, 0, 7, 34, 48, 50, 48, 45, 43, 46, 48, 47, 46, 50, 51, 52, 54, 56, 56, 54, 18, 0, 0, 0, 0, 5, 28, 27, 32, 43, 53, 56, 54, 51, 50, 49, 48, 46, 47, 49, 50, 51, 50, 50, 46, 45, 53, 20, 0, 0, 0, 0, 31, 38, 42, 50, 55, 57, 56, 53, 49, 47, 46, 46, 45, 45, 46, 46, 51, 51, 44, 38, 64, 32, 0, 0, 0, 0, 0, 23, 29, 40, 49, 56, 59, 55, 49, 46, 47, 47, 47, 47, 47, 52, 56, 52, 43, 38, 52, 46, 45, 48, 51, 50, 44, 35, 41, 57, 69, 57, 32, 17, 14, 22, 32, 43, 53, 67, 79, 75, 71, 74, 73, 66, 61, 53, 49, 49, 50, 43, 35, 22, 36, 53, 56, 42, 19, 0, 1, 9, 19, 23, 37, 68, 85, 81, 78, 81, 77, 72, 68, 59, 54, 55, 53, 50, 42, 26, 34, 39, 45, 41, 30, 19, 21, 26, 26, 23, 40, 70, 91, 84, 78, 80, 81, 74, 79, 76, 72, 70, 64, 59, 50, 31, 19, 22, 29, 29, 34, 42, 47, 44, 36, 28, 37, 58, 72, 67, 61, 66, 80, 80, 80, 86, 95, 92, 73, 54, 36, 17, 6, 7, 17, 33, 50, 58, 53, 51, 45, 36, 37, 53, 68, 59, 46, 56, 76, 85, 89, 95, 107, 100, 59, 25, 0, 0, 3, 16, 24, 45, 65, 70, 65, 60, 47, 31, 34, 49, 69, 64, 49, 53, 72, 85, 130, 126, 124, 90, 28, 0, 0, 0, 13, 25, 25, 42, 67, 68, 69, 65, 35, 16, 19, 51, 80, 74, 58, 53, 65, 82, 158, 147, 135, 73, 0, 0, 0, 0, 17, 26, 22, 39, 67, 63, 56, 50, 25, 5, 11, 50, 85, 83, 65, 54, 61, 75, 166, 158, 143, 80, 0, 0, 0, 0, 2, 19, 23, 46, 69, 60, 55, 41, 23, 11, 20, 56, 78, 77, 67, 53, 51, 60, 157, 159, 152, 91, 14, 0, 0, 0, 1, 15, 33, 61, 77, 65, 64, 49, 35, 23, 25, 58, 77, 81, 72, 57, 46, 52, 143, 154, 167, 115, 54, 5, 0, 0, 0, 3, 33, 62, 69, 61, 70, 54, 38, 23, 17, 54, 80, 86, 77, 67, 53, 58, 126, 148, 180, 145, 90, 45, 21, 3, 1, 3, 20, 45, 48, 42, 59, 53, 35, 16, 11, 34, 62, 75, 68, 63, 58, 70, 105, 139, 192, 177, 115, 68, 32, 0, 0, 0, 0, 8, 29, 41, 60, 52, 27, 6, 0, 13, 41, 56, 53, 56, 62, 73, 99, 122, 184, 193, 145, 98, 59, 14, 0, 0, 0, 1, 19, 46, 80, 77, 44, 5, 0, 0, 0, 16, 37, 49, 55, 69, 101, 110, 157, 191, 160, 120, 83, 48, 3, 0, 3, 20, 21, 52, 105, 107, 68, 18, 0, 0, 0, 5, 35, 50, 56, 69, 92, 97, 131, 164, 147, 106, 77, 70, 36, 11, 8, 3, 6, 49, 102, 114, 65, 6, 0, 0, 0, 17, 59, 76, 82, 95, 78, 86, 109, 136, 109, 62, 57, 74, 63, 34, 13, 3, 10, 59, 110, 111, 52, 0, 0, 0, 0, 43, 90, 110, 118, 122, 75, 82, 88, 95, 59, 0, 14, 72, 83, 50, 8, 0, 0, 48, 101, 107, 51, 0, 0, 0, 12, 54, 97, 127, 133, 119, 74, 81, 77, 70, 22, 0, 0, 56, 68, 35, 0, 0, 0, 0, 43, 64, 23, 0, 0, 0, 6, 33, 73, 104, 109, 93, 51, 62, 76, 68, 5, 0, 0, 40, 54, 31, 0, 0, 0, 0, 0, 15, 9, 0, 0, 0, 0, 9, 30, 58, 63, 51, 24, 41, 66, 69, 3, 0, 9, 20, 25, 12, 0, 0, 0, 0, 0, 0, 9, 6, 1, 0, 0, 4, 15, 29, 33, 28, 40, 38, 62, 58, 13, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 5, 5, 3, 3, 7, 11, 19, 27, 25, 19, 60, 52, 51, 38, 8, 0, 0, 0, 0, 0, 12, 16, 13, 9, 8, 9, 8, 4, 5, 8, 14, 20, 28, 29, 20, 12, 77, 69, 48, 8, 0, 0, 0, 11, 5, 15, 26, 31, 30, 22, 14, 8, 5, 4, 8, 16, 23, 28, 28, 22, 12, 11, 80, 81, 58, 0, 0, 0, 0, 16, 9, 15, 22, 29, 29, 21, 11, 5, 5, 8, 17, 27, 30, 26, 15, 6, 5, 21, 75, 84, 74, 0, 0, 0, 0, 3, 1, 4, 11, 20, 24, 19, 11, 4, 6, 14, 26, 35, 32, 18, 0, 0, 6, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 104, 76, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 143, 138, 123, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 161, 157, 168, 103, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 154, 154, 173, 139, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 127, 133, 156, 143, 64, 0, 0, 0, 0, 0, 0, 0, 6, 55, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 100, 105, 133, 128, 69, 33, 69, 93, 84, 46, 15, 19, 45, 85, 83, 6, 0, 0, 0, 11, 68, 105, 96, 45, 0, 0, 88, 92, 120, 116, 83, 83, 137, 175, 172, 115, 66, 35, 43, 78, 98, 72, 42, 45, 92, 140, 176, 203, 206, 175, 120, 82, 85, 99, 122, 115, 98, 119, 171, 205, 174, 105, 27, 0, 0, 21, 88, 138, 167, 190, 213, 231, 245, 259, 270, 263, 242, 223, 77, 98, 118, 109, 108, 119, 128, 111, 88, 68, 30, 0, 10, 63, 133, 192, 232, 250, 262, 276, 287, 297, 306, 310, 307, 304, 95, 93, 102, 102, 93, 86, 82, 78, 115, 151, 153, 144, 150, 174, 210, 243, 264, 277, 289, 302, 312, 321, 328, 331, 330, 331, 159, 125, 107, 87, 66, 84, 107, 150, 210, 249, 264, 262, 257, 258, 263, 271, 282, 295, 308, 320, 328, 335, 338, 338, 339, 345, 252, 198, 141, 72, 51, 102, 171, 228, 264, 280, 287, 287, 281, 276, 276, 283, 295, 309, 323, 331, 334, 335, 336, 341, 350, 361, 320, 264, 164, 51, 20, 100, 196, 257, 271, 275, 282, 286, 286, 282, 283, 291, 304, 319, 330, 333, 329, 325, 330, 345, 366, 377, 350, 299, 183, 48, 6, 82, 186, 247, 257, 264, 272, 277, 278, 277, 281, 291, 306, 322, 332, 329, 320, 315, 322, 347, 377, 384, 73, 80, 83, 81, 78, 75, 73, 76, 78, 73, 60, 35, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 37, 68, 82, 84, 82, 78, 65, 58, 55, 53, 50, 34, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 57, 76, 82, 82, 80, 63, 43, 22, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 57, 77, 87, 87, 71, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 48, 73, 92, 92, 78, 45, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66, 67, 79, 90, 88, 86, 72, 51, 39, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 106, 92, 81, 63, 61, 83, 96, 96, 84, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 120, 100, 73, 32, 10, 24, 50, 76, 84, 60, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 107, 89, 66, 8, 0, 0, 0, 1, 54, 57, 28, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 84, 71, 65, 12, 0, 0, 0, 0, 17, 34, 20, 11, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 56, 63, 28, 0, 0, 0, 0, 10, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 47, 67, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 50, 76, 58, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 57, 78, 71, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 47, 64, 72, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 42, 27, 43, 64, 55, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 23, 7, 20, 45, 52, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 25, 29, 19, 5, 11, 44, 63, 40, 23, 30, 22, 7, 18, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 19, 6, 28, 21, 20, 66, 91, 51, 30, 46, 33, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 44, 56, 101, 83, 19, 0, 4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 49, 88, 111, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 14, 84, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 15, 19, 20, 0, 0, 44, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 10, 14, 19, 24, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 10, 13, 17, 22, 21, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 8, 16, 19, 15, 22, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 14, 18, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 38, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 108, 133, 104, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 33, 4, 0, 0, 0, 0, 20, 69, 129, 184, 217, 228, 211, 158, 89, 39, 0, 0, 0, 0, 0, 0, 0, 0, 16, 67, 65, 30, 24, 56, 97, 141, 187, 230, 264, 288, 302, 309, 306, 285, 252, 228, 75, 6, 0, 0, 0, 0, 0, 0, 39, 113, 125, 112, 128, 170, 219, 266, 299, 319, 334, 345, 355, 362, 365, 362, 354, 349, 171, 101, 50, 0, 0, 0, 0, 7, 156, 227, 237, 234, 247, 274, 305, 332, 352, 365, 374, 380, 385, 389, 390, 390, 390, 391, 245, 203, 149, 49, 0, 0, 0, 154, 286, 327, 332, 331, 335, 342, 352, 362, 373, 384, 393, 399, 403, 404, 403, 404, 409, 413, 316, 289, 239, 115, 0, 0, 91, 272, 351, 358, 353, 352, 353, 356, 362, 371, 383, 396, 408, 415, 415, 412, 411, 419, 430, 433, 371, 341, 277, 157, 26, 60, 196, 327, 369, 365, 359, 357, 358, 361, 368, 377, 388, 402, 415, 422, 418, 413, 420, 435, 442, 435, 404, 363, 285, 181, 104, 147, 259, 346, 368, 368, 365, 364, 364, 366, 372, 379, 387, 398, 408, 414, 416, 420, 427, 435, 432, 411, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 24, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 5, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 4, 2, 7, 21, 21, 3, 0, 0, 0, 0, 0, 14, 17, 0, 0, 0, 0, 0, 54, 20, 1, 0, 0, 0, 0, 5, 34, 31, 33, 44, 37, 14, 0, 0, 0, 0, 0, 27, 36, 11, 0, 0, 0, 0, 72, 40, 10, 0, 0, 0, 0, 0, 40, 46, 48, 61, 50, 27, 17, 2, 0, 0, 1, 35, 43, 14, 0, 0, 0, 4, 72, 43, 6, 0, 0, 0, 0, 0, 28, 45, 50, 75, 66, 41, 33, 13, 0, 0, 3, 41, 42, 15, 0, 0, 0, 0, 64, 42, 7, 0, 0, 0, 0, 0, 9, 37, 50, 72, 69, 48, 44, 16, 0, 0, 0, 43, 41, 14, 0, 0, 0, 0, 64, 60, 21, 0, 0, 0, 0, 0, 0, 9, 30, 54, 46, 33, 32, 9, 0, 0, 0, 45, 47, 21, 0, 0, 0, 0, 85, 101, 63, 0, 0, 0, 0, 0, 0, 0, 0, 6, 5, 6, 13, 0, 0, 0, 0, 18, 32, 15, 0, 0, 0, 0, 106, 139, 121, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 113, 149, 156, 90, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 108, 134, 165, 125, 54, 17, 0, 0, 0, 0, 0, 0, 0, 10, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 98, 116, 151, 137, 76, 39, 23, 0, 0, 0, 0, 0, 17, 46, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 84, 100, 135, 133, 80, 53, 70, 73, 39, 1, 4, 14, 44, 85, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 76, 96, 131, 130, 72, 51, 109, 154, 122, 47, 0, 0, 0, 39, 50, 8, 0, 0, 0, 2, 16, 21, 22, 6, 0, 0, 51, 91, 132, 126, 68, 45, 97, 132, 91, 13, 0, 0, 0, 0, 23, 30, 9, 2, 15, 24, 30, 38, 43, 38, 22, 13, 14, 70, 120, 105, 38, 10, 46, 71, 44, 0, 0, 0, 0, 0, 0, 36, 42, 33, 30, 30, 32, 35, 45, 49, 44, 40, 0, 34, 83, 67, 4, 0, 0, 6, 3, 0, 0, 0, 0, 0, 0, 25, 35, 29, 27, 29, 29, 31, 36, 43, 45, 45, 0, 5, 40, 20, 0, 0, 0, 6, 5, 0, 0, 0, 0, 0, 0, 14, 22, 22, 24, 27, 31, 33, 37, 42, 42, 41, 0, 0, 0, 0, 0, 0, 11, 25, 10, 13, 20, 22, 20, 18, 20, 24, 24, 24, 26, 29, 31, 34, 38, 40, 39, 37, 19, 3, 0, 0, 0, 0, 30, 34, 19, 24, 34, 39, 38, 32, 27, 25, 25, 25, 26, 28, 28, 29, 33, 39, 36, 31, 46, 14, 0, 0, 0, 0, 17, 22, 7, 12, 23, 33, 36, 32, 27, 25, 25, 27, 28, 26, 24, 24, 28, 31, 32, 30, 52, 20, 0, 0, 0, 0, 0, 10, 0, 0, 4, 13, 19, 21, 21, 20, 25, 31, 32, 29, 26, 23, 20, 23, 31, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 0, 0, 0, 0, 0, 0, 3, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 30, 41, 54, 57, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 19, 33, 44, 57, 70, 80, 93, 102, 102, 91, 76, 71, 0, 0, 0, 0, 0, 0, 0, 1, 42, 49, 42, 44, 55, 65, 72, 76, 77, 85, 96, 105, 112, 116, 119, 119, 116, 115, 0, 0, 0, 0, 0, 0, 0, 64, 93, 96, 92, 89, 88, 87, 88, 90, 93, 101, 109, 116, 119, 120, 120, 124, 125, 128, 39, 0, 0, 0, 0, 0, 50, 101, 105, 100, 97, 95, 90, 88, 90, 94, 102, 110, 117, 121, 122, 123, 126, 128, 132, 133, 91, 30, 0, 0, 0, 0, 80, 108, 98, 91, 93, 93, 92, 91, 95, 102, 110, 117, 121, 122, 124, 126, 130, 135, 136, 130, 120, 71, 0, 0, 0, 13, 83, 101, 90, 89, 92, 95, 96, 97, 101, 108, 115, 119, 121, 120, 120, 122, 134, 147, 148, 139, 136, 101, 53, 0, 0, 31, 75, 86, 76, 81, 87, 92, 96, 96, 100, 107, 114, 118, 118, 117, 115, 118, 129, 146, 154, 149, 191, 190, 185, 181, 178, 175, 180, 188, 185, 183, 186, 197, 198, 181, 147, 103, 63, 29, 13, 18, 32, 55, 77, 103, 123, 128, 201, 190, 182, 182, 182, 176, 180, 189, 186, 176, 165, 157, 143, 120, 84, 43, 7, 0, 0, 0, 0, 3, 32, 65, 93, 109, 175, 174, 173, 179, 184, 177, 168, 162, 155, 129, 95, 76, 62, 47, 19, 0, 0, 0, 0, 0, 0, 0, 0, 26, 60, 87, 120, 135, 157, 175, 184, 178, 160, 141, 116, 79, 34, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 63, 74, 103, 133, 163, 177, 167, 142, 117, 88, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 51, 80, 111, 147, 178, 167, 128, 89, 64, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 21, 49, 82, 133, 189, 202, 154, 98, 64, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 30, 60, 108, 159, 187, 170, 123, 69, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 42, 69, 98, 125, 147, 141, 113, 70, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 47, 78, 97, 108, 111, 103, 71, 38, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 60, 76, 79, 74, 75, 55, 33, 27, 19, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 35, 48, 45, 33, 42, 54, 56, 56, 49, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 23, 7, 32, 60, 83, 86, 66, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 34, 71, 66, 35, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 8, 0, 0, 0, 0, 0, 0, 21, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 49, 74, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 34, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 48, 0, 0, 0, 0, 0, 0, 0, 0, 15, 48, 78, 87, 71, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 14, 40, 43, 37, 41, 53, 74, 86, 67, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 19, 4, 0, 29, 60, 80, 77, 44, 19, 17, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 32, 25, 28, 40, 71, 69, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 42, 47, 51, 53, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 46, 69, 68, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 73, 72, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 30, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 39, 27, 20, 22, 16, 0, 0, 0, 49, 153, 256, 340, 376, 308, 162, 10, 0, 0, 0, 0, 17, 47, 46, 24, 0, 65, 33, 24, 31, 42, 51, 62, 81, 124, 206, 281, 345, 373, 339, 203, 13, 0, 0, 0, 0, 0, 0, 0, 16, 7, 0, 63, 0, 0, 18, 39, 70, 130, 204, 251, 263, 251, 247, 219, 139, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 52, 119, 186, 184, 120, 61, 39, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 48, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 93, 135, 73, 59, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 161, 279, 283, 252, 160, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 104, 106, 0, 0, 0, 0, 0, 0, 0, 46, 150, 256, 281, 207, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 157, 114, 0, 0, 0, 0, 0, 0, 12, 41, 56, 126, 131, 16, 0, 0, 0, 0, 37, 13, 0, 0, 0, 0, 0, 16, 110, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 199, 258, 163, 39, 0, 0, 0, 0, 39, 91, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 293, 429, 383, 225, 57, 0, 0, 0, 49, 123, 155, 128, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 119, 333, 471, 430, 283, 110, 0, 0, 0, 21, 187, 265, 288, 247, 122, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 181, 326, 312, 161, 6, 0, 0, 0, 0, 40, 240, 356, 392, 304, 124, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 71, 105, 0, 0, 0, 0, 0, 0, 0, 96, 268, 370, 365, 230, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 105, 245, 336, 322, 243, 95, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 73, 162, 238, 290, 281, 193, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 110, 146, 114, 149, 271, 385, 394, 349, 271, 195, 113, 30, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 0, 0, 235, 481, 519, 506, 556, 658, 698, 603, 426, 231, 76, 0, 0, 0, 0, 0, 0, 0, 0, 15, 114, 0, 0, 0, 0, 229, 696, 839, 734, 596, 551, 569, 548, 439, 285, 133, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 248, 13, 0, 0, 18, 579, 902, 805, 531, 331, 262, 253, 231, 176, 108, 48, 8, 0, 0, 0, 0, 0, 0, 5, 2, 0, 264, 59, 0, 0, 240, 696, 782, 519, 226, 83, 52, 50, 43, 30, 16, 6, 0, 0, 0, 0, 0, 11, 29, 27, 5, 0, 202, 86, 0, 75, 426, 668, 565, 275, 68, 11, 16, 22, 18, 10, 2, 0, 0, 0, 0, 7, 25, 44, 54, 33, 6, 22, 134, 136, 190, 385, 613, 650, 441, 182, 39, 9, 14, 18, 15, 5, 0, 0, 0, 3, 21, 40, 53, 51, 30, 0, 2, 79, 98, 169, 332, 553, 682, 602, 382, 175, 68, 46, 43, 39, 25, 6, 0, 0, 0, 10, 35, 53, 46, 9, 0, 0, 4, 119, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 51, 66, 67, 54, 35, 8, 0, 0, 14, 30, 43, 45, 40, 26, 30, 19, 5, 0, 0, 0, 0, 11, 19, 24, 34, 56, 73, 80, 67, 45, 21, 0, 0, 0, 0, 0, 20, 36, 42, 37, 64, 37, 7, 0, 0, 0, 7, 26, 46, 53, 44, 35, 41, 45, 36, 26, 14, 0, 0, 0, 0, 0, 6, 20, 36, 37, 48, 27, 0, 0, 0, 0, 0, 5, 17, 23, 3, 0, 0, 15, 21, 20, 17, 0, 0, 0, 0, 0, 8, 17, 25, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 18, 27, 26, 9, 0, 0, 0, 0, 3, 5, 11, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 19, 22, 1, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 74, 67, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 68, 96, 69, 19, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 4, 3, 0, 0, 0, 0, 0, 0, 0, 7, 37, 72, 57, 16, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 6, 30, 26, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 15, 4, 0, 0, 15, 13, 2, 2, 2, 7, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 12, 40, 53, 57, 63, 60, 41, 21, 12, 7, 14, 26, 22, 0, 0, 10, 19, 17, 5, 0, 0, 0, 0, 0, 0, 0, 5, 49, 93, 107, 88, 53, 21, 6, 0, 0, 10, 44, 56, 39, 36, 33, 29, 22, 3, 0, 0, 0, 0, 0, 0, 0, 0, 9, 53, 72, 44, 0, 0, 0, 0, 0, 0, 36, 58, 59, 54, 40, 26, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 22, 1, 0, 0, 0, 0, 0, 8, 41, 64, 66, 58, 32, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 53, 66, 68, 59, 40, 28, 19, 8, 3, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 43, 55, 41, 25, 7, 13, 29, 33, 32, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 56, 66, 62, 45, 22, 9, 9, 8, 0, 0, 0, 0, 0, 7, 14, 19, 0, 0, 0, 0, 0, 0, 0, 0, 27, 84, 120, 134, 126, 99, 64, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 27, 0, 0, 0, 0, 0, 30, 66, 73, 76, 83, 78, 56, 31, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 73, 42, 0, 0, 0, 4, 37, 28, 9, 4, 8, 10, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 78, 66, 23, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 61, 74, 49, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 77, 79, 67, 32, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 60, 90, 95, 64, 26, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 19, 26, 29, 28, 22, 24, 30, 37, 3, 5, 3, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 12, 24, 41, 57, 67, 64, 57, 46, 35, 36, 17, 16, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 29, 41, 64, 86, 96, 97, 90, 67, 43, 34, 16, 28, 21, 11, 1, 0, 0, 0, 0, 0, 0, 0, 13, 26, 37, 41, 47, 58, 77, 96, 101, 94, 85, 74, 54, 35, 6, 28, 33, 24, 0, 0, 0, 0, 0, 0, 0, 30, 62, 75, 71, 59, 50, 51, 60, 72, 79, 71, 66, 72, 67, 47, 29, 42, 50, 31, 0, 0, 0, 0, 0, 0, 1, 45, 80, 91, 77, 52, 25, 19, 26, 43, 62, 65, 67, 77, 82, 64, 70, 80, 68, 27, 0, 0, 0, 0, 0, 0, 0, 31, 66, 79, 66, 39, 2, 0, 0, 23, 67, 83, 88, 88, 89, 77, 100, 96, 76, 24, 0, 0, 0, 0, 0, 0, 0, 15, 48, 58, 59, 36, 0, 0, 0, 28, 73, 97, 105, 99, 93, 84, 103, 99, 75, 19, 0, 0, 0, 0, 0, 0, 0, 4, 38, 51, 61, 41, 4, 0, 0, 35, 65, 86, 97, 98, 93, 88, 86, 91, 65, 22, 0, 0, 0, 0, 0, 0, 0, 2, 41, 57, 73, 56, 23, 0, 0, 30, 57, 77, 87, 93, 93, 91, 54, 72, 62, 42, 0, 0, 0, 0, 0, 0, 0, 0, 33, 63, 92, 73, 34, 5, 3, 34, 64, 86, 88, 90, 92, 102, 29, 60, 77, 63, 47, 2, 0, 0, 0, 0, 0, 0, 17, 53, 82, 64, 25, 0, 4, 42, 72, 85, 85, 86, 99, 120, 22, 63, 95, 94, 82, 48, 0, 0, 0, 0, 0, 0, 0, 30, 66, 57, 14, 0, 0, 22, 57, 67, 68, 77, 100, 112, 37, 65, 111, 114, 101, 81, 27, 0, 0, 0, 0, 0, 0, 26, 66, 65, 22, 0, 0, 0, 8, 22, 37, 55, 72, 83, 58, 70, 106, 122, 109, 91, 46, 0, 0, 0, 0, 0, 0, 37, 75, 71, 23, 0, 0, 0, 0, 0, 15, 42, 57, 64, 69, 70, 98, 109, 94, 71, 38, 0, 0, 0, 0, 0, 0, 29, 72, 65, 21, 0, 0, 0, 0, 0, 24, 50, 60, 64, 66, 66, 86, 86, 50, 7, 0, 0, 0, 0, 0, 0, 0, 12, 61, 61, 6, 0, 0, 0, 0, 4, 52, 73, 81, 76, 58, 61, 70, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 40, 0, 0, 0, 0, 0, 32, 73, 90, 90, 75, 40, 48, 53, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 2, 23, 48, 62, 53, 32, 2, 31, 48, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 10, 19, 17, 19, 25, 32, 25, 8, 0, 15, 61, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 37, 36, 33, 30, 26, 26, 29, 29, 24, 0, 0, 46, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 36, 43, 39, 34, 30, 28, 32, 35, 34, 25, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 22, 31, 35, 38, 43, 46, 45, 40, 34, 32, 29, 32, 38, 38, 27, 12, 0, 0, 0, 0, 0, 0, 0, 0, 21, 44, 59, 64, 63, 58, 52, 46, 40, 36, 35, 37, 39, 43, 41, 31, 15, 5, 21, 0, 0, 0, 0, 0, 0, 20, 38, 51, 57, 59, 59, 53, 45, 39, 37, 39, 43, 48, 52, 46, 31, 14, 3, 7, 40, 16, 0, 0, 0, 0, 0, 17, 34, 41, 46, 53, 56, 52, 43, 36, 37, 44, 53, 60, 57, 40, 17, 0, 0, 19, 197, 211, 210, 205, 203, 194, 174, 145, 125, 133, 152, 173, 181, 177, 142, 81, 12, 0, 0, 0, 0, 0, 4, 31, 64, 97, 158, 175, 192, 206, 211, 203, 179, 145, 127, 124, 129, 135, 130, 113, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 47, 93, 115, 156, 197, 212, 206, 188, 157, 128, 88, 72, 71, 66, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 53, 119, 180, 203, 198, 188, 161, 119, 62, 26, 14, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 79, 147, 167, 154, 151, 139, 99, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 107, 106, 73, 54, 49, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 79, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 73, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 74, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 106, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 85, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 131, 140, 149, 154, 155, 156, 159, 163, 174, 179, 157, 99, 33, 0, 0, 0, 10, 41, 58, 56, 36, 18, 8, 17, 46, 75, 111, 128, 143, 148, 147, 145, 139, 135, 132, 131, 101, 31, 0, 0, 0, 0, 33, 78, 105, 112, 93, 60, 29, 11, 14, 43, 59, 99, 133, 148, 147, 135, 111, 72, 40, 31, 29, 0, 0, 0, 0, 7, 51, 84, 114, 129, 111, 78, 45, 7, 0, 13, 38, 90, 138, 155, 152, 139, 112, 57, 20, 18, 41, 38, 19, 6, 10, 29, 48, 75, 107, 124, 94, 46, 16, 0, 0, 0, 105, 143, 171, 171, 159, 157, 148, 123, 107, 106, 121, 121, 96, 57, 23, 17, 26, 56, 93, 113, 75, 10, 0, 0, 0, 0, 193, 220, 217, 192, 170, 183, 213, 227, 225, 199, 176, 154, 116, 59, 3, 0, 0, 28, 94, 128, 101, 38, 0, 0, 6, 0, 249, 283, 263, 199, 156, 167, 216, 267, 285, 246, 205, 175, 125, 62, 2, 0, 2, 60, 130, 161, 141, 92, 35, 13, 20, 7, 268, 313, 283, 183, 106, 72, 116, 204, 280, 268, 229, 210, 157, 93, 41, 32, 48, 98, 140, 162, 141, 97, 49, 21, 21, 24, 245, 305, 279, 155, 25, 0, 0, 61, 201, 250, 247, 242, 202, 138, 92, 80, 69, 98, 116, 134, 105, 65, 35, 18, 17, 39, 203, 263, 248, 146, 23, 0, 0, 1, 144, 226, 250, 258, 232, 179, 126, 106, 76, 76, 79, 96, 68, 35, 14, 15, 28, 59, 153, 210, 210, 150, 65, 5, 0, 48, 154, 215, 221, 233, 212, 178, 140, 113, 75, 66, 75, 93, 74, 48, 28, 36, 60, 93, 124, 192, 215, 164, 118, 92, 84, 115, 148, 158, 150, 147, 127, 118, 118, 99, 66, 54, 62, 86, 78, 57, 39, 51, 77, 112, 111, 179, 238, 200, 173, 153, 126, 97, 62, 41, 35, 30, 23, 41, 83, 88, 53, 29, 22, 35, 41, 24, 14, 28, 66, 112, 101, 139, 217, 222, 193, 181, 134, 21, 0, 0, 0, 0, 0, 37, 91, 87, 33, 0, 0, 0, 0, 0, 0, 0, 44, 106, 94, 99, 159, 205, 190, 184, 134, 0, 0, 0, 0, 0, 59, 102, 133, 105, 34, 0, 0, 0, 0, 0, 0, 0, 73, 130, 100, 81, 113, 161, 158, 162, 154, 70, 0, 0, 28, 86, 127, 156, 172, 115, 45, 0, 0, 0, 0, 0, 0, 56, 116, 147, 110, 82, 92, 131, 117, 117, 144, 144, 105, 87, 118, 127, 124, 139, 148, 73, 0, 0, 0, 0, 0, 0, 0, 70, 112, 131, 106, 84, 95, 129, 106, 96, 121, 156, 142, 102, 77, 42, 21, 31, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 23, 69, 85, 115, 156, 118, 92, 74, 75, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 69, 145, 177, 122, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 126, 156, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 14, 8, 4, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 1, 13, 15, 10, 4, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 34, 13, 10, 14, 17, 16, 10, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 47, 19, 1, 1, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 36, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 20, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 8, 12, 11, 9, 22, 47, 37, 0, 0, 0, 0, 0, 0, 22, 124, 193, 195, 176, 164, 175, 186, 196, 199, 191, 162, 70, 58, 33, 10, 2, 12, 24, 8, 0, 0, 0, 0, 0, 29, 129, 234, 267, 226, 170, 158, 174, 190, 202, 220, 241, 227, 176, 154, 82, 24, 4, 0, 0, 0, 0, 0, 0, 18, 66, 141, 242, 316, 315, 221, 140, 133, 159, 173, 181, 223, 268, 278, 262, 224, 116, 41, 13, 0, 0, 0, 28, 58, 57, 68, 130, 215, 296, 346, 328, 222, 129, 114, 148, 165, 183, 231, 285, 301, 273, 226, 115, 59, 43, 5, 0, 0, 26, 70, 59, 69, 139, 225, 295, 344, 349, 262, 151, 106, 132, 173, 205, 237, 277, 303, 227, 169, 81, 74, 93, 42, 0, 0, 0, 10, 1, 22, 105, 193, 272, 343, 373, 299, 155, 72, 102, 181, 227, 238, 253, 281, 168, 95, 27, 48, 92, 47, 0, 0, 0, 0, 0, 0, 58, 150, 258, 354, 392, 289, 105, 6, 62, 179, 243, 241, 228, 251, 134, 45, 0, 0, 54, 55, 0, 0, 0, 0, 0, 0, 4, 106, 238, 360, 388, 227, 0, 0, 21, 178, 258, 253, 229, 235, 91, 0, 0, 0, 0, 39, 0, 0, 0, 0, 0, 0, 0, 71, 215, 346, 361, 149, 0, 0, 21, 197, 284, 289, 259, 247, 27, 0, 0, 0, 0, 53, 102, 114, 113, 27, 0, 0, 0, 32, 188, 329, 321, 92, 0, 0, 39, 215, 311, 327, 300, 272, 0, 0, 15, 47, 39, 109, 198, 235, 160, 0, 0, 0, 0, 15, 169, 312, 289, 81, 0, 0, 60, 228, 327, 345, 318, 287, 0, 0, 44, 126, 117, 166, 259, 262, 104, 0, 0, 0, 0, 57, 193, 301, 250, 75, 0, 0, 57, 211, 312, 333, 310, 285, 0, 0, 16, 158, 176, 192, 234, 202, 12, 0, 0, 0, 35, 149, 243, 285, 212, 80, 0, 0, 33, 179, 293, 333, 321, 289, 0, 0, 0, 134, 192, 180, 167, 126, 3, 0, 0, 46, 141, 227, 278, 264, 180, 85, 3, 0, 27, 175, 300, 348, 330, 277, 0, 0, 0, 81, 187, 155, 103, 73, 64, 103, 145, 162, 168, 217, 259, 230, 136, 53, 0, 0, 71, 215, 328, 360, 322, 241, 0, 0, 0, 25, 157, 116, 35, 42, 133, 230, 248, 182, 97, 103, 166, 151, 77, 10, 0, 25, 152, 292, 372, 372, 303, 195, 0, 0, 0, 5, 121, 41, 0, 0, 121, 250, 256, 126, 0, 0, 0, 40, 33, 17, 43, 107, 210, 323, 379, 361, 274, 176, 0, 0, 0, 33, 97, 0, 0, 0, 0, 112, 100, 0, 0, 0, 0, 0, 22, 74, 113, 153, 201, 258, 304, 290, 223, 157, 0, 0, 0, 62, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 77, 105, 116, 116, 125, 143, 142, 115, 87, 0, 0, 0, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 47, 31, 3, 0, 0, 0, 0, 0, 0, 0, 51, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 78, 154, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 133, 193, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 96, 120, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 11, 0, 0, 0, 0, 0, 0, 0, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 26, 3, 0, 0, 0, 0, 0, 0, 0, 19, 27, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 30, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 42, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 47, 52, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 10, 12, 23, 42, 49, 41, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 43, 81, 88, 73, 59, 53, 44, 32, 26, 15, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 60, 63, 54, 56, 77, 103, 122, 121, 103, 81, 59, 49, 48, 49, 46, 40, 36, 39, 45, 0, 0, 0, 0, 0, 0, 73, 133, 137, 105, 85, 92, 103, 103, 93, 79, 68, 61, 59, 58, 58, 59, 59, 58, 60, 64, 7, 0, 0, 0, 0, 31, 122, 164, 141, 107, 97, 99, 99, 94, 82, 70, 63, 62, 63, 63, 62, 62, 64, 67, 68, 69, 25, 0, 0, 0, 6, 104, 157, 146, 108, 84, 78, 77, 74, 70, 67, 65, 64, 64, 64, 64, 65, 68, 74, 74, 73, 71, 43, 0, 0, 0, 72, 153, 148, 107, 77, 67, 69, 67, 65, 64, 64, 64, 65, 66, 66, 68, 73, 79, 79, 74, 69, 66, 61, 5, 0, 11, 112, 168, 136, 93, 68, 70, 73, 72, 68, 64, 63, 63, 65, 67, 70, 73, 77, 78, 75, 67, 64, 77, 79, 41, 20, 62, 123, 150, 124, 87, 66, 67, 72, 76, 74, 68, 63, 61, 64, 69, 73, 74, 72, 67, 59, 57, 72, 100, 36, 39, 37, 35, 36, 34, 23, 15, 30, 47, 49, 29, 11, 9, 10, 6, 0, 5, 20, 24, 15, 5, 0, 0, 0, 10, 13, 29, 37, 38, 38, 32, 14, 0, 0, 15, 25, 15, 5, 7, 4, 0, 0, 0, 17, 25, 24, 16, 3, 0, 0, 0, 0, 11, 34, 42, 41, 35, 16, 0, 0, 2, 28, 36, 24, 11, 0, 0, 0, 0, 4, 16, 18, 14, 5, 0, 0, 0, 0, 10, 33, 43, 40, 42, 38, 25, 18, 32, 55, 60, 44, 20, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 26, 28, 42, 42, 34, 47, 74, 83, 66, 46, 45, 48, 35, 3, 0, 0, 0, 0, 0, 14, 14, 1, 0, 0, 0, 0, 36, 48, 57, 36, 5, 19, 66, 96, 73, 44, 42, 46, 33, 4, 0, 0, 0, 0, 0, 41, 42, 20, 6, 1, 0, 0, 36, 63, 74, 37, 0, 0, 13, 78, 79, 53, 53, 59, 47, 18, 0, 0, 0, 0, 8, 51, 54, 29, 5, 0, 2, 0, 13, 64, 87, 43, 0, 0, 0, 5, 47, 45, 58, 77, 70, 41, 12, 0, 0, 0, 17, 50, 48, 24, 0, 0, 0, 4, 0, 47, 93, 70, 0, 0, 0, 0, 0, 18, 51, 84, 85, 55, 22, 0, 0, 0, 7, 44, 36, 12, 0, 0, 0, 3, 0, 24, 75, 84, 32, 0, 0, 0, 0, 0, 32, 73, 89, 57, 20, 0, 0, 0, 6, 58, 47, 11, 0, 0, 0, 0, 0, 25, 58, 70, 55, 2, 0, 0, 0, 0, 16, 50, 65, 51, 17, 0, 0, 0, 12, 67, 56, 17, 0, 0, 0, 0, 9, 48, 65, 56, 55, 23, 0, 0, 0, 0, 5, 23, 23, 19, 1, 0, 0, 0, 4, 56, 50, 15, 0, 0, 0, 0, 29, 65, 68, 40, 38, 27, 0, 0, 0, 0, 0, 11, 5, 0, 0, 0, 0, 0, 0, 31, 33, 5, 0, 0, 0, 0, 31, 62, 59, 29, 15, 24, 0, 0, 0, 0, 0, 15, 6, 0, 0, 0, 0, 0, 0, 6, 16, 0, 0, 0, 0, 0, 24, 50, 52, 19, 0, 18, 17, 0, 0, 0, 1, 25, 26, 16, 1, 0, 0, 0, 0, 2, 13, 4, 0, 0, 0, 4, 15, 40, 53, 12, 0, 12, 44, 40, 10, 0, 0, 20, 38, 37, 18, 0, 10, 10, 10, 13, 8, 0, 0, 0, 0, 4, 8, 33, 48, 19, 0, 12, 65, 86, 49, 0, 0, 7, 50, 62, 32, 1, 0, 3, 17, 20, 13, 0, 0, 0, 0, 0, 3, 24, 32, 10, 0, 32, 95, 119, 74, 14, 0, 9, 50, 79, 67, 27, 0, 0, 15, 23, 10, 0, 0, 0, 0, 0, 0, 25, 24, 0, 0, 32, 114, 152, 100, 16, 0, 0, 0, 20, 53, 59, 48, 42, 39, 28, 16, 0, 0, 0, 0, 0, 0, 8, 9, 0, 0, 17, 70, 87, 41, 0, 0, 0, 0, 0, 19, 43, 41, 31, 22, 12, 6, 7, 5, 2, 9, 21, 0, 0, 0, 0, 0, 0, 34, 54, 26, 0, 0, 0, 0, 10, 15, 16, 9, 2, 1, 0, 0, 0, 1, 4, 6, 8, 0, 0, 0, 0, 0, 11, 75, 73, 55, 40, 31, 30, 30, 25, 16, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 109, 82, 43, 20, 14, 10, 6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 88, 107, 51, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 70, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 53, 57, 59, 64, 60, 54, 49, 41, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 82, 80, 76, 85, 103, 106, 98, 91, 80, 65, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 122, 129, 89, 67, 83, 107, 115, 117, 115, 107, 90, 52, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 96, 147, 170, 142, 85, 55, 68, 91, 98, 107, 122, 122, 109, 57, 44, 10, 0, 0, 0, 0, 0, 0, 0, 0, 21, 96, 147, 172, 173, 141, 85, 43, 45, 72, 95, 111, 126, 132, 122, 46, 33, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 84, 133, 154, 159, 129, 64, 11, 14, 58, 107, 132, 142, 142, 129, 36, 25, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 98, 139, 155, 118, 28, 0, 0, 35, 118, 159, 162, 148, 135, 29, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 125, 161, 110, 0, 0, 0, 6, 112, 167, 179, 163, 141, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 123, 170, 103, 0, 0, 0, 0, 107, 169, 192, 178, 153, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 115, 173, 92, 0, 0, 0, 0, 112, 180, 204, 193, 168, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 97, 164, 79, 0, 0, 0, 23, 134, 199, 211, 196, 182, 0, 0, 2, 53, 58, 50, 42, 0, 0, 0, 0, 0, 0, 0, 90, 137, 46, 0, 0, 0, 22, 121, 178, 190, 180, 180, 0, 0, 18, 98, 119, 118, 74, 0, 0, 0, 0, 0, 0, 4, 107, 123, 30, 0, 0, 0, 0, 73, 134, 161, 170, 170, 0, 0, 12, 103, 136, 131, 73, 0, 0, 0, 0, 0, 0, 62, 144, 132, 40, 0, 0, 0, 0, 8, 87, 135, 146, 129, 0, 0, 0, 77, 126, 105, 41, 0, 0, 0, 0, 0, 3, 79, 145, 128, 44, 0, 0, 0, 0, 0, 86, 135, 126, 89, 0, 0, 0, 48, 76, 46, 0, 0, 0, 0, 0, 0, 0, 18, 85, 79, 4, 0, 0, 0, 0, 37, 136, 165, 134, 80, 0, 0, 0, 27, 21, 0, 0, 0, 0, 28, 24, 0, 0, 0, 0, 10, 0, 0, 0, 0, 7, 116, 192, 199, 152, 98, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 83, 143, 186, 193, 158, 113, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 34, 68, 86, 98, 109, 116, 107, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 55, 67, 65, 53, 45, 46, 43, 35, 23, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 61, 52, 38, 25, 13, 6, 3, 0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 44, 47, 35, 20, 6, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 1, 15, 25, 35, 44, 46, 42, 33, 20, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 28, 35, 43, 46, 43, 36, 27, 19, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 26, 24, 28, 33, 35, 29, 20, 11, 8, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 18, 11, 14, 24, 30, 24, 12, 1, 0, 6, 12, 12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 59, 70, 74, 74, 74, 88, 102, 103, 78, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 35, 56, 68, 72, 71, 73, 83, 86, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 44, 60, 67, 61, 44, 31, 27, 6, 0, 0, 0, 0, 0, 0, 0, 4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 16, 43, 59, 67, 56, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 11, 0, 0, 0, 0, 0, 0, 0, 0, 13, 42, 62, 77, 68, 43, 16, 11, 16, 0, 0, 0, 0, 0, 0, 0, 7, 13, 0, 0, 0, 0, 0, 0, 0, 21, 54, 52, 62, 93, 112, 107, 89, 83, 86, 64, 11, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 88, 111, 72, 48, 85, 141, 168, 161, 147, 137, 103, 33, 0, 0, 0, 0, 0, 2, 34, 8, 0, 0, 0, 0, 0, 0, 120, 142, 82, 32, 47, 123, 183, 203, 193, 177, 133, 60, 0, 0, 0, 0, 0, 26, 52, 12, 0, 0, 0, 0, 0, 0, 121, 143, 71, 0, 0, 14, 86, 157, 191, 202, 163, 94, 20, 0, 0, 0, 0, 60, 57, 0, 0, 0, 0, 0, 0, 0, 92, 115, 58, 0, 0, 0, 0, 66, 156, 203, 183, 114, 46, 0, 0, 0, 20, 62, 31, 0, 0, 0, 0, 0, 0, 0, 37, 65, 43, 0, 0, 0, 0, 56, 135, 179, 178, 111, 50, 6, 0, 6, 31, 51, 11, 0, 0, 0, 0, 0, 0, 0, 4, 15, 12, 8, 0, 0, 9, 78, 140, 143, 107, 57, 27, 0, 0, 1, 21, 40, 9, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 7, 11, 0, 7, 52, 86, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 1, 30, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 43, 0, 0, 0, 28, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 56, 0, 0, 0, 5, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 67, 0, 0, 0, 0, 16, 0, 0, 0, 0, 15, 44, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 66, 14, 0, 0, 6, 17, 0, 0, 0, 0, 9, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 12, 0, 19, 69, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 23, 71, 103, 88, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 101, 106, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 94, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 79, 86, 80, 74, 72, 70, 51, 21, 0, 16, 59, 97, 125, 140, 118, 64, 0, 0, 0, 0, 0, 0, 0, 0, 7, 25, 68, 72, 74, 76, 81, 78, 64, 44, 28, 44, 74, 101, 117, 108, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 29, 48, 71, 83, 88, 91, 89, 68, 52, 47, 54, 51, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 58, 79, 86, 100, 97, 58, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 58, 56, 54, 44, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 80, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 78, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 19, 10, 5, 5, 2, 0, 0, 0, 1, 40, 78, 116, 130, 99, 38, 0, 0, 0, 0, 0, 0, 7, 21, 22, 5, 50, 30, 15, 10, 11, 13, 26, 49, 65, 76, 85, 100, 113, 108, 65, 0, 0, 0, 0, 0, 0, 0, 0, 5, 20, 14, 50, 16, 2, 5, 6, 11, 37, 79, 94, 77, 44, 30, 32, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 14, 0, 0, 0, 0, 0, 0, 7, 33, 36, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 83, 105, 92, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 130, 183, 199, 129, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 20, 0, 0, 0, 0, 0, 0, 0, 6, 48, 103, 149, 166, 89, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 56, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 92, 115, 78, 30, 0, 0, 0, 1, 24, 15, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 112, 189, 222, 191, 115, 44, 0, 0, 29, 72, 85, 66, 56, 36, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 102, 216, 264, 220, 136, 46, 0, 0, 0, 40, 108, 145, 152, 141, 101, 61, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 71, 165, 174, 93, 1, 0, 0, 0, 0, 7, 93, 159, 194, 172, 105, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 38, 0, 0, 0, 0, 0, 0, 34, 112, 162, 173, 122, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 88, 136, 137, 101, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 36, 63, 72, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 54, 112, 169, 206, 177, 107, 43, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 87, 190, 217, 230, 270, 318, 324, 262, 156, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 86, 0, 0, 0, 0, 99, 279, 334, 281, 220, 211, 224, 220, 177, 109, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 139, 54, 0, 0, 0, 204, 334, 292, 178, 101, 76, 78, 79, 65, 41, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 111, 65, 0, 0, 68, 220, 259, 179, 79, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 53, 50, 91, 184, 241, 193, 102, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 7, 46, 122, 222, 302, 287, 182, 80, 26, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 8, 0, 0, 0, 5, 1, 41, 135, 248, 318, 285, 179, 88, 48, 33, 27, 19, 7, 0, 0, 0, 0, 0, 0, 6, 9, 0, 0, 0, 0, 12, 52, 63, 68, 69, 71, 74, 66, 46, 39, 41, 57, 72, 81, 83, 70, 40, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 40, 57, 69, 76, 75, 63, 38, 27, 33, 55, 68, 65, 58, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 39, 68, 81, 84, 76, 59, 48, 53, 59, 53, 34, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 58, 82, 89, 90, 84, 72, 59, 39, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 75, 80, 86, 85, 59, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 48, 41, 47, 53, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 112, 166, 186, 157, 102, 57, 36, 38, 59, 84, 99, 96, 79, 51, 34, 16, 0, 0, 0, 0, 0, 8, 28, 52, 89, 145, 202, 227, 200, 132, 64, 20, 0, 0, 7, 38, 73, 100, 106, 82, 101, 53, 1, 0, 0, 0, 7, 68, 128, 157, 149, 154, 168, 168, 129, 84, 43, 22, 1, 0, 20, 45, 75, 108, 121, 101, 80, 29, 0, 0, 0, 0, 8, 69, 109, 106, 71, 56, 65, 77, 79, 77, 66, 50, 24, 29, 59, 96, 113, 116, 118, 107, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 49, 82, 105, 110, 94, 56, 47, 77, 120, 134, 112, 104, 105, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 64, 114, 142, 137, 97, 42, 14, 38, 78, 101, 89, 80, 97, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 61, 109, 124, 89, 39, 0, 0, 0, 37, 66, 75, 68, 77, 0, 0, 0, 0, 62, 110, 96, 22, 0, 0, 0, 0, 0, 23, 52, 60, 39, 2, 0, 0, 17, 55, 71, 79, 69, 58, 0, 0, 0, 27, 130, 209, 237, 161, 62, 0, 0, 0, 0, 0, 0, 16, 12, 0, 0, 29, 67, 92, 92, 89, 72, 48, 0, 0, 7, 57, 140, 211, 243, 183, 61, 0, 0, 0, 0, 0, 0, 2, 10, 15, 40, 66, 86, 99, 100, 88, 65, 39, 0, 0, 12, 42, 81, 132, 152, 95, 5, 0, 0, 0, 1, 5, 5, 23, 31, 46, 63, 62, 63, 72, 76, 66, 48, 23, 0, 0, 0, 0, 13, 41, 51, 28, 5, 13, 64, 114, 116, 91, 61, 56, 63, 87, 98, 78, 67, 73, 79, 71, 54, 30, 0, 0, 0, 0, 0, 0, 29, 76, 124, 186, 227, 241, 204, 155, 95, 80, 103, 144, 160, 133, 114, 123, 125, 110, 83, 51, 0, 0, 0, 0, 0, 0, 39, 154, 277, 350, 332, 266, 188, 121, 69, 78, 136, 212, 248, 235, 217, 204, 177, 142, 98, 40, 0, 0, 0, 0, 0, 0, 42, 165, 292, 328, 255, 151, 69, 22, 10, 46, 116, 212, 281, 315, 307, 250, 180, 112, 51, 0, 0, 0, 0, 0, 0, 0, 4, 72, 154, 164, 100, 26, 0, 0, 0, 41, 124, 220, 298, 337, 290, 196, 104, 41, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 72, 203, 287, 318, 287, 206, 122, 57, 23, 10, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 110, 232, 278, 244, 173, 104, 58, 31, 31, 40, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 92, 149, 185, 175, 157, 153, 169, 159, 122, 78, 47, 26, 17, 32, 57, 84, 29, 0, 0, 0, 0, 0, 0, 29, 120, 204, 292, 367, 386, 337, 252, 162, 97, 62, 45, 27, 17, 9, 5, 15, 32, 45, 140, 33, 0, 0, 0, 0, 152, 272, 314, 313, 328, 353, 350, 296, 209, 117, 60, 29, 19, 11, 4, 0, 0, 0, 0, 1, 203, 123, 1, 0, 0, 151, 302, 348, 290, 219, 188, 189, 184, 156, 114, 70, 41, 24, 16, 7, 0, 0, 0, 0, 0, 0, 179, 147, 64, 38, 101, 222, 288, 254, 161, 83, 54, 51, 53, 49, 41, 32, 25, 18, 10, 3, 0, 0, 0, 1, 0, 0, 105, 112, 113, 158, 222, 247, 228, 143, 67, 22, 10, 12, 18, 22, 23, 21, 16, 11, 7, 6, 6, 8, 11, 4, 0, 0, 42, 82, 165, 278, 348, 312, 218, 111, 53, 27, 19, 15, 14, 16, 16, 13, 8, 5, 7, 13, 21, 23, 12, 0, 0, 0, 19, 71, 186, 329, 407, 355, 231, 123, 74, 57, 46, 36, 26, 21, 16, 8, 2, 0, 6, 17, 25, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 84, 74, 47, 18, 0, 0, 10, 28, 45, 40, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 91, 138, 133, 94, 50, 9, 0, 0, 0, 10, 43, 70, 61, 12, 3, 0, 0, 0, 0, 0, 0, 0, 18, 31, 16, 41, 88, 118, 106, 82, 57, 14, 0, 0, 3, 35, 64, 103, 108, 65, 22, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 16, 55, 81, 95, 89, 44, 0, 0, 41, 88, 111, 127, 134, 101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 104, 137, 140, 99, 31, 10, 55, 108, 131, 126, 127, 119, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 144, 180, 173, 125, 31, 0, 6, 60, 91, 92, 91, 113, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 133, 161, 141, 83, 0, 0, 0, 14, 53, 64, 64, 85, 0, 0, 0, 0, 0, 102, 90, 0, 0, 0, 0, 0, 0, 0, 63, 96, 95, 36, 0, 0, 0, 39, 69, 66, 56, 57, 0, 0, 0, 0, 38, 213, 272, 162, 9, 0, 0, 0, 0, 0, 2, 45, 64, 18, 0, 0, 31, 91, 107, 84, 61, 40, 0, 0, 0, 0, 21, 177, 279, 206, 57, 0, 0, 0, 0, 0, 0, 24, 58, 32, 0, 9, 65, 110, 120, 94, 61, 31, 0, 0, 0, 0, 0, 57, 160, 128, 23, 0, 0, 0, 0, 0, 0, 37, 75, 58, 21, 13, 49, 82, 95, 79, 49, 11, 0, 0, 0, 0, 0, 0, 37, 77, 44, 13, 35, 69, 67, 53, 41, 70, 109, 104, 66, 33, 49, 87, 106, 90, 56, 9, 0, 0, 0, 0, 0, 0, 2, 116, 175, 189, 201, 212, 187, 141, 89, 87, 137, 164, 148, 113, 111, 148, 163, 134, 80, 18, 0, 0, 0, 0, 0, 0, 0, 169, 317, 363, 322, 254, 186, 130, 71, 62, 126, 208, 252, 241, 225, 236, 217, 164, 90, 0, 0, 0, 0, 0, 0, 0, 0, 150, 306, 345, 267, 159, 78, 44, 21, 29, 85, 193, 294, 335, 326, 285, 211, 124, 33, 0, 0, 0, 0, 0, 0, 0, 0, 46, 154, 187, 121, 34, 0, 0, 0, 41, 106, 208, 311, 362, 330, 246, 139, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 47, 16, 0, 0, 0, 0, 75, 201, 298, 345, 334, 267, 187, 111, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 12, 0, 0, 0, 111, 252, 321, 303, 242, 168, 128, 101, 75, 53, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 159, 200, 197, 169, 148, 160, 213, 226, 184, 126, 89, 76, 79, 90, 101, 114, 32, 0, 0, 0, 0, 0, 0, 0, 72, 224, 349, 419, 434, 377, 278, 185, 130, 98, 77, 59, 47, 43, 44, 56, 75, 89, 191, 52, 0, 0, 0, 0, 99, 210, 287, 346, 398, 428, 418, 354, 252, 150, 87, 56, 44, 33, 24, 15, 9, 7, 10, 10, 281, 190, 51, 0, 0, 113, 251, 315, 293, 254, 236, 233, 220, 186, 139, 92, 61, 44, 33, 22, 11, 1, 0, 0, 0, 0, 258, 250, 170, 97, 89, 176, 238, 230, 159, 91, 61, 60, 65, 63, 57, 49, 41, 34, 25, 12, 1, 0, 0, 0, 0, 0, 159, 223, 245, 243, 223, 213, 173, 121, 66, 24, 9, 12, 23, 30, 33, 33, 28, 22, 15, 6, 0, 0, 0, 0, 0, 0, 66, 160, 275, 359, 380, 294, 178, 102, 59, 30, 16, 10, 16, 23, 25, 22, 16, 10, 7, 9, 11, 9, 4, 0, 0, 0, 14, 110, 251, 398, 453, 368, 232, 139, 95, 69, 50, 34, 26, 23, 20, 13, 4, 0, 0, 9, 17, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 23, 23, 19, 9, 0, 0, 2, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 38, 48, 57, 58, 46, 27, 11, 3, 11, 0, 13, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 23, 43, 51, 57, 63, 64, 55, 39, 24, 12, 14, 19, 33, 27, 14, 4, 0, 0, 0, 0, 0, 0, 0, 2, 20, 34, 36, 43, 51, 65, 71, 65, 51, 40, 34, 29, 19, 47, 54, 46, 28, 15, 4, 0, 0, 0, 0, 16, 31, 39, 48, 45, 37, 44, 57, 69, 67, 55, 45, 44, 44, 41, 28, 88, 84, 66, 32, 6, 0, 0, 0, 0, 4, 25, 43, 55, 55, 49, 39, 46, 52, 60, 60, 52, 47, 48, 53, 49, 40, 123, 111, 82, 21, 0, 0, 0, 0, 0, 15, 35, 52, 58, 53, 47, 45, 54, 46, 42, 45, 50, 56, 60, 64, 58, 48, 145, 128, 90, 6, 0, 0, 0, 0, 5, 38, 50, 62, 59, 59, 53, 59, 59, 38, 22, 25, 39, 54, 64, 64, 64, 55, 142, 116, 79, 0, 0, 0, 0, 0, 19, 51, 60, 70, 64, 64, 67, 71, 66, 39, 18, 24, 41, 58, 65, 66, 70, 69, 119, 95, 74, 25, 0, 0, 0, 0, 27, 41, 43, 54, 61, 62, 73, 79, 70, 36, 17, 30, 46, 58, 68, 73, 79, 79, 103, 86, 80, 60, 0, 0, 0, 0, 28, 10, 4, 16, 34, 48, 73, 82, 67, 32, 22, 37, 51, 63, 72, 77, 76, 82, 102, 99, 97, 85, 51, 13, 0, 0, 0, 0, 0, 0, 3, 36, 71, 72, 38, 6, 3, 29, 47, 57, 59, 62, 66, 82, 109, 118, 123, 107, 92, 58, 13, 0, 0, 0, 0, 0, 0, 33, 69, 63, 10, 0, 0, 0, 8, 23, 28, 45, 67, 91, 124, 130, 137, 125, 114, 85, 27, 0, 0, 0, 0, 0, 17, 47, 76, 66, 7, 0, 0, 0, 0, 0, 12, 46, 65, 79, 133, 136, 141, 132, 127, 103, 44, 0, 0, 0, 0, 24, 34, 53, 75, 65, 6, 0, 0, 0, 0, 0, 25, 56, 64, 63, 134, 132, 141, 136, 128, 114, 71, 16, 0, 2, 29, 44, 45, 56, 66, 47, 0, 0, 0, 0, 0, 3, 54, 74, 70, 60, 127, 124, 132, 139, 128, 99, 73, 50, 43, 47, 53, 44, 39, 57, 50, 24, 0, 0, 0, 0, 0, 40, 73, 89, 75, 54, 118, 123, 133, 139, 124, 78, 51, 54, 37, 13, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 21, 42, 66, 75, 65, 38, 91, 113, 135, 146, 121, 45, 8, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 22, 40, 52, 63, 57, 46, 28, 51, 96, 136, 151, 86, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 23, 29, 43, 55, 59, 63, 69, 68, 59, 48, 9, 74, 142, 148, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 55, 65, 67, 70, 72, 77, 82, 86, 84, 82, 0, 52, 128, 120, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 51, 69, 77, 78, 80, 82, 84, 87, 93, 94, 95, 8, 39, 81, 42, 0, 0, 0, 0, 9, 36, 50, 55, 59, 64, 71, 78, 80, 81, 81, 84, 85, 86, 89, 94, 97, 92, 50, 45, 29, 0, 0, 0, 0, 25, 58, 78, 85, 88, 88, 85, 82, 82, 81, 81, 83, 85, 87, 88, 93, 99, 96, 84, 85, 57, 0, 0, 0, 0, 0, 45, 60, 75, 83, 87, 87, 85, 83, 81, 82, 85, 88, 90, 91, 94, 97, 97, 90, 79, 99, 72, 0, 0, 0, 0, 0, 44, 53, 57, 61, 68, 75, 80, 82, 82, 85, 89, 93, 96, 97, 99, 97, 93, 85, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 8, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 14, 32, 37, 35, 33, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 15, 30, 42, 47, 48, 51, 45, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 15, 14, 17, 27, 39, 43, 43, 37, 40, 40, 30, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 36, 36, 26, 21, 18, 11, 20, 34, 29, 23, 29, 30, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 28, 42, 38, 20, 3, 0, 0, 0, 26, 35, 31, 34, 38, 34, 12, 3, 0, 0, 0, 0, 0, 0, 0, 17, 12, 15, 27, 40, 41, 13, 0, 0, 0, 0, 31, 44, 42, 44, 48, 43, 26, 2, 4, 9, 0, 0, 0, 0, 0, 18, 22, 23, 27, 39, 42, 19, 1, 0, 0, 23, 50, 49, 42, 44, 52, 49, 31, 0, 4, 17, 6, 0, 0, 0, 0, 0, 0, 11, 30, 44, 43, 27, 16, 3, 8, 38, 50, 42, 32, 28, 40, 43, 30, 4, 0, 8, 10, 0, 0, 0, 0, 0, 0, 0, 30, 53, 50, 37, 29, 15, 13, 43, 53, 45, 27, 20, 25, 28, 25, 11, 5, 8, 3, 0, 0, 0, 0, 0, 0, 0, 19, 45, 50, 46, 30, 11, 10, 38, 55, 49, 33, 24, 24, 26, 25, 24, 23, 22, 7, 10, 0, 0, 0, 0, 12, 15, 16, 26, 28, 32, 25, 6, 5, 28, 47, 47, 29, 24, 30, 28, 27, 33, 50, 36, 21, 16, 14, 4, 0, 0, 2, 15, 16, 6, 0, 15, 24, 8, 0, 13, 36, 38, 23, 17, 17, 14, 6, 42, 62, 51, 29, 22, 29, 28, 0, 0, 0, 0, 0, 0, 0, 6, 22, 6, 0, 0, 2, 9, 6, 2, 0, 0, 0, 48, 63, 63, 42, 20, 23, 44, 15, 0, 0, 0, 0, 0, 0, 11, 17, 19, 8, 0, 0, 0, 0, 0, 0, 0, 0, 47, 62, 69, 47, 9, 11, 16, 10, 0, 0, 0, 0, 2, 12, 18, 22, 30, 28, 3, 0, 0, 0, 0, 9, 5, 3, 43, 60, 60, 42, 0, 0, 0, 0, 0, 0, 0, 0, 6, 34, 42, 31, 7, 0, 0, 0, 0, 0, 0, 1, 15, 16, 42, 51, 40, 17, 0, 0, 0, 9, 0, 0, 0, 0, 25, 60, 69, 48, 11, 0, 0, 9, 14, 8, 0, 1, 5, 7, 33, 45, 34, 3, 0, 0, 22, 59, 51, 24, 0, 0, 1, 23, 42, 52, 43, 30, 33, 40, 41, 38, 35, 29, 30, 30, 6, 34, 38, 1, 0, 0, 47, 65, 47, 16, 0, 0, 0, 0, 9, 37, 57, 59, 57, 55, 53, 52, 53, 54, 55, 55, 0, 0, 18, 4, 5, 22, 35, 25, 13, 1, 0, 0, 0, 0, 21, 40, 54, 59, 58, 55, 53, 53, 57, 61, 61, 58, 0, 0, 0, 0, 24, 39, 30, 17, 25, 33, 42, 45, 48, 51, 55, 58, 59, 57, 55, 54, 56, 59, 63, 64, 60, 53, 0, 0, 0, 0, 31, 50, 46, 37, 48, 59, 66, 67, 64, 63, 61, 60, 59, 58, 58, 60, 65, 71, 69, 60, 52, 52, 23, 0, 0, 0, 23, 60, 68, 55, 55, 62, 67, 68, 65, 62, 61, 60, 61, 62, 64, 68, 73, 72, 62, 53, 52, 60, 54, 14, 0, 0, 0, 38, 61, 56, 53, 59, 65, 67, 65, 62, 59, 58, 61, 66, 70, 70, 67, 60, 53, 53, 63, 69, 30, 36, 38, 38, 38, 33, 22, 13, 15, 28, 43, 64, 80, 84, 64, 20, 0, 0, 0, 0, 0, 0, 5, 20, 16, 11, 42, 41, 40, 41, 42, 41, 46, 52, 69, 74, 73, 76, 79, 71, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 49, 39, 36, 36, 38, 40, 49, 67, 87, 77, 52, 33, 22, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 11, 17, 25, 28, 29, 31, 39, 37, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 28, 54, 91, 104, 89, 36, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 22, 44, 72, 122, 148, 126, 60, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 29, 44, 44, 57, 74, 88, 71, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 10, 0, 0, 0, 0, 0, 0, 0, 11, 27, 21, 25, 16, 3, 0, 0, 0, 17, 20, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 74, 88, 55, 12, 0, 0, 6, 15, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 89, 126, 137, 120, 72, 27, 1, 0, 29, 47, 36, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 71, 152, 167, 134, 70, 19, 0, 0, 0, 30, 71, 76, 54, 28, 22, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 96, 87, 43, 0, 0, 0, 0, 0, 0, 36, 71, 70, 48, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 50, 50, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 52, 36, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 53, 85, 87, 59, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 50, 66, 105, 148, 169, 155, 106, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 0, 0, 0, 72, 131, 119, 86, 72, 72, 71, 52, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 25, 0, 0, 39, 110, 119, 63, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 25, 7, 2, 50, 77, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 36, 52, 64, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 71, 112, 105, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 108, 107, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 23, 26, 31, 36, 33, 32, 30, 43, 54, 44, 24, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 14, 22, 30, 33, 29, 17, 6, 23, 44, 41, 7, 0, 0, 0, 0, 0, 0, 0, 12, 2, 0, 0, 0, 0, 0, 0, 8, 27, 35, 33, 31, 20, 5, 3, 9, 12, 0, 0, 0, 0, 0, 0, 0, 0, 5, 1, 0, 0, 0, 0, 0, 0, 3, 34, 42, 36, 34, 29, 12, 0, 0, 5, 1, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 22, 48, 50, 37, 32, 42, 37, 22, 13, 17, 18, 0, 0, 0, 0, 0, 0, 6, 15, 0, 0, 0, 0, 0, 0, 30, 66, 82, 65, 36, 45, 81, 100, 78, 54, 47, 35, 4, 0, 0, 0, 0, 0, 9, 31, 11, 0, 0, 0, 0, 0, 51, 105, 113, 68, 22, 22, 74, 132, 121, 89, 74, 57, 18, 0, 0, 0, 0, 0, 18, 53, 37, 0, 0, 0, 0, 0, 49, 126, 139, 74, 0, 0, 11, 94, 121, 102, 93, 82, 40, 0, 0, 0, 0, 0, 30, 59, 36, 0, 0, 0, 0, 0, 33, 129, 151, 82, 0, 0, 0, 37, 84, 96, 105, 108, 69, 24, 0, 0, 0, 0, 39, 58, 21, 0, 0, 0, 0, 0, 26, 111, 137, 87, 6, 0, 0, 0, 50, 80, 112, 126, 88, 44, 7, 0, 0, 0, 34, 47, 3, 0, 0, 0, 0, 0, 18, 90, 111, 83, 32, 0, 0, 0, 29, 61, 100, 111, 86, 45, 2, 0, 0, 0, 29, 37, 0, 0, 0, 0, 0, 0, 11, 73, 85, 70, 42, 0, 0, 0, 19, 56, 81, 71, 53, 30, 0, 0, 0, 0, 18, 14, 0, 0, 0, 0, 0, 0, 1, 49, 71, 64, 54, 24, 0, 0, 0, 33, 47, 20, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 51, 49, 53, 49, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 21, 37, 56, 38, 0, 0, 0, 0, 0, 0, 0, 2, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 24, 47, 30, 0, 0, 0, 0, 10, 12, 5, 19, 13, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 38, 46, 15, 0, 0, 7, 16, 14, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 2, 1, 0, 0, 0, 38, 60, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 39, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 40, 39, 35, 33, 29, 29, 42, 53, 51, 23, 0, 0, 0, 0, 0, 0, 0, 12, 6, 0, 0, 0, 0, 0, 0, 3, 27, 39, 36, 30, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 27, 26, 21, 8, 0, 0, 0, 0, 0, 7, 37, 42, 36, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 42, 47, 44, 32, 7, 0, 0, 0, 1, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 61, 55, 49, 52, 63, 64, 46, 26, 26, 29, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 90, 92, 69, 46, 52, 89, 117, 107, 71, 41, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 85, 93, 69, 18, 0, 22, 63, 86, 75, 45, 20, 4, 0, 0, 0, 0, 0, 0, 16, 7, 0, 0, 0, 3, 7, 0, 41, 65, 56, 0, 0, 0, 0, 0, 0, 24, 26, 27, 17, 2, 0, 0, 0, 15, 9, 0, 0, 0, 0, 0, 10, 14, 0, 16, 33, 0, 0, 0, 0, 0, 0, 0, 27, 41, 40, 25, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 5, 22, 36, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 6, 19, 14, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 42, 45, 28, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 39, 41, 23, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 14, 22, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 24, 30, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 22, 22, 0, 0, 0, 0, 5, 30, 42, 21, 0, 0, 0, 35, 51, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 86, 106, 98, 58, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 3, 58, 90, 92, 74, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 39, 41, 32, 14, 0, 0, 0, 0, 0, 0, 14, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 42, 47, 45, 41, 37, 32, 25, 18, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 22, 30, 35, 35, 35, 36, 38, 38, 36, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 12, 11, 10, 11, 18, 25, 29, 31, 33, 35, 38, 39, 37, 36, 37, 42, 0, 0, 0, 0, 0, 0, 0, 0, 18, 35, 38, 35, 31, 29, 29, 31, 32, 34, 35, 38, 39, 34, 29, 29, 34, 43, 0, 0, 0, 0, 0, 0, 0, 11, 28, 31, 33, 35, 32, 30, 31, 33, 35, 35, 33, 30, 27, 25, 25, 28, 34, 30, 7, 0, 0, 0, 0, 0, 0, 8, 16, 24, 32, 37, 35, 31, 31, 33, 34, 33, 28, 21, 18, 21, 29, 43, 44, 24, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 23, 30, 30, 30, 31, 35, 35, 30, 23, 19, 24, 37, 51, 52, 36, 287, 287, 289, 293, 297, 290, 263, 221, 202, 214, 244, 268, 280, 281, 281, 267, 254, 240, 234, 242, 263, 288, 303, 313, 315, 317, 291, 298, 302, 303, 304, 303, 286, 248, 234, 246, 281, 301, 310, 302, 280, 241, 209, 177, 163, 168, 199, 237, 268, 292, 314, 320, 327, 329, 322, 309, 304, 310, 318, 312, 312, 311, 318, 319, 310, 289, 253, 213, 179, 152, 144, 148, 173, 206, 241, 266, 293, 313, 324, 337, 338, 314, 296, 300, 317, 325, 314, 286, 266, 258, 247, 236, 223, 208, 180, 162, 165, 178, 198, 217, 232, 250, 265, 294, 231, 288, 318, 299, 265, 242, 239, 240, 216, 196, 195, 200, 208, 219, 228, 227, 214, 200, 206, 221, 242, 253, 245, 238, 244, 271, 137, 237, 288, 270, 208, 141, 107, 95, 97, 114, 143, 170, 198, 226, 244, 252, 236, 211, 197, 204, 222, 242, 236, 224, 229, 247, 73, 200, 275, 268, 175, 61, 0, 0, 6, 46, 97, 139, 177, 219, 240, 231, 194, 157, 135, 142, 168, 207, 223, 217, 214, 229, 41, 183, 270, 287, 202, 87, 0, 0, 0, 14, 57, 95, 140, 182, 200, 173, 125, 80, 74, 96, 132, 187, 222, 219, 205, 206, 33, 172, 262, 308, 273, 191, 122, 75, 37, 17, 29, 50, 99, 141, 161, 121, 74, 41, 58, 94, 140, 198, 233, 233, 206, 194, 31, 170, 265, 321, 319, 261, 209, 150, 91, 20, 3, 12, 63, 116, 138, 101, 61, 53, 77, 107, 155, 213, 244, 248, 222, 205, 0, 146, 247, 317, 337, 283, 218, 142, 66, 1, 0, 10, 54, 110, 140, 114, 91, 89, 94, 99, 138, 191, 226, 240, 236, 230, 0, 51, 169, 269, 313, 279, 200, 101, 22, 0, 30, 64, 113, 158, 179, 158, 143, 133, 116, 110, 136, 173, 205, 227, 245, 261, 0, 0, 46, 186, 269, 272, 211, 122, 68, 78, 111, 157, 199, 229, 241, 227, 213, 186, 150, 133, 150, 175, 213, 247, 279, 297, 0, 0, 0, 86, 205, 262, 247, 232, 226, 239, 240, 250, 249, 251, 261, 281, 299, 275, 229, 189, 184, 195, 239, 283, 307, 309, 0, 0, 0, 0, 123, 210, 250, 289, 311, 301, 267, 237, 210, 197, 216, 267, 311, 303, 278, 246, 223, 224, 260, 288, 297, 295, 0, 0, 0, 0, 45, 126, 182, 237, 257, 237, 192, 142, 104, 109, 155, 220, 260, 254, 245, 231, 207, 195, 224, 246, 263, 273, 0, 0, 0, 0, 0, 5, 50, 100, 131, 128, 84, 20, 0, 0, 78, 192, 241, 239, 211, 173, 139, 135, 171, 208, 237, 255, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 110, 185, 181, 122, 60, 15, 12, 53, 111, 160, 190, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 287, 294, 301, 304, 303, 296, 283, 277, 279, 277, 256, 228, 195, 156, 123, 112, 100, 90, 82, 81, 83, 90, 108, 135, 170, 203, 254, 277, 293, 302, 305, 298, 282, 261, 249, 240, 205, 163, 122, 94, 80, 71, 62, 61, 57, 57, 57, 64, 70, 86, 123, 170, 207, 256, 287, 300, 304, 296, 276, 238, 204, 176, 148, 111, 76, 56, 47, 40, 45, 55, 53, 42, 37, 37, 32, 41, 79, 133, 171, 234, 278, 298, 301, 291, 263, 220, 185, 158, 132, 94, 59, 41, 27, 22, 35, 57, 66, 51, 37, 22, 8, 10, 45, 98, 171, 236, 275, 288, 286, 278, 257, 226, 198, 168, 140, 102, 56, 25, 8, 7, 28, 65, 84, 71, 45, 23, 3, 2, 19, 64, 162, 237, 275, 263, 247, 246, 249, 233, 205, 175, 143, 98, 46, 15, 0, 1, 35, 75, 101, 89, 59, 33, 13, 4, 10, 37, 148, 230, 263, 242, 205, 194, 209, 213, 200, 182, 153, 110, 61, 25, 0, 6, 42, 88, 109, 98, 64, 36, 21, 9, 8, 19, 134, 227, 258, 230, 170, 140, 159, 176, 179, 175, 164, 126, 82, 52, 10, 11, 38, 86, 104, 82, 48, 23, 13, 6, 3, 14, 124, 217, 249, 226, 158, 119, 113, 143, 164, 167, 170, 142, 98, 70, 24, 7, 26, 77, 88, 57, 25, 13, 10, 3, 4, 16, 105, 183, 223, 222, 161, 117, 100, 125, 150, 157, 156, 137, 100, 76, 30, 8, 27, 66, 65, 37, 12, 5, 8, 11, 16, 32, 76, 135, 185, 202, 170, 122, 100, 117, 140, 146, 134, 119, 100, 76, 30, 15, 34, 62, 59, 37, 11, 0, 4, 17, 32, 56, 39, 89, 139, 179, 172, 131, 103, 103, 114, 119, 97, 81, 80, 72, 47, 40, 48, 69, 65, 40, 11, 0, 3, 24, 55, 85, 3, 39, 81, 138, 160, 132, 100, 75, 72, 76, 68, 59, 61, 64, 59, 64, 66, 68, 55, 37, 7, 0, 0, 33, 78, 119, 0, 0, 12, 72, 126, 130, 99, 54, 36, 37, 48, 55, 59, 66, 77, 84, 70, 58, 43, 24, 0, 0, 9, 56, 108, 156, 0, 0, 0, 10, 73, 107, 89, 50, 32, 39, 61, 70, 70, 66, 83, 93, 83, 52, 16, 0, 0, 0, 32, 84, 138, 192, 0, 0, 0, 0, 29, 76, 84, 56, 49, 57, 78, 93, 91, 66, 63, 71, 57, 21, 0, 0, 0, 0, 43, 99, 153, 202, 0, 0, 0, 0, 1, 61, 73, 65, 64, 66, 71, 66, 57, 39, 25, 21, 2, 0, 0, 0, 0, 0, 7, 74, 126, 153, 0, 0, 0, 0, 0, 44, 53, 35, 14, 13, 14, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 13, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 63, 44, 28, 53, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 120, 108, 72, 46, 0, 0, 0, 0, 0, 26, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 107, 115, 62, 0, 0, 0, 0, 0, 0, 43, 46, 30, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 105, 70, 0, 0, 0, 0, 0, 0, 57, 55, 38, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 61, 0, 0, 20, 120, 104, 0, 0, 0, 0, 0, 0, 73, 84, 45, 35, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 91, 57, 0, 59, 163, 160, 45, 0, 0, 0, 0, 0, 88, 141, 68, 10, 11, 0, 0, 0, 0, 86, 0, 0, 0, 0, 52, 104, 44, 97, 206, 213, 110, 0, 0, 0, 0, 0, 128, 198, 89, 0, 3, 28, 0, 0, 0, 156, 82, 0, 0, 0, 0, 41, 19, 93, 235, 260, 168, 16, 0, 0, 0, 0, 200, 240, 89, 0, 0, 28, 18, 0, 0, 182, 164, 0, 0, 0, 0, 0, 0, 39, 236, 287, 199, 42, 0, 0, 0, 0, 282, 268, 71, 0, 0, 0, 9, 0, 27, 163, 171, 46, 0, 0, 0, 0, 0, 0, 211, 284, 201, 44, 0, 0, 0, 59, 327, 270, 54, 0, 0, 0, 0, 0, 108, 148, 104, 75, 0, 0, 0, 0, 0, 0, 182, 225, 162, 24, 0, 0, 0, 71, 297, 242, 46, 0, 0, 0, 0, 29, 200, 166, 38, 42, 0, 0, 0, 0, 0, 53, 162, 138, 86, 0, 0, 0, 0, 28, 228, 206, 36, 0, 0, 0, 0, 72, 241, 212, 29, 0, 0, 0, 0, 0, 0, 121, 140, 52, 0, 0, 0, 0, 0, 0, 157, 176, 32, 0, 0, 0, 0, 68, 247, 253, 49, 0, 0, 0, 0, 0, 0, 55, 43, 0, 0, 0, 0, 0, 0, 0, 95, 148, 29, 0, 0, 0, 0, 39, 223, 272, 76, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 85, 116, 0, 0, 0, 0, 0, 0, 183, 270, 101, 0, 0, 74, 118, 0, 0, 0, 0, 0, 22, 0, 0, 0, 32, 62, 102, 57, 0, 0, 0, 0, 0, 0, 139, 235, 86, 0, 0, 124, 250, 67, 0, 0, 0, 0, 163, 169, 81, 57, 87, 115, 93, 0, 0, 0, 0, 0, 0, 0, 110, 173, 0, 0, 0, 176, 359, 172, 0, 0, 0, 0, 226, 314, 257, 152, 101, 84, 31, 0, 0, 0, 0, 0, 0, 0, 69, 82, 0, 0, 0, 210, 452, 300, 0, 0, 0, 0, 186, 307, 293, 176, 74, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 268, 524, 395, 93, 0, 0, 5, 108, 185, 188, 109, 38, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 433, 585, 415, 166, 23, 11, 35, 58, 81, 81, 49, 19, 4, 0, 0, 0, 6, 18, 22, 29, 0, 0, 0, 0, 0, 245, 598, 539, 298, 122, 58, 49, 46, 38, 36, 32, 16, 1, 0, 0, 0, 3, 20, 32, 25, 16, 0, 0, 0, 0, 0, 456, 620, 394, 142, 59, 66, 70, 57, 42, 31, 23, 10, 0, 0, 0, 3, 16, 31, 25, 0, 0, 0, 0, 0, 0, 0, 484, 529, 255, 55, 37, 74, 87, 72, 49, 29, 17, 8, 0, 0, 0, 11, 29, 34, 2, 0, 0, 25, 0, 0, 0, 0, 366, 371, 152, 12, 19, 60, 81, 72, 45, 20, 7, 8, 12, 14, 17, 21, 23, 2, 0, 0, 27, 83, 0, 0, 0, 8, 215, 217, 83, 0, 0, 33, 58, 57, 28, 0, 0, 11, 37, 53, 49, 22, 0, 0, 0, 15, 132, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 87, 74, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 38, 59, 86, 91, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 51, 29, 18, 22, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 30, 46, 53, 44, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 35, 29, 14, 0, 5, 23, 39, 32, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 37, 42, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 116, 137, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 18, 0, 0, 0, 0, 0, 0, 0, 0, 68, 180, 240, 188, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 78, 84, 55, 21, 0, 0, 0, 0, 0, 0, 0, 4, 87, 121, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 90, 66, 33, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 69, 48, 21, 0, 0, 0, 28, 68, 67, 36, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 99, 198, 224, 174, 111, 43, 9, 36, 86, 101, 87, 61, 32, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 75, 194, 302, 330, 274, 187, 101, 25, 16, 80, 157, 178, 164, 143, 109, 71, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 148, 297, 351, 282, 175, 77, 2, 0, 0, 65, 169, 233, 251, 218, 153, 84, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 88, 187, 184, 95, 8, 0, 0, 0, 0, 27, 134, 228, 271, 225, 130, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 80, 156, 209, 219, 159, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66, 167, 208, 189, 131, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 44, 54, 67, 103, 133, 140, 95, 31, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 39, 110, 197, 288, 329, 284, 198, 109, 38, 4, 0, 0, 0, 0, 0, 0, 0, 0, 87, 13, 0, 0, 0, 0, 138, 242, 287, 308, 351, 404, 405, 339, 226, 97, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 194, 95, 0, 0, 0, 191, 363, 401, 337, 252, 216, 219, 208, 172, 116, 54, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 212, 149, 23, 0, 100, 292, 377, 315, 179, 76, 33, 25, 27, 25, 18, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 138, 121, 59, 67, 188, 273, 270, 164, 60, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 89, 121, 205, 295, 282, 201, 99, 30, 5, 1, 1, 3, 3, 0, 0, 0, 0, 0, 0, 1, 8, 10, 0, 0, 0, 19, 81, 187, 327, 399, 337, 210, 106, 44, 21, 10, 3, 2, 0, 0, 0, 0, 0, 0, 12, 22, 20, 1, 0, 0, 0, 3, 58, 166, 301, 367, 320, 210, 127, 80, 64, 51, 38, 27, 13, 1, 0, 0, 0, 0, 16, 23, 10, 0, 0, 0, 0, 334, 349, 357, 358, 358, 350, 329, 297, 272, 270, 280, 275, 249, 222, 188, 150, 101, 64, 46, 55, 79, 103, 123, 143, 171, 207, 278, 308, 338, 359, 366, 361, 333, 280, 231, 215, 216, 207, 194, 171, 135, 87, 30, 0, 0, 0, 0, 19, 52, 84, 120, 160, 221, 264, 317, 355, 369, 362, 333, 279, 225, 187, 175, 165, 145, 114, 72, 26, 0, 0, 0, 0, 0, 0, 0, 24, 73, 119, 181, 225, 292, 345, 360, 353, 331, 295, 240, 178, 133, 99, 71, 39, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 87, 136, 189, 262, 317, 328, 316, 300, 269, 220, 148, 81, 37, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 61, 59, 138, 230, 278, 273, 239, 217, 200, 164, 98, 38, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 79, 201, 253, 210, 129, 81, 73, 84, 57, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 41, 178, 245, 201, 96, 10, 0, 8, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 151, 237, 220, 134, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 124, 215, 235, 176, 76, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 97, 175, 206, 173, 95, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 116, 152, 142, 83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 76, 93, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 28, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 67, 0, 0, 0, 0, 0, 0, 0, 15, 4, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 22, 65, 125, 0, 0, 0, 0, 0, 0, 0, 13, 25, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 75, 128, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 6, 46, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 10, 76, 77, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 2, 82, 59, 0, 0, 1, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 29, 0, 0, 0, 0, 0, 0, 0, 0, 94, 44, 0, 0, 14, 55, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 74, 69, 0, 0, 0, 0, 0, 0, 0, 0, 106, 35, 0, 0, 0, 53, 37, 0, 0, 0, 0, 0, 0, 0, 0, 23, 110, 81, 0, 0, 0, 0, 0, 0, 0, 0, 116, 20, 0, 0, 0, 0, 42, 17, 8, 8, 0, 0, 0, 0, 0, 44, 138, 74, 0, 0, 0, 0, 0, 0, 0, 0, 88, 1, 0, 0, 0, 0, 15, 60, 80, 61, 0, 0, 0, 0, 0, 50, 139, 45, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 0, 7, 106, 125, 75, 0, 0, 0, 0, 0, 42, 111, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 129, 109, 0, 0, 0, 0, 0, 0, 22, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 76, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 29, 9, 0, 0, 0, 0, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 44, 37, 1, 3, 0, 0, 0, 83, 31, 0, 0, 0, 53, 88, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 58, 25, 0, 10, 0, 0, 39, 129, 67, 0, 0, 0, 89, 129, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 60, 65, 21, 0, 20, 0, 0, 119, 196, 107, 0, 0, 0, 7, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 37, 36, 5, 0, 44, 9, 68, 179, 236, 80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 78, 68, 139, 218, 183, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 104, 148, 225, 231, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 0, 0, 1, 7, 85, 204, 281, 192, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 0, 0, 6, 22, 33, 49, 194, 265, 118, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 0, 0, 0, 21, 42, 38, 19, 127, 169, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 35, 40, 9, 0, 42, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 35, 39, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 12, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 28, 22, 18, 22, 34, 36, 41, 43, 42, 29, 14, 13, 0, 0, 0, 0, 0, 0, 0, 2, 32, 31, 19, 20, 38, 55, 65, 66, 61, 56, 60, 66, 70, 73, 74, 70, 66, 68, 10, 0, 0, 0, 0, 0, 0, 51, 74, 61, 47, 49, 60, 72, 80, 81, 81, 79, 82, 84, 84, 84, 86, 88, 88, 85, 37, 15, 0, 0, 0, 0, 26, 85, 96, 83, 78, 77, 78, 81, 84, 85, 86, 87, 88, 89, 87, 88, 93, 97, 93, 86, 48, 36, 0, 0, 0, 0, 65, 99, 94, 88, 88, 89, 89, 87, 86, 86, 88, 90, 92, 93, 95, 101, 105, 105, 96, 88, 71, 48, 17, 0, 0, 39, 90, 98, 86, 84, 86, 87, 88, 87, 86, 87, 90, 96, 101, 106, 110, 112, 109, 103, 96, 96, 98, 61, 28, 7, 24, 73, 97, 95, 82, 81, 82, 84, 86, 85, 85, 86, 91, 100, 108, 114, 115, 109, 100, 91, 93, 103, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 1, 0, 0, 0, 45, 69, 54, 38, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 11, 0, 0, 0, 64, 98, 80, 62, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 4, 0, 0, 0, 25, 44, 27, 25, 34, 1, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 20, 17, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 44, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 48, 73, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 72, 61, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 12, 23, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 57, 22, 0, 0, 36, 71, 53, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 81, 105, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 124, 105, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 127, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 418, 425, 426, 424, 422, 414, 383, 324, 278, 268, 302, 339, 359, 349, 334, 300, 254, 205, 181, 194, 231, 268, 298, 323, 351, 378, 388, 413, 429, 433, 432, 423, 384, 317, 256, 240, 273, 318, 340, 331, 299, 237, 152, 68, 24, 41, 104, 175, 234, 279, 316, 350, 371, 410, 427, 436, 438, 435, 406, 348, 289, 261, 277, 299, 305, 290, 249, 164, 54, 0, 0, 0, 3, 80, 158, 221, 281, 324, 341, 389, 414, 422, 430, 428, 413, 375, 319, 268, 241, 230, 223, 210, 175, 101, 2, 0, 0, 0, 0, 53, 118, 186, 252, 302, 247, 312, 361, 382, 383, 358, 329, 293, 239, 174, 117, 99, 108, 126, 118, 77, 14, 0, 0, 0, 24, 73, 121, 174, 226, 281, 63, 178, 272, 316, 286, 197, 116, 68, 37, 1, 0, 0, 32, 82, 111, 109, 61, 4, 0, 0, 34, 82, 122, 159, 205, 254, 0, 22, 183, 258, 198, 40, 0, 0, 0, 0, 0, 0, 5, 77, 123, 129, 75, 0, 0, 0, 0, 55, 94, 122, 167, 225, 0, 0, 119, 237, 181, 0, 0, 0, 0, 0, 0, 0, 0, 54, 105, 92, 11, 0, 0, 0, 0, 21, 64, 82, 121, 182, 0, 0, 76, 255, 250, 90, 0, 0, 0, 0, 0, 0, 0, 0, 44, 9, 0, 0, 0, 0, 0, 18, 61, 66, 83, 134, 0, 0, 45, 260, 324, 228, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 68, 67, 64, 91, 0, 0, 2, 225, 321, 274, 148, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 61, 57, 46, 64, 0, 0, 0, 139, 254, 239, 125, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 48, 47, 48, 77, 0, 0, 0, 0, 133, 165, 84, 0, 0, 0, 0, 0, 0, 0, 13, 20, 0, 0, 0, 0, 0, 13, 53, 67, 87, 135, 0, 0, 0, 0, 0, 54, 48, 0, 0, 0, 0, 0, 0, 21, 51, 72, 55, 0, 0, 0, 9, 65, 113, 141, 174, 210, 0, 0, 0, 0, 0, 0, 4, 42, 33, 24, 28, 28, 9, 0, 15, 65, 94, 75, 51, 47, 82, 138, 183, 213, 236, 257, 0, 0, 0, 0, 0, 0, 0, 16, 74, 82, 33, 0, 0, 0, 0, 10, 78, 100, 102, 101, 121, 154, 178, 196, 216, 234, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 74, 94, 90, 79, 82, 85, 95, 115, 149, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 26, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 153, 158, 162, 163, 161, 157, 150, 144, 128, 108, 88, 65, 42, 22, 25, 38, 42, 40, 32, 31, 38, 55, 69, 84, 102, 120, 142, 154, 161, 163, 162, 156, 146, 124, 91, 68, 44, 18, 2, 0, 7, 24, 37, 24, 4, 0, 7, 19, 32, 54, 81, 106, 133, 153, 162, 164, 164, 153, 138, 108, 86, 57, 30, 8, 0, 0, 10, 29, 48, 22, 0, 0, 0, 0, 0, 24, 55, 89, 134, 158, 165, 166, 166, 154, 131, 99, 79, 45, 17, 0, 0, 0, 13, 29, 40, 23, 0, 0, 0, 0, 0, 2, 31, 70, 121, 157, 160, 162, 164, 150, 119, 85, 64, 45, 15, 0, 0, 0, 9, 25, 45, 34, 9, 0, 0, 0, 0, 0, 19, 52, 99, 134, 134, 138, 150, 131, 92, 58, 48, 36, 9, 0, 0, 0, 0, 18, 48, 49, 14, 0, 0, 0, 0, 0, 10, 40, 81, 109, 102, 97, 104, 80, 34, 3, 10, 13, 0, 0, 0, 0, 0, 19, 54, 58, 10, 0, 0, 0, 0, 0, 0, 24, 61, 84, 70, 69, 73, 52, 13, 0, 0, 2, 0, 0, 0, 0, 0, 24, 62, 48, 0, 0, 0, 0, 0, 0, 0, 10, 36, 51, 39, 33, 25, 32, 5, 8, 5, 8, 0, 0, 0, 0, 0, 30, 66, 27, 0, 0, 0, 0, 0, 0, 0, 3, 19, 35, 31, 26, 9, 21, 27, 47, 40, 16, 0, 0, 0, 0, 0, 28, 56, 1, 0, 0, 0, 0, 1, 5, 3, 11, 0, 25, 40, 48, 37, 38, 57, 73, 56, 3, 0, 0, 0, 0, 0, 25, 43, 0, 0, 0, 0, 0, 4, 21, 24, 32, 0, 0, 29, 62, 70, 66, 79, 73, 18, 0, 0, 0, 0, 0, 0, 21, 21, 0, 0, 0, 0, 0, 0, 21, 37, 53, 0, 0, 0, 56, 75, 66, 60, 25, 0, 0, 0, 0, 0, 0, 13, 26, 5, 0, 0, 0, 0, 0, 0, 23, 57, 78, 0, 0, 0, 28, 60, 53, 32, 0, 0, 0, 0, 0, 0, 1, 34, 35, 9, 0, 0, 0, 0, 0, 0, 35, 77, 94, 0, 0, 0, 0, 35, 31, 0, 0, 0, 0, 0, 0, 0, 22, 37, 24, 0, 0, 0, 0, 0, 0, 3, 63, 99, 114, 0, 0, 0, 0, 8, 12, 0, 0, 0, 0, 6, 0, 0, 15, 17, 0, 0, 0, 0, 0, 0, 0, 30, 93, 117, 119, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 91, 98, 91, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 44, 41, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 22, 43, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 11, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 9, 14, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 8, 9, 12, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 9, 14, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 19, 31, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 10, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 14, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 22, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 1, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 10, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 8, 0, 45, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 0, 45, 8, 0, 4, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 37, 5, 0, 12, 32, 4, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 19, 4, 0, 0, 37, 7, 0, 19, 48, 22, 0, 0, 0, 0, 8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 9, 29, 40, 26, 0, 0, 48, 20, 11, 31, 66, 37, 0, 0, 0, 0, 11, 5, 0, 0, 0, 0, 0, 0, 8, 29, 44, 58, 61, 48, 23, 0, 60, 44, 39, 55, 68, 26, 0, 0, 0, 0, 0, 0, 0, 0, 3, 11, 20, 38, 49, 58, 68, 74, 79, 74, 60, 51, 65, 73, 75, 82, 57, 0, 0, 0, 0, 0, 0, 0, 0, 7, 32, 49, 57, 64, 72, 78, 83, 89, 91, 89, 86, 85, 58, 84, 107, 104, 28, 0, 0, 0, 0, 11, 12, 12, 19, 35, 50, 63, 70, 77, 84, 88, 91, 94, 94, 95, 99, 103, 55, 81, 115, 103, 0, 0, 0, 0, 44, 59, 60, 57, 57, 61, 65, 69, 74, 82, 89, 94, 96, 96, 95, 98, 105, 109, 60, 78, 102, 76, 0, 0, 0, 37, 74, 79, 73, 68, 65, 67, 70, 74, 79, 86, 93, 96, 96, 96, 98, 104, 110, 109, 71, 76, 75, 38, 0, 0, 6, 53, 74, 77, 76, 73, 70, 71, 75, 80, 84, 88, 92, 94, 95, 98, 103, 109, 112, 102, 81, 66, 53, 12, 0, 0, 28, 57, 68, 69, 66, 67, 70, 76, 83, 87, 88, 87, 87, 89, 93, 101, 108, 112, 111, 93, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 37, 32, 26, 35, 43, 33, 5, 0, 2, 20, 23, 18, 12, 18, 22, 11, 22, 9, 0, 0, 0, 0, 0, 0, 15, 57, 72, 54, 33, 32, 25, 8, 0, 0, 16, 39, 39, 30, 20, 19, 25, 21, 36, 9, 0, 0, 0, 0, 0, 4, 24, 53, 58, 33, 12, 7, 3, 0, 0, 3, 42, 69, 72, 55, 43, 32, 24, 22, 19, 0, 0, 0, 0, 0, 0, 0, 1, 7, 14, 17, 12, 7, 1, 3, 12, 21, 51, 76, 79, 65, 50, 37, 25, 19, 4, 0, 1, 6, 0, 0, 0, 0, 0, 0, 5, 31, 36, 25, 18, 24, 32, 31, 49, 73, 73, 51, 31, 24, 15, 12, 29, 23, 34, 26, 0, 0, 0, 21, 37, 34, 43, 64, 63, 46, 34, 33, 29, 10, 26, 63, 67, 43, 13, 4, 11, 6, 71, 74, 77, 49, 0, 0, 24, 92, 117, 91, 69, 76, 68, 50, 34, 17, 0, 0, 9, 66, 87, 60, 18, 0, 8, 12, 102, 116, 116, 69, 20, 19, 68, 145, 179, 124, 78, 83, 72, 52, 29, 0, 0, 0, 24, 95, 125, 89, 44, 9, 8, 12, 113, 145, 152, 89, 23, 5, 47, 124, 161, 109, 76, 95, 87, 66, 33, 5, 0, 0, 56, 124, 140, 93, 54, 20, 7, 7, 108, 154, 169, 106, 24, 0, 12, 59, 93, 67, 77, 123, 121, 97, 56, 29, 4, 11, 76, 135, 133, 85, 47, 17, 3, 9, 104, 148, 161, 103, 33, 8, 0, 4, 27, 51, 102, 165, 167, 137, 88, 51, 19, 26, 84, 126, 117, 74, 36, 10, 6, 20, 97, 129, 147, 102, 41, 18, 0, 0, 18, 85, 155, 203, 188, 146, 94, 52, 25, 46, 94, 119, 111, 79, 42, 27, 29, 41, 85, 118, 136, 101, 58, 34, 3, 4, 53, 139, 200, 200, 164, 116, 76, 41, 25, 54, 87, 110, 111, 84, 58, 49, 44, 40, 76, 108, 142, 114, 85, 59, 41, 34, 79, 147, 175, 146, 96, 59, 53, 49, 36, 50, 71, 93, 107, 83, 62, 43, 22, 19, 76, 97, 136, 132, 99, 74, 74, 59, 65, 86, 82, 57, 40, 37, 49, 57, 43, 41, 46, 77, 93, 72, 37, 9, 0, 0, 79, 92, 124, 136, 106, 70, 81, 79, 61, 43, 19, 0, 17, 42, 62, 74, 63, 57, 48, 52, 58, 39, 10, 0, 0, 1, 82, 95, 124, 125, 74, 41, 65, 85, 79, 34, 7, 0, 25, 62, 90, 91, 85, 80, 60, 41, 26, 19, 10, 12, 19, 33, 86, 102, 118, 102, 34, 0, 29, 70, 67, 43, 31, 33, 73, 112, 124, 114, 67, 40, 22, 0, 0, 0, 5, 28, 49, 65, 103, 109, 102, 82, 14, 0, 23, 97, 120, 100, 83, 87, 112, 137, 134, 107, 43, 0, 0, 0, 0, 0, 0, 3, 22, 33, 118, 125, 102, 76, 8, 0, 65, 150, 154, 115, 78, 65, 71, 73, 59, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 109, 138, 122, 70, 7, 20, 109, 153, 109, 45, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 113, 109, 44, 17, 53, 115, 89, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 65, 66, 22, 28, 74, 88, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 28, 19, 43, 83, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 12, 45, 75, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 15, 24, 27, 33, 33, 15, 0, 0, 0, 0, 0, 0, 0, 20, 50, 53, 47, 45, 50, 48, 43, 40, 40, 43, 2, 8, 15, 19, 22, 25, 33, 17, 0, 0, 0, 0, 0, 0, 0, 39, 63, 60, 51, 54, 63, 63, 62, 55, 54, 53, 32, 31, 26, 22, 23, 25, 33, 23, 4, 0, 1, 5, 0, 4, 38, 74, 84, 76, 64, 70, 74, 70, 63, 61, 61, 61, 49, 52, 43, 34, 30, 29, 26, 20, 7, 2, 8, 17, 35, 52, 78, 98, 96, 78, 70, 73, 83, 81, 65, 58, 65, 68, 42, 54, 57, 50, 33, 6, 0, 0, 0, 1, 19, 41, 70, 81, 95, 111, 113, 85, 70, 73, 85, 83, 73, 61, 67, 71, 38, 45, 62, 57, 30, 0, 0, 0, 0, 0, 19, 48, 80, 91, 92, 109, 108, 78, 53, 49, 69, 84, 85, 78, 70, 73, 50, 46, 56, 50, 11, 0, 0, 0, 0, 0, 0, 30, 68, 86, 85, 93, 83, 56, 26, 18, 50, 85, 101, 96, 74, 67, 71, 43, 30, 33, 5, 0, 0, 0, 0, 0, 0, 6, 50, 67, 76, 90, 70, 32, 0, 0, 37, 82, 110, 109, 85, 63, 73, 27, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 31, 53, 77, 92, 75, 28, 0, 0, 34, 84, 117, 121, 101, 73, 62, 22, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 38, 77, 101, 89, 31, 0, 0, 36, 85, 119, 128, 112, 90, 45, 17, 30, 21, 23, 29, 28, 12, 0, 0, 0, 0, 0, 18, 77, 113, 97, 35, 0, 0, 46, 90, 120, 129, 118, 107, 24, 11, 53, 54, 60, 67, 75, 37, 0, 0, 0, 0, 0, 18, 80, 110, 79, 16, 0, 0, 41, 79, 106, 114, 113, 121, 18, 15, 59, 90, 80, 86, 85, 29, 0, 0, 0, 0, 0, 37, 86, 103, 62, 2, 0, 0, 7, 46, 80, 108, 122, 125, 32, 25, 61, 103, 97, 91, 83, 36, 0, 0, 0, 0, 27, 64, 104, 111, 75, 11, 0, 0, 0, 17, 71, 109, 113, 106, 50, 36, 62, 102, 108, 85, 70, 30, 0, 0, 0, 18, 39, 75, 116, 99, 57, 0, 0, 0, 0, 1, 61, 93, 96, 93, 63, 41, 56, 93, 102, 66, 35, 28, 18, 12, 22, 26, 16, 51, 96, 70, 7, 0, 0, 0, 0, 16, 74, 101, 99, 84, 66, 40, 48, 77, 76, 23, 0, 0, 27, 42, 33, 2, 0, 0, 45, 49, 0, 0, 0, 0, 0, 46, 103, 118, 100, 76, 60, 42, 49, 61, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 22, 69, 116, 127, 102, 69, 34, 28, 44, 51, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 36, 52, 72, 95, 107, 94, 68, 6, 16, 48, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 37, 48, 57, 65, 67, 74, 85, 91, 84, 71, 0, 22, 68, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 70, 79, 78, 76, 76, 76, 79, 84, 83, 77, 14, 48, 95, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 43, 68, 84, 88, 85, 81, 79, 77, 78, 80, 79, 73, 44, 71, 99, 50, 0, 0, 0, 0, 17, 50, 67, 72, 75, 80, 84, 87, 88, 86, 83, 82, 79, 76, 78, 81, 79, 68, 69, 85, 85, 0, 0, 0, 0, 25, 69, 83, 88, 90, 93, 91, 88, 85, 83, 82, 82, 82, 82, 84, 84, 82, 75, 59, 86, 92, 71, 0, 0, 0, 0, 56, 81, 84, 85, 85, 88, 88, 84, 80, 80, 84, 88, 91, 93, 90, 82, 74, 64, 58, 93, 90, 54, 0, 0, 0, 0, 58, 74, 73, 72, 75, 82, 84, 81, 77, 78, 84, 93, 100, 99, 92, 77, 60, 56, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 53, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66, 76, 76, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 67, 83, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 60, 63, 19, 0, 0, 0, 0, 20, 42, 58, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 25, 90, 138, 171, 170, 134, 46, 0, 0, 0, 22, 28, 25, 0, 0, 0, 0, 0, 24, 0, 0, 2, 67, 136, 187, 192, 187, 215, 251, 279, 290, 281, 239, 177, 122, 106, 62, 34, 0, 0, 0, 0, 24, 129, 191, 188, 169, 185, 234, 291, 339, 351, 337, 338, 355, 376, 394, 404, 404, 385, 366, 357, 130, 72, 0, 0, 0, 2, 158, 309, 387, 385, 358, 355, 378, 409, 427, 432, 433, 433, 442, 454, 467, 479, 487, 489, 488, 488, 217, 130, 44, 5, 20, 145, 318, 451, 497, 471, 436, 420, 425, 438, 453, 463, 471, 480, 489, 498, 506, 515, 522, 528, 531, 533, 310, 200, 109, 81, 127, 264, 417, 509, 511, 487, 469, 463, 460, 462, 470, 480, 491, 502, 512, 523, 532, 540, 544, 549, 553, 551, 409, 278, 181, 155, 221, 345, 480, 520, 502, 486, 482, 480, 475, 474, 480, 491, 504, 519, 533, 544, 551, 557, 566, 574, 577, 576, 495, 373, 274, 237, 292, 402, 505, 510, 487, 480, 483, 482, 480, 479, 485, 498, 516, 534, 549, 557, 561, 565, 573, 582, 595, 600, 550, 468, 384, 334, 365, 449, 510, 500, 478, 477, 479, 478, 476, 477, 485, 500, 520, 539, 553, 555, 552, 549, 555, 578, 605, 620, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 43, 36, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 48, 63, 57, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 8, 17, 0, 0, 8, 19, 26, 26, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 0, 0, 16, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 15, 8, 13, 25, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 9, 35, 60, 50, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 59, 52, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 62, 67, 67, 67, 61, 46, 32, 36, 57, 62, 58, 51, 40, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 30, 52, 67, 71, 62, 46, 29, 31, 48, 54, 41, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 59, 74, 71, 63, 46, 31, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 73, 79, 78, 60, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 54, 64, 75, 66, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 28, 29, 62, 83, 57, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 16, 0, 0, 23, 69, 69, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 23, 0, 0, 0, 0, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 31, 61, 81, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 85, 65, 7, 0, 0, 34, 83, 134, 163, 126, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 125, 143, 103, 23, 0, 0, 0, 71, 152, 210, 211, 119, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 70, 159, 178, 139, 32, 0, 0, 0, 54, 142, 210, 234, 184, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 158, 193, 148, 26, 0, 0, 0, 34, 127, 194, 226, 217, 126, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 115, 177, 122, 0, 0, 0, 0, 27, 121, 181, 217, 224, 176, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 134, 82, 0, 0, 0, 0, 51, 138, 179, 207, 211, 175, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 91, 53, 0, 0, 0, 0, 104, 171, 188, 190, 177, 132, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 34, 0, 0, 0, 10, 145, 197, 194, 161, 123, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 4, 0, 0, 0, 26, 152, 196, 176, 115, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 32, 149, 190, 163, 79, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 136, 176, 143, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 69, 153, 184, 123, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 152, 226, 214, 107, 0, 0, 0, 0, 0, 27, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 82, 190, 286, 324, 274, 130, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 118, 168, 272, 365, 425, 428, 365, 232, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 167, 283, 360, 436, 493, 513, 489, 445, 369, 277, 199, 171, 0, 0, 0, 0, 0, 0, 0, 0, 2, 34, 4, 0, 58, 194, 338, 446, 511, 543, 553, 546, 533, 517, 493, 459, 428, 422, 0, 0, 0, 0, 0, 0, 0, 8, 224, 304, 302, 303, 348, 431, 513, 571, 596, 597, 591, 582, 572, 562, 554, 546, 541, 541, 63, 0, 0, 0, 0, 0, 0, 255, 440, 494, 487, 488, 515, 557, 599, 625, 634, 627, 615, 601, 587, 575, 569, 567, 562, 554, 239, 111, 0, 0, 0, 0, 196, 441, 560, 590, 592, 597, 609, 622, 633, 639, 638, 629, 616, 601, 586, 577, 574, 573, 562, 543, 393, 240, 31, 0, 0, 101, 390, 551, 605, 605, 608, 615, 620, 624, 625, 626, 625, 622, 612, 602, 592, 590, 590, 586, 568, 538, 505, 353, 137, 0, 31, 273, 502, 597, 610, 603, 606, 613, 614, 611, 608, 608, 611, 618, 620, 617, 613, 608, 599, 586, 565, 544, 568, 462, 288, 163, 225, 419, 575, 622, 615, 603, 603, 605, 606, 600, 592, 591, 598, 615, 630, 635, 625, 603, 577, 556, 556, 569, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 14, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 75, 76, 63, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 57, 51, 33, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 17, 27, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 30, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 33, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 20, 1, 0, 0, 0, 10, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 80, 81, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 63, 96, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 47, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 87, 83, 88, 90, 89, 92, 102, 112, 101, 68, 35, 13, 0, 0, 16, 67, 110, 125, 123, 112, 104, 106, 114, 118, 122, 120, 91, 94, 94, 89, 84, 84, 86, 80, 56, 23, 1, 0, 0, 11, 52, 108, 147, 142, 121, 104, 105, 112, 115, 120, 132, 139, 115, 128, 113, 93, 83, 76, 65, 49, 36, 30, 33, 30, 40, 69, 109, 151, 172, 146, 112, 97, 99, 100, 100, 105, 128, 150, 162, 173, 135, 97, 84, 75, 59, 55, 71, 87, 89, 79, 82, 111, 142, 165, 171, 142, 104, 85, 83, 82, 80, 96, 118, 147, 197, 200, 145, 104, 98, 98, 79, 72, 93, 116, 105, 85, 86, 109, 130, 140, 160, 156, 124, 97, 89, 86, 87, 94, 113, 134, 185, 188, 131, 103, 120, 127, 101, 73, 79, 91, 79, 62, 66, 88, 108, 130, 170, 185, 146, 106, 92, 100, 106, 102, 105, 115, 151, 164, 113, 87, 106, 120, 89, 44, 42, 63, 60, 52, 54, 79, 107, 141, 187, 197, 143, 88, 73, 101, 119, 110, 99, 101, 132, 148, 93, 49, 53, 69, 52, 23, 30, 60, 61, 49, 50, 76, 112, 148, 197, 176, 91, 31, 40, 91, 125, 118, 101, 102, 103, 124, 79, 31, 25, 44, 49, 50, 80, 96, 71, 47, 45, 73, 111, 144, 179, 130, 27, 0, 18, 88, 129, 129, 114, 116, 57, 85, 76, 40, 27, 51, 93, 132, 157, 137, 74, 34, 35, 69, 103, 136, 163, 98, 2, 0, 24, 96, 138, 147, 143, 144, 1, 46, 85, 83, 61, 77, 146, 190, 188, 123, 33, 4, 24, 62, 97, 137, 159, 95, 15, 0, 41, 105, 150, 169, 171, 168, 0, 0, 84, 126, 109, 118, 172, 212, 175, 60, 0, 0, 19, 66, 107, 154, 165, 107, 39, 19, 49, 100, 147, 171, 179, 177, 0, 0, 37, 127, 144, 142, 155, 154, 81, 0, 0, 0, 50, 106, 142, 168, 152, 97, 51, 30, 41, 81, 127, 156, 178, 188, 0, 0, 0, 84, 144, 147, 121, 83, 25, 0, 3, 55, 113, 156, 178, 170, 129, 83, 48, 14, 15, 59, 117, 163, 195, 199, 0, 0, 0, 19, 109, 134, 108, 72, 56, 80, 125, 143, 150, 166, 180, 171, 127, 76, 35, 3, 16, 77, 142, 189, 213, 196, 0, 0, 0, 0, 67, 90, 76, 63, 90, 155, 186, 161, 120, 106, 125, 125, 87, 39, 6, 0, 33, 96, 163, 210, 210, 173, 0, 0, 0, 0, 31, 49, 20, 28, 80, 154, 172, 118, 39, 5, 18, 32, 14, 0, 0, 0, 21, 81, 139, 182, 176, 139, 0, 0, 0, 0, 12, 0, 0, 0, 1, 74, 84, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 66, 67, 50, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 12, 43, 92, 143, 179, 181, 143, 77, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 25, 110, 169, 194, 214, 245, 276, 300, 314, 311, 292, 269, 254, 0, 0, 0, 0, 0, 0, 0, 46, 112, 126, 108, 95, 108, 151, 214, 268, 299, 321, 341, 360, 378, 392, 402, 404, 404, 405, 0, 0, 0, 0, 0, 0, 33, 143, 226, 260, 256, 244, 245, 263, 295, 326, 352, 374, 393, 408, 420, 429, 436, 442, 447, 453, 126, 0, 0, 0, 0, 19, 137, 237, 304, 344, 356, 353, 347, 345, 352, 367, 385, 403, 420, 433, 444, 451, 456, 462, 467, 470, 287, 115, 0, 0, 0, 94, 212, 301, 352, 378, 387, 384, 376, 371, 376, 389, 406, 424, 439, 450, 456, 463, 472, 481, 489, 491, 408, 247, 74, 0, 14, 131, 250, 319, 351, 368, 380, 386, 383, 380, 386, 400, 419, 438, 451, 457, 459, 464, 474, 493, 512, 515, 469, 357, 205, 93, 79, 164, 266, 318, 334, 348, 359, 365, 366, 370, 380, 399, 423, 445, 456, 455, 446, 441, 456, 490, 526, 540, 
    
    
    others => 0);
end ifmap_package;
