library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    160, 18, 64, 
    260, 81, 188, 
    257, 0, 0, 
    
    -- channel=1
    71, 0, 28, 
    0, 0, 186, 
    0, 0, 0, 
    
    -- channel=2
    0, 49, 0, 
    0, 146, 0, 
    0, 0, 0, 
    
    -- channel=3
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=4
    260, 0, 0, 
    2, 0, 0, 
    0, 0, 0, 
    
    -- channel=5
    168, 0, 56, 
    0, 0, 0, 
    0, 0, 2, 
    
    -- channel=6
    0, 0, 0, 
    0, 0, 0, 
    0, 83, 55, 
    
    -- channel=7
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=8
    0, 0, 15, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=9
    168, 378, 308, 
    55, 275, 130, 
    183, 53, 0, 
    
    -- channel=10
    0, 45, 121, 
    0, 333, 98, 
    0, 0, 0, 
    
    -- channel=11
    0, 0, 126, 
    16, 53, 0, 
    106, 0, 209, 
    
    -- channel=12
    0, 0, 0, 
    0, 176, 176, 
    0, 160, 51, 
    
    -- channel=13
    119, 210, 129, 
    198, 0, 0, 
    8, 169, 87, 
    
    -- channel=14
    0, 101, 200, 
    0, 161, 60, 
    0, 88, 122, 
    
    -- channel=15
    0, 0, 0, 
    6, 0, 92, 
    0, 0, 0, 
    
    -- channel=16
    0, 44, 230, 
    0, 119, 72, 
    0, 255, 36, 
    
    -- channel=17
    0, 0, 25, 
    0, 54, 0, 
    0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=19
    0, 0, 0, 
    0, 0, 0, 
    0, 93, 77, 
    
    -- channel=20
    181, 108, 170, 
    0, 0, 0, 
    0, 0, 63, 
    
    -- channel=21
    0, 27, 48, 
    21, 0, 0, 
    0, 281, 179, 
    
    -- channel=22
    0, 18, 0, 
    170, 0, 189, 
    182, 38, 0, 
    
    -- channel=23
    0, 40, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=24
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=25
    192, 292, 324, 
    335, 208, 104, 
    23, 0, 64, 
    
    -- channel=26
    0, 0, 9, 
    87, 22, 0, 
    207, 93, 0, 
    
    -- channel=27
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=28
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=29
    168, 1, 184, 
    30, 40, 150, 
    144, 21, 99, 
    
    -- channel=30
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=31
    0, 0, 0, 
    0, 0, 0, 
    0, 283, 158, 
    
    -- channel=32
    0, 0, 108, 
    0, 0, 0, 
    0, 121, 248, 
    
    -- channel=33
    67, 4, 255, 
    103, 18, 17, 
    0, 0, 28, 
    
    -- channel=34
    0, 105, 65, 
    0, 134, 78, 
    49, 0, 0, 
    
    -- channel=35
    145, 108, 81, 
    23, 38, 70, 
    0, 176, 253, 
    
    -- channel=36
    224, 0, 120, 
    0, 16, 0, 
    0, 0, 0, 
    
    -- channel=37
    0, 89, 171, 
    193, 251, 239, 
    106, 143, 219, 
    
    -- channel=38
    59, 83, 20, 
    16, 0, 0, 
    123, 70, 171, 
    
    -- channel=39
    98, 90, 316, 
    162, 109, 140, 
    122, 291, 81, 
    
    -- channel=40
    151, 161, 0, 
    0, 0, 0, 
    60, 0, 7, 
    
    -- channel=41
    0, 0, 0, 
    0, 0, 0, 
    260, 0, 0, 
    
    -- channel=42
    0, 0, 30, 
    79, 162, 303, 
    140, 0, 0, 
    
    -- channel=43
    347, 314, 353, 
    131, 161, 114, 
    312, 18, 0, 
    
    -- channel=44
    0, 136, 112, 
    220, 224, 173, 
    318, 205, 174, 
    
    -- channel=45
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=46
    200, 31, 191, 
    70, 75, 78, 
    27, 38, 0, 
    
    -- channel=47
    30, 115, 315, 
    159, 54, 30, 
    6, 170, 165, 
    
    -- channel=48
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=49
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=50
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=51
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=52
    106, 67, 118, 
    257, 102, 124, 
    0, 0, 0, 
    
    -- channel=53
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=54
    0, 89, 105, 
    0, 49, 0, 
    0, 0, 0, 
    
    -- channel=55
    61, 0, 0, 
    16, 49, 114, 
    237, 0, 0, 
    
    -- channel=56
    0, 0, 0, 
    0, 0, 0, 
    112, 300, 383, 
    
    -- channel=57
    208, 0, 0, 
    0, 0, 50, 
    0, 103, 8, 
    
    -- channel=58
    57, 33, 222, 
    109, 68, 118, 
    132, 321, 235, 
    
    -- channel=59
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=60
    178, 120, 110, 
    63, 127, 146, 
    0, 0, 0, 
    
    -- channel=61
    0, 0, 28, 
    401, 0, 30, 
    52, 135, 328, 
    
    -- channel=62
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 88, 
    
    -- channel=63
    74, 70, 0, 
    0, 0, 0, 
    243, 215, 197, 
    
    
    others => 0);
end gold_package_package;
