-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;


-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity ifmap_36k_layer0_entity9 is
    generic (
        DEVICE: string := "7SERIES"
        );

    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic_vector(2-1 downto 0);;
        DI   : in std_logic_vector(16-1 downto 0);
        ADDR : in std_logic_vector(11-1 downto 0);
        DO   : out std_logic_vector(16-1 downto 0)
    );
 end ifmap_36k_layer0_entity9;

  architecture a1 of bram is

    begin

    BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
    generic map (
       BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
       DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
       DO_REG => 0,                     -- Optional output register (0 or 1)
       INIT => X"000000000000000000",   -- Initial values on output port
       INIT_FILE => "NONE",
       WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       SRVAL => X"000000000000000000",  -- Set/Reset value for port output
       WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
       -- The following INIT_xx declarations specify the initial contents of the RAM
       INIT_00 => X"00a000b900d100d900e600f600f900f600f800f300e600dd00da00dd00d800c7",
       INIT_01 => X"00bc00bb00b800b400a600900079008b006a00660066004f005e0065005b005e",
       INIT_02 => X"00e100ef00f200e600e800f500f300eb00ed00e600d800cd00c900cb00c800ba",
       INIT_03 => X"00af00ab00a1007f008e008d007a00870076005200250034005f006b00610064",
       INIT_04 => X"00fc00f900f100dc00d900e200df00d600d500cf00c300b800b300b600b300a7",
       INIT_05 => X"009f0098009400810080008c0080007200570028000400260063007300690069",
       INIT_06 => X"00e900e100de00d300d300cb00c800c000bb00b700ae00a400a000a500a00099",
       INIT_07 => X"0091008d008c008a007d007d007f0069003b0025001a0037007000780070006d",
       INIT_08 => X"00cf00c300cf00c900be00b400b300ab00a3009f00990092009100970093008d",
       INIT_09 => X"00870088008300870081007a0084005a003a003d00300056007500780072006d",
       INIT_0A => X"00b600ab00aa00a20099009c009f00970090008d008c008a008b008d008a008a",
       INIT_0B => X"0087008c0086008a008c008900660045004b003e00430074008100800070006e",
       INIT_0C => X"008d00880088008600880086008c008500870089008b008d008f0092008e0091",
       INIT_0D => X"00910091008a008f008e006b002f00210048004b006c007f00840084006f0070",
       INIT_0E => X"0076007d0080008100880083008a00840088008c009000930096009e009a0099",
       INIT_0F => X"009200950093009400800042000d0011005000750080007a007b008000720070",
       INIT_10 => X"0073007e00840085008b0087008f0089008b0091009500980094009a00a300aa",
       INIT_11 => X"009e00a2009d00940073002c000e001e0069008b0088007e0077007a0074006f",
       INIT_12 => X"0076008000880088008d00880091008d008d0093009a00a5009d009a00a200a7",
       INIT_13 => X"009b00930091008a00630038002e0037006d007c007a007e007300740075006e",
       INIT_14 => X"007d0084008b0089008e00880090008c008b0090009600990083008b00900098",
       INIT_15 => X"00a600ba00d300d60080005c0045002a0055005f006300730070006f0071006b",
       INIT_16 => X"00850089008e008a008d0088008e008a0089008f00880084008e00b600c900cb",
       INIT_17 => X"00d200ce00cf00c000a200bd0092002a001b002800670072006d006a006c0068",
       INIT_18 => X"008c008b008f008b008f008c008a008900870085009000a400ab00a000890073",
       INIT_19 => X"006a005d004b003b006f00dc00c9005f000d0007003e00740063006500690064",
       INIT_1A => X"0090008a008f008c009200920082008700820091008c006e005e005c00310013",
       INIT_1B => X"001d003200190012007800d100d2009d0026000600130044004500520063005f",
       INIT_1C => X"0091008b0092008e0090008e007900800085007f0054004400560052002e0016",
       INIT_1D => X"00130032001e004100af00c900cd00cb006600100012001600230038004f0058",
       INIT_1E => X"008f008b00940090008a0084008b00830075004200480056006a004e00280022",
       INIT_1F => X"00240046007300b600cb00c500cd00c3006c003d002500120018004f00640053",
       INIT_20 => X"008e008b00930090008500720084007900510059003c0045005500440053009b",
       INIT_21 => X"00c000db00ed00eb00d700d700d300720030005d003500140041008b008f0054",
       INIT_22 => X"008f008d008e008900740045003a00430051004b001d001c00240019008c00f2",
       INIT_23 => X"00ec00eb00e300dc00db00df0095003a00390054004e004e008500a100a7005b",
       INIT_24 => X"008f008c00880086008d0047002d00340043002100170016002f0029009b00d9",
       INIT_25 => X"00c700be00bf00d000dc00df00ad0067005d0073008700950098009400a50059",
       INIT_26 => X"008f008c007e00b500bd004c0021002b003900150010001700390042009e00c2",
       INIT_27 => X"00b600b300c400c900c200ce00de00b30097009c009500970096009200880042",
       INIT_28 => X"008c0085009a00ea00b5005a0026002a0034000b000b000b0014003100a000ba",
       INIT_29 => X"00b000b900b900730045005a00a100c400b700aa00a0009900930088004d0026",
       INIT_2A => X"0082008000a300a3008b006a002d002e001c00030009000f001e003600a200b4",
       INIT_2B => X"00ac00be00710015001400150030009500bb00ab008e00850080004300150027",
       INIT_2C => X"007c00840067001a0048006c0034003000120007000b003b005a006300a500b0",
       INIT_2D => X"00b100a9002a001d002f0026000e00460095008800750075003c000e00150030",
       INIT_2E => X"0079007c0049001e003b00720044001f000d000e00180048004f006c00bb00bb",
       INIT_2F => X"00bf008b001b002b001e001b001c001b006c0084007b005900160015002a003b",
       INIT_30 => X"006d00660047003f003c0071004d001c0010001f003000470046008800bd00b3",
       INIT_31 => X"00b40074001f003600350029001b000e00480085007c003c001200220032003b",
       INIT_32 => X"00570051003d003c003a0069004b00150014002e004c00600061009100a400a3",
       INIT_33 => X"00aa00710020003900470031002500110029006c00600021000c001d00280032",
       INIT_34 => X"004900490040003c0039005f0057002f003d0062008900a500a900b000b700b6",
       INIT_35 => X"00b6007c002200360060005c0033001b00110046003b000c00060012001d0028",
       INIT_36 => X"004900490045004e004100590045002f0034003c004a0056005b006000620060",
       INIT_37 => X"006200530020003c003b003e001d001400040011000a00030007000a00110021",
       INIT_38 => X"004b005300480036002d0027000f0004000300020005000700070008000a000b",
       INIT_39 => X"000b000d000800420043002f0038000f00020002000100030006000a000f0020",
       INIT_3A => X"005000590051002f0015000a00100019000e000a000e000e000e000e000e000c",
       INIT_3B => X"000a000900060017003e0048002a000700030004000500050007000b00150021",
       INIT_3C => X"0049004f00490037002e002f003b003a001a00110019001c001f0020001d001c",
       INIT_3D => X"001800150010000c00140016000800060008000700080008000b000f001b001f",
       INIT_3E => X"00450048004c004e005800530048003800200026002b002a002f003300320031",
       INIT_3F => X"002c0026001e001c002200220013000c000e0010000f000d0012001a001e001d",

       -- The next set of INIT_xx are valid when configured as 36Kb
       INIT_40 => X"002500310039003a0042004e0050005100560052004900420041004300430038",
       INIT_41 => X"0032003200400073003400380032002700160022002e0024001d001200150013",
       INIT_42 => X"00430048004d00440043004a004800420044004000390034003200360037002e",
       INIT_43 => X"0029002a0027002900280023001e00210022002e001e001b001c001500160012",
       INIT_44 => X"004800440048003e003a003d003800310030002d002b00280026002a002b0026",
       INIT_45 => X"00220023001e001c00230021001f002200300022000d000e0015001400130011",
       INIT_46 => X"00380036003d003c003e0030002b00240023002300220020001f002100220020",
       INIT_47 => X"001d001e001b001d0020001c001d0025002a0012000b000f0016001300100011",
       INIT_48 => X"003900390042003b003400240020001b001c001d001c001a001a001a001c001e",
       INIT_49 => X"001c001c001c001c001c00300043002a00190012000d0019001b001f00130011",
       INIT_4A => X"003b003a002f0021001a001a0019001600170019001a001900180018001b001f",
       INIT_4B => X"001d001e0021001e0021005d005e003c0029001b001e002c002b002d00180013",
       INIT_4C => X"0022001c001700140016001700160015001600160019001a00180019001d0023",
       INIT_4D => X"0020001f0023001e003300590037002500380028002b002d0024001e00170015",
       INIT_4E => X"0011001100100012001600170016001600180017001a001b0019001b001d0027",
       INIT_4F => X"0028002d00330030004100400012000b00220025001f00200019001600160015",
       INIT_50 => X"0011001200120012001500160017001700190018001c001e002500380033003b",
       INIT_51 => X"003b003a00370036003d002800110010001a00190018001b001a001700150014",
       INIT_52 => X"001300120012001200150014001600180018001900200031003e004c00390034",
       INIT_53 => X"0031002e0032003a003800310030002c00290023001900190019001800140014",
       INIT_54 => X"00140012001300120015001500150017001900190024003500310042003e004a",
       INIT_55 => X"0068008900a600b8007c0068004b00210038003d002600190018001900120013",
       INIT_56 => X"001500120014001300180018001600180019001d001f00300055009700b200be",
       INIT_57 => X"00cd00cd00ca00c500b200d00098001600180025004600280015001600110011",
       INIT_58 => X"0014001400160015001800180019001a00190020004200700090009b008c0075",
       INIT_59 => X"006400580047003d007500e800d5004e000f000a00320046001a001500110010",
       INIT_5A => X"0014001600190016001700170019001a001a00480067005b0050005600340012",
       INIT_5B => X"00110022000f0010007c00dd00e0009b002400070016003b0021001300120010",
       INIT_5C => X"00180017001b0016001800190013001500370055003a0029003d004e00320018",
       INIT_5D => X"000b002b001e004900bf00d800d100cd0067000e00100017001b001600140012",
       INIT_5E => X"001a0016001a001700190025003c0034004c00340038003b0050004d002e0026",
       INIT_5F => X"00230049007c00c400df00d800d900d2007600390015000e001f0047003e0011",
       INIT_60 => X"0019001400190017002100350060005c0049005d003e004200510047005a00a2",
       INIT_61 => X"00c400df00f500f500e300e400de00790025003b001100090048008c00750013",
       INIT_62 => X"001900150018001a0028002c00350045005800520025002900310020009400fb",
       INIT_63 => X"00f600f200e900e200e100e2008b001f000b001900280043008500a200970022",
       INIT_64 => X"0016001300160026005d0046002e0036004b00260018001b0038003100a300e3",
       INIT_65 => X"00d600cd00cb00da00e500e400a3004a0039005a008000950097009600a00033",
       INIT_66 => X"0013000f0026007c00af005a0024002a003f0017000b00150040004f00aa00d0",
       INIT_67 => X"00c700c500d300d600ce00d900e300b1009800a800a700a2009a00970088002a",
       INIT_68 => X"0012000a006500dc00be006f002f002e0039000a0009000e001f004200b100cc",
       INIT_69 => X"00c200ca00c6007c004f006600ac00d300c800b800b100a9009c008c004a0011",
       INIT_6A => X"000e0014008400a50096008000370034001e0003000a0016002d004800b400c6",
       INIT_6B => X"00be00cd007b0019001a001e003800a300ca00b8009e009300880044000d0011",
       INIT_6C => X"000a00230053002100530082003e00350013000700100048006c007500b700c2",
       INIT_6D => X"00c300b7002f001e0031002b0014004f00a10094008400810040000a00090018",
       INIT_6E => X"000a00210037002300460088004e0024000f0011002200580061007e00cd00cd",
       INIT_6F => X"00d000980020002b0020001f0020001f00750091008a00630017000c00190021",
       INIT_70 => X"000a001500360041004700880057002100150027003f00570056009a00cf00c5",
       INIT_71 => X"00c60081002500380037002c001c000f004d0093008b0043000e0014001c001f",
       INIT_72 => X"0007000e002f003e004500800056001c001e003c005e006f006f00a200b600b4",
       INIT_73 => X"00bc007f0029003c004b00350023000f002c007a006f00260007000d00100016",
       INIT_74 => X"000b00110027003b004600750068003d00510079009f00b700b900c300c900c7",
       INIT_75 => X"00c60088002a003c006600620034001c0015004f0045001000030007000c0016",
       INIT_76 => X"00130014001d0043004900670055003c00450050005b0064006800710071006d",
       INIT_77 => X"006d00590025004100400042001f001700080014000e000500060006000b0018",
       INIT_78 => X"0017001c001d0025002c002c00160007000a000a000c000c000d001000110010",
       INIT_79 => X"000f000f000900430044003000380010000400030003000400060009000e0019",
       INIT_7A => X"002100250027002000170012001900200017001500170017001700150013000f",
       INIT_7B => X"000b000a00070018003e00470029000800040005000500060009000e0018001d",
       INIT_7C => X"0023002500290032003c00430051004d002c0024002d00300031002c00270023",
       INIT_7D => X"001d001b0015001000170019000a0009000b0009000a000b000e0014001f001e",
       INIT_7E => X"002a002a003b0057006d006f006600520037003e00450047004a004800460043",
       INIT_7F => X"003b0033002b0029002f002c0018001200140016001500130016001c0020001e",

       -- The next set of INITP_xx are for the parity bits
       INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

       -- The next set of INIT_xx are valid when configured as 36Kb
       INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000")
    port map (
       DO => DO,      -- Output data, width defined by READ_WIDTH parameter
       ADDR => ADDR,  -- Input address, width defined by read/write port depth
       CLK => CLK,    -- 1-bit input clock
       DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
       EN => EN,      -- 1-bit input RAM enable
       REGCE => REGCE, -- 1-bit input output register enable
       RST => RST,    -- 1-bit input reset
       WE => WE       -- Input write enable, width defined by write port depth
    );


-- End of BRAM_SINGLE_MACRO_inst instantiation
