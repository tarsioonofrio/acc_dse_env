library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    5, 0, 6, 10, 1, 0, 3, 3, 6, 7, 3, 0, 0, 0, 0, 4, 9, 16, 24, 37, 37, 32, 27, 21, 20, 20, 20, 21, 28, 32, 
    4, 0, 2, 6, 0, 0, 1, 3, 0, 0, 0, 7, 6, 2, 4, 10, 31, 38, 47, 52, 60, 58, 47, 48, 29, 24, 21, 19, 22, 27, 
    2, 0, 0, 4, 0, 0, 3, 2, 0, 0, 0, 21, 23, 9, 27, 50, 61, 56, 36, 40, 50, 60, 65, 57, 50, 30, 19, 17, 23, 26, 
    12, 5, 4, 5, 0, 0, 6, 2, 0, 0, 0, 56, 58, 50, 64, 90, 78, 24, 8, 23, 35, 52, 52, 58, 58, 55, 27, 12, 21, 28, 
    62, 41, 4, 0, 0, 0, 2, 1, 0, 0, 10, 57, 68, 84, 81, 76, 49, 0, 0, 17, 34, 44, 45, 46, 73, 88, 46, 6, 13, 29, 
    95, 86, 0, 0, 0, 0, 0, 1, 7, 15, 25, 24, 43, 74, 55, 43, 45, 0, 0, 10, 51, 49, 32, 49, 90, 88, 68, 14, 3, 27, 
    108, 58, 0, 0, 2, 0, 0, 0, 30, 39, 15, 0, 24, 70, 53, 42, 53, 25, 0, 0, 59, 61, 44, 60, 79, 88, 80, 39, 0, 15, 
    99, 18, 0, 0, 13, 1, 0, 0, 0, 43, 0, 0, 34, 77, 66, 54, 65, 51, 0, 0, 36, 63, 65, 55, 59, 69, 86, 74, 12, 0, 
    58, 0, 0, 20, 26, 19, 0, 0, 0, 28, 0, 0, 53, 65, 72, 56, 82, 60, 0, 0, 12, 55, 68, 46, 46, 59, 82, 93, 50, 8, 
    49, 0, 0, 31, 29, 28, 0, 0, 0, 48, 17, 0, 51, 57, 55, 69, 91, 39, 0, 0, 14, 57, 84, 46, 30, 57, 74, 94, 70, 35, 
    47, 0, 0, 30, 26, 24, 28, 0, 0, 51, 3, 0, 22, 58, 48, 44, 98, 9, 0, 0, 45, 74, 89, 47, 32, 48, 64, 76, 69, 52, 
    48, 0, 0, 49, 24, 16, 61, 0, 0, 31, 0, 0, 0, 57, 42, 29, 86, 0, 0, 0, 63, 85, 77, 55, 41, 40, 47, 56, 54, 54, 
    32, 0, 26, 90, 17, 3, 69, 10, 0, 0, 0, 0, 0, 49, 36, 39, 85, 0, 0, 6, 60, 70, 69, 53, 43, 28, 19, 42, 48, 40, 
    17, 0, 41, 103, 19, 0, 58, 26, 0, 0, 0, 0, 37, 47, 32, 47, 83, 0, 0, 6, 62, 60, 70, 55, 28, 17, 12, 40, 44, 27, 
    11, 0, 21, 98, 33, 0, 43, 42, 0, 0, 0, 21, 80, 37, 43, 54, 58, 0, 0, 0, 37, 66, 80, 57, 26, 23, 28, 40, 31, 4, 
    14, 0, 0, 86, 63, 0, 23, 51, 11, 0, 0, 63, 70, 43, 46, 43, 24, 0, 0, 11, 21, 66, 84, 71, 41, 29, 37, 30, 3, 0, 
    12, 0, 0, 69, 85, 0, 0, 50, 38, 21, 34, 39, 42, 20, 41, 47, 0, 2, 60, 44, 17, 78, 117, 78, 50, 17, 6, 3, 0, 10, 
    3, 0, 0, 41, 90, 15, 0, 29, 36, 82, 31, 7, 19, 0, 28, 73, 0, 3, 45, 32, 67, 105, 99, 59, 25, 0, 0, 0, 0, 11, 
    0, 0, 0, 18, 84, 31, 0, 33, 46, 82, 48, 0, 0, 0, 9, 82, 39, 19, 51, 71, 113, 109, 81, 47, 5, 0, 0, 9, 19, 22, 
    0, 0, 0, 13, 86, 24, 0, 0, 61, 66, 18, 0, 0, 0, 5, 68, 56, 68, 86, 104, 98, 83, 68, 39, 26, 15, 19, 47, 54, 50, 
    0, 0, 0, 17, 84, 0, 0, 0, 3, 51, 7, 0, 0, 0, 30, 75, 80, 85, 101, 82, 63, 52, 44, 49, 44, 42, 55, 71, 76, 74, 
    0, 0, 0, 11, 47, 0, 0, 0, 24, 78, 80, 44, 45, 61, 72, 95, 97, 92, 82, 61, 54, 52, 54, 60, 59, 54, 50, 60, 68, 64, 
    2, 0, 0, 13, 0, 0, 0, 0, 82, 147, 108, 73, 75, 75, 79, 81, 76, 75, 70, 61, 61, 60, 60, 55, 52, 49, 48, 57, 60, 54, 
    49, 14, 0, 14, 0, 0, 0, 61, 148, 125, 77, 63, 65, 66, 65, 63, 65, 67, 63, 56, 58, 59, 49, 42, 39, 46, 49, 54, 49, 39, 
    68, 39, 7, 6, 0, 0, 0, 132, 147, 73, 61, 61, 66, 67, 65, 65, 64, 62, 56, 53, 49, 47, 43, 42, 49, 58, 51, 41, 30, 19, 
    76, 62, 44, 19, 0, 0, 47, 153, 100, 58, 51, 64, 72, 65, 62, 62, 61, 57, 53, 56, 50, 44, 46, 59, 69, 64, 43, 25, 28, 38, 
    75, 69, 60, 40, 0, 0, 85, 137, 74, 56, 51, 55, 65, 66, 63, 63, 59, 57, 56, 56, 59, 54, 57, 65, 66, 49, 29, 33, 73, 73, 
    75, 65, 64, 57, 15, 0, 78, 133, 73, 61, 48, 48, 56, 61, 63, 58, 55, 53, 54, 60, 62, 61, 60, 52, 39, 22, 27, 68, 105, 75, 
    81, 65, 59, 64, 53, 40, 80, 101, 82, 68, 58, 58, 57, 61, 58, 47, 42, 41, 48, 58, 63, 66, 53, 25, 0, 4, 46, 81, 96, 79, 
    78, 67, 58, 62, 64, 62, 71, 81, 85, 68, 65, 69, 72, 72, 61, 48, 41, 31, 37, 59, 67, 64, 39, 6, 0, 8, 63, 96, 93, 77, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 41, 44, 40, 25, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 31, 52, 69, 72, 65, 55, 49, 28, 21, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 6, 1, 17, 29, 57, 61, 62, 90, 105, 102, 80, 62, 47, 30, 15, 0, 0, 0, 
    2, 17, 0, 0, 0, 0, 0, 0, 0, 0, 29, 96, 55, 48, 72, 75, 57, 45, 73, 114, 130, 127, 111, 93, 82, 65, 39, 10, 0, 0, 
    56, 59, 20, 0, 0, 0, 0, 0, 0, 0, 10, 48, 58, 66, 57, 53, 60, 66, 86, 108, 124, 126, 108, 101, 111, 90, 40, 14, 0, 0, 
    99, 72, 0, 0, 0, 0, 0, 0, 0, 7, 23, 36, 64, 88, 81, 78, 84, 71, 88, 110, 117, 104, 93, 103, 110, 95, 65, 19, 0, 0, 
    127, 99, 9, 0, 0, 0, 0, 0, 17, 43, 52, 46, 90, 110, 100, 96, 102, 80, 70, 106, 129, 101, 90, 98, 97, 86, 66, 36, 10, 0, 
    177, 100, 61, 53, 5, 0, 2, 13, 61, 70, 48, 72, 120, 124, 96, 91, 89, 91, 56, 62, 122, 117, 97, 78, 82, 93, 80, 47, 13, 12, 
    208, 147, 104, 94, 29, 0, 5, 65, 127, 171, 122, 103, 121, 120, 98, 89, 93, 79, 38, 63, 124, 125, 119, 94, 85, 92, 100, 79, 34, 2, 
    203, 153, 149, 114, 28, 0, 0, 61, 155, 190, 134, 102, 124, 118, 110, 100, 89, 83, 33, 98, 153, 151, 138, 98, 96, 105, 100, 88, 60, 13, 
    207, 141, 154, 139, 39, 0, 0, 14, 68, 152, 118, 114, 138, 143, 109, 103, 103, 72, 44, 143, 188, 157, 131, 92, 90, 106, 108, 100, 79, 34, 
    200, 122, 160, 160, 65, 0, 0, 8, 40, 120, 84, 98, 164, 171, 121, 107, 129, 93, 67, 160, 184, 146, 121, 103, 92, 101, 103, 97, 85, 47, 
    186, 126, 193, 169, 69, 13, 22, 23, 41, 99, 92, 133, 200, 195, 149, 117, 119, 96, 85, 157, 172, 145, 111, 95, 85, 80, 90, 96, 76, 34, 
    189, 138, 202, 184, 103, 43, 54, 39, 42, 59, 119, 168, 167, 151, 132, 137, 118, 66, 61, 146, 151, 134, 136, 118, 99, 95, 90, 84, 51, 3, 
    203, 163, 200, 200, 144, 86, 77, 65, 66, 76, 135, 219, 192, 127, 122, 120, 94, 55, 59, 109, 127, 129, 110, 83, 82, 89, 78, 60, 15, 0, 
    217, 187, 208, 223, 176, 121, 113, 102, 69, 70, 132, 133, 131, 107, 101, 117, 92, 50, 64, 107, 124, 131, 119, 101, 73, 72, 47, 10, 0, 0, 
    226, 205, 212, 229, 194, 126, 122, 147, 101, 80, 108, 74, 84, 76, 94, 122, 97, 85, 90, 48, 66, 127, 112, 73, 39, 23, 0, 0, 0, 0, 
    211, 210, 207, 216, 205, 150, 128, 159, 163, 114, 63, 71, 100, 93, 134, 141, 96, 102, 109, 100, 107, 100, 88, 69, 38, 9, 0, 0, 0, 0, 
    190, 203, 194, 203, 209, 166, 123, 141, 158, 182, 122, 95, 121, 111, 168, 184, 116, 94, 130, 146, 152, 115, 99, 102, 95, 92, 72, 77, 79, 77, 
    188, 211, 193, 197, 210, 174, 124, 181, 186, 140, 138, 115, 124, 161, 211, 212, 173, 125, 117, 129, 133, 133, 124, 130, 150, 158, 171, 182, 179, 175, 
    212, 231, 203, 203, 205, 146, 105, 202, 283, 255, 200, 207, 229, 248, 267, 264, 241, 215, 185, 155, 157, 171, 193, 209, 219, 228, 235, 234, 235, 232, 
    256, 275, 226, 212, 205, 129, 138, 239, 313, 331, 294, 237, 237, 240, 243, 249, 233, 212, 212, 213, 220, 222, 230, 242, 244, 244, 246, 253, 255, 251, 
    263, 270, 253, 226, 211, 164, 196, 285, 334, 300, 237, 204, 198, 196, 197, 201, 213, 218, 223, 229, 237, 242, 243, 242, 245, 246, 246, 253, 257, 258, 
    267, 235, 227, 242, 195, 157, 229, 324, 320, 257, 218, 214, 216, 212, 212, 213, 219, 221, 224, 230, 239, 244, 246, 249, 252, 260, 265, 269, 271, 268, 
    293, 255, 224, 226, 202, 181, 275, 334, 274, 218, 224, 219, 225, 221, 212, 211, 215, 219, 225, 236, 248, 255, 255, 263, 275, 281, 282, 286, 283, 280, 
    301, 274, 244, 214, 201, 236, 305, 322, 240, 216, 224, 229, 226, 217, 217, 216, 219, 224, 233, 245, 254, 269, 277, 279, 275, 276, 277, 285, 292, 301, 
    301, 281, 260, 239, 205, 245, 325, 303, 243, 232, 225, 227, 231, 220, 216, 217, 224, 233, 239, 250, 259, 258, 263, 269, 270, 268, 277, 302, 314, 288, 
    289, 277, 263, 254, 230, 221, 287, 289, 230, 232, 231, 237, 240, 233, 224, 213, 215, 224, 237, 248, 253, 254, 251, 248, 251, 262, 294, 312, 289, 240, 
    292, 265, 256, 255, 245, 226, 224, 236, 222, 212, 212, 225, 234, 239, 230, 218, 225, 236, 240, 244, 245, 241, 235, 228, 241, 272, 300, 306, 289, 247, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 21, 13, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 27, 33, 29, 13, 11, 11, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 12, 0, 4, 22, 29, 20, 12, 26, 24, 9, 0, 0, 0, 
    0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 10, 19, 20, 7, 0, 11, 16, 10, 16, 24, 28, 17, 0, 0, 0, 
    25, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 23, 19, 22, 25, 20, 0, 3, 11, 11, 14, 13, 20, 15, 5, 0, 0, 
    53, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 13, 18, 20, 32, 14, 0, 0, 2, 12, 14, 6, 16, 15, 13, 0, 0, 
    83, 46, 2, 0, 0, 0, 0, 0, 0, 9, 13, 0, 0, 10, 4, 20, 13, 39, 0, 0, 7, 3, 28, 22, 7, 18, 22, 19, 9, 0, 
    100, 50, 19, 0, 0, 0, 0, 0, 0, 20, 18, 0, 0, 11, 6, 14, 6, 47, 0, 0, 31, 21, 41, 25, 15, 17, 26, 21, 17, 0, 
    108, 43, 14, 4, 0, 0, 0, 0, 0, 16, 9, 0, 0, 13, 8, 5, 4, 49, 0, 0, 42, 32, 37, 22, 22, 22, 28, 20, 17, 0, 
    102, 24, 18, 41, 0, 0, 0, 0, 0, 6, 0, 0, 0, 29, 16, 6, 15, 54, 0, 10, 44, 33, 30, 26, 25, 21, 17, 14, 11, 0, 
    91, 17, 28, 53, 0, 0, 0, 0, 0, 1, 0, 0, 33, 43, 20, 12, 21, 40, 0, 14, 38, 25, 26, 30, 19, 14, 8, 2, 0, 0, 
    81, 24, 34, 46, 40, 0, 0, 0, 0, 0, 0, 9, 50, 34, 26, 22, 13, 14, 0, 3, 24, 30, 33, 37, 24, 17, 7, 0, 0, 0, 
    79, 42, 41, 41, 69, 0, 0, 0, 0, 0, 14, 45, 48, 30, 16, 23, 11, 0, 0, 6, 9, 13, 22, 28, 24, 18, 6, 0, 0, 0, 
    79, 61, 53, 48, 81, 43, 0, 0, 0, 0, 30, 16, 10, 12, 0, 30, 12, 0, 0, 9, 0, 18, 39, 34, 15, 2, 0, 0, 0, 0, 
    70, 69, 63, 55, 70, 63, 15, 18, 10, 0, 26, 0, 0, 0, 0, 36, 27, 0, 0, 0, 0, 33, 32, 29, 0, 0, 0, 0, 0, 0, 
    51, 63, 60, 52, 61, 76, 35, 31, 29, 13, 31, 0, 21, 0, 0, 40, 35, 0, 4, 9, 34, 40, 32, 32, 0, 0, 0, 0, 0, 0, 
    31, 55, 51, 42, 55, 83, 36, 17, 46, 43, 40, 10, 18, 0, 18, 43, 42, 17, 30, 50, 62, 55, 52, 51, 46, 21, 0, 0, 0, 0, 
    31, 63, 50, 39, 62, 87, 19, 0, 35, 39, 37, 34, 37, 48, 64, 70, 72, 49, 54, 61, 68, 67, 72, 78, 90, 77, 73, 68, 75, 75, 
    70, 90, 64, 45, 59, 62, 0, 21, 55, 88, 110, 104, 108, 119, 121, 123, 127, 102, 93, 90, 100, 107, 117, 128, 136, 138, 138, 132, 138, 138, 
    137, 131, 91, 56, 64, 44, 0, 45, 96, 155, 158, 131, 129, 131, 129, 130, 134, 124, 126, 133, 138, 141, 146, 152, 151, 155, 155, 155, 158, 160, 
    176, 159, 116, 80, 91, 34, 11, 67, 140, 159, 137, 122, 121, 120, 120, 125, 135, 137, 143, 149, 152, 156, 156, 157, 152, 155, 156, 158, 165, 166, 
    186, 168, 135, 105, 94, 20, 28, 108, 167, 144, 134, 131, 134, 135, 131, 132, 137, 140, 143, 149, 155, 158, 158, 157, 160, 163, 169, 172, 173, 162, 
    196, 180, 155, 128, 103, 39, 59, 141, 150, 131, 137, 136, 141, 138, 133, 132, 135, 139, 144, 151, 160, 165, 166, 170, 177, 180, 186, 178, 173, 175, 
    199, 188, 168, 148, 128, 80, 88, 159, 136, 135, 141, 136, 141, 138, 135, 135, 140, 143, 150, 155, 168, 175, 175, 178, 181, 185, 180, 180, 188, 200, 
    196, 191, 178, 163, 150, 124, 116, 172, 139, 144, 144, 138, 142, 138, 139, 138, 141, 144, 151, 158, 166, 170, 173, 176, 174, 173, 177, 198, 200, 198, 
    192, 189, 177, 171, 158, 148, 133, 160, 144, 150, 146, 146, 148, 144, 142, 133, 134, 141, 147, 152, 160, 165, 166, 161, 155, 158, 176, 193, 190, 178, 
    185, 179, 168, 169, 158, 149, 138, 138, 144, 144, 140, 149, 149, 148, 145, 138, 139, 142, 141, 148, 157, 153, 154, 145, 144, 150, 173, 192, 194, 169, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    152, 163, 164, 157, 154, 159, 157, 158, 156, 154, 151, 150, 160, 170, 171, 168, 159, 148, 147, 144, 138, 138, 136, 141, 136, 133, 134, 139, 138, 130, 
    150, 160, 165, 156, 155, 160, 158, 161, 158, 154, 137, 131, 152, 166, 162, 160, 146, 143, 133, 112, 95, 92, 107, 118, 129, 138, 136, 137, 137, 130, 
    148, 150, 160, 157, 162, 164, 164, 163, 163, 165, 133, 118, 139, 153, 147, 147, 156, 137, 95, 72, 57, 51, 54, 69, 81, 103, 126, 134, 135, 134, 
    143, 145, 157, 161, 164, 167, 167, 164, 162, 161, 200, 184, 144, 142, 151, 136, 116, 80, 73, 67, 64, 51, 49, 51, 43, 72, 108, 126, 128, 129, 
    124, 135, 163, 165, 159, 166, 165, 160, 160, 148, 208, 178, 129, 103, 93, 72, 49, 59, 76, 68, 72, 77, 73, 50, 61, 51, 66, 105, 127, 126, 
    95, 78, 102, 137, 158, 167, 170, 163, 156, 148, 162, 138, 105, 77, 48, 46, 38, 57, 89, 87, 78, 82, 72, 78, 74, 50, 41, 72, 118, 127, 
    77, 38, 38, 92, 147, 164, 165, 163, 139, 137, 128, 97, 92, 79, 58, 66, 56, 46, 97, 127, 97, 68, 75, 92, 69, 50, 29, 47, 103, 124, 
    71, 19, 33, 86, 134, 157, 165, 144, 104, 68, 65, 86, 105, 89, 63, 61, 61, 56, 79, 110, 104, 71, 62, 65, 65, 46, 33, 24, 73, 123, 
    95, 27, 62, 103, 135, 150, 163, 145, 136, 91, 86, 105, 104, 91, 56, 55, 56, 59, 54, 75, 92, 76, 61, 61, 58, 53, 50, 27, 35, 95, 
    91, 60, 94, 115, 129, 145, 121, 177, 196, 157, 111, 122, 96, 82, 74, 60, 48, 49, 47, 72, 88, 96, 83, 67, 68, 60, 55, 38, 16, 47, 
    66, 85, 100, 123, 131, 155, 106, 149, 166, 155, 132, 140, 109, 76, 87, 61, 50, 26, 44, 111, 106, 113, 82, 57, 72, 71, 65, 47, 25, 29, 
    62, 67, 87, 129, 142, 161, 137, 98, 136, 142, 111, 118, 134, 93, 78, 76, 73, 22, 61, 131, 108, 104, 71, 57, 64, 80, 65, 51, 37, 47, 
    54, 64, 99, 100, 115, 151, 153, 94, 133, 131, 89, 104, 158, 139, 94, 74, 88, 36, 85, 122, 111, 86, 52, 51, 48, 54, 56, 56, 50, 75, 
    49, 78, 122, 65, 74, 122, 142, 95, 110, 102, 107, 84, 131, 126, 104, 103, 95, 41, 96, 134, 102, 85, 76, 70, 60, 53, 68, 78, 81, 93, 
    55, 88, 121, 63, 48, 89, 119, 80, 114, 101, 140, 169, 137, 107, 110, 108, 88, 59, 102, 136, 111, 86, 65, 51, 62, 65, 78, 104, 102, 95, 
    67, 85, 109, 89, 39, 88, 103, 74, 92, 93, 151, 184, 121, 106, 90, 83, 83, 53, 100, 160, 145, 91, 79, 65, 67, 81, 83, 94, 89, 108, 
    85, 81, 103, 113, 37, 66, 94, 99, 49, 95, 129, 112, 96, 79, 64, 60, 77, 72, 106, 83, 92, 117, 94, 62, 53, 71, 90, 93, 110, 141, 
    109, 92, 102, 116, 57, 42, 92, 110, 76, 68, 71, 84, 95, 81, 75, 42, 61, 111, 104, 49, 77, 99, 64, 46, 33, 46, 88, 108, 134, 145, 
    126, 101, 105, 115, 82, 41, 72, 65, 77, 97, 53, 93, 89, 69, 97, 56, 32, 95, 114, 116, 101, 57, 50, 29, 47, 64, 107, 132, 143, 139, 
    125, 104, 108, 111, 98, 64, 81, 59, 23, 48, 13, 46, 30, 58, 109, 78, 27, 47, 71, 88, 59, 22, 4, 0, 25, 41, 90, 110, 103, 101, 
    112, 102, 101, 109, 98, 56, 57, 111, 80, 29, 26, 58, 74, 117, 135, 117, 81, 63, 48, 15, 0, 2, 0, 2, 7, 28, 55, 62, 53, 52, 
    109, 112, 99, 108, 89, 33, 60, 139, 148, 111, 98, 87, 102, 111, 114, 105, 64, 49, 24, 5, 0, 0, 7, 10, 2, 6, 11, 21, 16, 5, 
    63, 104, 108, 104, 108, 69, 115, 138, 156, 141, 60, 33, 35, 29, 31, 33, 14, 10, 10, 7, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 34, 81, 108, 102, 86, 132, 150, 158, 75, 13, 4, 0, 2, 0, 5, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 31, 97, 73, 92, 134, 157, 93, 25, 3, 0, 4, 4, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 8, 4, 0, 0, 
    0, 0, 0, 36, 57, 113, 146, 123, 34, 7, 4, 3, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 11, 
    0, 0, 0, 0, 20, 125, 162, 87, 33, 10, 4, 3, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 8, 28, 
    0, 0, 0, 0, 0, 75, 147, 70, 27, 21, 10, 15, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 76, 26, 8, 4, 2, 13, 19, 20, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 7, 0, 0, 0, 0, 0, 7, 14, 21, 21, 15, 9, 5, 1, 0, 0, 0, 5, 21, 18, 7, 0, 0, 
    
    -- channel=5
    12, 11, 12, 17, 11, 7, 11, 6, 8, 8, 8, 10, 9, 9, 12, 10, 9, 6, 6, 9, 9, 10, 11, 9, 9, 4, 8, 8, 10, 11, 
    12, 8, 9, 17, 9, 8, 8, 12, 10, 4, 0, 0, 7, 9, 9, 5, 1, 0, 6, 2, 2, 6, 5, 13, 15, 12, 10, 7, 8, 6, 
    7, 4, 5, 10, 9, 9, 9, 12, 13, 19, 0, 0, 5, 5, 1, 7, 5, 26, 8, 0, 0, 0, 0, 0, 7, 11, 11, 7, 7, 8, 
    4, 2, 5, 5, 10, 9, 13, 13, 13, 31, 0, 21, 18, 8, 8, 9, 35, 23, 0, 0, 0, 1, 0, 0, 0, 0, 10, 10, 4, 8, 
    0, 19, 23, 13, 6, 9, 11, 11, 4, 0, 7, 52, 16, 0, 22, 21, 9, 0, 0, 0, 0, 4, 19, 0, 0, 2, 6, 12, 7, 9, 
    0, 21, 23, 7, 6, 11, 12, 7, 7, 0, 4, 25, 6, 3, 5, 0, 0, 0, 0, 0, 0, 17, 12, 0, 18, 5, 0, 5, 6, 9, 
    0, 13, 0, 0, 5, 11, 8, 3, 0, 0, 17, 0, 0, 3, 3, 0, 0, 0, 2, 6, 6, 6, 0, 14, 11, 12, 0, 0, 7, 9, 
    0, 23, 0, 0, 4, 9, 4, 0, 0, 0, 0, 0, 0, 7, 6, 3, 7, 0, 4, 9, 12, 0, 0, 10, 11, 1, 0, 0, 8, 8, 
    21, 0, 0, 0, 10, 6, 35, 0, 0, 0, 0, 0, 5, 16, 8, 0, 0, 16, 5, 0, 0, 3, 0, 0, 0, 3, 1, 0, 0, 7, 
    46, 0, 0, 0, 21, 0, 25, 0, 11, 21, 24, 0, 2, 18, 0, 8, 0, 24, 0, 0, 0, 0, 15, 16, 0, 0, 3, 3, 0, 0, 
    25, 0, 0, 7, 22, 4, 0, 7, 17, 43, 35, 15, 0, 0, 10, 1, 0, 26, 0, 0, 3, 5, 28, 5, 7, 4, 8, 4, 0, 0, 
    32, 0, 0, 21, 31, 14, 0, 3, 0, 22, 32, 0, 0, 1, 2, 5, 0, 17, 0, 0, 14, 21, 24, 0, 0, 7, 11, 1, 3, 0, 
    41, 0, 0, 31, 29, 11, 10, 5, 0, 40, 0, 0, 0, 27, 6, 0, 10, 15, 0, 0, 18, 14, 5, 0, 0, 5, 0, 0, 2, 5, 
    28, 0, 0, 20, 9, 2, 2, 0, 0, 20, 0, 0, 0, 46, 23, 0, 15, 13, 0, 0, 30, 16, 7, 15, 2, 0, 0, 0, 9, 21, 
    12, 0, 8, 3, 7, 0, 3, 4, 0, 9, 0, 0, 34, 16, 14, 26, 22, 0, 0, 17, 9, 3, 10, 13, 5, 0, 0, 8, 30, 9, 
    6, 0, 5, 0, 12, 0, 13, 0, 12, 0, 0, 61, 45, 21, 12, 12, 9, 0, 0, 22, 34, 16, 8, 9, 3, 3, 4, 20, 13, 0, 
    6, 0, 0, 6, 2, 7, 0, 0, 0, 0, 19, 28, 17, 17, 0, 2, 16, 0, 0, 28, 4, 6, 34, 18, 4, 13, 15, 16, 0, 4, 
    13, 0, 0, 15, 6, 0, 0, 21, 0, 0, 32, 0, 11, 4, 0, 0, 4, 3, 29, 0, 0, 33, 26, 16, 0, 0, 0, 0, 0, 11, 
    10, 0, 0, 11, 8, 1, 0, 2, 19, 0, 15, 0, 19, 0, 0, 0, 0, 3, 29, 5, 20, 24, 14, 13, 0, 0, 0, 0, 3, 1, 
    0, 0, 0, 3, 15, 24, 1, 0, 0, 9, 0, 0, 0, 0, 0, 6, 0, 0, 0, 25, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 31, 0, 0, 0, 0, 0, 0, 0, 0, 17, 25, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 17, 16, 0, 0, 29, 0, 5, 2, 0, 20, 31, 31, 31, 29, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 25, 11, 4, 26, 0, 0, 0, 0, 49, 40, 0, 1, 2, 9, 18, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 13, 0, 36, 0, 0, 0, 48, 63, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 26, 0, 0, 9, 75, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 6, 0, 0, 55, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 11, 59, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 24, 59, 10, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 0, 0, 23, 32, 0, 1, 0, 1, 5, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 5, 8, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 
    
    -- channel=6
    52, 55, 56, 51, 53, 52, 52, 52, 52, 51, 48, 47, 53, 60, 60, 60, 55, 51, 49, 52, 52, 53, 53, 51, 52, 49, 48, 53, 55, 53, 
    54, 58, 59, 49, 51, 51, 51, 50, 51, 45, 34, 22, 40, 55, 51, 50, 51, 48, 50, 35, 26, 25, 39, 48, 51, 59, 52, 50, 52, 52, 
    51, 51, 53, 53, 53, 55, 53, 55, 53, 35, 20, 0, 21, 44, 46, 50, 66, 54, 28, 1, 0, 0, 0, 14, 26, 31, 49, 52, 51, 52, 
    44, 49, 53, 56, 56, 58, 57, 56, 57, 42, 60, 42, 40, 52, 65, 68, 42, 26, 9, 0, 0, 0, 0, 0, 5, 18, 43, 52, 49, 44, 
    47, 46, 74, 67, 55, 55, 56, 54, 58, 64, 57, 46, 42, 34, 23, 24, 13, 13, 5, 0, 0, 0, 0, 0, 2, 14, 23, 44, 52, 44, 
    32, 19, 39, 53, 54, 57, 58, 55, 52, 57, 52, 35, 18, 5, 2, 7, 6, 4, 10, 0, 0, 0, 9, 13, 11, 18, 24, 29, 48, 48, 
    0, 0, 7, 8, 39, 55, 51, 43, 39, 32, 34, 11, 0, 0, 5, 14, 15, 11, 15, 26, 3, 0, 13, 21, 21, 11, 16, 25, 44, 51, 
    0, 0, 0, 0, 19, 49, 40, 13, 0, 0, 0, 0, 0, 2, 3, 10, 14, 26, 21, 15, 0, 0, 0, 5, 13, 10, 10, 15, 32, 57, 
    0, 0, 0, 0, 16, 50, 25, 14, 0, 0, 0, 0, 0, 0, 0, 1, 20, 11, 13, 0, 0, 0, 0, 4, 7, 2, 10, 17, 21, 41, 
    0, 0, 0, 0, 7, 48, 33, 37, 24, 0, 0, 0, 0, 0, 4, 0, 11, 1, 2, 0, 0, 0, 0, 9, 14, 6, 0, 6, 10, 24, 
    0, 0, 0, 0, 10, 47, 58, 26, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 9, 14, 7, 5, 0, 16, 
    0, 0, 0, 0, 28, 49, 56, 31, 33, 2, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 4, 13, 14, 17, 10, 0, 0, 10, 
    0, 0, 0, 0, 11, 46, 55, 39, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 27, 40, 33, 20, 0, 0, 0, 0, 0, 0, 10, 7, 0, 4, 0, 0, 0, 11, 11, 11, 2, 0, 9, 13, 23, 
    0, 0, 0, 0, 0, 2, 11, 22, 19, 13, 0, 11, 1, 3, 13, 10, 14, 11, 16, 0, 1, 0, 0, 0, 9, 12, 15, 27, 28, 31, 
    0, 0, 0, 0, 0, 0, 3, 4, 0, 34, 26, 23, 26, 13, 14, 4, 8, 3, 23, 40, 42, 8, 9, 29, 27, 27, 24, 13, 19, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 24, 25, 0, 0, 0, 0, 0, 15, 10, 3, 13, 33, 36, 30, 33, 22, 25, 16, 26, 38, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 16, 0, 8, 11, 22, 35, 18, 19, 4, 20, 26, 37, 44, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 9, 16, 0, 0, 0, 0, 0, 7, 34, 45, 41, 31, 25, 19, 11, 11, 23, 29, 35, 44, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 27, 18, 9, 0, 0, 0, 0, 3, 16, 14, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 14, 13, 11, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=7
    91, 92, 86, 88, 92, 94, 95, 94, 97, 96, 93, 87, 89, 96, 97, 99, 103, 97, 93, 85, 82, 79, 80, 82, 83, 80, 81, 81, 83, 83, 
    92, 95, 87, 89, 93, 97, 96, 96, 100, 108, 98, 91, 95, 100, 102, 102, 91, 92, 88, 87, 81, 74, 73, 66, 75, 74, 82, 86, 88, 87, 
    98, 100, 91, 88, 94, 95, 94, 96, 101, 137, 102, 95, 99, 100, 87, 74, 71, 83, 89, 88, 80, 76, 70, 72, 71, 76, 83, 85, 85, 86, 
    96, 98, 90, 90, 95, 94, 93, 96, 98, 120, 77, 69, 78, 73, 64, 55, 72, 89, 80, 77, 70, 65, 67, 65, 61, 65, 77, 83, 81, 85, 
    69, 83, 85, 90, 98, 97, 96, 98, 100, 105, 78, 82, 77, 74, 78, 67, 78, 88, 77, 70, 63, 59, 64, 58, 52, 55, 71, 78, 72, 78, 
    58, 81, 97, 92, 95, 97, 98, 98, 101, 96, 94, 97, 81, 76, 81, 68, 69, 86, 83, 66, 61, 65, 63, 50, 46, 51, 56, 73, 69, 72, 
    57, 97, 96, 92, 96, 102, 104, 109, 92, 100, 110, 106, 80, 66, 70, 61, 60, 69, 79, 63, 59, 64, 59, 52, 52, 50, 48, 63, 71, 71, 
    67, 112, 92, 78, 96, 104, 129, 140, 118, 112, 124, 91, 69, 58, 64, 57, 50, 57, 82, 71, 69, 66, 62, 64, 59, 57, 46, 52, 71, 71, 
    89, 107, 85, 69, 92, 90, 146, 135, 102, 82, 97, 70, 61, 64, 55, 60, 40, 64, 101, 79, 85, 64, 63, 69, 60, 60, 48, 46, 63, 69, 
    99, 100, 81, 67, 95, 81, 113, 111, 66, 56, 86, 73, 58, 67, 57, 60, 39, 86, 116, 78, 87, 53, 59, 68, 64, 60, 58, 48, 59, 59, 
    102, 94, 78, 66, 90, 78, 82, 107, 61, 44, 85, 85, 65, 74, 71, 74, 39, 112, 111, 67, 74, 51, 61, 66, 64, 58, 61, 51, 57, 50, 
    108, 98, 59, 65, 83, 80, 67, 112, 56, 64, 100, 116, 78, 83, 82, 76, 42, 117, 100, 65, 71, 55, 62, 58, 61, 63, 68, 58, 60, 49, 
    116, 95, 46, 67, 89, 83, 64, 107, 66, 95, 108, 106, 74, 79, 81, 69, 47, 114, 89, 65, 75, 66, 66, 67, 68, 76, 77, 61, 60, 59, 
    116, 88, 51, 66, 96, 88, 74, 110, 87, 132, 119, 90, 82, 75, 70, 59, 50, 102, 83, 66, 68, 61, 51, 60, 67, 71, 70, 53, 61, 68, 
    111, 88, 68, 56, 102, 89, 86, 89, 101, 110, 83, 51, 55, 65, 58, 62, 57, 94, 72, 73, 72, 64, 59, 67, 66, 62, 55, 50, 67, 76, 
    104, 91, 80, 47, 86, 87, 80, 80, 104, 87, 56, 48, 58, 67, 62, 74, 77, 81, 56, 73, 64, 51, 48, 48, 52, 55, 56, 69, 83, 82, 
    97, 91, 85, 54, 75, 90, 76, 73, 94, 62, 68, 62, 75, 94, 68, 81, 89, 75, 73, 97, 69, 42, 38, 54, 50, 61, 62, 74, 79, 79, 
    92, 91, 87, 65, 62, 90, 65, 74, 83, 50, 91, 58, 81, 102, 65, 72, 88, 63, 81, 79, 48, 46, 47, 67, 61, 77, 73, 78, 80, 85, 
    89, 92, 91, 72, 58, 93, 85, 65, 70, 41, 75, 64, 101, 109, 73, 68, 75, 56, 53, 43, 37, 44, 51, 63, 63, 78, 83, 86, 95, 95, 
    87, 95, 95, 71, 49, 96, 112, 91, 87, 92, 110, 106, 127, 111, 82, 75, 79, 55, 57, 52, 60, 65, 71, 73, 76, 85, 92, 93, 101, 101, 
    88, 97, 98, 72, 59, 126, 131, 105, 99, 89, 99, 88, 79, 67, 59, 50, 56, 50, 62, 73, 74, 71, 70, 63, 71, 76, 88, 89, 95, 91, 
    78, 88, 96, 80, 83, 149, 129, 107, 72, 59, 53, 54, 47, 44, 45, 45, 56, 56, 68, 68, 65, 64, 61, 59, 62, 63, 67, 63, 66, 65, 
    64, 82, 85, 66, 95, 138, 116, 89, 57, 54, 66, 61, 56, 56, 55, 55, 57, 54, 60, 61, 58, 59, 58, 61, 60, 62, 63, 61, 61, 62, 
    64, 77, 82, 59, 115, 137, 100, 57, 54, 63, 63, 57, 53, 51, 50, 51, 51, 53, 58, 60, 59, 61, 65, 65, 62, 61, 62, 61, 68, 74, 
    59, 66, 66, 68, 127, 125, 72, 48, 65, 66, 55, 51, 49, 49, 52, 55, 58, 60, 62, 63, 65, 66, 66, 61, 57, 55, 63, 69, 77, 74, 
    58, 61, 60, 69, 126, 101, 52, 66, 75, 62, 57, 49, 50, 52, 52, 54, 57, 59, 61, 59, 61, 61, 59, 55, 55, 62, 76, 76, 64, 55, 
    57, 58, 57, 60, 94, 88, 29, 76, 69, 63, 61, 56, 57, 54, 52, 50, 53, 54, 56, 55, 57, 58, 55, 54, 59, 73, 73, 59, 36, 51, 
    56, 57, 52, 52, 64, 67, 30, 64, 61, 58, 57, 55, 59, 55, 57, 57, 58, 58, 56, 54, 54, 53, 54, 62, 72, 79, 67, 54, 40, 63, 
    50, 56, 49, 49, 53, 61, 46, 64, 58, 59, 53, 51, 51, 49, 55, 56, 59, 63, 62, 58, 55, 53, 61, 74, 83, 77, 61, 51, 46, 51, 
    49, 54, 48, 48, 49, 55, 53, 54, 54, 56, 49, 52, 49, 46, 48, 50, 57, 65, 60, 54, 56, 54, 67, 73, 79, 66, 50, 44, 50, 45, 
    
    -- channel=8
    451, 464, 459, 450, 460, 466, 465, 464, 463, 450, 441, 450, 476, 504, 507, 499, 476, 443, 406, 372, 355, 352, 367, 375, 381, 392, 404, 415, 408, 388, 
    461, 477, 472, 462, 468, 473, 471, 470, 461, 435, 426, 434, 460, 489, 484, 463, 427, 368, 325, 278, 259, 260, 281, 309, 333, 360, 389, 409, 408, 392, 
    458, 472, 475, 473, 477, 480, 477, 476, 469, 433, 416, 384, 414, 436, 419, 387, 333, 280, 230, 174, 143, 139, 175, 200, 255, 303, 351, 383, 396, 390, 
    421, 426, 450, 470, 485, 488, 484, 484, 485, 484, 433, 352, 359, 363, 321, 279, 244, 209, 166, 119, 93, 80, 88, 118, 160, 214, 288, 341, 371, 381, 
    350, 343, 402, 453, 482, 492, 488, 491, 493, 487, 457, 354, 302, 264, 225, 188, 162, 161, 149, 122, 107, 93, 98, 104, 104, 140, 215, 292, 345, 365, 
    232, 230, 338, 421, 470, 496, 494, 484, 471, 437, 388, 320, 250, 177, 141, 126, 121, 147, 160, 141, 126, 126, 133, 119, 100, 94, 145, 238, 320, 356, 
    132, 109, 252, 365, 446, 488, 482, 452, 420, 362, 319, 275, 210, 146, 121, 114, 106, 144, 184, 175, 142, 141, 149, 136, 105, 91, 108, 186, 286, 343, 
    73, 73, 190, 297, 407, 465, 432, 387, 309, 260, 243, 230, 176, 132, 117, 121, 111, 122, 180, 207, 157, 132, 136, 134, 112, 88, 90, 144, 244, 317, 
    50, 70, 172, 260, 371, 437, 395, 340, 231, 158, 175, 196, 157, 125, 116, 106, 107, 109, 157, 195, 158, 132, 111, 117, 121, 100, 84, 95, 181, 278, 
    67, 86, 158, 245, 355, 411, 396, 332, 243, 158, 174, 186, 153, 136, 120, 110, 97, 97, 167, 182, 147, 135, 108, 122, 120, 107, 88, 75, 109, 214, 
    51, 104, 158, 227, 345, 406, 366, 328, 272, 181, 194, 213, 170, 141, 140, 113, 90, 96, 190, 178, 140, 132, 107, 121, 131, 113, 90, 71, 78, 157, 
    36, 109, 152, 203, 333, 414, 358, 302, 277, 190, 229, 242, 196, 139, 145, 135, 87, 100, 194, 176, 132, 122, 105, 112, 125, 120, 105, 86, 89, 149, 
    42, 117, 115, 157, 299, 399, 369, 307, 275, 203, 226, 236, 199, 141, 138, 144, 103, 109, 186, 159, 116, 108, 99, 96, 110, 117, 112, 104, 121, 179, 
    57, 128, 90, 95, 215, 337, 338, 295, 271, 217, 218, 193, 165, 160, 150, 138, 118, 143, 199, 161, 130, 113, 96, 93, 102, 114, 133, 145, 172, 247, 
    60, 117, 85, 61, 121, 239, 265, 275, 249, 252, 234, 155, 137, 158, 160, 155, 146, 177, 244, 203, 148, 124, 111, 106, 116, 125, 154, 189, 241, 310, 
    57, 94, 83, 46, 70, 158, 203, 216, 243, 263, 231, 199, 160, 161, 159, 143, 152, 214, 259, 231, 195, 137, 102, 105, 122, 136, 170, 223, 293, 346, 
    58, 74, 83, 48, 36, 109, 154, 158, 190, 224, 186, 196, 177, 169, 151, 121, 156, 201, 225, 244, 223, 149, 120, 110, 137, 176, 231, 292, 356, 390, 
    89, 76, 85, 61, 28, 75, 136, 125, 128, 155, 160, 186, 161, 165, 130, 93, 146, 189, 172, 170, 160, 135, 104, 92, 135, 197, 294, 346, 385, 404, 
    132, 100, 102, 85, 40, 47, 94, 110, 107, 94, 132, 166, 153, 175, 120, 65, 124, 184, 186, 152, 103, 90, 73, 75, 125, 203, 321, 367, 380, 385, 
    155, 115, 121, 108, 58, 43, 84, 59, 59, 67, 83, 111, 118, 134, 100, 51, 62, 125, 139, 115, 61, 26, 18, 19, 64, 122, 198, 223, 225, 217, 
    126, 96, 115, 107, 60, 63, 142, 98, 11, 15, 32, 54, 71, 87, 67, 37, 18, 22, 26, 12, 0, 0, 0, 0, 0, 0, 40, 53, 42, 38, 
    55, 54, 83, 86, 52, 86, 172, 161, 97, 9, 3, 35, 40, 46, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 49, 76, 66, 131, 186, 155, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 21, 50, 86, 171, 189, 110, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 73, 161, 149, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 46, 129, 82, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 83, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 2, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 12, 0, 0, 0, 0, 6, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 7, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 4, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 30, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 8, 0, 8, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 23, 0, 0, 15, 14, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 25, 0, 0, 8, 15, 0, 0, 0, 0, 0, 2, 8, 0, 0, 14, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 0, 0, 13, 4, 0, 0, 0, 0, 1, 3, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 38, 38, 0, 21, 0, 29, 10, 0, 25, 9, 0, 0, 0, 0, 3, 7, 14, 0, 13, 8, 0, 0, 0, 0, 
    22, 0, 0, 0, 0, 0, 24, 62, 36, 16, 0, 3, 0, 0, 2, 1, 0, 5, 8, 10, 19, 30, 20, 21, 16, 17, 20, 18, 10, 15, 
    29, 10, 1, 10, 18, 0, 0, 10, 7, 0, 0, 0, 0, 0, 0, 0, 2, 26, 21, 21, 22, 20, 21, 24, 21, 23, 23, 27, 24, 23, 
    11, 12, 14, 6, 9, 0, 6, 0, 0, 0, 0, 0, 0, 0, 4, 12, 12, 20, 16, 20, 24, 21, 23, 28, 28, 25, 27, 32, 25, 30, 
    5, 5, 9, 6, 4, 0, 0, 0, 0, 2, 16, 22, 20, 20, 16, 15, 18, 21, 21, 23, 28, 29, 31, 32, 32, 30, 30, 31, 34, 45, 
    27, 4, 1, 28, 8, 8, 0, 0, 0, 9, 21, 19, 18, 19, 20, 20, 22, 25, 26, 28, 34, 35, 33, 26, 26, 27, 27, 40, 46, 39, 
    36, 25, 8, 19, 2, 18, 0, 0, 0, 13, 20, 21, 18, 19, 23, 23, 25, 25, 28, 28, 26, 32, 28, 26, 23, 28, 38, 44, 25, 16, 
    37, 37, 30, 5, 0, 13, 26, 0, 6, 15, 24, 29, 23, 20, 19, 20, 22, 25, 26, 25, 22, 24, 27, 29, 33, 43, 36, 22, 10, 17, 
    31, 34, 37, 23, 0, 0, 28, 0, 4, 16, 18, 29, 29, 24, 22, 24, 24, 25, 22, 27, 24, 21, 25, 35, 47, 40, 29, 29, 27, 19, 
    29, 30, 33, 33, 9, 0, 36, 2, 8, 13, 12, 15, 17, 23, 25, 26, 25, 29, 31, 25, 21, 24, 30, 38, 45, 37, 37, 30, 38, 15, 
    31, 23, 30, 29, 32, 14, 25, 20, 17, 16, 16, 13, 12, 10, 10, 14, 22, 28, 29, 23, 23, 25, 25, 29, 29, 32, 24, 21, 36, 22, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    119, 122, 120, 113, 117, 121, 121, 116, 117, 120, 120, 120, 123, 122, 118, 117, 118, 123, 120, 113, 104, 98, 100, 96, 95, 93, 88, 83, 79, 71, 
    110, 116, 115, 113, 119, 124, 125, 119, 119, 119, 132, 136, 126, 119, 121, 123, 128, 114, 105, 102, 97, 94, 88, 90, 89, 85, 88, 88, 84, 76, 
    106, 118, 117, 116, 120, 127, 125, 122, 126, 137, 171, 167, 135, 126, 131, 128, 97, 79, 94, 99, 91, 81, 80, 73, 80, 87, 88, 91, 91, 82, 
    115, 122, 122, 122, 124, 126, 123, 121, 133, 201, 201, 158, 134, 125, 98, 76, 59, 81, 111, 128, 115, 98, 74, 62, 71, 69, 74, 86, 94, 88, 
    123, 109, 99, 116, 127, 122, 119, 121, 131, 207, 194, 147, 116, 95, 64, 42, 54, 91, 136, 166, 153, 121, 94, 95, 63, 48, 58, 74, 86, 89, 
    92, 70, 85, 119, 129, 122, 118, 121, 127, 144, 132, 120, 106, 72, 53, 49, 72, 111, 153, 176, 160, 124, 118, 101, 65, 26, 28, 60, 80, 90, 
    71, 27, 82, 135, 133, 124, 128, 127, 141, 121, 115, 146, 145, 107, 85, 71, 74, 119, 158, 164, 146, 127, 113, 85, 62, 27, 14, 36, 62, 87, 
    100, 80, 120, 149, 139, 129, 131, 161, 175, 166, 167, 190, 171, 123, 95, 85, 73, 79, 128, 167, 151, 124, 100, 81, 59, 37, 11, 23, 49, 73, 
    140, 162, 189, 175, 144, 137, 159, 237, 249, 221, 205, 209, 182, 121, 97, 77, 59, 38, 95, 175, 180, 143, 101, 77, 76, 62, 21, 0, 31, 63, 
    199, 216, 229, 194, 153, 127, 211, 281, 307, 266, 236, 212, 191, 145, 99, 79, 47, 29, 122, 213, 221, 168, 109, 89, 85, 83, 49, 5, 9, 44, 
    218, 230, 253, 201, 158, 114, 173, 235, 279, 254, 225, 223, 213, 179, 118, 96, 51, 63, 190, 251, 241, 163, 105, 98, 96, 91, 66, 29, 14, 26, 
    201, 236, 271, 198, 150, 124, 106, 166, 207, 203, 224, 272, 255, 206, 157, 129, 64, 107, 230, 265, 230, 146, 97, 85, 93, 87, 86, 65, 47, 25, 
    205, 250, 250, 182, 143, 135, 101, 139, 152, 171, 240, 317, 289, 215, 178, 167, 93, 136, 230, 259, 203, 136, 105, 81, 83, 96, 108, 97, 82, 40, 
    233, 270, 226, 165, 131, 140, 112, 126, 139, 204, 275, 346, 291, 226, 192, 155, 96, 153, 226, 233, 201, 146, 98, 73, 77, 108, 128, 115, 84, 62, 
    259, 275, 240, 173, 133, 147, 129, 143, 134, 239, 320, 282, 225, 190, 169, 139, 98, 141, 209, 216, 187, 149, 109, 92, 95, 117, 129, 98, 72, 81, 
    281, 284, 274, 194, 160, 146, 151, 150, 159, 245, 286, 227, 179, 140, 136, 123, 97, 156, 191, 171, 156, 143, 86, 64, 79, 91, 98, 81, 91, 103, 
    296, 299, 302, 217, 177, 162, 171, 139, 174, 180, 155, 155, 136, 130, 138, 125, 112, 152, 141, 163, 174, 118, 62, 37, 50, 68, 73, 91, 113, 112, 
    308, 305, 308, 240, 176, 174, 187, 166, 153, 133, 113, 122, 119, 147, 155, 142, 139, 135, 110, 133, 124, 64, 22, 10, 30, 71, 93, 116, 119, 116, 
    307, 307, 303, 261, 186, 170, 181, 215, 179, 91, 107, 113, 144, 218, 202, 150, 151, 146, 144, 107, 51, 26, 0, 28, 42, 92, 128, 139, 130, 124, 
    302, 306, 299, 275, 197, 162, 186, 227, 228, 139, 134, 145, 219, 282, 258, 181, 142, 134, 119, 69, 29, 14, 24, 67, 85, 132, 155, 152, 148, 137, 
    301, 309, 304, 275, 193, 183, 288, 312, 260, 215, 194, 206, 266, 290, 274, 209, 138, 88, 54, 42, 45, 44, 64, 81, 109, 140, 163, 162, 154, 144, 
    283, 296, 303, 269, 196, 241, 376, 435, 389, 283, 220, 228, 242, 243, 230, 182, 142, 101, 77, 68, 82, 99, 110, 112, 125, 134, 145, 139, 132, 127, 
    254, 267, 287, 282, 229, 310, 414, 464, 385, 238, 171, 154, 149, 145, 144, 124, 108, 101, 102, 102, 108, 113, 118, 121, 127, 135, 139, 136, 135, 126, 
    190, 229, 265, 259, 262, 367, 447, 416, 257, 148, 111, 99, 97, 90, 93, 94, 92, 91, 98, 104, 109, 114, 117, 131, 138, 140, 140, 140, 136, 141, 
    131, 166, 216, 203, 269, 394, 442, 311, 177, 119, 109, 111, 103, 96, 96, 96, 94, 93, 100, 107, 113, 124, 138, 150, 149, 149, 146, 146, 161, 185, 
    128, 125, 155, 183, 279, 397, 387, 233, 145, 118, 114, 112, 105, 96, 94, 94, 97, 102, 108, 121, 129, 137, 148, 151, 148, 140, 149, 176, 203, 201, 
    132, 116, 115, 157, 274, 357, 312, 201, 131, 119, 120, 115, 108, 104, 102, 99, 102, 107, 118, 125, 133, 145, 146, 135, 126, 129, 169, 196, 184, 155, 
    140, 120, 113, 122, 216, 293, 231, 167, 127, 111, 118, 120, 117, 110, 104, 103, 112, 119, 126, 126, 125, 128, 125, 121, 128, 162, 188, 180, 137, 118, 
    138, 121, 117, 112, 134, 196, 157, 129, 102, 100, 114, 121, 121, 109, 106, 108, 118, 125, 133, 137, 126, 115, 111, 128, 162, 202, 199, 164, 96, 100, 
    136, 124, 115, 113, 106, 116, 107, 93, 75, 76, 86, 96, 106, 104, 104, 111, 126, 141, 151, 142, 122, 111, 116, 151, 203, 226, 207, 154, 98, 90, 
    
    -- channel=12
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 13, 11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 23, 16, 5, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 19, 17, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 1, 0, 0, 0, 0, 0, 5, 12, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 0, 13, 18, 5, 14, 14, 9, 2, 0, 0, 0, 0, 9, 11, 9, 3, 0, 0, 0, 0, 0, 0, 0, 
    16, 19, 0, 0, 0, 0, 0, 9, 23, 23, 16, 26, 25, 9, 7, 0, 0, 0, 0, 18, 19, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 28, 14, 0, 0, 0, 0, 14, 39, 39, 30, 26, 31, 12, 2, 1, 0, 0, 0, 27, 27, 17, 2, 0, 0, 0, 0, 0, 0, 0, 
    39, 35, 25, 0, 0, 0, 0, 20, 35, 32, 16, 22, 32, 22, 5, 3, 0, 0, 7, 31, 35, 18, 5, 0, 0, 0, 0, 0, 0, 0, 
    36, 42, 39, 0, 0, 0, 0, 0, 10, 16, 24, 29, 37, 28, 13, 6, 0, 0, 20, 41, 37, 17, 2, 0, 0, 0, 2, 0, 0, 0, 
    34, 41, 46, 6, 0, 0, 0, 0, 0, 2, 26, 42, 37, 22, 17, 21, 3, 0, 24, 42, 30, 18, 10, 0, 0, 1, 4, 0, 0, 0, 
    41, 45, 47, 23, 0, 0, 0, 0, 0, 10, 41, 74, 53, 31, 16, 11, 4, 6, 20, 35, 32, 11, 0, 0, 0, 0, 1, 0, 0, 0, 
    49, 48, 52, 38, 0, 0, 0, 0, 0, 17, 33, 34, 33, 16, 15, 8, 0, 0, 14, 22, 23, 21, 13, 2, 0, 0, 0, 0, 0, 0, 
    61, 54, 56, 45, 17, 0, 2, 1, 0, 16, 36, 27, 15, 3, 11, 2, 0, 0, 0, 0, 3, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    67, 63, 63, 52, 37, 10, 7, 3, 14, 8, 4, 15, 6, 6, 20, 7, 0, 0, 7, 18, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    67, 64, 64, 53, 39, 20, 19, 11, 12, 15, 0, 0, 0, 4, 27, 21, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    61, 61, 58, 55, 42, 28, 32, 48, 16, 0, 0, 0, 7, 28, 34, 28, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    56, 55, 53, 56, 39, 18, 26, 59, 68, 31, 24, 26, 40, 47, 52, 39, 17, 15, 13, 5, 0, 0, 5, 13, 0, 0, 0, 0, 0, 0, 
    58, 58, 56, 58, 42, 27, 49, 56, 58, 55, 30, 26, 41, 44, 50, 40, 13, 5, 12, 13, 12, 10, 16, 24, 28, 34, 40, 42, 43, 42, 
    51, 56, 60, 58, 41, 36, 65, 86, 87, 55, 42, 47, 53, 54, 57, 53, 40, 29, 26, 22, 27, 34, 40, 43, 50, 52, 51, 50, 53, 52, 
    59, 47, 54, 57, 28, 43, 76, 104, 98, 71, 57, 53, 54, 51, 55, 51, 41, 39, 41, 40, 43, 45, 49, 52, 54, 56, 55, 55, 55, 52, 
    67, 57, 50, 51, 40, 61, 93, 103, 77, 56, 42, 38, 38, 33, 35, 36, 35, 37, 42, 45, 47, 49, 50, 55, 53, 54, 56, 58, 58, 63, 
    56, 51, 49, 35, 41, 72, 104, 87, 65, 46, 43, 43, 40, 37, 38, 39, 39, 39, 42, 47, 49, 54, 57, 57, 54, 56, 57, 62, 67, 70, 
    59, 50, 50, 42, 40, 77, 101, 73, 54, 43, 41, 44, 43, 37, 37, 38, 41, 43, 46, 53, 53, 53, 58, 61, 62, 61, 67, 73, 72, 64, 
    63, 55, 49, 50, 53, 63, 86, 59, 44, 41, 45, 45, 44, 43, 40, 40, 42, 46, 50, 55, 59, 61, 60, 58, 60, 65, 75, 74, 67, 56, 
    67, 58, 54, 50, 61, 64, 60, 54, 41, 35, 39, 41, 43, 43, 42, 45, 50, 52, 53, 56, 56, 55, 54, 54, 61, 73, 80, 80, 67, 49, 
    65, 58, 56, 51, 50, 61, 53, 49, 40, 38, 41, 40, 39, 36, 37, 39, 45, 50, 57, 59, 54, 50, 49, 52, 63, 80, 84, 73, 49, 46, 
    62, 57, 53, 51, 44, 41, 41, 38, 34, 32, 36, 39, 43, 36, 31, 34, 41, 47, 52, 52, 49, 46, 43, 51, 64, 76, 80, 67, 49, 45, 
    
    -- channel=13
    19, 24, 31, 36, 32, 32, 33, 29, 25, 31, 37, 40, 34, 23, 21, 17, 17, 11, 8, 0, 0, 0, 0, 8, 17, 15, 7, 0, 0, 0, 
    10, 19, 27, 36, 35, 38, 37, 33, 36, 70, 80, 71, 45, 24, 29, 34, 16, 12, 0, 5, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    18, 29, 34, 37, 36, 35, 36, 31, 41, 129, 157, 157, 76, 35, 26, 4, 0, 0, 27, 67, 69, 54, 12, 0, 0, 0, 0, 0, 0, 0, 
    22, 32, 32, 34, 30, 29, 28, 25, 29, 86, 125, 132, 51, 0, 0, 0, 0, 9, 77, 126, 128, 106, 81, 44, 3, 0, 0, 0, 3, 2, 
    0, 0, 0, 10, 31, 30, 29, 26, 26, 53, 41, 57, 34, 0, 0, 0, 0, 49, 117, 158, 142, 114, 93, 71, 34, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 29, 27, 29, 32, 26, 24, 28, 53, 66, 53, 30, 14, 22, 59, 125, 174, 151, 100, 75, 64, 19, 0, 0, 0, 0, 9, 
    57, 34, 10, 43, 41, 29, 37, 63, 45, 46, 55, 106, 131, 98, 55, 28, 28, 32, 80, 134, 147, 98, 51, 31, 14, 0, 0, 0, 0, 0, 
    157, 135, 123, 126, 70, 32, 92, 175, 226, 200, 175, 172, 175, 117, 66, 23, 5, 6, 45, 96, 152, 126, 66, 32, 19, 11, 0, 0, 0, 0, 
    229, 215, 211, 172, 97, 21, 117, 243, 361, 343, 285, 221, 198, 141, 76, 44, 0, 0, 64, 139, 205, 156, 104, 60, 36, 34, 0, 0, 0, 0, 
    239, 232, 258, 202, 122, 35, 69, 189, 305, 334, 298, 259, 230, 169, 102, 60, 0, 18, 112, 211, 260, 165, 104, 52, 54, 53, 26, 0, 0, 0, 
    247, 217, 255, 219, 137, 58, 53, 116, 183, 248, 254, 264, 272, 222, 129, 102, 30, 74, 148, 252, 258, 147, 84, 42, 41, 48, 46, 18, 2, 0, 
    259, 228, 240, 196, 107, 61, 37, 92, 113, 205, 219, 287, 309, 277, 178, 128, 70, 122, 177, 253, 234, 127, 66, 28, 23, 35, 54, 52, 42, 0, 
    280, 254, 251, 170, 72, 51, 26, 60, 67, 184, 244, 302, 287, 265, 208, 151, 82, 130, 180, 246, 228, 143, 88, 54, 40, 56, 83, 84, 60, 14, 
    308, 275, 269, 181, 92, 54, 47, 66, 68, 217, 321, 353, 288, 200, 171, 141, 85, 114, 162, 227, 202, 132, 73, 46, 50, 81, 97, 79, 54, 10, 
    335, 304, 305, 216, 149, 85, 97, 63, 91, 175, 275, 303, 226, 148, 113, 92, 68, 114, 132, 190, 191, 144, 73, 39, 37, 63, 70, 48, 32, 17, 
    362, 330, 336, 254, 179, 125, 135, 113, 91, 113, 167, 143, 121, 99, 70, 80, 82, 89, 68, 98, 107, 110, 59, 1, 0, 22, 39, 41, 41, 41, 
    381, 351, 348, 282, 207, 147, 158, 166, 132, 66, 88, 79, 102, 116, 93, 95, 91, 111, 95, 57, 41, 44, 0, 0, 0, 0, 25, 53, 52, 41, 
    367, 355, 346, 298, 221, 170, 139, 179, 179, 89, 82, 56, 127, 170, 170, 137, 97, 92, 126, 104, 44, 0, 0, 0, 0, 43, 52, 74, 61, 39, 
    332, 348, 337, 304, 235, 201, 191, 190, 168, 90, 72, 63, 156, 227, 256, 205, 109, 49, 44, 25, 0, 0, 0, 0, 7, 62, 69, 69, 52, 31, 
    297, 349, 331, 294, 219, 206, 261, 351, 316, 199, 169, 186, 265, 331, 333, 271, 189, 72, 6, 0, 0, 0, 0, 21, 40, 64, 77, 70, 56, 40, 
    283, 358, 337, 295, 228, 248, 325, 457, 485, 362, 267, 240, 267, 285, 270, 217, 157, 88, 38, 9, 16, 36, 69, 82, 82, 86, 87, 79, 76, 59, 
    236, 324, 343, 320, 286, 338, 415, 504, 435, 333, 200, 131, 127, 124, 120, 104, 87, 59, 56, 62, 73, 79, 89, 100, 106, 107, 111, 111, 110, 101, 
    138, 218, 288, 293, 313, 378, 458, 471, 359, 204, 107, 80, 74, 74, 71, 64, 66, 60, 61, 67, 79, 89, 95, 111, 124, 133, 132, 128, 128, 127, 
    116, 126, 194, 237, 309, 387, 452, 389, 247, 120, 93, 89, 88, 82, 77, 70, 65, 65, 67, 76, 88, 99, 116, 135, 149, 154, 151, 148, 160, 173, 
    129, 109, 117, 167, 297, 409, 426, 316, 163, 96, 103, 99, 93, 83, 77, 72, 71, 73, 82, 95, 112, 130, 141, 145, 142, 134, 143, 164, 194, 213, 
    134, 109, 100, 116, 260, 382, 387, 269, 139, 99, 109, 103, 92, 79, 78, 82, 86, 91, 102, 107, 117, 131, 142, 139, 121, 119, 144, 177, 197, 193, 
    136, 113, 107, 111, 176, 283, 278, 225, 113, 105, 113, 114, 115, 96, 85, 80, 88, 99, 109, 116, 118, 116, 117, 119, 121, 139, 161, 177, 143, 123, 
    148, 122, 112, 115, 124, 143, 139, 130, 64, 67, 88, 106, 120, 116, 109, 104, 109, 117, 122, 118, 113, 106, 103, 116, 149, 187, 206, 182, 113, 87, 
    153, 125, 114, 116, 111, 99, 64, 64, 42, 35, 45, 60, 73, 85, 99, 112, 131, 148, 154, 143, 123, 103, 107, 139, 201, 246, 239, 182, 120, 77, 
    149, 128, 110, 112, 99, 90, 65, 47, 36, 30, 31, 40, 33, 31, 42, 65, 101, 139, 160, 155, 130, 103, 117, 154, 218, 252, 233, 167, 105, 71, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 5, 12, 19, 19, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 10, 10, 0, 0, 0, 0, 13, 21, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 15, 0, 0, 10, 18, 18, 20, 40, 30, 12, 0, 0, 0, 0, 0, 11, 22, 1, 0, 0, 
    1, 12, 9, 0, 0, 0, 0, 0, 0, 70, 64, 0, 0, 0, 12, 0, 12, 59, 52, 27, 19, 14, 4, 0, 0, 0, 30, 34, 0, 0, 
    0, 13, 46, 0, 0, 0, 0, 0, 0, 0, 12, 4, 0, 0, 0, 0, 9, 69, 73, 22, 6, 21, 37, 17, 0, 0, 16, 53, 21, 0, 
    0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 14, 10, 69, 112, 50, 0, 5, 41, 25, 1, 0, 0, 47, 45, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 7, 32, 21, 48, 115, 88, 0, 0, 5, 21, 2, 0, 0, 18, 64, 25, 
    0, 20, 12, 0, 0, 0, 38, 52, 0, 0, 0, 32, 0, 0, 0, 14, 16, 23, 87, 71, 1, 0, 0, 8, 9, 0, 0, 0, 48, 60, 
    7, 77, 24, 0, 0, 0, 105, 193, 88, 0, 22, 30, 0, 0, 0, 0, 0, 20, 100, 44, 0, 0, 0, 22, 19, 0, 0, 0, 0, 46, 
    35, 123, 47, 0, 0, 0, 59, 209, 164, 34, 57, 57, 0, 0, 0, 0, 0, 30, 142, 49, 4, 0, 0, 37, 38, 11, 0, 0, 0, 0, 
    24, 130, 58, 0, 0, 0, 0, 119, 140, 41, 69, 90, 0, 0, 0, 0, 0, 47, 161, 54, 0, 0, 0, 30, 48, 34, 16, 0, 0, 0, 
    17, 125, 27, 0, 2, 0, 0, 64, 102, 39, 56, 92, 34, 0, 0, 11, 0, 75, 148, 45, 0, 0, 0, 12, 28, 33, 26, 0, 0, 0, 
    28, 122, 0, 0, 7, 3, 0, 14, 69, 81, 62, 42, 41, 34, 23, 10, 0, 85, 144, 47, 0, 0, 0, 14, 23, 31, 32, 0, 0, 0, 
    33, 105, 3, 0, 0, 26, 0, 0, 54, 135, 116, 17, 8, 54, 58, 26, 0, 64, 121, 58, 10, 0, 0, 33, 56, 49, 39, 6, 0, 0, 
    32, 93, 37, 0, 0, 56, 0, 0, 49, 159, 160, 78, 33, 42, 44, 29, 1, 41, 81, 85, 47, 0, 0, 29, 69, 63, 32, 0, 0, 0, 
    32, 87, 70, 0, 0, 80, 42, 0, 6, 88, 89, 64, 14, 20, 13, 14, 25, 17, 2, 64, 84, 24, 9, 36, 51, 49, 14, 0, 0, 0, 
    45, 77, 80, 0, 0, 72, 92, 0, 0, 0, 44, 50, 5, 27, 0, 0, 64, 26, 0, 0, 30, 19, 10, 22, 10, 11, 7, 0, 0, 0, 
    63, 66, 79, 22, 0, 41, 90, 39, 4, 0, 38, 65, 43, 63, 0, 0, 40, 70, 50, 28, 0, 12, 20, 46, 19, 7, 3, 0, 0, 0, 
    81, 49, 73, 42, 0, 37, 84, 0, 0, 0, 7, 25, 48, 64, 0, 0, 0, 28, 60, 51, 20, 6, 17, 53, 56, 53, 29, 0, 1, 4, 
    103, 37, 65, 40, 0, 53, 138, 7, 0, 0, 0, 44, 95, 101, 66, 8, 0, 0, 0, 4, 15, 9, 18, 31, 54, 67, 55, 32, 31, 36, 
    148, 66, 67, 26, 0, 55, 150, 94, 6, 0, 56, 141, 166, 163, 149, 98, 64, 32, 13, 14, 31, 53, 63, 62, 69, 75, 75, 60, 56, 59, 
    192, 145, 108, 46, 4, 106, 136, 96, 66, 41, 76, 108, 112, 108, 107, 84, 65, 60, 64, 67, 66, 71, 77, 78, 72, 73, 81, 72, 70, 70, 
    140, 178, 170, 87, 76, 153, 126, 63, 23, 32, 48, 52, 52, 50, 56, 61, 62, 63, 69, 77, 74, 72, 73, 76, 70, 66, 71, 69, 66, 65, 
    60, 126, 177, 113, 122, 159, 93, 5, 21, 60, 61, 63, 62, 63, 63, 61, 60, 60, 64, 70, 69, 67, 72, 80, 81, 82, 86, 79, 71, 73, 
    53, 77, 123, 138, 193, 182, 40, 0, 23, 65, 70, 63, 60, 65, 64, 60, 59, 62, 67, 74, 80, 83, 85, 84, 88, 94, 101, 96, 93, 102, 
    62, 68, 77, 121, 234, 230, 34, 0, 39, 62, 72, 58, 46, 56, 66, 70, 73, 73, 76, 79, 86, 99, 97, 82, 77, 83, 102, 109, 103, 113, 
    61, 76, 78, 85, 186, 245, 89, 20, 70, 77, 86, 72, 52, 46, 54, 65, 72, 73, 77, 76, 75, 85, 90, 85, 74, 83, 93, 87, 65, 93, 
    55, 79, 86, 74, 96, 162, 101, 50, 68, 90, 102, 98, 89, 69, 61, 63, 64, 64, 61, 61, 65, 71, 78, 85, 85, 83, 64, 48, 29, 74, 
    53, 76, 87, 78, 63, 71, 69, 51, 48, 71, 83, 89, 97, 93, 96, 99, 92, 82, 65, 49, 52, 60, 77, 101, 112, 93, 61, 49, 48, 63, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 0, 5, 20, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 88, 103, 63, 55, 45, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    58, 50, 14, 0, 0, 0, 0, 0, 0, 111, 110, 49, 27, 2, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 7, 3, 0, 0, 
    56, 36, 0, 0, 2, 0, 0, 0, 0, 56, 34, 0, 0, 0, 0, 0, 0, 0, 20, 41, 47, 48, 45, 30, 17, 15, 18, 1, 0, 0, 
    13, 0, 0, 18, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 16, 26, 29, 37, 34, 22, 10, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 15, 18, 15, 23, 27, 27, 25, 17, 
    0, 0, 9, 1, 0, 0, 0, 3, 4, 3, 14, 8, 20, 41, 36, 23, 16, 47, 54, 28, 30, 52, 66, 62, 50, 46, 36, 22, 14, 7, 
    0, 44, 47, 41, 42, 44, 42, 41, 38, 33, 34, 32, 47, 52, 40, 28, 31, 59, 57, 41, 51, 65, 66, 56, 44, 38, 31, 20, 12, 5, 
    90, 91, 87, 84, 85, 84, 79, 73, 64, 58, 53, 53, 59, 58, 50, 45, 54, 68, 70, 69, 72, 71, 68, 60, 50, 45, 36, 20, 5, 0, 
    117, 89, 88, 102, 112, 114, 111, 106, 102, 99, 94, 92, 97, 99, 94, 88, 93, 100, 102, 98, 90, 81, 72, 58, 38, 27, 23, 9, 0, 0, 
    113, 76, 46, 70, 97, 107, 110, 113, 113, 113, 102, 78, 95, 110, 108, 102, 106, 111, 103, 90, 76, 58, 37, 18, 7, 12, 22, 14, 0, 0, 
    114, 89, 44, 45, 83, 100, 110, 117, 115, 113, 99, 20, 2, 54, 64, 61, 64, 62, 52, 38, 21, 10, 5, 8, 19, 32, 32, 5, 0, 0, 
    118, 105, 73, 64, 93, 113, 120, 124, 119, 112, 104, 14, 0, 0, 22, 16, 11, 10, 10, 13, 15, 22, 36, 51, 47, 26, 6, 0, 0, 0, 
    125, 113, 95, 93, 104, 118, 124, 123, 116, 110, 108, 46, 0, 0, 37, 41, 37, 43, 55, 67, 77, 77, 63, 42, 15, 0, 0, 0, 0, 0, 
    137, 121, 107, 105, 107, 115, 121, 117, 112, 109, 110, 81, 7, 3, 66, 89, 97, 108, 112, 105, 86, 52, 17, 0, 2, 0, 0, 0, 0, 0, 
    143, 132, 109, 109, 108, 113, 116, 113, 111, 110, 109, 98, 38, 24, 91, 130, 134, 122, 95, 60, 26, 3, 0, 3, 11, 0, 0, 0, 0, 0, 
    141, 131, 106, 105, 106, 108, 109, 109, 109, 109, 108, 103, 66, 55, 111, 144, 118, 69, 23, 0, 0, 2, 10, 8, 0, 0, 0, 0, 0, 0, 
    127, 107, 94, 93, 94, 96, 98, 98, 98, 98, 96, 93, 73, 64, 88, 85, 43, 5, 0, 0, 8, 18, 13, 1, 0, 0, 0, 0, 0, 0, 
    96, 76, 72, 74, 74, 74, 74, 73, 72, 71, 67, 60, 46, 32, 27, 15, 1, 0, 0, 7, 21, 18, 4, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=17
    250, 248, 248, 248, 248, 248, 248, 248, 248, 248, 249, 249, 249, 249, 247, 245, 245, 248, 252, 254, 252, 251, 248, 248, 248, 249, 248, 248, 248, 249, 
    254, 252, 252, 252, 252, 252, 252, 252, 251, 252, 252, 252, 252, 252, 250, 248, 248, 252, 256, 264, 254, 256, 250, 250, 252, 252, 251, 251, 252, 253, 
    253, 250, 250, 250, 250, 250, 250, 251, 250, 250, 251, 251, 250, 250, 250, 250, 252, 259, 265, 269, 257, 257, 252, 250, 250, 251, 251, 250, 251, 252, 
    254, 251, 251, 251, 251, 251, 252, 251, 250, 250, 250, 251, 252, 251, 255, 258, 260, 265, 273, 255, 236, 238, 234, 247, 251, 250, 251, 250, 251, 252, 
    251, 248, 249, 249, 250, 251, 251, 251, 249, 249, 252, 254, 254, 254, 263, 273, 284, 285, 280, 249, 225, 239, 240, 246, 253, 251, 251, 252, 253, 252, 
    256, 254, 254, 253, 251, 251, 251, 249, 247, 249, 252, 261, 252, 256, 272, 272, 269, 269, 264, 248, 240, 248, 254, 253, 258, 255, 255, 255, 256, 254, 
    264, 261, 261, 258, 256, 254, 250, 249, 249, 250, 254, 260, 245, 251, 267, 263, 242, 236, 244, 235, 222, 214, 226, 255, 268, 263, 262, 261, 259, 256, 
    262, 268, 267, 258, 251, 254, 250, 250, 252, 253, 259, 247, 225, 246, 255, 245, 242, 245, 249, 243, 237, 230, 228, 253, 274, 269, 265, 260, 263, 259, 
    297, 293, 291, 277, 256, 255, 248, 247, 253, 256, 264, 246, 224, 245, 258, 251, 244, 257, 268, 272, 277, 282, 284, 284, 283, 279, 273, 262, 265, 262, 
    211, 204, 204, 208, 232, 252, 245, 244, 249, 258, 266, 255, 244, 255, 263, 264, 263, 271, 281, 293, 300, 294, 279, 258, 243, 233, 221, 243, 265, 264, 
    183, 172, 166, 164, 209, 249, 245, 241, 249, 266, 278, 265, 266, 266, 265, 264, 269, 269, 284, 283, 261, 237, 218, 206, 198, 186, 176, 218, 263, 266, 
    257, 248, 245, 242, 246, 249, 239, 239, 253, 274, 290, 277, 278, 277, 275, 273, 272, 273, 282, 267, 244, 239, 238, 236, 235, 206, 201, 241, 263, 266, 
    265, 263, 265, 264, 270, 257, 224, 207, 242, 274, 237, 190, 191, 190, 192, 199, 198, 216, 253, 263, 262, 263, 261, 257, 258, 242, 244, 265, 263, 264, 
    196, 189, 187, 196, 208, 217, 220, 236, 272, 280, 209, 144, 140, 135, 129, 130, 154, 209, 255, 268, 272, 270, 261, 249, 252, 261, 262, 249, 241, 253, 
    143, 129, 126, 165, 184, 172, 186, 236, 266, 260, 212, 171, 161, 172, 212, 243, 258, 267, 266, 256, 243, 227, 212, 197, 194, 200, 204, 201, 198, 223, 
    99, 107, 159, 197, 170, 128, 148, 190, 216, 228, 230, 233, 235, 263, 279, 263, 244, 228, 220, 208, 193, 180, 178, 183, 183, 187, 200, 212, 219, 238, 
    47, 102, 217, 240, 175, 155, 172, 196, 222, 249, 267, 277, 282, 299, 280, 237, 214, 222, 232, 235, 237, 236, 238, 242, 239, 243, 258, 267, 265, 251, 
    67, 168, 278, 286, 268, 268, 275, 286, 294, 300, 302, 293, 291, 311, 307, 296, 278, 279, 296, 296, 299, 302, 297, 285, 274, 268, 252, 230, 215, 201, 
    139, 236, 273, 273, 284, 295, 294, 292, 290, 292, 295, 289, 286, 283, 264, 254, 255, 261, 242, 223, 235, 246, 235, 214, 198, 193, 185, 177, 181, 190, 
    217, 239, 228, 228, 230, 232, 232, 234, 231, 230, 235, 240, 243, 230, 212, 207, 216, 226, 211, 198, 202, 202, 193, 187, 184, 186, 184, 178, 174, 175, 
    150, 149, 151, 163, 172, 174, 175, 177, 179, 187, 200, 214, 228, 228, 225, 224, 223, 219, 212, 205, 199, 188, 180, 177, 176, 171, 160, 149, 148, 160, 
    61, 56, 66, 71, 81, 82, 82, 82, 83, 91, 107, 126, 150, 180, 187, 186, 186, 181, 172, 165, 159, 156, 149, 140, 133, 127, 128, 130, 140, 156, 
    62, 40, 55, 70, 63, 48, 40, 38, 32, 30, 36, 53, 64, 95, 119, 122, 129, 131, 121, 113, 105, 101, 99, 96, 97, 110, 133, 141, 139, 149, 
    62, 45, 41, 64, 79, 68, 55, 44, 32, 25, 22, 28, 50, 63, 53, 42, 40, 39, 37, 35, 37, 47, 64, 94, 126, 139, 134, 128, 139, 162, 
    39, 32, 20, 25, 44, 48, 47, 42, 29, 19, 17, 0, 9, 51, 36, 0, 0, 0, 2, 22, 44, 72, 100, 111, 103, 100, 118, 143, 159, 183, 
    55, 31, 15, 11, 11, 16, 21, 21, 18, 14, 15, 0, 0, 0, 0, 0, 0, 0, 1, 33, 56, 62, 61, 66, 83, 112, 140, 156, 173, 200, 
    86, 41, 15, 12, 12, 15, 18, 17, 15, 13, 15, 0, 0, 0, 0, 0, 0, 0, 0, 15, 28, 34, 53, 88, 123, 141, 148, 164, 189, 212, 
    108, 52, 16, 16, 18, 21, 21, 17, 14, 14, 17, 6, 0, 0, 0, 0, 0, 0, 9, 18, 40, 72, 102, 125, 137, 141, 151, 169, 194, 218, 
    117, 57, 18, 18, 21, 25, 23, 19, 16, 17, 21, 18, 0, 0, 0, 1, 1, 0, 11, 42, 84, 119, 135, 137, 140, 148, 159, 176, 194, 216, 
    106, 53, 27, 22, 24, 27, 25, 22, 19, 20, 23, 23, 14, 1, 6, 5, 7, 25, 52, 80, 112, 134, 138, 139, 145, 160, 172, 186, 203, 222, 
    
    -- channel=18
    60, 58, 58, 58, 58, 58, 58, 58, 58, 58, 59, 59, 59, 58, 57, 56, 56, 57, 61, 64, 63, 61, 58, 58, 58, 59, 58, 59, 58, 58, 
    61, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 59, 58, 57, 57, 59, 62, 77, 68, 71, 62, 59, 60, 60, 60, 60, 59, 60, 
    61, 59, 59, 59, 59, 59, 59, 60, 59, 59, 59, 59, 60, 59, 59, 58, 59, 67, 71, 97, 73, 76, 59, 57, 59, 59, 59, 60, 59, 59, 
    61, 59, 59, 59, 59, 59, 60, 60, 59, 58, 59, 60, 61, 59, 60, 65, 72, 82, 86, 101, 67, 68, 57, 56, 59, 59, 59, 59, 59, 59, 
    61, 58, 59, 58, 58, 58, 59, 59, 58, 57, 58, 62, 65, 61, 68, 84, 96, 101, 99, 98, 77, 78, 69, 59, 60, 59, 60, 60, 60, 60, 
    68, 62, 63, 61, 59, 59, 58, 58, 57, 57, 54, 71, 68, 60, 74, 90, 96, 95, 97, 98, 92, 89, 75, 60, 65, 62, 62, 62, 62, 61, 
    73, 70, 71, 67, 63, 60, 58, 57, 57, 58, 53, 80, 60, 57, 70, 79, 78, 75, 84, 83, 78, 73, 67, 61, 72, 68, 68, 67, 65, 63, 
    95, 94, 94, 86, 69, 62, 58, 57, 59, 60, 55, 77, 48, 53, 60, 69, 68, 66, 78, 73, 72, 71, 75, 79, 87, 84, 82, 73, 68, 64, 
    126, 120, 116, 98, 62, 63, 59, 57, 59, 62, 61, 69, 49, 56, 61, 66, 66, 69, 79, 84, 96, 106, 111, 111, 107, 104, 95, 70, 69, 66, 
    82, 74, 75, 64, 42, 64, 60, 56, 61, 65, 69, 71, 65, 68, 71, 72, 73, 77, 84, 105, 115, 112, 105, 94, 86, 92, 75, 54, 68, 68, 
    62, 50, 50, 46, 48, 67, 69, 66, 62, 71, 96, 97, 97, 94, 93, 89, 92, 85, 85, 96, 84, 71, 67, 57, 61, 71, 45, 51, 71, 70, 
    104, 95, 92, 86, 80, 76, 81, 67, 59, 89, 138, 125, 125, 122, 119, 111, 101, 74, 73, 77, 70, 66, 73, 68, 69, 68, 51, 76, 82, 75, 
    124, 120, 120, 105, 90, 80, 69, 53, 60, 95, 126, 92, 94, 90, 77, 64, 51, 44, 66, 77, 84, 86, 93, 89, 84, 84, 86, 101, 95, 82, 
    101, 98, 84, 64, 80, 81, 61, 67, 82, 95, 91, 58, 51, 32, 24, 34, 46, 66, 88, 98, 107, 106, 106, 99, 97, 97, 98, 97, 90, 76, 
    83, 59, 30, 54, 83, 62, 44, 67, 75, 72, 60, 46, 41, 40, 71, 94, 98, 101, 101, 97, 96, 88, 78, 72, 72, 68, 65, 64, 69, 69, 
    70, 15, 17, 70, 57, 26, 19, 40, 45, 53, 55, 67, 67, 76, 99, 93, 85, 77, 75, 70, 69, 63, 60, 64, 65, 63, 69, 78, 90, 95, 
    27, 0, 50, 80, 50, 37, 37, 53, 64, 75, 81, 96, 86, 96, 98, 88, 84, 77, 96, 100, 97, 97, 101, 108, 106, 109, 117, 116, 112, 101, 
    15, 54, 107, 114, 106, 110, 110, 115, 119, 120, 118, 122, 114, 135, 133, 132, 120, 124, 145, 139, 133, 141, 142, 142, 131, 123, 113, 98, 87, 81, 
    63, 115, 129, 131, 136, 142, 140, 139, 139, 137, 135, 136, 132, 138, 125, 122, 115, 121, 123, 113, 116, 124, 119, 112, 101, 95, 90, 85, 78, 75, 
    113, 127, 123, 124, 127, 131, 130, 129, 125, 124, 127, 130, 131, 126, 114, 112, 114, 117, 115, 111, 114, 113, 108, 103, 102, 101, 94, 81, 69, 63, 
    88, 89, 87, 93, 100, 105, 105, 105, 104, 108, 117, 126, 135, 138, 135, 132, 129, 129, 126, 121, 118, 113, 107, 101, 96, 81, 67, 59, 52, 53, 
    43, 39, 37, 41, 48, 49, 51, 54, 55, 59, 71, 86, 94, 111, 119, 120, 118, 119, 113, 105, 100, 94, 84, 69, 54, 41, 45, 48, 43, 44, 
    32, 29, 32, 22, 23, 21, 22, 25, 24, 24, 31, 47, 32, 52, 67, 71, 74, 76, 67, 60, 50, 38, 29, 25, 31, 38, 45, 41, 33, 36, 
    25, 25, 32, 23, 24, 20, 20, 22, 21, 16, 19, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 31, 40, 33, 28, 31, 32, 38, 
    17, 18, 20, 17, 14, 12, 14, 17, 16, 11, 12, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 16, 16, 10, 10, 23, 36, 39, 47, 
    21, 21, 12, 10, 4, 1, 5, 10, 11, 9, 8, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 21, 33, 40, 44, 57, 
    27, 29, 9, 9, 8, 7, 9, 9, 9, 8, 8, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 23, 34, 37, 43, 51, 62, 
    36, 32, 7, 8, 9, 11, 12, 10, 9, 9, 10, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 24, 28, 33, 38, 46, 53, 62, 
    41, 22, 4, 3, 6, 10, 11, 9, 6, 6, 9, 10, 6, 0, 0, 0, 0, 0, 0, 0, 0, 18, 30, 31, 30, 34, 41, 47, 53, 61, 
    34, 8, 0, 0, 0, 4, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 27, 31, 32, 33, 39, 45, 51, 57, 65, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=20
    138, 139, 139, 139, 139, 139, 139, 139, 138, 139, 140, 140, 140, 139, 139, 140, 140, 140, 137, 138, 137, 137, 139, 139, 140, 139, 139, 138, 139, 139, 
    139, 139, 139, 139, 139, 139, 139, 139, 139, 140, 140, 140, 140, 140, 140, 140, 142, 142, 136, 146, 149, 149, 147, 140, 140, 139, 139, 139, 140, 140, 
    140, 139, 139, 139, 139, 139, 139, 139, 139, 139, 138, 138, 139, 139, 139, 138, 136, 135, 135, 133, 139, 133, 134, 137, 138, 138, 138, 138, 139, 139, 
    139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 138, 138, 138, 138, 137, 141, 147, 143, 141, 102, 117, 120, 132, 138, 139, 139, 139, 139, 139, 139, 
    144, 142, 142, 142, 140, 139, 140, 139, 138, 139, 138, 139, 141, 138, 134, 135, 137, 130, 121, 89, 113, 138, 149, 143, 139, 141, 140, 140, 140, 140, 
    139, 135, 135, 138, 140, 141, 141, 139, 138, 140, 136, 144, 145, 140, 138, 121, 99, 88, 84, 73, 79, 97, 122, 137, 138, 139, 138, 138, 140, 140, 
    123, 128, 127, 131, 138, 142, 142, 141, 140, 141, 140, 135, 134, 142, 133, 111, 93, 83, 78, 66, 56, 52, 77, 120, 136, 137, 136, 138, 139, 140, 
    168, 174, 173, 169, 152, 142, 143, 143, 142, 140, 149, 116, 122, 141, 133, 115, 105, 107, 100, 92, 85, 91, 108, 144, 157, 162, 162, 149, 140, 140, 
    110, 114, 123, 139, 140, 141, 147, 144, 140, 140, 150, 114, 121, 134, 139, 126, 119, 127, 117, 123, 133, 141, 140, 138, 134, 139, 150, 145, 139, 140, 
    21, 22, 22, 44, 107, 138, 148, 150, 146, 143, 147, 134, 138, 140, 141, 135, 131, 133, 124, 123, 116, 96, 83, 69, 59, 69, 80, 114, 135, 140, 
    67, 72, 67, 68, 118, 127, 140, 155, 143, 136, 161, 176, 174, 175, 173, 172, 171, 157, 138, 109, 86, 73, 69, 69, 61, 45, 53, 108, 136, 139, 
    131, 144, 150, 155, 154, 133, 113, 101, 105, 109, 108, 111, 114, 123, 132, 137, 128, 122, 128, 113, 106, 110, 109, 122, 116, 78, 102, 137, 148, 146, 
    100, 105, 123, 122, 121, 141, 114, 96, 120, 109, 35, 16, 22, 21, 10, 15, 36, 96, 135, 143, 151, 158, 154, 157, 160, 146, 155, 145, 143, 145, 
    58, 47, 31, 42, 97, 129, 128, 142, 153, 119, 25, 0, 0, 0, 17, 60, 105, 149, 158, 152, 144, 141, 123, 109, 114, 118, 107, 82, 81, 101, 
    59, 41, 0, 46, 72, 69, 100, 124, 124, 101, 60, 50, 49, 66, 99, 118, 124, 115, 98, 77, 54, 45, 36, 34, 38, 45, 46, 45, 50, 93, 
    23, 20, 58, 69, 26, 24, 58, 75, 90, 98, 104, 113, 119, 130, 108, 71, 61, 53, 46, 46, 35, 28, 33, 45, 48, 61, 85, 104, 106, 120, 
    0, 34, 133, 101, 71, 76, 100, 110, 124, 131, 138, 134, 138, 154, 135, 114, 93, 91, 106, 119, 109, 104, 108, 113, 115, 117, 119, 116, 102, 86, 
    0, 89, 129, 114, 116, 123, 129, 130, 132, 133, 137, 118, 123, 122, 118, 114, 98, 101, 91, 85, 93, 98, 94, 80, 76, 72, 64, 63, 65, 68, 
    94, 126, 113, 105, 105, 101, 98, 98, 93, 91, 90, 78, 80, 58, 48, 43, 59, 65, 41, 36, 52, 55, 51, 35, 32, 39, 47, 57, 62, 67, 
    106, 101, 91, 87, 86, 83, 83, 86, 88, 87, 88, 86, 81, 64, 58, 55, 64, 64, 53, 51, 50, 44, 40, 36, 37, 41, 44, 47, 54, 63, 
    20, 32, 27, 19, 23, 29, 35, 43, 54, 61, 68, 67, 62, 60, 63, 65, 59, 54, 47, 40, 35, 32, 30, 30, 27, 21, 22, 38, 60, 73, 
    1, 2, 18, 7, 0, 0, 0, 0, 7, 13, 19, 21, 0, 0, 0, 8, 16, 16, 9, 6, 6, 5, 2, 0, 2, 23, 51, 65, 68, 75, 
    24, 11, 34, 51, 39, 20, 9, 4, 4, 3, 1, 19, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 64, 87, 79, 64, 69, 76, 
    16, 14, 15, 54, 68, 57, 39, 25, 14, 8, 1, 8, 76, 76, 37, 16, 11, 9, 13, 20, 35, 61, 84, 96, 92, 76, 64, 69, 78, 83, 
    5, 9, 4, 25, 44, 42, 34, 23, 12, 10, 7, 0, 78, 153, 148, 134, 125, 118, 115, 113, 116, 115, 102, 74, 53, 61, 76, 79, 80, 93, 
    11, 6, 7, 9, 20, 25, 22, 15, 10, 9, 10, 0, 38, 122, 148, 144, 136, 132, 128, 118, 95, 69, 54, 55, 68, 82, 85, 83, 92, 100, 
    29, 10, 8, 8, 11, 15, 14, 11, 9, 9, 9, 7, 19, 89, 126, 130, 131, 122, 96, 64, 46, 44, 58, 79, 84, 80, 79, 87, 101, 104, 
    52, 16, 8, 7, 8, 10, 10, 9, 8, 8, 8, 6, 6, 63, 114, 115, 95, 68, 52, 47, 55, 68, 82, 87, 83, 77, 80, 86, 96, 102, 
    53, 20, 11, 8, 6, 6, 6, 6, 5, 4, 4, 1, 0, 29, 74, 63, 39, 35, 56, 75, 83, 88, 85, 82, 85, 86, 87, 91, 98, 104, 
    44, 28, 21, 16, 13, 10, 6, 4, 4, 3, 1, 3, 0, 14, 37, 42, 47, 57, 76, 92, 96, 90, 82, 80, 84, 89, 90, 96, 105, 112, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 4, 4, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 1, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 12, 22, 6, 0, 5, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 0, 0, 3, 2, 0, 0, 0, 0, 2, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 1, 0, 7, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 26, 25, 15, 2, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 15, 11, 2, 0, 0, 
    15, 20, 31, 33, 3, 0, 0, 0, 0, 0, 6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 12, 17, 26, 31, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 4, 2, 0, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 11, 5, 2, 23, 33, 30, 30, 28, 23, 20, 9, 0, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 21, 22, 11, 13, 0, 0, 0, 0, 0, 23, 27, 27, 28, 31, 27, 32, 7, 6, 3, 0, 0, 0, 0, 7, 0, 0, 0, 8, 3, 
    19, 21, 26, 33, 24, 29, 18, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 6, 11, 14, 21, 30, 33, 8, 5, 26, 22, 9, 
    12, 6, 8, 0, 0, 33, 15, 0, 15, 40, 12, 0, 0, 0, 0, 0, 0, 0, 12, 19, 24, 27, 26, 15, 13, 16, 18, 7, 0, 0, 
    31, 17, 0, 0, 1, 0, 0, 3, 19, 29, 1, 0, 0, 0, 0, 0, 2, 10, 10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 6, 1, 26, 32, 7, 4, 0, 3, 14, 9, 0, 2, 12, 7, 2, 10, 17, 18, 17, 
    0, 0, 14, 21, 3, 1, 5, 7, 12, 14, 17, 11, 0, 17, 22, 30, 4, 0, 15, 18, 9, 13, 15, 18, 17, 18, 16, 11, 8, 0, 
    0, 13, 26, 17, 16, 22, 22, 19, 16, 14, 18, 7, 3, 10, 3, 1, 0, 10, 7, 0, 0, 13, 17, 12, 2, 0, 0, 0, 0, 2, 
    30, 48, 40, 35, 33, 35, 35, 38, 35, 32, 30, 27, 29, 24, 14, 2, 7, 19, 14, 7, 11, 13, 13, 7, 0, 0, 2, 3, 0, 0, 
    11, 17, 8, 3, 9, 18, 20, 22, 26, 28, 30, 31, 32, 31, 28, 25, 21, 21, 23, 23, 17, 13, 8, 3, 3, 1, 0, 0, 0, 0, 
    3, 7, 0, 0, 0, 0, 0, 0, 2, 5, 10, 5, 0, 0, 6, 10, 10, 15, 13, 7, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 2, 12, 10, 9, 1, 0, 0, 2, 2, 7, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 6, 0, 0, 
    10, 0, 0, 6, 25, 27, 20, 14, 10, 6, 0, 24, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 23, 5, 0, 0, 0, 
    0, 1, 0, 0, 13, 19, 18, 17, 11, 6, 0, 0, 0, 25, 51, 44, 37, 30, 26, 18, 15, 22, 30, 27, 6, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 4, 9, 10, 9, 5, 3, 4, 0, 0, 0, 29, 39, 40, 38, 30, 29, 31, 25, 9, 0, 0, 0, 0, 0, 0, 0, 
    2, 10, 2, 3, 2, 4, 7, 5, 4, 3, 4, 0, 0, 0, 20, 29, 25, 27, 27, 21, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 17, 0, 1, 1, 2, 3, 2, 3, 2, 3, 0, 0, 0, 12, 28, 29, 23, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 26, 10, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    21, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 14, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 22, 22, 19, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 8, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 8, 4, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 51, 42, 36, 36, 32, 30, 27, 25, 20, 14, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 34, 29, 16, 19, 29, 36, 42, 47, 49, 48, 43, 30, 24, 23, 23, 19, 14, 15, 10, 7, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 24, 24, 14, 0, 0, 11, 26, 36, 42, 41, 33, 11, 0, 0, 5, 10, 9, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 45, 38, 40, 27, 21, 23, 29, 37, 43, 41, 22, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    31, 48, 49, 51, 55, 51, 48, 46, 45, 46, 48, 27, 24, 9, 0, 0, 0, 0, 0, 0, 0, 2, 24, 27, 11, 0, 0, 0, 0, 0, 
    16, 39, 51, 49, 51, 52, 50, 49, 47, 47, 49, 50, 44, 59, 45, 36, 35, 35, 36, 43, 50, 45, 27, 2, 0, 0, 0, 0, 0, 0, 
    13, 29, 48, 47, 48, 49, 49, 49, 48, 47, 48, 52, 49, 58, 56, 53, 53, 53, 57, 53, 35, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 27, 45, 47, 47, 47, 46, 47, 47, 48, 47, 47, 44, 50, 58, 58, 68, 64, 44, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 33, 39, 43, 44, 43, 44, 46, 46, 46, 45, 45, 43, 48, 64, 60, 47, 24, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 30, 32, 33, 35, 35, 36, 36, 36, 36, 34, 33, 32, 30, 29, 21, 6, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 21, 23, 23, 24, 23, 20, 17, 17, 16, 14, 12, 11, 5, 0, 0, 0, 0, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=23
    117, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 115, 114, 116, 117, 116, 117, 114, 116, 117, 118, 117, 116, 116, 117, 116, 116, 
    117, 117, 117, 117, 117, 117, 117, 117, 117, 116, 116, 116, 117, 116, 115, 116, 116, 115, 101, 111, 101, 112, 113, 116, 117, 117, 116, 117, 117, 117, 
    117, 117, 117, 117, 117, 117, 116, 116, 117, 117, 117, 117, 117, 117, 118, 118, 116, 110, 88, 111, 105, 117, 118, 115, 116, 117, 117, 118, 117, 117, 
    118, 117, 117, 117, 117, 117, 116, 117, 117, 117, 117, 116, 118, 115, 112, 108, 102, 96, 85, 112, 110, 117, 114, 114, 116, 117, 117, 118, 118, 118, 
    114, 112, 114, 115, 117, 117, 117, 118, 117, 117, 114, 114, 118, 112, 103, 99, 99, 94, 87, 97, 93, 103, 110, 111, 117, 118, 118, 118, 118, 118, 
    118, 116, 117, 118, 118, 118, 118, 118, 116, 117, 102, 113, 116, 107, 102, 105, 110, 105, 100, 99, 100, 112, 123, 116, 120, 121, 121, 120, 120, 119, 
    125, 120, 121, 122, 121, 119, 119, 116, 115, 116, 95, 118, 119, 111, 106, 114, 117, 110, 113, 114, 120, 129, 134, 123, 123, 124, 123, 123, 122, 120, 
    74, 76, 90, 110, 114, 118, 117, 115, 115, 117, 99, 126, 122, 117, 114, 119, 120, 112, 117, 115, 112, 108, 104, 94, 96, 101, 114, 118, 123, 121, 
    81, 81, 97, 124, 112, 115, 115, 114, 116, 118, 112, 129, 123, 120, 118, 120, 119, 113, 107, 96, 85, 82, 82, 80, 80, 93, 119, 119, 122, 122, 
    122, 120, 130, 140, 112, 108, 108, 109, 110, 112, 113, 118, 115, 116, 117, 119, 119, 115, 103, 103, 106, 109, 113, 104, 93, 114, 131, 125, 123, 124, 
    106, 104, 111, 111, 97, 93, 100, 105, 94, 74, 75, 67, 68, 72, 78, 83, 102, 108, 109, 122, 127, 122, 121, 108, 98, 126, 126, 119, 122, 123, 
    65, 62, 67, 76, 83, 94, 117, 127, 95, 54, 68, 59, 58, 61, 71, 90, 119, 121, 119, 122, 119, 106, 106, 99, 96, 110, 96, 99, 109, 115, 
    48, 50, 70, 75, 84, 97, 115, 116, 85, 59, 83, 79, 90, 107, 121, 132, 131, 108, 95, 87, 80, 68, 69, 70, 71, 71, 64, 80, 100, 104, 
    48, 70, 87, 72, 69, 84, 91, 91, 84, 85, 106, 110, 121, 116, 101, 87, 72, 60, 60, 56, 59, 60, 67, 73, 81, 84, 88, 100, 118, 110, 
    61, 94, 83, 72, 81, 97, 93, 104, 110, 116, 120, 121, 121, 94, 81, 80, 81, 84, 90, 90, 97, 100, 102, 104, 111, 115, 114, 111, 112, 97, 
    106, 114, 92, 104, 124, 128, 121, 128, 126, 123, 114, 123, 119, 107, 112, 116, 123, 116, 116, 112, 111, 109, 104, 103, 100, 93, 85, 76, 77, 78, 
    123, 101, 84, 109, 111, 110, 103, 105, 103, 102, 98, 113, 100, 92, 89, 90, 87, 73, 73, 74, 70, 67, 58, 59, 58, 57, 65, 71, 77, 81, 
    98, 71, 74, 84, 80, 79, 76, 74, 74, 76, 76, 87, 72, 72, 70, 76, 69, 55, 66, 70, 62, 57, 54, 61, 64, 68, 74, 75, 74, 75, 
    30, 35, 43, 48, 48, 50, 50, 51, 55, 60, 65, 69, 63, 69, 70, 72, 63, 55, 60, 56, 49, 48, 50, 54, 54, 55, 58, 62, 66, 73, 
    7, 11, 7, 8, 4, 2, 2, 6, 11, 14, 20, 22, 22, 25, 29, 32, 30, 28, 27, 24, 25, 29, 32, 35, 40, 47, 55, 63, 69, 75, 
    25, 32, 25, 19, 10, 4, 0, 1, 1, 1, 4, 4, 0, 0, 3, 10, 10, 10, 12, 14, 20, 26, 31, 40, 52, 58, 60, 65, 68, 80, 
    26, 40, 46, 36, 31, 24, 18, 15, 13, 11, 18, 31, 19, 19, 18, 19, 14, 14, 18, 23, 33, 46, 57, 62, 60, 49, 49, 62, 76, 96, 
    23, 33, 45, 32, 24, 20, 17, 17, 17, 16, 21, 61, 55, 55, 61, 57, 52, 52, 51, 54, 59, 59, 50, 37, 31, 36, 54, 78, 92, 108, 
    29, 31, 38, 25, 14, 10, 12, 14, 19, 20, 21, 58, 52, 32, 36, 39, 38, 35, 32, 27, 20, 12, 9, 20, 43, 64, 76, 90, 103, 114, 
    33, 31, 29, 21, 14, 11, 13, 17, 21, 21, 22, 42, 32, 0, 0, 0, 0, 0, 0, 0, 0, 8, 34, 59, 74, 81, 87, 102, 110, 116, 
    34, 35, 24, 21, 16, 13, 14, 19, 22, 22, 22, 28, 26, 0, 0, 0, 0, 0, 0, 0, 24, 52, 69, 75, 77, 85, 96, 109, 111, 116, 
    34, 36, 24, 23, 21, 18, 19, 22, 23, 23, 24, 24, 23, 0, 0, 0, 0, 0, 11, 46, 67, 77, 79, 79, 84, 94, 101, 108, 112, 116, 
    36, 39, 31, 29, 28, 27, 25, 25, 25, 25, 27, 26, 24, 0, 0, 0, 2, 39, 62, 73, 77, 81, 82, 88, 94, 99, 106, 112, 117, 118, 
    50, 51, 44, 42, 41, 40, 38, 37, 35, 35, 38, 39, 41, 27, 16, 36, 59, 71, 75, 74, 76, 83, 90, 95, 98, 101, 107, 115, 118, 116, 
    69, 67, 63, 59, 58, 58, 58, 57, 56, 57, 59, 61, 67, 66, 63, 68, 71, 75, 80, 79, 80, 89, 96, 99, 101, 104, 109, 113, 115, 114, 
    
    -- channel=24
    137, 139, 139, 139, 139, 139, 139, 139, 139, 140, 139, 139, 139, 140, 141, 142, 144, 142, 136, 129, 129, 133, 139, 142, 141, 139, 139, 139, 140, 139, 
    139, 140, 140, 140, 140, 140, 141, 140, 141, 141, 141, 141, 141, 142, 145, 147, 148, 142, 135, 125, 133, 131, 141, 142, 142, 141, 141, 141, 141, 140, 
    138, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 141, 142, 143, 140, 129, 112, 111, 131, 133, 142, 140, 139, 140, 139, 140, 140, 140, 
    140, 141, 141, 141, 141, 141, 140, 139, 140, 141, 139, 138, 138, 140, 140, 134, 122, 105, 78, 84, 115, 119, 133, 138, 139, 141, 141, 140, 140, 140, 
    140, 142, 141, 141, 143, 142, 141, 140, 141, 141, 139, 135, 135, 135, 125, 114, 101, 82, 61, 62, 99, 117, 131, 139, 140, 144, 142, 141, 141, 141, 
    135, 134, 136, 140, 143, 144, 143, 141, 141, 142, 141, 132, 141, 137, 106, 82, 67, 54, 38, 41, 69, 106, 132, 140, 135, 140, 140, 140, 140, 141, 
    113, 112, 116, 129, 140, 144, 146, 143, 141, 141, 134, 129, 152, 138, 106, 77, 56, 42, 24, 17, 26, 59, 106, 126, 124, 131, 132, 134, 137, 140, 
    107, 111, 114, 124, 140, 145, 148, 146, 142, 143, 126, 122, 153, 143, 114, 95, 87, 69, 50, 42, 40, 53, 84, 110, 120, 126, 128, 135, 136, 139, 
    94, 106, 120, 141, 153, 144, 149, 148, 143, 141, 126, 119, 140, 141, 125, 111, 107, 98, 87, 79, 75, 79, 89, 98, 109, 123, 138, 146, 135, 139, 
    11, 25, 52, 113, 145, 142, 155, 152, 144, 141, 130, 122, 126, 127, 124, 119, 113, 105, 89, 73, 68, 64, 57, 52, 52, 70, 124, 145, 133, 138, 
    1, 11, 23, 67, 109, 130, 145, 152, 149, 138, 121, 127, 123, 125, 124, 124, 115, 111, 84, 60, 51, 41, 34, 26, 12, 36, 95, 121, 124, 131, 
    60, 72, 79, 84, 97, 99, 109, 131, 117, 79, 68, 95, 96, 104, 112, 117, 128, 130, 99, 79, 75, 73, 71, 68, 51, 62, 93, 105, 119, 127, 
    51, 67, 82, 105, 109, 95, 92, 98, 69, 0, 0, 1, 2, 16, 38, 65, 99, 119, 113, 110, 109, 107, 107, 117, 113, 104, 103, 105, 119, 128, 
    0, 7, 47, 74, 88, 123, 137, 118, 75, 0, 0, 0, 0, 1, 16, 43, 85, 110, 113, 109, 106, 102, 99, 109, 115, 106, 85, 78, 97, 113, 
    0, 17, 38, 38, 72, 126, 152, 137, 105, 58, 26, 22, 37, 54, 63, 82, 94, 85, 69, 51, 37, 34, 33, 33, 39, 44, 39, 35, 58, 77, 
    39, 86, 44, 17, 46, 88, 112, 112, 104, 93, 91, 89, 99, 77, 51, 46, 37, 26, 7, 0, 0, 0, 0, 0, 6, 23, 33, 36, 45, 60, 
    58, 95, 57, 25, 36, 57, 72, 78, 82, 88, 92, 100, 107, 75, 42, 18, 19, 17, 7, 7, 4, 0, 4, 12, 23, 34, 47, 51, 48, 51, 
    36, 49, 39, 34, 33, 33, 38, 39, 40, 42, 39, 41, 45, 34, 33, 26, 18, 6, 5, 17, 12, 1, 0, 0, 10, 13, 17, 23, 24, 29, 
    23, 15, 6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 22, 36, 
    41, 24, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 36, 52, 
    23, 27, 15, 0, 0, 0, 0, 4, 16, 16, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 29, 57, 76, 
    9, 31, 21, 0, 0, 0, 0, 8, 22, 27, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 29, 58, 87, 100, 
    41, 60, 75, 57, 24, 14, 16, 21, 29, 32, 27, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 37, 61, 77, 93, 107, 118, 
    65, 70, 94, 109, 91, 74, 59, 48, 48, 50, 50, 79, 82, 19, 0, 0, 0, 0, 5, 22, 45, 62, 77, 93, 109, 117, 107, 107, 120, 127, 
    57, 64, 74, 95, 101, 92, 78, 66, 60, 60, 59, 102, 188, 206, 178, 173, 166, 160, 158, 154, 150, 151, 148, 140, 130, 126, 120, 119, 125, 126, 
    48, 55, 66, 73, 81, 79, 71, 66, 63, 65, 64, 91, 182, 268, 295, 299, 281, 254, 227, 205, 182, 166, 155, 143, 134, 132, 130, 128, 126, 120, 
    50, 51, 67, 68, 70, 68, 64, 65, 65, 65, 65, 83, 159, 251, 294, 293, 270, 234, 200, 173, 156, 150, 148, 145, 138, 133, 133, 133, 130, 119, 
    58, 60, 74, 72, 71, 67, 64, 65, 66, 67, 64, 76, 134, 214, 246, 235, 214, 190, 171, 158, 152, 149, 145, 144, 137, 132, 130, 130, 129, 120, 
    78, 84, 89, 85, 80, 74, 71, 72, 72, 71, 67, 72, 105, 159, 180, 170, 158, 160, 171, 177, 167, 154, 146, 143, 141, 134, 131, 128, 126, 118, 
    99, 113, 112, 104, 98, 90, 85, 83, 82, 80, 80, 86, 103, 132, 146, 149, 157, 177, 191, 192, 171, 153, 147, 142, 143, 139, 135, 131, 129, 119, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 1, 4, 0, 0, 0, 0, 0, 0, 
    1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 11, 17, 20, 24, 22, 9, 2, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 3, 0, 0, 3, 2, 0, 6, 14, 16, 20, 15, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 11, 0, 0, 0, 3, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    25, 24, 10, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 6, 0, 0, 0, 7, 0, 0, 
    28, 33, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 13, 14, 23, 25, 25, 27, 22, 12, 0, 2, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 16, 8, 7, 7, 0, 9, 20, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 12, 1, 9, 8, 0, 2, 13, 25, 26, 22, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 4, 0, 0, 0, 0, 0, 15, 42, 26, 42, 52, 45, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 49, 11, 0, 0, 0, 0, 0, 18, 35, 30, 32, 21, 0, 0, 0, 0, 0, 0, 3, 4, 14, 16, 15, 16, 24, 26, 16, 0, 0, 
    26, 44, 31, 32, 21, 13, 14, 7, 14, 11, 6, 0, 2, 11, 13, 11, 20, 29, 31, 39, 39, 35, 30, 27, 19, 8, 0, 0, 0, 0, 
    18, 10, 37, 26, 24, 14, 10, 0, 0, 0, 0, 0, 0, 3, 5, 8, 8, 0, 0, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 8, 3, 6, 0, 3, 11, 0, 0, 0, 0, 6, 6, 6, 5, 0, 0, 2, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 3, 2, 1, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 11, 16, 5, 0, 0, 0, 
    0, 0, 8, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 15, 21, 21, 12, 0, 0, 0, 0, 3, 
    0, 0, 0, 8, 2, 0, 0, 0, 0, 0, 0, 13, 51, 38, 22, 18, 22, 22, 20, 21, 23, 19, 5, 0, 0, 0, 0, 0, 1, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 34, 19, 13, 14, 10, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 3, 2, 3, 4, 3, 4, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=27
    432, 430, 431, 431, 431, 431, 431, 431, 432, 432, 432, 432, 432, 432, 430, 429, 429, 430, 433, 431, 431, 431, 432, 433, 432, 431, 431, 432, 432, 432, 
    435, 433, 433, 433, 433, 433, 434, 433, 434, 434, 434, 434, 434, 435, 433, 432, 432, 433, 435, 421, 420, 422, 426, 434, 434, 433, 433, 434, 435, 434, 
    434, 433, 433, 433, 433, 433, 433, 432, 432, 432, 433, 432, 433, 433, 431, 432, 434, 430, 407, 391, 391, 411, 425, 432, 432, 432, 432, 434, 435, 434, 
    435, 434, 434, 434, 434, 434, 433, 432, 432, 433, 433, 433, 433, 435, 436, 430, 418, 402, 352, 354, 366, 399, 421, 431, 433, 433, 434, 435, 436, 436, 
    430, 431, 431, 431, 434, 435, 434, 433, 434, 435, 436, 432, 431, 434, 430, 410, 387, 365, 326, 333, 351, 377, 404, 428, 437, 435, 435, 437, 438, 438, 
    427, 430, 432, 433, 436, 437, 435, 435, 436, 437, 438, 420, 422, 428, 401, 364, 348, 338, 317, 313, 326, 359, 398, 428, 440, 438, 439, 440, 440, 440, 
    432, 432, 434, 438, 440, 439, 438, 437, 437, 439, 423, 403, 414, 416, 391, 357, 343, 340, 324, 309, 312, 352, 411, 438, 444, 442, 443, 443, 443, 443, 
    390, 391, 393, 403, 427, 439, 438, 436, 437, 440, 402, 395, 413, 416, 401, 387, 387, 382, 375, 369, 373, 385, 412, 419, 420, 415, 418, 433, 446, 444, 
    316, 322, 339, 373, 417, 434, 430, 432, 436, 439, 404, 408, 421, 431, 420, 415, 423, 421, 427, 419, 404, 387, 372, 361, 357, 358, 381, 421, 445, 446, 
    240, 249, 290, 373, 417, 422, 417, 419, 425, 432, 419, 419, 424, 431, 431, 433, 438, 436, 428, 397, 362, 339, 315, 299, 286, 288, 358, 420, 445, 447, 
    285, 287, 314, 379, 399, 401, 391, 388, 409, 416, 384, 367, 373, 378, 385, 393, 399, 412, 399, 368, 346, 331, 319, 303, 274, 289, 369, 421, 439, 445, 
    340, 342, 354, 361, 361, 354, 352, 380, 394, 345, 280, 256, 266, 275, 288, 309, 358, 409, 413, 402, 397, 389, 384, 363, 331, 359, 391, 405, 417, 433, 
    257, 265, 276, 311, 337, 318, 335, 382, 360, 242, 160, 132, 136, 159, 209, 274, 359, 411, 422, 415, 402, 381, 367, 357, 348, 357, 349, 351, 370, 403, 
    120, 134, 195, 257, 269, 290, 345, 377, 340, 231, 170, 150, 172, 221, 264, 306, 350, 367, 362, 340, 317, 289, 274, 281, 290, 289, 279, 291, 333, 381, 
    44, 108, 220, 224, 203, 251, 311, 344, 342, 306, 285, 284, 321, 359, 356, 338, 322, 304, 282, 255, 234, 217, 212, 217, 231, 247, 263, 284, 330, 354, 
    55, 219, 279, 230, 216, 257, 303, 346, 375, 389, 394, 399, 417, 396, 347, 314, 288, 279, 273, 256, 247, 249, 255, 255, 271, 293, 305, 306, 315, 311, 
    150, 326, 331, 301, 298, 327, 353, 383, 404, 419, 417, 422, 428, 389, 341, 306, 308, 317, 311, 304, 311, 313, 304, 292, 290, 292, 289, 280, 270, 267, 
    262, 344, 356, 357, 360, 370, 377, 383, 385, 383, 366, 374, 367, 348, 326, 310, 314, 301, 289, 296, 300, 287, 259, 241, 231, 221, 217, 215, 218, 224, 
    244, 267, 274, 282, 289, 292, 292, 290, 293, 295, 291, 293, 270, 251, 239, 250, 245, 212, 197, 204, 199, 182, 157, 147, 149, 157, 165, 175, 194, 210, 
    145, 142, 143, 148, 150, 152, 155, 161, 168, 177, 187, 192, 183, 175, 173, 182, 182, 164, 148, 138, 128, 119, 114, 117, 123, 134, 146, 163, 185, 209, 
    16, 12, 27, 44, 43, 36, 38, 48, 59, 72, 87, 102, 111, 114, 118, 120, 120, 108, 94, 84, 79, 77, 80, 89, 102, 122, 143, 160, 180, 207, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 31, 33, 37, 34, 25, 20, 22, 30, 43, 61, 91, 126, 142, 144, 155, 183, 217, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 21, 16, 10, 9, 14, 24, 42, 73, 107, 131, 138, 134, 142, 168, 199, 249, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 76, 71, 56, 50, 54, 59, 72, 93, 109, 116, 116, 123, 137, 159, 189, 231, 287, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 83, 127, 118, 94, 90, 90, 91, 90, 88, 85, 82, 95, 124, 156, 181, 219, 268, 315, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 59, 48, 50, 48, 43, 34, 31, 47, 82, 122, 153, 177, 204, 246, 288, 327, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 45, 90, 135, 160, 174, 192, 222, 264, 300, 332, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 69, 115, 149, 165, 174, 184, 205, 233, 272, 309, 340, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 90, 132, 159, 168, 173, 186, 201, 220, 246, 280, 316, 345, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 33, 66, 104, 138, 163, 168, 169, 179, 195, 215, 236, 261, 294, 324, 345, 
    
    -- channel=28
    90, 89, 89, 89, 89, 89, 89, 89, 89, 90, 90, 90, 90, 90, 88, 88, 88, 90, 92, 90, 91, 89, 89, 89, 89, 89, 89, 89, 90, 90, 
    91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 89, 88, 90, 91, 93, 82, 85, 83, 87, 91, 91, 91, 91, 91, 91, 91, 
    91, 90, 90, 90, 90, 90, 90, 90, 90, 90, 91, 90, 90, 90, 89, 91, 94, 94, 92, 81, 82, 87, 89, 91, 91, 91, 91, 91, 91, 91, 
    91, 91, 91, 91, 91, 91, 91, 90, 90, 91, 91, 91, 90, 91, 91, 88, 86, 87, 79, 77, 74, 79, 85, 90, 91, 90, 91, 91, 91, 91, 
    88, 89, 89, 89, 90, 91, 91, 91, 91, 91, 93, 90, 89, 93, 96, 93, 87, 84, 75, 70, 66, 67, 77, 88, 91, 90, 91, 91, 91, 91, 
    90, 92, 91, 90, 89, 90, 90, 91, 91, 91, 95, 85, 87, 92, 92, 90, 88, 87, 81, 79, 78, 78, 80, 88, 92, 91, 91, 92, 92, 92, 
    94, 94, 94, 92, 90, 90, 91, 91, 91, 92, 93, 83, 83, 88, 91, 82, 79, 83, 80, 78, 78, 85, 91, 92, 93, 93, 93, 92, 92, 92, 
    67, 67, 67, 72, 85, 89, 90, 91, 92, 92, 86, 82, 83, 85, 87, 86, 85, 85, 85, 84, 81, 79, 81, 80, 79, 77, 79, 89, 93, 92, 
    78, 77, 73, 70, 83, 86, 87, 90, 92, 92, 85, 85, 86, 90, 88, 88, 91, 93, 97, 90, 84, 81, 79, 78, 77, 71, 72, 85, 92, 92, 
    70, 73, 78, 84, 84, 83, 81, 83, 87, 90, 85, 84, 86, 89, 91, 93, 95, 98, 102, 97, 91, 89, 83, 82, 77, 66, 78, 86, 92, 93, 
    54, 54, 62, 77, 81, 82, 73, 72, 87, 86, 66, 59, 61, 63, 65, 69, 72, 86, 93, 91, 83, 77, 73, 70, 67, 65, 80, 87, 91, 93, 
    62, 60, 62, 64, 70, 76, 80, 87, 95, 91, 70, 60, 60, 59, 60, 65, 79, 92, 92, 88, 83, 81, 78, 72, 68, 74, 79, 80, 84, 89, 
    62, 62, 59, 72, 70, 59, 68, 81, 85, 72, 55, 44, 44, 53, 67, 75, 82, 85, 86, 82, 75, 70, 66, 62, 58, 63, 67, 70, 72, 82, 
    30, 38, 52, 57, 46, 47, 63, 74, 76, 61, 50, 43, 44, 49, 45, 45, 56, 66, 72, 71, 67, 62, 61, 63, 64, 67, 68, 72, 77, 86, 
    0, 19, 54, 45, 37, 44, 63, 75, 78, 69, 61, 56, 62, 73, 73, 72, 74, 77, 76, 75, 70, 64, 60, 59, 60, 63, 65, 68, 73, 73, 
    0, 42, 61, 56, 47, 51, 67, 79, 81, 80, 80, 77, 86, 90, 90, 85, 75, 75, 71, 66, 63, 62, 61, 57, 59, 59, 56, 57, 62, 65, 
    27, 61, 67, 60, 54, 57, 66, 77, 83, 87, 89, 90, 91, 79, 66, 59, 64, 65, 59, 57, 62, 63, 61, 56, 55, 59, 63, 65, 65, 63, 
    56, 78, 86, 84, 83, 85, 90, 94, 94, 92, 89, 92, 92, 88, 82, 77, 80, 83, 82, 82, 81, 78, 74, 71, 66, 62, 58, 52, 48, 48, 
    46, 64, 71, 78, 84, 85, 86, 86, 89, 90, 90, 92, 88, 84, 79, 78, 74, 68, 64, 64, 62, 57, 49, 46, 42, 38, 35, 35, 40, 46, 
    29, 30, 34, 37, 39, 39, 39, 40, 40, 42, 48, 54, 52, 49, 46, 49, 50, 46, 42, 40, 38, 34, 32, 34, 33, 34, 35, 36, 37, 41, 
    3, 1, 12, 19, 18, 15, 12, 12, 11, 15, 23, 33, 37, 37, 36, 38, 39, 36, 33, 31, 28, 25, 25, 29, 33, 34, 34, 28, 29, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 28, 31, 27, 24, 22, 20, 18, 18, 19, 22, 26, 30, 32, 26, 20, 21, 27, 35, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 31, 28, 26, 25, 23, 20, 21, 25, 24, 14, 9, 13, 21, 25, 28, 41, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 6, 7, 5, 3, 0, 0, 0, 4, 14, 19, 21, 25, 35, 49, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 11, 14, 22, 33, 45, 57, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 18, 27, 37, 49, 61, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 12, 19, 23, 30, 42, 52, 63, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 11, 15, 21, 26, 34, 46, 56, 66, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 13, 14, 17, 22, 28, 36, 46, 57, 67, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 15, 16, 20, 26, 33, 40, 49, 57, 66, 
    
    -- channel=29
    510, 507, 507, 507, 507, 507, 507, 507, 507, 507, 508, 508, 509, 509, 508, 507, 505, 506, 505, 508, 507, 509, 506, 506, 506, 507, 507, 508, 508, 509, 
    511, 508, 508, 508, 508, 508, 507, 506, 506, 506, 506, 506, 507, 507, 505, 502, 499, 497, 471, 469, 454, 481, 489, 503, 506, 506, 506, 507, 508, 508, 
    511, 508, 509, 509, 509, 509, 508, 507, 506, 507, 507, 506, 507, 507, 508, 506, 498, 483, 433, 418, 409, 457, 484, 504, 509, 507, 508, 509, 510, 510, 
    512, 509, 509, 509, 509, 509, 508, 508, 508, 510, 510, 507, 508, 504, 491, 473, 453, 431, 392, 384, 391, 450, 487, 506, 511, 509, 510, 511, 513, 514, 
    501, 499, 503, 506, 509, 511, 510, 510, 512, 514, 508, 502, 501, 496, 470, 425, 384, 363, 338, 334, 333, 382, 446, 491, 511, 509, 509, 511, 513, 516, 
    489, 498, 502, 503, 508, 512, 513, 515, 517, 518, 490, 482, 474, 479, 461, 419, 389, 372, 358, 340, 326, 346, 411, 474, 512, 511, 511, 513, 515, 517, 
    500, 509, 511, 509, 509, 511, 513, 515, 518, 519, 479, 466, 453, 479, 468, 447, 442, 439, 439, 428, 430, 439, 464, 490, 512, 511, 512, 514, 516, 518, 
    334, 344, 377, 430, 474, 505, 509, 510, 512, 513, 482, 475, 462, 487, 493, 487, 486, 490, 499, 492, 485, 469, 448, 423, 411, 418, 452, 486, 512, 518, 
    201, 201, 240, 333, 422, 490, 497, 501, 506, 506, 492, 496, 491, 500, 504, 508, 511, 508, 492, 457, 413, 368, 330, 301, 278, 287, 354, 436, 504, 517, 
    334, 332, 356, 397, 434, 464, 458, 467, 479, 477, 472, 476, 481, 489, 496, 504, 511, 507, 478, 434, 384, 356, 347, 329, 299, 304, 351, 438, 502, 515, 
    432, 440, 467, 482, 462, 422, 395, 401, 406, 362, 310, 270, 285, 303, 328, 355, 408, 453, 475, 468, 450, 447, 451, 441, 417, 414, 430, 474, 499, 511, 
    300, 306, 331, 370, 393, 400, 403, 411, 401, 296, 170, 76, 83, 101, 141, 214, 324, 423, 489, 503, 498, 481, 472, 459, 454, 457, 439, 437, 446, 473, 
    133, 136, 176, 225, 287, 342, 398, 446, 424, 313, 195, 109, 132, 184, 254, 328, 402, 446, 454, 426, 393, 354, 327, 307, 310, 325, 313, 307, 341, 394, 
    64, 117, 161, 190, 213, 236, 306, 380, 389, 357, 326, 306, 333, 366, 393, 395, 378, 349, 313, 266, 226, 196, 186, 184, 198, 222, 249, 275, 323, 366, 
    30, 167, 255, 256, 199, 213, 273, 347, 389, 423, 443, 458, 476, 459, 408, 336, 295, 283, 279, 266, 255, 243, 249, 261, 280, 307, 341, 361, 369, 362, 
    62, 250, 393, 384, 341, 361, 397, 441, 469, 494, 488, 497, 496, 488, 445, 387, 370, 368, 385, 391, 395, 390, 379, 370, 361, 352, 344, 329, 316, 296, 
    167, 344, 420, 429, 428, 445, 456, 468, 473, 472, 452, 440, 414, 401, 377, 371, 361, 341, 333, 327, 338, 336, 303, 272, 251, 240, 229, 227, 234, 240, 
    278, 353, 352, 350, 355, 364, 366, 366, 362, 357, 347, 343, 313, 287, 258, 262, 272, 258, 230, 213, 219, 215, 188, 168, 157, 162, 173, 187, 207, 227, 
    192, 209, 209, 216, 222, 231, 238, 249, 257, 265, 272, 283, 275, 265, 245, 244, 240, 227, 209, 188, 171, 155, 142, 137, 138, 142, 151, 168, 192, 218, 
    0, 0, 2, 20, 31, 41, 48, 62, 78, 100, 123, 151, 169, 180, 180, 180, 170, 154, 140, 122, 105, 96, 92, 95, 106, 118, 135, 157, 185, 214, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 16, 27, 33, 32, 23, 16, 19, 27, 44, 71, 108, 140, 160, 173, 187, 218, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 40, 92, 144, 177, 181, 176, 173, 189, 237, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 142, 128, 86, 70, 72, 81, 100, 128, 156, 172, 173, 166, 157, 157, 178, 217, 274, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 207, 267, 241, 225, 216, 207, 192, 173, 153, 130, 111, 107, 125, 163, 205, 247, 306, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 88, 186, 196, 187, 172, 142, 105, 71, 52, 57, 82, 119, 152, 185, 226, 274, 327, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 112, 125, 93, 59, 26, 6, 7, 36, 80, 121, 147, 162, 189, 240, 292, 341, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 45, 0, 0, 0, 20, 60, 100, 130, 144, 153, 169, 200, 246, 295, 344, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 84, 118, 135, 139, 148, 166, 190, 223, 263, 308, 351, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 47, 89, 120, 134, 132, 134, 150, 175, 205, 238, 280, 324, 361, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 78, 96, 115, 124, 130, 129, 138, 161, 184, 212, 244, 282, 322, 357, 
    
    -- channel=30
    80, 83, 83, 83, 83, 83, 83, 83, 84, 84, 84, 84, 84, 83, 81, 82, 84, 83, 84, 87, 86, 82, 81, 82, 83, 82, 83, 84, 84, 82, 
    83, 85, 85, 85, 85, 85, 85, 86, 87, 87, 87, 87, 87, 86, 83, 84, 87, 89, 90, 104, 109, 100, 95, 88, 86, 86, 86, 87, 87, 85, 
    82, 84, 84, 84, 84, 84, 84, 84, 85, 84, 84, 84, 86, 85, 81, 81, 84, 90, 81, 111, 124, 108, 103, 88, 83, 84, 84, 85, 85, 84, 
    83, 85, 85, 85, 85, 85, 84, 84, 85, 84, 83, 84, 86, 86, 86, 91, 94, 95, 62, 94, 116, 106, 102, 88, 83, 83, 84, 85, 84, 84, 
    87, 89, 88, 88, 85, 84, 83, 84, 85, 85, 84, 85, 90, 87, 84, 96, 109, 104, 72, 97, 133, 140, 126, 96, 83, 85, 86, 86, 86, 85, 
    94, 89, 88, 90, 86, 83, 83, 84, 85, 86, 82, 88, 104, 87, 62, 60, 74, 75, 64, 78, 110, 144, 149, 110, 82, 83, 85, 86, 85, 85, 
    91, 82, 81, 85, 85, 84, 85, 86, 86, 88, 64, 81, 114, 82, 46, 39, 47, 40, 29, 25, 31, 70, 115, 105, 83, 83, 84, 85, 84, 85, 
    154, 149, 138, 124, 100, 86, 89, 90, 88, 89, 43, 62, 105, 78, 48, 50, 65, 52, 42, 40, 38, 58, 100, 120, 122, 123, 116, 100, 88, 85, 
    175, 180, 185, 182, 133, 90, 91, 92, 89, 89, 48, 58, 87, 84, 66, 64, 81, 77, 81, 94, 106, 117, 131, 140, 150, 163, 169, 132, 93, 86, 
    20, 32, 67, 135, 123, 92, 103, 104, 97, 93, 79, 84, 94, 94, 89, 87, 90, 87, 81, 84, 87, 79, 71, 64, 64, 102, 158, 137, 95, 87, 
    0, 4, 20, 78, 85, 83, 112, 127, 116, 111, 141, 168, 168, 162, 157, 149, 137, 112, 58, 30, 25, 13, 11, 3, 0, 32, 108, 112, 98, 90, 
    141, 151, 152, 141, 104, 67, 78, 108, 87, 60, 126, 193, 199, 201, 203, 192, 179, 138, 69, 45, 52, 51, 61, 57, 21, 56, 101, 114, 123, 111, 
    173, 188, 203, 188, 145, 91, 74, 84, 33, 0, 0, 60, 70, 69, 70, 83, 120, 122, 104, 108, 122, 123, 132, 145, 131, 133, 132, 144, 164, 147, 
    106, 94, 114, 124, 129, 155, 161, 131, 54, 0, 0, 0, 0, 0, 1, 51, 112, 136, 140, 142, 150, 145, 140, 151, 157, 140, 109, 110, 142, 140, 
    103, 70, 43, 26, 65, 138, 158, 132, 77, 3, 0, 0, 15, 41, 65, 106, 124, 113, 94, 67, 55, 52, 44, 40, 49, 50, 35, 36, 82, 105, 
    138, 131, 10, 0, 0, 37, 57, 65, 64, 50, 46, 64, 83, 47, 15, 25, 34, 27, 13, 0, 0, 0, 0, 5, 25, 50, 66, 73, 98, 109, 
    147, 160, 42, 0, 5, 33, 52, 77, 96, 100, 91, 112, 124, 81, 49, 41, 59, 71, 87, 97, 87, 83, 90, 106, 122, 130, 136, 129, 113, 103, 
    153, 154, 126, 127, 134, 141, 147, 155, 160, 156, 131, 142, 146, 142, 150, 148, 148, 132, 148, 179, 169, 148, 136, 142, 141, 119, 105, 97, 87, 83, 
    173, 161, 164, 173, 178, 176, 173, 167, 165, 159, 144, 138, 111, 97, 103, 120, 114, 76, 78, 110, 111, 96, 81, 79, 80, 75, 78, 87, 88, 81, 
    190, 185, 180, 177, 177, 179, 178, 174, 168, 164, 162, 153, 127, 108, 102, 109, 106, 90, 90, 98, 96, 89, 88, 91, 90, 85, 84, 87, 82, 78, 
    94, 122, 118, 112, 123, 137, 146, 155, 165, 173, 185, 190, 183, 174, 168, 156, 142, 130, 125, 118, 107, 100, 96, 91, 81, 64, 55, 66, 74, 74, 
    0, 37, 38, 3, 0, 10, 28, 46, 64, 79, 103, 116, 105, 97, 112, 120, 111, 98, 92, 84, 76, 69, 57, 46, 46, 46, 47, 60, 68, 67, 
    0, 37, 70, 33, 0, 0, 0, 0, 0, 9, 36, 68, 20, 0, 0, 0, 7, 10, 12, 11, 15, 21, 31, 47, 63, 64, 55, 58, 59, 68, 
    2, 27, 84, 95, 54, 18, 1, 0, 0, 2, 24, 121, 112, 0, 0, 0, 0, 0, 0, 0, 23, 50, 71, 81, 80, 63, 48, 53, 62, 76, 
    0, 0, 36, 64, 57, 33, 14, 1, 0, 2, 7, 121, 217, 158, 80, 64, 64, 65, 70, 80, 92, 96, 76, 46, 37, 43, 48, 60, 73, 83, 
    0, 0, 5, 18, 25, 15, 3, 0, 0, 1, 0, 49, 152, 172, 124, 110, 116, 110, 96, 76, 54, 38, 28, 23, 30, 45, 57, 73, 79, 82, 
    0, 0, 0, 3, 10, 6, 0, 0, 0, 0, 0, 10, 79, 115, 73, 54, 60, 52, 30, 7, 0, 6, 26, 36, 37, 46, 64, 84, 87, 85, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 60, 108, 69, 29, 16, 7, 4, 3, 9, 21, 33, 36, 35, 42, 59, 78, 85, 86, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 63, 31, 0, 0, 0, 18, 31, 31, 30, 34, 40, 44, 47, 57, 72, 80, 82, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 30, 37, 29, 29, 35, 43, 52, 57, 65, 80, 88, 84, 
    
    -- channel=31
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=32
    0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 87, 64, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 56, 73, 88, 67, 43, 65, 47, 0, 0, 0, 0, 0, 0, 0, 
    34, 54, 13, 0, 19, 13, 0, 0, 0, 0, 0, 0, 0, 0, 26, 71, 68, 53, 48, 46, 38, 54, 28, 0, 0, 0, 15, 40, 0, 0, 
    56, 66, 44, 36, 51, 36, 25, 27, 34, 28, 23, 30, 24, 15, 51, 69, 51, 38, 49, 55, 36, 44, 11, 0, 0, 0, 35, 64, 29, 32, 
    51, 60, 36, 23, 44, 54, 38, 27, 36, 42, 29, 27, 23, 29, 53, 56, 38, 34, 48, 53, 12, 0, 0, 8, 23, 0, 3, 77, 44, 49, 
    31, 47, 18, 7, 52, 61, 29, 0, 11, 37, 22, 9, 20, 41, 52, 45, 36, 28, 33, 32, 0, 0, 0, 0, 37, 0, 0, 89, 70, 46, 
    18, 47, 37, 31, 62, 61, 16, 0, 6, 26, 29, 18, 26, 45, 45, 39, 32, 20, 20, 10, 0, 0, 0, 0, 37, 13, 0, 86, 104, 44, 
    30, 58, 49, 51, 68, 41, 13, 7, 6, 12, 18, 12, 12, 22, 14, 5, 2, 0, 0, 0, 0, 0, 0, 0, 21, 50, 32, 82, 116, 58, 
    32, 41, 38, 30, 29, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 5, 64, 89, 82, 82, 57, 
    20, 12, 17, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 11, 47, 35, 0, 0, 0, 0, 0, 50, 74, 18, 10, 42, 
    17, 11, 20, 18, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 18, 12, 0, 10, 48, 29, 0, 0, 0, 0, 1, 27, 27, 0, 0, 32, 
    31, 38, 48, 36, 6, 0, 0, 0, 5, 10, 13, 13, 11, 8, 6, 3, 0, 0, 18, 0, 0, 0, 0, 0, 4, 14, 10, 0, 18, 22, 
    59, 48, 29, 2, 0, 0, 0, 16, 21, 15, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 13, 27, 40, 53, 48, 7, 
    54, 14, 0, 0, 0, 14, 21, 18, 8, 0, 0, 0, 0, 3, 16, 31, 7, 0, 0, 0, 0, 0, 18, 34, 40, 60, 74, 74, 63, 28, 
    18, 0, 2, 11, 13, 16, 26, 10, 0, 0, 0, 0, 27, 57, 68, 72, 16, 0, 0, 6, 14, 27, 47, 63, 67, 72, 76, 68, 63, 68, 
    9, 12, 15, 14, 17, 26, 37, 31, 26, 13, 1, 5, 47, 88, 78, 60, 7, 0, 7, 35, 45, 57, 70, 69, 68, 77, 76, 65, 78, 109, 
    0, 13, 18, 18, 45, 65, 67, 58, 55, 20, 0, 0, 44, 74, 54, 38, 15, 9, 41, 55, 59, 65, 72, 73, 78, 83, 78, 78, 102, 111, 
    0, 17, 20, 20, 60, 84, 61, 44, 37, 8, 0, 20, 58, 69, 56, 50, 43, 41, 51, 59, 64, 70, 75, 76, 78, 84, 83, 93, 100, 97, 
    1, 16, 22, 23, 55, 69, 45, 35, 38, 28, 38, 62, 76, 72, 58, 53, 51, 51, 61, 72, 78, 77, 64, 64, 87, 93, 89, 92, 93, 90, 
    24, 38, 50, 55, 71, 73, 63, 61, 64, 64, 65, 65, 61, 55, 53, 61, 68, 68, 76, 79, 74, 72, 66, 75, 98, 97, 87, 88, 90, 88, 
    66, 76, 83, 83, 86, 83, 73, 68, 66, 61, 60, 61, 63, 64, 71, 77, 69, 66, 70, 74, 78, 83, 79, 86, 98, 90, 84, 85, 84, 87, 
    88, 91, 85, 80, 80, 75, 66, 64, 69, 71, 72, 74, 75, 72, 76, 70, 42, 49, 84, 87, 84, 86, 85, 91, 90, 85, 83, 80, 85, 97, 
    89, 87, 80, 78, 78, 76, 72, 73, 76, 77, 74, 71, 68, 68, 76, 65, 31, 62, 105, 93, 83, 87, 92, 90, 86, 82, 81, 79, 96, 116, 
    89, 87, 81, 78, 77, 77, 73, 72, 69, 68, 67, 68, 72, 76, 87, 74, 38, 72, 109, 91, 84, 94, 91, 89, 86, 82, 79, 88, 114, 127, 
    83, 82, 77, 75, 75, 74, 71, 70, 70, 73, 78, 82, 89, 94, 104, 89, 46, 74, 107, 91, 91, 91, 90, 90, 89, 81, 81, 104, 130, 119, 
    
    -- channel=33
    291, 278, 253, 250, 281, 290, 290, 285, 281, 280, 271, 263, 266, 267, 270, 267, 256, 266, 268, 269, 266, 257, 262, 265, 267, 258, 264, 268, 258, 251, 
    291, 279, 247, 240, 274, 283, 280, 273, 273, 276, 265, 256, 263, 269, 270, 269, 257, 263, 268, 279, 261, 242, 255, 264, 265, 255, 263, 267, 253, 252, 
    281, 271, 238, 227, 262, 272, 267, 255, 259, 266, 252, 246, 252, 260, 260, 263, 253, 261, 273, 281, 250, 230, 249, 259, 262, 251, 260, 266, 248, 249, 
    271, 258, 229, 217, 248, 256, 256, 245, 250, 258, 244, 236, 242, 252, 252, 256, 249, 257, 282, 267, 196, 204, 249, 260, 260, 247, 253, 262, 243, 244, 
    262, 250, 219, 202, 234, 241, 242, 226, 235, 249, 236, 230, 238, 243, 238, 249, 246, 255, 275, 256, 200, 212, 246, 251, 253, 241, 243, 250, 237, 241, 
    248, 240, 202, 182, 213, 221, 220, 207, 220, 234, 223, 220, 233, 234, 218, 235, 234, 254, 271, 211, 169, 215, 249, 244, 235, 224, 226, 232, 221, 219, 
    227, 220, 178, 156, 185, 195, 193, 187, 202, 209, 202, 205, 225, 224, 200, 215, 231, 248, 270, 235, 194, 213, 226, 226, 232, 212, 206, 209, 196, 189, 
    222, 212, 171, 160, 193, 196, 191, 186, 194, 194, 190, 198, 214, 217, 230, 247, 234, 206, 181, 169, 155, 141, 117, 95, 153, 192, 208, 209, 181, 176, 
    203, 198, 176, 170, 198, 192, 181, 191, 192, 192, 194, 207, 218, 223, 247, 248, 213, 190, 187, 187, 178, 168, 145, 105, 108, 132, 158, 189, 159, 172, 
    168, 170, 167, 157, 162, 158, 158, 161, 165, 177, 183, 195, 207, 216, 236, 229, 205, 195, 200, 196, 183, 159, 133, 143, 161, 149, 138, 152, 136, 149, 
    148, 157, 152, 141, 158, 160, 150, 152, 164, 174, 182, 188, 198, 213, 222, 205, 186, 185, 185, 178, 151, 130, 137, 143, 134, 126, 156, 175, 156, 149, 
    152, 161, 159, 168, 193, 180, 155, 152, 182, 197, 192, 207, 228, 238, 231, 217, 207, 202, 196, 187, 152, 144, 185, 197, 175, 120, 136, 180, 167, 148, 
    170, 187, 175, 166, 189, 182, 167, 188, 225, 239, 234, 227, 235, 237, 224, 209, 203, 200, 199, 187, 157, 160, 187, 199, 208, 157, 134, 176, 156, 128, 
    192, 194, 181, 172, 171, 172, 183, 193, 203, 222, 235, 232, 230, 233, 228, 217, 210, 204, 198, 186, 162, 169, 176, 177, 190, 183, 154, 163, 155, 112, 
    198, 190, 182, 180, 178, 175, 186, 208, 228, 240, 251, 261, 265, 263, 253, 250, 250, 238, 227, 210, 183, 178, 177, 176, 183, 192, 171, 117, 105, 104, 
    218, 215, 215, 206, 219, 237, 251, 264, 272, 278, 283, 286, 284, 282, 269, 253, 246, 239, 229, 194, 156, 150, 162, 178, 187, 194, 177, 108, 90, 105, 
    234, 223, 231, 236, 240, 257, 266, 271, 277, 280, 282, 283, 281, 276, 263, 239, 220, 212, 203, 169, 136, 150, 172, 187, 194, 194, 178, 148, 171, 190, 
    230, 235, 235, 226, 212, 226, 258, 274, 280, 281, 278, 268, 254, 240, 226, 214, 204, 210, 217, 197, 178, 188, 193, 195, 194, 188, 179, 172, 176, 172, 
    236, 218, 199, 197, 216, 233, 250, 268, 267, 259, 245, 234, 228, 226, 224, 228, 223, 208, 219, 215, 203, 204, 204, 202, 196, 192, 189, 176, 156, 147, 
    212, 193, 215, 248, 265, 265, 250, 243, 232, 230, 237, 243, 245, 250, 241, 232, 222, 204, 213, 217, 209, 206, 210, 208, 202, 193, 171, 149, 128, 117, 
    239, 245, 251, 253, 247, 246, 240, 225, 227, 245, 246, 250, 247, 241, 221, 197, 174, 174, 206, 214, 213, 214, 213, 203, 175, 159, 150, 128, 115, 114, 
    239, 249, 251, 247, 245, 249, 243, 231, 225, 231, 227, 231, 238, 219, 173, 145, 131, 145, 197, 217, 211, 202, 183, 165, 154, 152, 137, 119, 119, 114, 
    203, 239, 249, 247, 248, 243, 220, 204, 197, 185, 188, 214, 226, 207, 169, 156, 160, 169, 186, 183, 176, 169, 163, 154, 142, 131, 116, 110, 106, 87, 
    187, 219, 229, 230, 234, 213, 175, 164, 168, 163, 169, 200, 217, 212, 197, 181, 168, 158, 156, 157, 161, 164, 152, 124, 112, 114, 108, 100, 89, 79, 
    180, 201, 210, 212, 219, 206, 177, 172, 181, 187, 194, 191, 177, 160, 151, 152, 153, 155, 158, 159, 146, 128, 117, 120, 125, 113, 101, 97, 92, 82, 
    169, 191, 200, 198, 197, 191, 181, 171, 164, 150, 140, 136, 138, 142, 148, 155, 155, 149, 146, 130, 117, 115, 112, 114, 118, 104, 92, 92, 92, 83, 
    137, 143, 146, 141, 138, 133, 128, 126, 126, 128, 131, 135, 142, 144, 142, 138, 126, 114, 122, 124, 115, 108, 101, 101, 102, 94, 90, 90, 84, 81, 
    91, 89, 90, 97, 104, 107, 108, 118, 127, 130, 132, 129, 126, 118, 112, 108, 107, 125, 144, 122, 101, 95, 93, 95, 93, 90, 88, 84, 80, 78, 
    83, 81, 81, 88, 95, 99, 101, 106, 110, 109, 107, 108, 115, 114, 108, 101, 102, 129, 147, 109, 90, 90, 91, 88, 89, 90, 88, 80, 80, 69, 
    84, 82, 82, 86, 89, 90, 90, 93, 98, 104, 108, 111, 114, 107, 96, 85, 88, 116, 131, 96, 85, 85, 82, 85, 88, 89, 85, 80, 75, 52, 
    
    -- channel=34
    122, 124, 125, 101, 109, 112, 112, 106, 97, 94, 93, 77, 76, 77, 70, 83, 70, 74, 70, 69, 76, 66, 64, 64, 75, 67, 64, 72, 70, 57, 
    116, 118, 117, 89, 99, 101, 103, 93, 84, 87, 85, 73, 72, 77, 66, 81, 69, 71, 67, 80, 87, 57, 59, 59, 73, 65, 60, 69, 69, 54, 
    107, 107, 107, 77, 88, 85, 90, 80, 70, 76, 75, 67, 61, 75, 60, 75, 67, 68, 73, 101, 88, 45, 56, 56, 70, 62, 57, 69, 66, 50, 
    95, 97, 100, 65, 77, 72, 79, 70, 57, 69, 67, 61, 54, 75, 58, 71, 70, 62, 73, 109, 74, 39, 60, 55, 67, 59, 53, 67, 61, 49, 
    86, 87, 95, 52, 67, 57, 64, 53, 44, 62, 59, 56, 47, 74, 63, 68, 72, 58, 82, 116, 67, 48, 72, 59, 65, 58, 45, 60, 54, 47, 
    73, 74, 88, 36, 49, 40, 46, 35, 30, 50, 46, 47, 41, 69, 56, 59, 72, 73, 93, 108, 73, 75, 96, 75, 65, 56, 36, 46, 44, 31, 
    64, 65, 73, 22, 35, 37, 35, 24, 22, 38, 34, 36, 39, 54, 42, 69, 93, 108, 110, 108, 95, 91, 101, 80, 56, 51, 34, 41, 44, 17, 
    71, 68, 69, 39, 54, 58, 42, 36, 34, 38, 35, 40, 52, 58, 60, 95, 99, 92, 80, 80, 74, 60, 68, 40, 39, 43, 41, 53, 50, 18, 
    77, 73, 78, 66, 69, 70, 57, 58, 53, 53, 55, 62, 75, 73, 83, 104, 97, 88, 88, 96, 94, 78, 62, 18, 38, 28, 22, 53, 48, 40, 
    74, 74, 77, 59, 60, 65, 64, 64, 54, 63, 69, 75, 83, 86, 100, 105, 95, 91, 92, 96, 95, 62, 43, 26, 47, 32, 0, 42, 42, 54, 
    71, 66, 72, 53, 66, 78, 76, 60, 55, 73, 77, 79, 88, 101, 109, 102, 94, 88, 83, 83, 77, 30, 22, 20, 27, 41, 0, 35, 59, 61, 
    71, 73, 87, 70, 86, 90, 75, 64, 76, 87, 94, 102, 110, 120, 119, 109, 100, 94, 85, 84, 67, 31, 37, 34, 26, 41, 3, 20, 74, 57, 
    86, 89, 92, 78, 92, 91, 88, 91, 100, 102, 108, 111, 110, 113, 110, 98, 91, 90, 82, 78, 55, 34, 44, 39, 35, 35, 32, 20, 74, 55, 
    99, 91, 89, 82, 83, 85, 85, 86, 92, 96, 102, 105, 106, 105, 105, 94, 90, 86, 77, 76, 56, 43, 40, 33, 38, 32, 59, 43, 52, 42, 
    103, 90, 86, 81, 77, 83, 90, 98, 104, 107, 113, 116, 118, 116, 117, 113, 107, 98, 91, 93, 65, 47, 36, 33, 42, 35, 62, 40, 4, 18, 
    117, 100, 96, 103, 109, 113, 120, 124, 125, 125, 127, 129, 130, 128, 124, 120, 107, 93, 84, 82, 45, 31, 35, 39, 51, 46, 52, 18, 0, 18, 
    119, 115, 122, 127, 123, 115, 121, 125, 130, 132, 135, 135, 132, 125, 113, 101, 87, 72, 67, 63, 37, 34, 47, 51, 60, 53, 53, 40, 39, 49, 
    132, 134, 123, 108, 101, 107, 119, 128, 139, 138, 132, 122, 110, 99, 88, 81, 85, 75, 73, 71, 58, 55, 56, 60, 61, 58, 62, 59, 61, 58, 
    131, 113, 94, 98, 107, 118, 123, 129, 127, 117, 108, 101, 95, 92, 92, 93, 101, 83, 78, 78, 70, 65, 62, 70, 72, 74, 73, 69, 64, 55, 
    115, 108, 113, 127, 130, 124, 119, 115, 103, 105, 107, 108, 103, 109, 112, 110, 111, 79, 75, 78, 75, 75, 78, 87, 83, 76, 72, 66, 51, 52, 
    127, 126, 129, 127, 120, 117, 117, 116, 110, 120, 114, 108, 103, 115, 109, 92, 89, 61, 73, 87, 89, 92, 89, 84, 74, 71, 70, 58, 46, 57, 
    118, 124, 129, 125, 120, 129, 128, 124, 118, 122, 101, 95, 94, 99, 82, 63, 68, 64, 84, 95, 90, 86, 81, 80, 73, 72, 67, 58, 56, 54, 
    102, 118, 125, 122, 118, 132, 119, 105, 99, 99, 82, 88, 95, 96, 85, 77, 81, 77, 79, 78, 79, 83, 85, 78, 63, 64, 60, 57, 52, 43, 
    97, 106, 112, 110, 107, 113, 94, 81, 83, 88, 89, 101, 107, 102, 92, 83, 79, 72, 72, 76, 82, 80, 74, 59, 55, 62, 58, 54, 49, 43, 
    94, 98, 108, 109, 109, 108, 98, 93, 99, 100, 96, 91, 82, 76, 73, 73, 79, 81, 79, 77, 70, 64, 65, 57, 63, 64, 55, 51, 51, 46, 
    96, 101, 110, 106, 104, 103, 98, 89, 81, 73, 68, 67, 70, 74, 76, 80, 85, 74, 66, 65, 60, 61, 60, 56, 62, 58, 52, 51, 51, 45, 
    77, 79, 79, 75, 74, 73, 70, 66, 66, 67, 69, 72, 76, 75, 70, 69, 65, 50, 63, 69, 61, 56, 52, 53, 56, 53, 50, 49, 44, 42, 
    50, 51, 50, 53, 57, 60, 61, 64, 68, 69, 68, 65, 64, 61, 56, 57, 56, 50, 76, 70, 52, 50, 50, 51, 52, 51, 49, 46, 36, 41, 
    43, 44, 43, 47, 51, 54, 54, 54, 56, 56, 57, 57, 61, 62, 56, 55, 53, 52, 78, 62, 47, 50, 48, 48, 51, 51, 50, 41, 36, 40, 
    42, 44, 42, 44, 47, 48, 47, 47, 51, 54, 56, 57, 59, 58, 51, 50, 48, 46, 72, 56, 47, 47, 44, 47, 51, 52, 46, 38, 40, 30, 
    
    -- channel=35
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=36
    77, 65, 57, 79, 90, 92, 99, 107, 108, 114, 113, 123, 129, 133, 136, 122, 129, 133, 135, 140, 147, 147, 143, 141, 132, 134, 139, 135, 134, 139, 
    87, 78, 64, 87, 103, 106, 105, 112, 119, 123, 118, 130, 134, 136, 141, 126, 131, 132, 134, 154, 162, 152, 145, 145, 134, 138, 145, 137, 135, 145, 
    90, 82, 71, 95, 111, 116, 112, 121, 130, 128, 124, 131, 134, 137, 148, 131, 134, 134, 135, 135, 122, 136, 144, 148, 137, 140, 149, 145, 134, 146, 
    98, 87, 78, 101, 115, 125, 120, 124, 136, 135, 128, 129, 136, 130, 153, 144, 145, 138, 137, 122, 107, 129, 141, 150, 138, 144, 156, 149, 136, 147, 
    109, 97, 82, 109, 121, 134, 127, 126, 144, 143, 132, 128, 138, 124, 146, 144, 138, 150, 139, 86, 85, 137, 160, 166, 144, 144, 157, 148, 144, 152, 
    111, 104, 80, 108, 118, 137, 136, 133, 150, 146, 136, 129, 147, 125, 106, 111, 118, 165, 174, 91, 93, 149, 177, 207, 179, 146, 151, 145, 154, 164, 
    129, 120, 81, 118, 132, 156, 153, 149, 163, 153, 145, 138, 154, 131, 111, 113, 106, 106, 93, 44, 42, 54, 62, 110, 149, 154, 164, 158, 164, 172, 
    140, 126, 86, 126, 149, 153, 153, 162, 172, 161, 159, 156, 157, 139, 140, 114, 83, 48, 32, 31, 27, 35, 28, 20, 73, 112, 138, 148, 142, 165, 
    104, 96, 79, 94, 96, 90, 109, 126, 128, 125, 132, 136, 123, 112, 119, 93, 64, 48, 48, 45, 48, 56, 30, 39, 76, 106, 98, 89, 79, 116, 
    56, 51, 47, 43, 39, 44, 67, 75, 65, 65, 76, 76, 59, 61, 70, 52, 41, 45, 45, 34, 39, 37, 12, 48, 46, 102, 119, 72, 59, 74, 
    26, 21, 28, 51, 53, 46, 42, 33, 41, 32, 33, 45, 46, 51, 50, 43, 44, 47, 44, 37, 28, 48, 72, 84, 50, 66, 144, 91, 71, 58, 
    21, 34, 30, 57, 69, 52, 30, 48, 76, 59, 41, 45, 50, 43, 33, 32, 30, 36, 41, 41, 30, 70, 114, 132, 115, 51, 131, 119, 65, 59, 
    33, 45, 28, 44, 45, 30, 28, 39, 47, 53, 40, 27, 29, 26, 21, 14, 10, 15, 28, 34, 45, 91, 116, 131, 140, 76, 96, 147, 77, 54, 
    24, 25, 18, 26, 5, 0, 0, 10, 22, 36, 39, 34, 39, 37, 34, 42, 48, 44, 56, 72, 95, 125, 125, 122, 125, 104, 63, 107, 57, 27, 
    24, 30, 24, 25, 28, 24, 27, 41, 49, 56, 58, 61, 62, 65, 61, 75, 86, 85, 86, 89, 99, 105, 110, 116, 108, 114, 65, 37, 13, 2, 
    32, 35, 45, 56, 77, 73, 61, 58, 61, 64, 68, 74, 79, 89, 85, 80, 84, 81, 73, 49, 54, 68, 91, 104, 100, 113, 77, 44, 82, 83, 
    35, 55, 73, 63, 47, 56, 64, 63, 67, 76, 81, 80, 76, 72, 69, 54, 61, 79, 78, 48, 57, 79, 86, 94, 92, 95, 79, 85, 130, 126, 
    47, 53, 32, 12, 8, 36, 61, 72, 75, 71, 63, 57, 54, 52, 58, 62, 69, 87, 90, 74, 81, 94, 87, 89, 86, 94, 98, 103, 107, 111, 
    12, 0, 9, 29, 52, 54, 59, 66, 53, 43, 46, 55, 65, 74, 84, 99, 101, 98, 93, 84, 85, 90, 92, 95, 103, 103, 91, 85, 71, 63, 
    17, 12, 33, 47, 55, 54, 49, 50, 53, 62, 70, 74, 74, 84, 96, 96, 87, 90, 87, 84, 88, 95, 107, 99, 86, 73, 67, 59, 39, 40, 
    49, 38, 41, 43, 43, 56, 65, 62, 76, 89, 86, 74, 69, 61, 50, 36, 20, 55, 89, 98, 99, 95, 85, 70, 61, 60, 54, 40, 48, 53, 
    46, 51, 51, 50, 49, 60, 71, 61, 59, 58, 63, 67, 73, 46, 20, 22, 20, 60, 88, 82, 71, 62, 59, 60, 55, 46, 33, 35, 50, 38, 
    40, 52, 49, 48, 47, 35, 26, 20, 19, 10, 37, 74, 93, 78, 58, 54, 46, 52, 53, 50, 54, 58, 56, 36, 27, 29, 27, 30, 26, 19, 
    37, 45, 44, 50, 60, 32, 16, 22, 36, 43, 71, 86, 80, 60, 45, 42, 40, 43, 51, 56, 51, 40, 34, 27, 30, 28, 27, 20, 16, 16, 
    46, 63, 67, 72, 80, 62, 51, 52, 51, 50, 51, 47, 41, 34, 33, 43, 50, 53, 48, 41, 29, 27, 27, 36, 38, 25, 18, 17, 17, 14, 
    48, 64, 64, 58, 54, 47, 41, 36, 32, 31, 31, 34, 41, 44, 45, 47, 40, 21, 17, 25, 31, 32, 23, 31, 29, 18, 15, 16, 14, 11, 
    25, 30, 28, 27, 26, 24, 24, 30, 34, 39, 41, 40, 34, 30, 29, 30, 24, 15, 23, 30, 30, 22, 20, 24, 19, 14, 14, 15, 12, 17, 
    18, 16, 15, 19, 21, 21, 22, 28, 29, 25, 22, 19, 18, 21, 25, 26, 28, 41, 36, 26, 21, 21, 23, 18, 15, 14, 15, 15, 16, 28, 
    21, 17, 16, 15, 15, 14, 13, 14, 15, 15, 16, 19, 22, 26, 30, 29, 34, 48, 31, 16, 20, 22, 16, 14, 14, 15, 17, 13, 27, 28, 
    16, 12, 12, 13, 14, 16, 17, 18, 21, 26, 28, 30, 31, 34, 37, 34, 36, 49, 27, 17, 22, 16, 15, 14, 13, 15, 14, 20, 32, 18, 
    
    -- channel=37
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 0, 1, 0, 0, 0, 1, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 4, 27, 4, 0, 0, 1, 0, 0, 0, 2, 0, 
    0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 3, 0, 0, 0, 16, 26, 0, 0, 0, 1, 0, 0, 2, 0, 0, 
    0, 1, 4, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 6, 3, 9, 5, 0, 2, 36, 7, 0, 0, 0, 3, 0, 0, 11, 0, 0, 
    0, 3, 11, 0, 0, 0, 4, 0, 0, 6, 2, 0, 0, 1, 6, 13, 15, 0, 0, 42, 1, 0, 9, 4, 4, 1, 0, 10, 0, 0, 
    0, 2, 13, 0, 0, 0, 7, 0, 0, 10, 5, 0, 0, 5, 0, 0, 2, 19, 51, 36, 0, 9, 47, 43, 27, 8, 0, 5, 5, 5, 
    8, 16, 16, 0, 0, 8, 14, 2, 4, 15, 5, 0, 13, 24, 0, 0, 0, 8, 40, 9, 0, 0, 7, 36, 33, 20, 7, 14, 21, 10, 
    28, 32, 13, 0, 13, 32, 22, 15, 23, 25, 16, 10, 23, 16, 0, 18, 24, 17, 0, 0, 0, 0, 0, 0, 0, 0, 8, 25, 34, 8, 
    24, 24, 6, 0, 15, 12, 6, 14, 21, 18, 14, 16, 22, 6, 15, 31, 20, 3, 0, 3, 0, 9, 23, 0, 0, 0, 0, 10, 2, 0, 
    3, 4, 7, 0, 0, 0, 0, 7, 0, 0, 0, 2, 0, 0, 2, 13, 0, 0, 0, 0, 7, 0, 0, 0, 0, 17, 0, 4, 0, 2, 
    0, 0, 2, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 9, 4, 0, 0, 0, 0, 4, 0, 0, 0, 0, 1, 0, 9, 8, 7, 
    0, 0, 0, 0, 9, 23, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 5, 29, 7, 
    0, 1, 0, 0, 12, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 28, 0, 5, 19, 36, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 17, 0, 0, 29, 32, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 12, 8, 12, 5, 0, 5, 5, 8, 8, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 3, 3, 0, 0, 9, 0, 0, 0, 0, 0, 14, 35, 4, 0, 0, 
    0, 0, 3, 5, 6, 0, 0, 0, 0, 0, 0, 1, 2, 4, 4, 0, 0, 0, 5, 0, 0, 0, 0, 0, 1, 9, 6, 0, 11, 39, 
    0, 9, 12, 0, 0, 0, 0, 0, 2, 3, 3, 1, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 2, 1, 2, 6, 21, 29, 
    5, 5, 0, 0, 0, 0, 0, 2, 7, 0, 0, 0, 0, 0, 0, 7, 16, 4, 1, 0, 0, 0, 0, 5, 4, 11, 17, 15, 17, 14, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 1, 14, 24, 36, 8, 0, 1, 0, 2, 6, 13, 19, 18, 13, 18, 1, 0, 
    1, 0, 0, 0, 0, 0, 4, 2, 0, 12, 10, 1, 0, 1, 16, 8, 3, 0, 0, 7, 8, 10, 21, 23, 11, 8, 17, 10, 0, 5, 
    0, 0, 0, 0, 0, 0, 15, 11, 5, 18, 5, 0, 1, 15, 5, 0, 0, 0, 0, 15, 16, 17, 8, 8, 9, 13, 10, 0, 11, 24, 
    0, 0, 0, 0, 0, 4, 7, 0, 0, 0, 0, 0, 22, 28, 8, 0, 0, 0, 7, 8, 5, 3, 6, 10, 4, 6, 0, 4, 13, 8, 
    0, 0, 0, 0, 6, 15, 0, 0, 0, 0, 0, 6, 20, 22, 15, 8, 4, 0, 0, 0, 7, 14, 18, 0, 0, 4, 7, 7, 3, 0, 
    0, 2, 9, 11, 26, 25, 7, 1, 0, 2, 11, 18, 14, 7, 0, 0, 0, 3, 7, 14, 10, 0, 1, 0, 8, 10, 5, 3, 2, 3, 
    3, 11, 21, 19, 19, 18, 14, 12, 11, 5, 2, 0, 0, 1, 1, 3, 8, 7, 0, 0, 0, 3, 1, 1, 13, 8, 0, 0, 2, 0, 
    1, 10, 15, 11, 9, 8, 6, 2, 2, 2, 1, 1, 3, 3, 3, 13, 13, 0, 0, 2, 7, 6, 0, 4, 7, 2, 0, 0, 0, 0, 
    2, 3, 0, 0, 0, 0, 0, 0, 0, 1, 3, 4, 0, 0, 0, 5, 0, 0, 5, 13, 4, 0, 4, 5, 3, 0, 0, 0, 0, 7, 
    2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 0, 0, 16, 10, 0, 5, 5, 2, 1, 0, 1, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 6, 9, 12, 16, 6, 0, 15, 2, 4, 5, 1, 1, 0, 1, 0, 0, 17, 20, 
    
    -- channel=38
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 16, 17, 31, 35, 34, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 9, 0, 0, 0, 0, 0, 
    4, 2, 0, 6, 16, 10, 10, 7, 6, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 11, 21, 
    15, 10, 11, 10, 1, 1, 9, 10, 11, 9, 10, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 25, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 11, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 7, 11, 13, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 2, 0, 0, 0, 0, 0, 0, 3, 1, 2, 7, 6, 10, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 7, 12, 12, 13, 22, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 4, 13, 18, 13, 13, 21, 26, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 4, 15, 13, 5, 2, 8, 19, 19, 20, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 14, 9, 0, 0, 0, 0, 0, 6, 15, 15, 8, 3, 9, 10, 14, 20, 19, 18, 20, 
    0, 0, 1, 7, 7, 9, 11, 12, 12, 9, 3, 0, 0, 0, 0, 6, 13, 18, 14, 6, 7, 12, 15, 18, 19, 19, 18, 18, 18, 18, 
    23, 27, 28, 24, 19, 16, 12, 6, 1, 3, 4, 8, 13, 16, 17, 18, 11, 0, 0, 5, 16, 17, 18, 19, 20, 19, 19, 18, 17, 19, 
    21, 21, 21, 20, 18, 16, 15, 16, 17, 20, 22, 21, 16, 9, 9, 8, 3, 1, 0, 12, 19, 16, 18, 20, 19, 19, 17, 17, 20, 23, 
    22, 22, 23, 23, 23, 23, 23, 21, 19, 14, 9, 7, 7, 8, 12, 14, 14, 13, 6, 14, 19, 19, 22, 21, 19, 19, 18, 17, 26, 32, 
    26, 23, 22, 20, 17, 14, 13, 11, 9, 8, 9, 12, 13, 16, 21, 24, 25, 20, 6, 15, 21, 21, 21, 20, 20, 20, 19, 22, 30, 41, 
    19, 16, 15, 14, 14, 14, 14, 15, 17, 18, 20, 24, 28, 33, 38, 41, 38, 30, 13, 20, 23, 21, 22, 21, 22, 20, 22, 28, 35, 44, 
    
    -- channel=39
    82, 80, 107, 102, 103, 101, 105, 107, 102, 100, 110, 110, 112, 118, 105, 120, 116, 119, 114, 103, 115, 116, 121, 113, 122, 123, 113, 114, 124, 115, 
    84, 82, 110, 103, 105, 101, 108, 112, 104, 102, 110, 110, 108, 120, 106, 120, 118, 117, 95, 90, 114, 114, 121, 112, 121, 123, 111, 112, 124, 113, 
    88, 84, 112, 102, 108, 101, 108, 115, 105, 106, 110, 112, 102, 119, 105, 115, 118, 111, 85, 97, 126, 115, 121, 110, 120, 122, 109, 113, 124, 112, 
    89, 82, 114, 101, 111, 103, 110, 121, 107, 110, 111, 115, 95, 111, 98, 102, 117, 99, 66, 101, 121, 109, 121, 108, 116, 119, 106, 115, 122, 109, 
    87, 75, 114, 95, 111, 102, 112, 120, 106, 111, 112, 116, 89, 101, 96, 96, 113, 92, 62, 103, 110, 91, 108, 102, 109, 118, 105, 113, 118, 104, 
    87, 72, 114, 94, 106, 99, 107, 113, 101, 111, 109, 112, 92, 109, 100, 92, 82, 56, 39, 62, 60, 43, 66, 81, 91, 114, 104, 105, 111, 95, 
    73, 63, 99, 78, 77, 82, 88, 94, 89, 101, 100, 98, 94, 107, 85, 74, 70, 67, 66, 77, 76, 61, 78, 88, 86, 91, 80, 79, 100, 80, 
    55, 51, 70, 53, 51, 63, 66, 66, 68, 78, 77, 73, 82, 89, 69, 70, 72, 73, 66, 66, 64, 52, 82, 83, 92, 83, 63, 64, 83, 64, 
    50, 48, 62, 59, 60, 69, 63, 65, 64, 69, 68, 67, 80, 79, 64, 67, 65, 61, 52, 54, 60, 56, 81, 63, 80, 89, 59, 78, 80, 66, 
    60, 59, 80, 77, 69, 64, 68, 75, 70, 76, 82, 84, 88, 78, 70, 71, 70, 67, 63, 66, 89, 92, 101, 77, 83, 110, 57, 71, 73, 63, 
    69, 62, 81, 68, 54, 63, 81, 89, 81, 81, 88, 85, 72, 62, 60, 63, 66, 73, 72, 77, 104, 99, 98, 87, 74, 115, 70, 53, 72, 62, 
    65, 54, 69, 55, 51, 60, 73, 71, 68, 69, 75, 77, 68, 63, 67, 72, 78, 85, 82, 90, 109, 94, 93, 88, 69, 94, 82, 36, 65, 59, 
    58, 52, 65, 56, 58, 69, 76, 78, 84, 83, 86, 89, 84, 82, 90, 94, 96, 99, 92, 97, 100, 87, 91, 86, 76, 65, 67, 26, 50, 56, 
    71, 67, 75, 81, 84, 92, 95, 94, 93, 92, 94, 94, 91, 87, 91, 91, 87, 84, 69, 75, 74, 76, 85, 83, 84, 54, 60, 51, 60, 65, 
    74, 74, 77, 84, 81, 80, 82, 82, 84, 87, 91, 91, 91, 84, 79, 78, 74, 68, 53, 72, 77, 84, 91, 85, 89, 61, 80, 103, 88, 80, 
    73, 67, 61, 61, 68, 72, 79, 82, 83, 83, 84, 82, 80, 76, 73, 79, 84, 78, 72, 95, 97, 92, 93, 85, 87, 71, 86, 95, 71, 70, 
    55, 45, 49, 66, 79, 82, 79, 74, 71, 69, 72, 77, 84, 90, 94, 94, 96, 88, 81, 97, 94, 87, 89, 85, 86, 77, 79, 72, 63, 79, 
    46, 60, 78, 92, 88, 78, 72, 65, 69, 77, 85, 93, 96, 97, 96, 88, 93, 90, 85, 90, 88, 85, 83, 80, 74, 63, 58, 52, 61, 81, 
    73, 83, 79, 74, 69, 67, 68, 78, 87, 94, 93, 91, 83, 76, 67, 60, 81, 84, 85, 88, 85, 80, 68, 62, 58, 52, 50, 53, 59, 64, 
    75, 76, 71, 73, 75, 74, 71, 80, 80, 82, 83, 84, 65, 53, 46, 45, 82, 86, 81, 81, 70, 60, 53, 56, 59, 56, 55, 58, 50, 40, 
    69, 74, 75, 75, 69, 61, 55, 57, 53, 68, 77, 82, 63, 59, 65, 67, 92, 80, 66, 61, 57, 57, 56, 60, 56, 51, 54, 51, 35, 29, 
    69, 68, 70, 69, 51, 47, 46, 50, 52, 77, 82, 80, 66, 67, 70, 64, 72, 61, 57, 63, 63, 60, 53, 53, 48, 50, 50, 42, 32, 33, 
    67, 68, 73, 73, 54, 60, 67, 69, 72, 83, 71, 56, 44, 45, 51, 53, 64, 64, 64, 59, 56, 54, 55, 57, 49, 46, 43, 37, 37, 37, 
    70, 69, 71, 67, 53, 60, 62, 56, 50, 50, 40, 40, 45, 55, 61, 61, 62, 56, 49, 49, 54, 56, 61, 50, 37, 39, 39, 38, 38, 39, 
    53, 44, 43, 39, 34, 38, 40, 41, 45, 51, 54, 56, 56, 57, 53, 48, 48, 49, 48, 54, 54, 50, 50, 38, 34, 38, 39, 38, 39, 39, 
    32, 27, 32, 34, 36, 41, 46, 49, 53, 56, 54, 51, 48, 47, 45, 50, 61, 59, 53, 50, 44, 42, 43, 36, 37, 40, 40, 40, 40, 34, 
    33, 33, 37, 39, 42, 45, 46, 44, 44, 46, 47, 49, 52, 52, 50, 58, 70, 51, 43, 45, 42, 39, 38, 36, 40, 41, 40, 42, 36, 27, 
    34, 36, 39, 41, 44, 45, 47, 47, 50, 52, 55, 56, 55, 50, 44, 54, 64, 39, 40, 45, 38, 35, 34, 36, 40, 41, 41, 40, 25, 21, 
    37, 41, 43, 47, 49, 51, 53, 53, 54, 53, 53, 51, 49, 45, 37, 47, 60, 36, 43, 42, 35, 32, 35, 36, 38, 41, 41, 31, 18, 22, 
    44, 47, 47, 48, 47, 47, 47, 47, 46, 44, 43, 39, 36, 31, 24, 36, 52, 32, 40, 37, 32, 33, 33, 35, 37, 42, 36, 21, 18, 27, 
    
    -- channel=40
    0, 0, 0, 14, 6, 9, 19, 34, 44, 49, 68, 92, 100, 105, 103, 98, 115, 115, 118, 119, 124, 140, 136, 126, 116, 126, 122, 116, 124, 133, 
    0, 0, 7, 45, 40, 40, 49, 70, 78, 79, 92, 110, 116, 118, 117, 108, 122, 123, 130, 122, 138, 159, 149, 136, 124, 136, 132, 121, 133, 145, 
    8, 5, 32, 72, 71, 73, 76, 99, 109, 103, 112, 126, 129, 127, 130, 117, 127, 126, 110, 100, 140, 165, 149, 141, 132, 146, 143, 128, 141, 151, 
    29, 25, 52, 95, 97, 103, 104, 131, 138, 124, 127, 136, 136, 135, 143, 131, 135, 133, 95, 68, 124, 156, 147, 146, 141, 158, 159, 141, 148, 153, 
    55, 45, 69, 118, 122, 131, 129, 156, 162, 144, 140, 147, 143, 134, 151, 146, 150, 133, 74, 65, 130, 151, 147, 153, 148, 168, 176, 160, 164, 164, 
    79, 61, 85, 137, 145, 155, 157, 181, 184, 166, 162, 164, 149, 126, 142, 136, 143, 130, 65, 50, 112, 147, 165, 174, 163, 172, 186, 180, 192, 198, 
    96, 75, 99, 149, 157, 167, 179, 199, 198, 187, 180, 177, 162, 139, 121, 92, 80, 74, 51, 26, 47, 79, 122, 183, 189, 184, 190, 188, 210, 233, 
    110, 91, 110, 151, 155, 170, 187, 198, 200, 197, 191, 179, 162, 150, 109, 51, 17, 0, 0, 0, 0, 0, 12, 101, 152, 180, 186, 179, 210, 230, 
    93, 81, 86, 110, 115, 125, 148, 156, 163, 165, 163, 145, 124, 112, 71, 21, 0, 0, 0, 0, 0, 0, 33, 70, 103, 142, 151, 130, 159, 163, 
    42, 36, 40, 52, 42, 52, 71, 81, 85, 81, 82, 68, 44, 27, 3, 0, 0, 0, 0, 0, 0, 23, 51, 82, 114, 153, 141, 86, 88, 81, 
    0, 0, 12, 29, 8, 0, 20, 33, 17, 4, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 66, 73, 75, 89, 161, 179, 96, 62, 50, 
    0, 0, 6, 34, 4, 0, 6, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 112, 131, 127, 94, 134, 182, 114, 60, 57, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 69, 121, 147, 161, 130, 116, 155, 120, 60, 66, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 38, 96, 133, 152, 156, 139, 102, 95, 107, 74, 62, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 14, 31, 66, 117, 146, 154, 145, 128, 87, 40, 66, 73, 52, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 26, 34, 27, 50, 98, 121, 128, 124, 107, 83, 57, 85, 87, 58, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 18, 34, 40, 26, 35, 74, 90, 96, 95, 89, 87, 90, 121, 136, 112, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 20, 36, 56, 49, 50, 71, 77, 77, 78, 82, 84, 91, 109, 118, 125, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 27, 36, 44, 64, 59, 56, 65, 71, 73, 73, 78, 81, 82, 80, 89, 115, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 16, 19, 28, 40, 56, 76, 64, 57, 61, 66, 65, 65, 72, 65, 54, 55, 62, 72, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 8, 0, 0, 3, 15, 44, 80, 66, 58, 58, 56, 56, 50, 47, 43, 41, 51, 49, 43, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 10, 0, 0, 0, 0, 20, 55, 58, 53, 49, 43, 36, 33, 37, 32, 36, 42, 42, 37, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 18, 5, 0, 0, 8, 21, 38, 39, 38, 33, 27, 22, 25, 25, 19, 22, 28, 30, 32, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 23, 21, 17, 17, 19, 19, 23, 25, 26, 28, 28, 21, 17, 13, 13, 18, 17, 18, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 19, 26, 24, 14, 9, 12, 18, 19, 21, 24, 24, 21, 18, 25, 27, 14, 11, 17, 16, 14, 18, 
    8, 11, 8, 10, 10, 6, 4, 9, 11, 18, 21, 21, 18, 19, 22, 22, 16, 18, 12, 15, 20, 21, 26, 26, 16, 13, 15, 15, 14, 19, 
    15, 17, 18, 16, 13, 12, 14, 17, 20, 25, 27, 26, 22, 22, 23, 22, 19, 12, 1, 12, 20, 20, 19, 18, 14, 14, 16, 17, 23, 27, 
    19, 20, 24, 25, 24, 23, 28, 28, 26, 24, 23, 20, 14, 15, 20, 29, 39, 27, 0, 10, 23, 18, 17, 17, 14, 15, 16, 24, 33, 37, 
    32, 30, 31, 29, 26, 24, 25, 22, 19, 14, 13, 16, 15, 22, 29, 40, 53, 36, 0, 13, 19, 17, 16, 16, 16, 16, 18, 31, 36, 48, 
    30, 28, 27, 24, 21, 19, 21, 23, 26, 27, 28, 30, 29, 35, 41, 50, 61, 39, 2, 12, 20, 17, 17, 16, 14, 16, 27, 32, 38, 55, 
    
    -- channel=41
    21, 8, 0, 18, 16, 7, 4, 8, 6, 2, 0, 2, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 6, 0, 11, 10, 5, 0, 1, 1, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 3, 0, 7, 5, 4, 0, 0, 1, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 11, 13, 13, 13, 15, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 1, 24, 12, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 10, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 6, 2, 0, 3, 7, 0, 15, 39, 8, 9, 0, 0, 20, 0, 0, 0, 
    18, 12, 1, 11, 6, 0, 13, 19, 21, 11, 8, 12, 6, 6, 10, 6, 8, 14, 16, 16, 16, 30, 22, 24, 0, 0, 25, 0, 0, 0, 
    14, 8, 0, 0, 1, 9, 2, 3, 20, 16, 5, 5, 12, 12, 11, 16, 14, 15, 18, 21, 2, 2, 0, 7, 8, 0, 1, 0, 0, 0, 
    8, 14, 0, 1, 6, 4, 3, 10, 13, 22, 19, 18, 26, 28, 32, 35, 30, 24, 23, 15, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 
    19, 24, 15, 30, 29, 28, 30, 29, 25, 28, 29, 26, 30, 30, 26, 28, 28, 15, 4, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    22, 32, 28, 28, 33, 28, 23, 24, 23, 21, 19, 19, 18, 16, 1, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 25, 28, 0, 
    18, 19, 5, 0, 7, 16, 15, 14, 14, 12, 8, 5, 0, 3, 0, 0, 2, 9, 10, 0, 5, 0, 0, 0, 0, 14, 16, 4, 16, 8, 
    0, 0, 0, 2, 4, 11, 12, 8, 2, 1, 1, 3, 6, 10, 15, 7, 5, 17, 24, 5, 5, 2, 0, 0, 0, 1, 0, 0, 0, 3, 
    0, 15, 30, 29, 11, 5, 1, 0, 0, 8, 13, 17, 20, 18, 16, 7, 0, 8, 11, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 28, 24, 14, 14, 5, 2, 12, 19, 20, 18, 13, 7, 0, 0, 0, 0, 4, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 14, 12, 8, 14, 15, 11, 12, 10, 10, 9, 4, 0, 0, 0, 0, 0, 7, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 17, 16, 15, 7, 3, 0, 0, 0, 0, 10, 9, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 13, 11, 9, 0, 0, 0, 0, 0, 0, 12, 12, 21, 15, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 10, 8, 11, 10, 1, 8, 14, 16, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    14, 13, 6, 7, 22, 14, 10, 7, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 2, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 1, 3, 4, 4, 2, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=42
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=43
    328, 296, 311, 353, 387, 400, 403, 408, 418, 410, 414, 424, 435, 441, 428, 427, 433, 445, 454, 447, 434, 438, 449, 442, 439, 447, 448, 439, 439, 450, 
    338, 301, 316, 361, 394, 401, 404, 414, 422, 412, 414, 422, 433, 441, 431, 431, 433, 447, 455, 420, 399, 424, 451, 446, 442, 450, 450, 439, 443, 454, 
    341, 305, 317, 360, 395, 399, 401, 411, 419, 410, 405, 413, 423, 432, 425, 427, 430, 441, 417, 363, 373, 416, 449, 445, 442, 450, 450, 432, 442, 451, 
    342, 305, 313, 354, 392, 397, 397, 411, 419, 406, 397, 407, 409, 419, 410, 411, 415, 428, 371, 300, 334, 406, 446, 442, 438, 443, 439, 427, 438, 446, 
    341, 298, 303, 343, 384, 389, 389, 408, 413, 399, 389, 402, 393, 391, 376, 379, 401, 397, 320, 279, 329, 386, 418, 420, 423, 427, 422, 420, 429, 435, 
    337, 283, 289, 329, 377, 380, 381, 401, 401, 389, 382, 397, 371, 348, 351, 352, 371, 338, 235, 218, 270, 309, 338, 342, 365, 399, 406, 407, 408, 407, 
    314, 257, 275, 312, 351, 347, 356, 378, 373, 368, 367, 380, 354, 336, 330, 303, 274, 240, 189, 172, 182, 199, 233, 277, 315, 356, 366, 360, 360, 367, 
    266, 224, 248, 274, 285, 292, 310, 326, 322, 326, 331, 334, 324, 330, 303, 247, 187, 154, 139, 122, 117, 94, 96, 186, 260, 310, 315, 282, 295, 306, 
    193, 174, 180, 194, 204, 221, 236, 245, 252, 261, 268, 264, 270, 285, 255, 204, 170, 160, 150, 141, 131, 109, 132, 165, 199, 228, 245, 214, 224, 224, 
    123, 120, 125, 144, 153, 154, 150, 162, 184, 193, 195, 203, 227, 234, 208, 183, 170, 161, 149, 138, 128, 142, 204, 207, 226, 224, 208, 188, 159, 149, 
    103, 114, 131, 147, 141, 118, 118, 157, 172, 176, 183, 194, 208, 200, 178, 161, 154, 153, 147, 133, 161, 215, 250, 232, 225, 259, 229, 205, 140, 121, 
    128, 126, 148, 159, 133, 110, 140, 182, 190, 190, 199, 210, 208, 192, 176, 165, 168, 175, 174, 170, 225, 291, 320, 296, 226, 258, 239, 190, 135, 106, 
    143, 127, 134, 131, 118, 120, 153, 196, 225, 222, 216, 222, 218, 204, 189, 190, 197, 209, 209, 216, 263, 300, 322, 319, 254, 240, 234, 141, 97, 85, 
    148, 139, 136, 122, 129, 151, 181, 209, 236, 249, 251, 255, 253, 249, 247, 248, 248, 253, 247, 241, 259, 272, 287, 293, 270, 216, 190, 103, 74, 74, 
    167, 163, 170, 179, 185, 206, 235, 258, 276, 290, 300, 305, 307, 298, 296, 292, 286, 277, 249, 225, 228, 252, 273, 275, 274, 206, 135, 103, 116, 115, 
    198, 212, 218, 227, 234, 258, 284, 300, 311, 318, 322, 322, 317, 300, 280, 271, 268, 257, 214, 194, 209, 244, 266, 269, 271, 220, 173, 189, 184, 149, 
    212, 208, 195, 199, 237, 269, 290, 303, 306, 302, 296, 290, 283, 275, 258, 256, 260, 250, 216, 212, 231, 252, 268, 265, 263, 243, 238, 254, 238, 200, 
    173, 154, 166, 193, 237, 270, 286, 284, 274, 268, 266, 265, 263, 265, 264, 262, 269, 272, 259, 258, 266, 267, 271, 262, 256, 239, 220, 203, 192, 197, 
    151, 162, 193, 226, 241, 255, 258, 247, 247, 257, 264, 271, 276, 277, 272, 251, 243, 260, 272, 273, 274, 275, 268, 249, 223, 195, 167, 133, 129, 172, 
    175, 205, 233, 250, 253, 247, 237, 236, 248, 263, 274, 282, 282, 256, 215, 186, 196, 234, 266, 271, 265, 256, 226, 196, 172, 143, 107, 82, 88, 109, 
    209, 231, 236, 237, 245, 237, 219, 224, 233, 237, 250, 265, 241, 187, 138, 118, 166, 224, 246, 238, 221, 199, 171, 143, 120, 93, 69, 69, 57, 24, 
    210, 228, 230, 233, 232, 208, 177, 170, 171, 190, 226, 249, 208, 150, 118, 106, 147, 184, 192, 182, 166, 147, 121, 97, 78, 60, 52, 46, 16, 0, 
    192, 215, 221, 222, 196, 155, 128, 127, 129, 173, 220, 232, 193, 146, 125, 119, 133, 142, 143, 135, 119, 99, 74, 67, 53, 35, 23, 7, 0, 0, 
    172, 198, 209, 208, 165, 127, 117, 124, 131, 154, 169, 166, 148, 129, 122, 116, 115, 114, 107, 93, 78, 67, 52, 49, 32, 15, 0, 0, 0, 0, 
    155, 172, 176, 172, 144, 120, 113, 113, 116, 118, 113, 103, 94, 91, 95, 96, 91, 82, 74, 61, 50, 40, 43, 39, 15, 0, 0, 0, 0, 0, 
    106, 109, 105, 99, 90, 81, 75, 73, 70, 68, 68, 71, 73, 74, 74, 64, 54, 60, 56, 43, 32, 21, 25, 16, 0, 0, 0, 0, 0, 0, 
    30, 26, 25, 24, 24, 26, 32, 40, 46, 49, 49, 49, 51, 50, 44, 34, 41, 59, 50, 28, 12, 7, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 17, 24, 27, 29, 30, 30, 32, 29, 22, 27, 58, 65, 37, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 9, 13, 16, 20, 25, 29, 24, 12, 17, 50, 50, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 8, 15, 18, 19, 17, 12, 0, 0, 0, 20, 24, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=44
    88, 80, 76, 87, 97, 100, 98, 97, 100, 96, 93, 93, 95, 95, 96, 93, 94, 97, 97, 95, 87, 90, 95, 97, 95, 96, 99, 96, 92, 97, 
    87, 77, 73, 84, 92, 96, 94, 93, 96, 93, 90, 90, 95, 94, 96, 93, 93, 97, 99, 82, 72, 85, 95, 97, 94, 95, 98, 94, 91, 97, 
    85, 75, 67, 79, 88, 90, 87, 85, 90, 88, 85, 86, 92, 89, 91, 92, 90, 97, 96, 79, 72, 83, 93, 96, 92, 93, 95, 91, 92, 96, 
    82, 72, 62, 73, 82, 85, 83, 82, 87, 84, 81, 81, 87, 85, 81, 82, 82, 96, 87, 53, 58, 81, 92, 94, 90, 87, 91, 88, 89, 93, 
    77, 69, 55, 66, 75, 78, 76, 77, 82, 79, 77, 79, 83, 79, 72, 75, 77, 83, 79, 60, 56, 66, 74, 82, 84, 80, 82, 84, 84, 88, 
    75, 64, 51, 62, 74, 72, 71, 72, 77, 74, 73, 76, 74, 72, 77, 72, 70, 57, 37, 35, 37, 42, 42, 42, 61, 72, 75, 75, 70, 73, 
    61, 51, 43, 48, 58, 53, 57, 61, 63, 63, 64, 69, 64, 60, 65, 65, 64, 64, 56, 51, 50, 55, 52, 46, 45, 54, 58, 56, 47, 52, 
    46, 38, 36, 37, 41, 42, 43, 45, 46, 47, 49, 53, 53, 59, 62, 59, 49, 40, 36, 30, 23, 13, 10, 37, 45, 55, 54, 41, 36, 37, 
    35, 30, 29, 36, 40, 39, 39, 39, 42, 42, 45, 48, 54, 61, 58, 48, 40, 35, 35, 32, 23, 19, 17, 17, 19, 29, 53, 42, 40, 36, 
    25, 25, 25, 33, 33, 30, 23, 31, 41, 40, 42, 50, 61, 64, 56, 49, 41, 37, 38, 35, 24, 28, 44, 45, 39, 14, 30, 38, 26, 27, 
    24, 25, 20, 23, 28, 22, 23, 36, 42, 48, 46, 48, 56, 55, 47, 37, 31, 30, 31, 24, 21, 28, 36, 40, 43, 30, 26, 45, 21, 21, 
    26, 25, 28, 30, 25, 22, 25, 32, 38, 45, 53, 56, 59, 58, 52, 46, 45, 44, 42, 34, 37, 47, 53, 47, 36, 40, 25, 38, 23, 12, 
    33, 29, 30, 31, 32, 30, 40, 55, 63, 63, 65, 69, 68, 64, 58, 58, 58, 58, 52, 44, 44, 49, 56, 57, 42, 43, 29, 11, 13, 10, 
    42, 40, 39, 37, 47, 54, 59, 61, 67, 71, 71, 71, 71, 70, 65, 61, 60, 57, 49, 35, 33, 35, 44, 50, 47, 44, 36, 10, 11, 12, 
    45, 42, 48, 47, 47, 56, 64, 69, 74, 78, 80, 81, 80, 76, 74, 68, 65, 60, 53, 37, 34, 39, 44, 48, 50, 42, 28, 17, 27, 26, 
    56, 56, 53, 52, 55, 70, 81, 86, 89, 89, 87, 83, 77, 70, 66, 63, 62, 62, 53, 41, 36, 42, 47, 50, 51, 42, 26, 14, 13, 18, 
    57, 51, 50, 57, 69, 74, 81, 85, 83, 80, 78, 77, 73, 70, 64, 61, 55, 51, 44, 38, 38, 45, 54, 53, 53, 48, 39, 34, 33, 25, 
    50, 50, 59, 63, 70, 75, 76, 77, 75, 75, 75, 72, 68, 65, 59, 55, 54, 55, 53, 51, 51, 53, 57, 53, 49, 41, 34, 29, 25, 24, 
    57, 53, 53, 57, 62, 70, 72, 70, 73, 69, 66, 63, 61, 58, 55, 47, 42, 50, 57, 57, 57, 57, 54, 45, 36, 32, 28, 18, 19, 24, 
    51, 58, 66, 72, 73, 70, 67, 62, 61, 60, 63, 66, 67, 56, 44, 38, 33, 43, 56, 55, 52, 48, 41, 38, 32, 24, 13, 6, 8, 10, 
    61, 68, 69, 68, 67, 60, 52, 52, 53, 51, 59, 66, 63, 51, 38, 32, 35, 41, 44, 43, 41, 39, 35, 25, 16, 9, 2, 0, 0, 0, 
    57, 62, 63, 63, 63, 52, 43, 44, 46, 46, 53, 60, 53, 39, 27, 17, 21, 29, 36, 38, 35, 27, 17, 10, 8, 4, 0, 0, 0, 0, 
    49, 58, 61, 62, 60, 50, 40, 40, 39, 45, 49, 47, 37, 24, 18, 18, 24, 28, 28, 24, 15, 11, 8, 9, 5, 0, 0, 0, 0, 0, 
    42, 52, 55, 53, 44, 35, 28, 25, 22, 23, 28, 33, 35, 32, 27, 23, 19, 15, 12, 10, 11, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 36, 36, 35, 28, 21, 19, 19, 22, 24, 23, 20, 18, 14, 11, 10, 8, 8, 10, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 21, 20, 21, 19, 17, 15, 13, 10, 6, 3, 3, 4, 4, 5, 6, 7, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 4, 1, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=45
    405, 369, 370, 402, 465, 482, 486, 495, 505, 502, 499, 500, 514, 526, 511, 514, 504, 524, 530, 515, 509, 504, 527, 524, 527, 528, 533, 526, 528, 533, 
    401, 364, 369, 398, 461, 477, 482, 488, 498, 493, 485, 488, 497, 517, 504, 513, 502, 513, 481, 441, 435, 464, 523, 524, 528, 528, 531, 526, 525, 527, 
    402, 359, 364, 388, 453, 464, 471, 478, 484, 484, 471, 475, 474, 498, 487, 503, 497, 495, 445, 387, 382, 438, 518, 520, 523, 520, 520, 520, 520, 522, 
    403, 353, 355, 373, 443, 453, 461, 466, 470, 474, 457, 465, 452, 459, 439, 454, 473, 459, 384, 334, 346, 428, 511, 510, 508, 501, 495, 503, 509, 513, 
    394, 334, 338, 348, 427, 438, 453, 458, 457, 458, 445, 456, 430, 415, 377, 382, 413, 413, 349, 288, 281, 357, 441, 460, 475, 473, 463, 478, 486, 492, 
    387, 324, 331, 342, 418, 429, 443, 449, 443, 443, 431, 440, 420, 411, 362, 333, 295, 245, 191, 158, 135, 140, 190, 268, 361, 430, 435, 440, 445, 446, 
    341, 292, 298, 309, 359, 372, 384, 401, 401, 403, 402, 406, 390, 385, 350, 298, 220, 161, 116, 114, 108, 77, 75, 105, 207, 314, 346, 342, 351, 349, 
    220, 197, 199, 194, 214, 227, 246, 272, 280, 288, 298, 303, 303, 305, 283, 244, 186, 162, 149, 141, 128, 110, 132, 137, 197, 235, 237, 212, 204, 206, 
    101, 96, 106, 106, 113, 126, 130, 150, 158, 170, 178, 188, 206, 216, 204, 184, 159, 151, 138, 119, 119, 120, 151, 163, 205, 239, 226, 194, 134, 124, 
    60, 72, 100, 116, 129, 105, 95, 118, 136, 148, 150, 171, 200, 206, 192, 169, 156, 147, 137, 121, 149, 200, 268, 249, 207, 235, 233, 229, 140, 101, 
    86, 98, 122, 130, 139, 121, 121, 164, 207, 207, 192, 200, 216, 207, 179, 156, 147, 146, 149, 156, 203, 270, 354, 354, 282, 253, 223, 217, 147, 83, 
    118, 122, 119, 95, 104, 98, 121, 168, 208, 227, 223, 217, 217, 211, 191, 171, 163, 171, 179, 202, 254, 303, 351, 356, 315, 268, 223, 174, 126, 46, 
    129, 119, 114, 93, 87, 102, 143, 186, 225, 251, 271, 276, 275, 272, 272, 268, 272, 272, 264, 273, 297, 317, 336, 326, 305, 248, 178, 90, 65, 10, 
    170, 163, 169, 176, 197, 223, 248, 285, 315, 328, 339, 349, 353, 344, 339, 337, 340, 328, 285, 261, 249, 269, 293, 302, 299, 235, 160, 59, 38, 34, 
    217, 225, 240, 256, 284, 316, 336, 349, 362, 370, 374, 374, 372, 360, 339, 317, 307, 291, 236, 197, 184, 220, 264, 284, 295, 248, 218, 188, 178, 165, 
    237, 240, 239, 234, 256, 300, 345, 364, 371, 368, 358, 342, 323, 303, 283, 272, 276, 275, 248, 223, 216, 248, 274, 277, 286, 260, 253, 256, 264, 252, 
    203, 187, 176, 188, 223, 278, 327, 344, 337, 319, 303, 290, 280, 277, 276, 275, 284, 291, 287, 284, 280, 291, 293, 284, 282, 263, 250, 229, 206, 212, 
    161, 157, 185, 238, 279, 295, 295, 290, 284, 278, 284, 294, 301, 306, 304, 294, 293, 289, 297, 303, 300, 304, 301, 284, 256, 223, 183, 134, 113, 142, 
    195, 202, 237, 274, 290, 288, 274, 269, 274, 292, 305, 311, 305, 288, 254, 216, 223, 245, 283, 300, 298, 294, 268, 228, 182, 138, 94, 62, 47, 55, 
    243, 257, 265, 270, 273, 277, 268, 262, 267, 285, 292, 292, 256, 200, 135, 88, 122, 186, 257, 275, 255, 226, 186, 145, 101, 67, 43, 29, 15, 1, 
    223, 260, 268, 266, 257, 239, 214, 198, 183, 205, 233, 262, 236, 172, 103, 74, 110, 148, 192, 191, 165, 139, 102, 74, 45, 18, 0, 0, 0, 0, 
    179, 232, 246, 243, 210, 165, 117, 106, 106, 143, 195, 249, 241, 195, 141, 108, 114, 114, 117, 112, 94, 71, 43, 20, 0, 0, 0, 0, 0, 0, 
    157, 203, 223, 227, 196, 151, 107, 107, 129, 159, 180, 189, 162, 130, 106, 90, 91, 86, 81, 63, 39, 18, 7, 0, 0, 0, 0, 0, 0, 0, 
    152, 190, 209, 205, 182, 155, 124, 110, 103, 103, 97, 89, 76, 67, 65, 63, 63, 54, 39, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    92, 109, 116, 101, 79, 68, 57, 48, 41, 33, 29, 33, 39, 43, 38, 24, 11, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=46
    60, 47, 110, 138, 109, 97, 103, 108, 100, 86, 98, 105, 96, 95, 72, 81, 102, 101, 98, 87, 92, 100, 94, 77, 82, 100, 85, 74, 95, 98, 
    68, 49, 109, 140, 113, 92, 97, 111, 99, 81, 99, 111, 102, 104, 80, 80, 100, 104, 102, 96, 122, 124, 100, 78, 84, 106, 86, 73, 103, 105, 
    62, 46, 106, 137, 113, 88, 89, 109, 93, 73, 90, 107, 98, 108, 90, 80, 99, 101, 72, 73, 141, 141, 105, 78, 82, 108, 90, 72, 103, 103, 
    55, 40, 103, 131, 109, 85, 81, 106, 90, 67, 81, 102, 88, 109, 111, 94, 108, 97, 34, 54, 148, 143, 109, 80, 79, 108, 92, 78, 104, 97, 
    57, 36, 103, 132, 108, 84, 72, 98, 84, 67, 78, 96, 71, 90, 120, 111, 126, 98, 11, 64, 173, 159, 134, 100, 78, 103, 91, 87, 109, 95, 
    54, 25, 99, 129, 103, 86, 77, 94, 76, 68, 79, 92, 55, 50, 84, 95, 139, 133, 45, 85, 188, 202, 213, 186, 120, 104, 86, 82, 111, 96, 
    64, 27, 100, 133, 110, 103, 102, 102, 80, 77, 88, 92, 60, 49, 53, 60, 98, 114, 82, 82, 116, 124, 174, 227, 189, 143, 105, 91, 127, 114, 
    104, 65, 122, 159, 138, 142, 147, 135, 113, 113, 119, 111, 99, 106, 69, 39, 36, 31, 26, 23, 25, 0, 26, 113, 151, 151, 116, 102, 150, 139, 
    116, 87, 111, 129, 111, 126, 143, 137, 126, 128, 136, 125, 123, 124, 78, 47, 52, 57, 51, 56, 66, 32, 34, 47, 76, 93, 43, 40, 115, 116, 
    82, 57, 61, 58, 40, 58, 84, 91, 77, 74, 89, 86, 91, 89, 62, 52, 62, 63, 49, 46, 58, 37, 36, 16, 47, 94, 3, 0, 40, 62, 
    52, 26, 50, 57, 24, 25, 52, 65, 31, 18, 45, 64, 67, 61, 53, 51, 54, 51, 31, 15, 53, 62, 19, 0, 0, 98, 56, 0, 10, 54, 
    57, 30, 69, 90, 52, 41, 72, 92, 62, 34, 49, 81, 79, 60, 57, 55, 54, 57, 43, 29, 81, 107, 81, 30, 0, 47, 88, 0, 0, 66, 
    72, 39, 56, 69, 56, 67, 93, 104, 97, 68, 49, 59, 55, 35, 26, 22, 18, 29, 29, 37, 82, 92, 91, 82, 9, 12, 86, 19, 3, 66, 
    54, 32, 30, 25, 19, 33, 50, 53, 56, 53, 43, 42, 40, 31, 35, 39, 28, 30, 35, 63, 99, 93, 83, 75, 49, 0, 31, 32, 8, 29, 
    47, 35, 23, 32, 28, 31, 52, 66, 68, 69, 72, 73, 71, 63, 76, 95, 93, 77, 60, 85, 112, 102, 90, 67, 59, 0, 0, 0, 0, 0, 
    75, 72, 66, 95, 117, 110, 99, 100, 101, 98, 98, 100, 101, 94, 87, 98, 103, 72, 18, 34, 67, 70, 75, 67, 64, 14, 0, 4, 0, 0, 
    98, 107, 104, 111, 135, 133, 113, 105, 108, 110, 109, 106, 98, 87, 67, 62, 74, 54, 0, 9, 47, 50, 60, 63, 63, 45, 47, 87, 78, 34, 
    98, 99, 82, 69, 85, 107, 117, 112, 110, 104, 93, 80, 66, 56, 50, 47, 70, 77, 45, 47, 68, 61, 56, 57, 63, 63, 71, 81, 94, 107, 
    45, 62, 70, 78, 81, 88, 98, 95, 84, 73, 67, 67, 69, 73, 85, 84, 99, 104, 76, 67, 75, 76, 66, 68, 77, 73, 67, 62, 77, 125, 
    38, 70, 95, 104, 100, 83, 70, 79, 86, 84, 85, 87, 86, 93, 107, 110, 137, 134, 88, 73, 81, 89, 80, 71, 68, 56, 43, 39, 48, 86, 
    99, 85, 82, 83, 88, 86, 82, 107, 126, 126, 114, 89, 53, 40, 56, 58, 108, 137, 104, 90, 92, 86, 69, 54, 49, 41, 36, 45, 40, 31, 
    130, 95, 88, 89, 86, 93, 105, 115, 116, 130, 126, 87, 22, 0, 3, 17, 70, 113, 100, 86, 74, 59, 50, 52, 49, 37, 42, 49, 32, 13, 
    128, 100, 92, 88, 52, 43, 65, 68, 57, 90, 117, 102, 64, 39, 44, 50, 66, 74, 64, 56, 54, 52, 42, 40, 33, 29, 34, 27, 17, 12, 
    108, 87, 81, 80, 33, 11, 35, 49, 56, 90, 114, 111, 95, 79, 68, 56, 53, 54, 52, 50, 48, 44, 36, 31, 19, 25, 28, 18, 13, 11, 
    115, 106, 102, 108, 84, 68, 78, 83, 85, 92, 87, 72, 58, 49, 49, 52, 62, 66, 54, 38, 31, 31, 49, 46, 22, 23, 28, 21, 17, 15, 
    125, 124, 116, 110, 98, 90, 84, 70, 52, 43, 42, 48, 57, 60, 57, 52, 52, 44, 28, 28, 33, 33, 45, 40, 23, 22, 25, 21, 18, 21, 
    74, 73, 71, 63, 52, 50, 54, 52, 49, 50, 51, 52, 55, 51, 38, 33, 40, 26, 11, 28, 33, 29, 32, 27, 22, 23, 23, 20, 20, 16, 
    23, 26, 35, 37, 35, 38, 48, 51, 47, 43, 39, 35, 32, 28, 20, 37, 71, 38, 4, 23, 32, 27, 26, 24, 23, 24, 23, 22, 16, 7, 
    18, 18, 24, 25, 24, 24, 26, 27, 24, 21, 23, 28, 32, 31, 26, 47, 84, 39, 0, 23, 31, 26, 25, 23, 25, 28, 26, 23, 4, 0, 
    15, 13, 16, 17, 16, 18, 20, 23, 28, 31, 35, 37, 39, 38, 33, 55, 91, 41, 3, 24, 27, 25, 24, 23, 25, 29, 30, 14, 0, 0, 
    
    -- channel=47
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=48
    0, 0, 0, 2, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 42, 6, 0, 4, 4, 10, 19, 10, 0, 2, 7, 2, 2, 5, 3, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 43, 3, 16, 28, 9, 19, 20, 12, 0, 7, 11, 2, 5, 10, 2, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 27, 28, 0, 22, 19, 0, 20, 21, 12, 1, 1, 1, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 42, 35, 0, 16, 17, 3, 23, 23, 12, 4, 6, 8, 0, 18, 8, 4, 0, 6, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 39, 24, 2, 7, 11, 5, 8, 14, 6, 3, 8, 5, 1, 21, 9, 2, 0, 0, 15, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 9, 18, 18, 10, 9, 6, 9, 11, 5, 3, 5, 4, 6, 19, 10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 15, 17, 3, 7, 2, 7, 0, 0, 0, 0, 0, 3, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17, 42, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 22, 38, 43, 25, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 30, 52, 40, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 28, 75, 56, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 80, 106, 48, 25, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 62, 126, 75, 43, 43, 31, 22, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 61, 149, 99, 57, 58, 45, 40, 40, 38, 35, 33, 37, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 83, 160, 122, 73, 62, 53, 48, 47, 49, 52, 61, 77, 73, 36, 16, 14, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 20, 94, 98, 87, 90, 64, 63, 45, 13, 16, 34, 65, 62, 49, 42, 43, 53, 16, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 34, 0, 10, 61, 51, 30, 6, 0, 0, 0, 45, 38, 0, 0, 27, 30, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 11, 0, 0, 0, 0, 0, 22, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 13, 19, 23, 25, 26, 28, 30, 28, 37, 49, 37, 27, 15, 7, 23, 36, 39, 26, 21, 24, 25, 20, 17, 24, 30, 31, 27, 20, 28, 
    32, 40, 51, 53, 53, 51, 52, 54, 50, 51, 56, 54, 51, 45, 34, 41, 50, 45, 45, 47, 47, 44, 43, 45, 46, 44, 48, 48, 46, 47, 
    29, 33, 39, 42, 44, 43, 44, 43, 41, 46, 47, 46, 44, 43, 41, 45, 56, 56, 52, 54, 58, 58, 53, 53, 53, 55, 61, 68, 62, 46, 
    55, 50, 56, 59, 63, 66, 61, 58, 61, 65, 65, 67, 66, 65, 62, 61, 69, 72, 70, 70, 71, 68, 68, 68, 68, 69, 74, 73, 51, 22, 
    73, 61, 68, 68, 71, 72, 64, 63, 70, 72, 71, 69, 65, 64, 60, 59, 63, 68, 69, 67, 63, 63, 66, 68, 68, 67, 58, 38, 10, 0, 
    74, 64, 70, 66, 68, 67, 60, 63, 70, 71, 67, 65, 66, 63, 59, 58, 64, 69, 66, 63, 61, 61, 62, 64, 62, 47, 22, 1, 0, 26, 
    74, 63, 70, 66, 68, 67, 62, 66, 66, 59, 54, 54, 58, 56, 48, 50, 56, 57, 56, 60, 60, 59, 61, 54, 36, 11, 0, 13, 55, 71, 
    74, 62, 65, 61, 64, 65, 64, 64, 63, 50, 42, 51, 56, 54, 46, 47, 52, 50, 52, 63, 67, 60, 54, 34, 6, 0, 24, 72, 82, 57, 
    
    -- channel=49
    204, 237, 248, 252, 238, 218, 206, 202, 207, 216, 223, 222, 221, 221, 219, 216, 214, 216, 219, 221, 222, 222, 222, 220, 218, 216, 218, 225, 234, 227, 
    220, 258, 269, 276, 248, 187, 161, 143, 151, 178, 185, 184, 180, 175, 172, 175, 179, 176, 176, 178, 185, 183, 190, 190, 204, 222, 232, 242, 249, 243, 
    219, 260, 268, 276, 258, 187, 144, 101, 110, 134, 131, 137, 136, 135, 128, 127, 134, 140, 140, 144, 149, 143, 167, 182, 214, 245, 244, 242, 244, 236, 
    222, 261, 271, 280, 262, 198, 143, 60, 67, 99, 88, 103, 103, 84, 88, 94, 112, 116, 120, 129, 129, 125, 143, 171, 226, 252, 245, 246, 247, 239, 
    221, 257, 266, 279, 252, 192, 143, 72, 98, 97, 76, 75, 69, 53, 71, 84, 100, 95, 101, 107, 100, 110, 106, 130, 196, 234, 243, 247, 249, 237, 
    219, 257, 266, 268, 223, 148, 97, 83, 123, 114, 113, 111, 102, 77, 92, 110, 134, 126, 125, 132, 122, 140, 132, 155, 191, 220, 251, 257, 256, 244, 
    218, 254, 263, 260, 216, 143, 73, 64, 118, 119, 126, 126, 119, 97, 99, 109, 122, 123, 125, 113, 115, 137, 129, 139, 154, 202, 249, 258, 259, 249, 
    221, 255, 258, 262, 245, 192, 135, 125, 146, 158, 156, 158, 169, 155, 147, 146, 148, 147, 146, 127, 129, 150, 157, 160, 151, 199, 251, 258, 258, 250, 
    225, 258, 257, 268, 265, 242, 229, 227, 215, 218, 221, 221, 226, 219, 215, 218, 222, 225, 223, 212, 208, 220, 224, 225, 223, 239, 254, 257, 259, 251, 
    233, 259, 254, 265, 267, 263, 260, 244, 228, 226, 224, 223, 216, 214, 215, 218, 228, 235, 231, 219, 217, 218, 221, 243, 257, 255, 254, 258, 262, 251, 
    235, 262, 255, 260, 258, 251, 247, 239, 228, 230, 223, 217, 218, 220, 223, 225, 223, 222, 226, 225, 221, 222, 225, 244, 259, 257, 255, 257, 258, 246, 
    236, 264, 258, 264, 251, 236, 232, 235, 240, 248, 252, 251, 250, 252, 255, 256, 256, 255, 255, 254, 250, 250, 253, 256, 257, 256, 252, 249, 251, 241, 
    233, 267, 254, 239, 209, 186, 210, 235, 237, 237, 240, 247, 251, 254, 256, 256, 254, 251, 250, 248, 247, 250, 252, 251, 252, 255, 254, 256, 259, 248, 
    234, 271, 250, 217, 183, 145, 128, 155, 191, 221, 235, 234, 239, 246, 251, 252, 251, 251, 251, 249, 247, 252, 257, 259, 258, 258, 256, 257, 260, 250, 
    234, 270, 262, 264, 253, 217, 153, 115, 123, 142, 182, 214, 225, 233, 244, 250, 252, 253, 252, 247, 244, 247, 249, 250, 250, 252, 252, 254, 258, 250, 
    231, 268, 259, 259, 256, 251, 237, 187, 138, 112, 117, 161, 205, 228, 231, 232, 235, 239, 245, 247, 246, 247, 252, 253, 255, 258, 257, 257, 260, 251, 
    227, 263, 254, 256, 254, 249, 252, 242, 185, 110, 86, 97, 120, 165, 206, 223, 224, 222, 224, 232, 236, 241, 247, 249, 252, 256, 255, 256, 260, 249, 
    223, 258, 249, 255, 256, 252, 247, 249, 221, 127, 78, 83, 78, 84, 108, 148, 185, 210, 223, 225, 219, 220, 228, 233, 239, 246, 249, 253, 256, 245, 
    220, 254, 244, 250, 252, 252, 244, 253, 222, 134, 90, 85, 79, 79, 74, 77, 93, 121, 157, 184, 197, 213, 227, 227, 223, 228, 229, 233, 243, 238, 
    220, 253, 245, 250, 252, 251, 248, 253, 206, 110, 76, 81, 69, 76, 76, 84, 97, 99, 96, 77, 85, 120, 158, 185, 201, 226, 241, 240, 242, 239, 
    222, 254, 246, 247, 251, 252, 253, 230, 168, 114, 82, 76, 85, 90, 92, 98, 105, 113, 118, 100, 80, 81, 99, 102, 113, 142, 170, 201, 231, 241, 
    217, 249, 245, 242, 246, 249, 248, 214, 166, 168, 168, 116, 83, 75, 80, 137, 188, 189, 141, 114, 141, 142, 116, 95, 121, 180, 201, 199, 216, 229, 
    211, 237, 236, 235, 237, 237, 237, 236, 236, 244, 247, 212, 179, 175, 179, 213, 249, 257, 230, 204, 217, 231, 224, 207, 216, 239, 251, 251, 251, 244, 
    210, 239, 236, 234, 235, 233, 230, 230, 228, 230, 231, 229, 227, 226, 227, 227, 227, 226, 229, 233, 230, 229, 233, 239, 236, 227, 218, 215, 219, 216, 
    131, 143, 144, 138, 137, 132, 127, 123, 117, 117, 119, 116, 115, 116, 127, 146, 157, 156, 155, 155, 157, 158, 161, 165, 169, 171, 167, 162, 167, 163, 
    130, 136, 136, 136, 138, 139, 140, 136, 135, 136, 133, 132, 133, 135, 134, 136, 141, 137, 133, 135, 135, 132, 131, 135, 137, 138, 137, 134, 139, 139, 
    121, 122, 125, 126, 127, 121, 111, 105, 105, 102, 100, 101, 98, 94, 95, 94, 95, 91, 84, 81, 80, 78, 77, 75, 75, 78, 82, 92, 107, 113, 
    74, 66, 71, 69, 71, 73, 67, 66, 68, 66, 63, 61, 64, 65, 65, 67, 72, 76, 72, 67, 66, 67, 68, 67, 70, 81, 93, 108, 121, 127, 
    78, 72, 77, 74, 76, 75, 71, 74, 75, 71, 68, 71, 70, 68, 68, 69, 75, 75, 72, 70, 69, 66, 67, 72, 81, 101, 119, 130, 144, 150, 
    69, 63, 69, 64, 65, 64, 62, 63, 62, 60, 55, 58, 62, 61, 59, 62, 64, 61, 58, 60, 64, 65, 72, 88, 106, 121, 134, 152, 153, 104, 
    
    -- channel=50
    66, 91, 86, 91, 95, 75, 61, 61, 64, 69, 69, 70, 65, 70, 66, 63, 66, 64, 67, 66, 64, 67, 65, 65, 63, 57, 56, 61, 68, 54, 
    79, 110, 108, 105, 93, 53, 30, 22, 21, 38, 42, 39, 35, 40, 36, 32, 37, 35, 37, 40, 36, 39, 50, 51, 61, 68, 74, 75, 76, 62, 
    80, 110, 107, 108, 101, 55, 33, 0, 0, 9, 5, 5, 8, 10, 4, 0, 4, 4, 6, 13, 11, 8, 34, 30, 55, 79, 76, 73, 73, 59, 
    84, 110, 109, 113, 106, 55, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 10, 8, 2, 22, 18, 58, 83, 77, 74, 77, 61, 
    82, 105, 108, 115, 99, 48, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 47, 70, 80, 81, 80, 61, 
    82, 106, 106, 109, 80, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 3, 0, 16, 3, 26, 40, 51, 78, 82, 85, 68, 
    81, 106, 105, 103, 85, 41, 0, 0, 3, 12, 19, 9, 10, 0, 0, 2, 13, 12, 9, 6, 0, 18, 4, 26, 19, 39, 84, 90, 89, 73, 
    81, 107, 104, 108, 97, 55, 7, 17, 30, 38, 36, 32, 43, 37, 32, 24, 25, 28, 23, 17, 11, 28, 31, 35, 26, 53, 85, 88, 90, 76, 
    79, 109, 102, 107, 103, 88, 79, 85, 74, 78, 78, 78, 82, 77, 74, 69, 75, 80, 78, 73, 65, 76, 77, 65, 67, 79, 89, 89, 92, 78, 
    76, 108, 97, 104, 109, 104, 100, 98, 83, 86, 85, 81, 79, 75, 75, 77, 81, 84, 81, 79, 73, 75, 79, 80, 90, 90, 91, 91, 94, 77, 
    73, 103, 91, 98, 109, 101, 88, 85, 80, 81, 79, 75, 75, 73, 74, 74, 75, 76, 77, 78, 74, 74, 80, 87, 92, 90, 88, 86, 89, 71, 
    71, 98, 99, 104, 107, 95, 84, 91, 92, 92, 92, 91, 91, 90, 90, 90, 90, 89, 90, 90, 88, 86, 87, 89, 89, 87, 85, 84, 86, 69, 
    68, 98, 97, 86, 75, 73, 76, 84, 87, 89, 90, 89, 88, 87, 87, 87, 86, 84, 85, 85, 85, 85, 86, 88, 89, 89, 89, 89, 90, 74, 
    67, 95, 82, 68, 51, 44, 43, 54, 72, 81, 84, 82, 80, 80, 83, 83, 83, 82, 83, 84, 83, 84, 89, 91, 90, 90, 90, 90, 93, 77, 
    65, 97, 90, 86, 72, 53, 32, 32, 49, 57, 64, 72, 76, 78, 81, 82, 83, 82, 82, 82, 81, 81, 84, 87, 86, 88, 89, 89, 94, 80, 
    63, 94, 84, 84, 81, 72, 53, 43, 56, 48, 44, 59, 69, 74, 76, 77, 77, 78, 79, 81, 82, 82, 85, 87, 87, 90, 90, 90, 96, 81, 
    60, 88, 77, 79, 79, 75, 69, 50, 65, 50, 20, 31, 42, 56, 66, 71, 74, 75, 76, 83, 84, 79, 82, 83, 85, 88, 90, 90, 94, 80, 
    55, 83, 72, 76, 77, 75, 72, 50, 75, 63, 17, 22, 19, 24, 35, 48, 60, 70, 77, 89, 86, 78, 80, 80, 81, 84, 85, 85, 90, 77, 
    54, 80, 69, 74, 76, 75, 65, 62, 85, 64, 27, 26, 17, 14, 11, 15, 26, 42, 60, 78, 83, 77, 79, 80, 77, 78, 81, 81, 83, 75, 
    55, 80, 72, 74, 76, 76, 68, 82, 72, 32, 19, 24, 18, 25, 17, 7, 7, 11, 30, 32, 34, 40, 58, 76, 68, 70, 76, 74, 78, 74, 
    58, 83, 74, 73, 77, 78, 72, 73, 36, 3, 16, 32, 20, 25, 6, 0, 5, 20, 41, 13, 7, 15, 26, 30, 13, 27, 51, 59, 70, 71, 
    59, 84, 75, 73, 78, 76, 69, 58, 40, 32, 41, 40, 13, 15, 13, 23, 48, 52, 52, 26, 30, 34, 32, 28, 30, 54, 69, 69, 75, 74, 
    69, 91, 86, 83, 86, 88, 87, 88, 91, 88, 89, 83, 71, 72, 75, 84, 99, 99, 92, 85, 90, 91, 89, 87, 94, 103, 108, 104, 100, 90, 
    81, 96, 95, 92, 95, 93, 91, 93, 92, 88, 94, 95, 95, 94, 91, 90, 98, 101, 101, 102, 102, 102, 104, 105, 105, 102, 100, 99, 97, 87, 
    46, 54, 51, 47, 48, 45, 43, 41, 38, 42, 45, 44, 46, 49, 56, 59, 67, 70, 68, 69, 70, 73, 73, 75, 77, 78, 77, 77, 75, 73, 
    49, 53, 50, 53, 57, 57, 56, 51, 49, 50, 50, 51, 52, 52, 54, 53, 54, 54, 52, 53, 54, 54, 53, 54, 55, 55, 53, 53, 60, 54, 
    47, 44, 44, 43, 42, 42, 37, 29, 29, 31, 33, 32, 31, 29, 29, 27, 24, 25, 24, 24, 22, 20, 19, 20, 20, 21, 25, 31, 31, 24, 
    21, 15, 18, 16, 16, 18, 13, 9, 12, 12, 14, 13, 12, 12, 11, 11, 13, 17, 16, 13, 13, 12, 14, 14, 15, 25, 33, 29, 29, 45, 
    23, 16, 22, 20, 19, 19, 15, 16, 17, 18, 15, 13, 12, 12, 10, 8, 13, 14, 12, 10, 12, 11, 12, 17, 28, 35, 31, 38, 60, 62, 
    14, 8, 16, 14, 13, 12, 11, 9, 8, 8, 3, 6, 8, 7, 5, 3, 7, 5, 6, 6, 12, 10, 13, 24, 28, 31, 48, 69, 61, 30, 
    
    -- channel=51
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=52
    96, 85, 96, 92, 73, 77, 85, 91, 91, 89, 90, 90, 90, 87, 88, 89, 85, 86, 87, 87, 90, 91, 92, 92, 92, 95, 103, 109, 112, 118, 
    85, 77, 87, 93, 80, 81, 108, 126, 118, 113, 118, 113, 120, 117, 113, 114, 113, 112, 109, 110, 113, 111, 116, 103, 87, 97, 110, 110, 109, 117, 
    84, 81, 89, 94, 90, 92, 107, 102, 111, 133, 141, 139, 140, 140, 135, 140, 144, 142, 143, 145, 142, 137, 142, 130, 108, 107, 114, 115, 113, 119, 
    83, 79, 86, 87, 94, 112, 100, 84, 100, 105, 94, 95, 101, 101, 99, 100, 91, 93, 93, 90, 92, 95, 84, 99, 105, 103, 105, 109, 109, 115, 
    83, 82, 85, 83, 94, 121, 122, 130, 123, 105, 104, 117, 124, 116, 117, 119, 119, 114, 117, 116, 114, 125, 101, 126, 140, 118, 106, 112, 113, 119, 
    79, 79, 86, 84, 96, 123, 112, 132, 128, 112, 122, 121, 111, 117, 122, 129, 128, 130, 140, 135, 137, 136, 114, 128, 138, 123, 112, 113, 113, 119, 
    76, 76, 86, 82, 93, 94, 69, 94, 92, 88, 90, 88, 83, 93, 93, 93, 83, 93, 95, 90, 99, 88, 105, 91, 82, 102, 107, 105, 104, 112, 
    75, 74, 84, 83, 91, 81, 86, 100, 95, 98, 94, 106, 102, 100, 100, 103, 97, 98, 106, 100, 107, 102, 124, 91, 78, 100, 104, 103, 100, 107, 
    81, 72, 82, 84, 86, 85, 93, 88, 88, 88, 88, 94, 85, 83, 85, 91, 94, 95, 94, 87, 94, 92, 97, 98, 101, 103, 100, 102, 101, 107, 
    91, 76, 83, 78, 83, 92, 87, 64, 65, 63, 63, 62, 60, 63, 65, 69, 69, 67, 64, 65, 72, 71, 70, 93, 103, 101, 101, 104, 102, 107, 
    105, 84, 92, 99, 112, 121, 106, 79, 77, 80, 78, 81, 82, 85, 88, 88, 86, 84, 86, 85, 88, 86, 86, 98, 100, 100, 99, 100, 98, 105, 
    109, 89, 94, 97, 93, 110, 143, 142, 120, 99, 91, 93, 95, 99, 98, 97, 96, 95, 94, 93, 94, 96, 97, 96, 98, 101, 102, 103, 103, 111, 
    111, 100, 80, 53, 30, 32, 83, 126, 144, 139, 118, 103, 98, 98, 99, 101, 100, 101, 100, 101, 102, 104, 104, 104, 104, 104, 106, 108, 107, 113, 
    113, 106, 92, 79, 73, 36, 10, 33, 82, 118, 132, 124, 110, 103, 104, 106, 107, 110, 108, 104, 104, 105, 103, 101, 99, 99, 100, 101, 100, 106, 
    112, 103, 105, 104, 110, 98, 56, 20, 29, 68, 104, 135, 150, 140, 121, 110, 106, 106, 106, 103, 102, 103, 103, 101, 100, 99, 98, 97, 96, 103, 
    113, 106, 110, 105, 110, 117, 119, 74, 29, 38, 62, 90, 125, 153, 159, 148, 129, 113, 105, 102, 104, 103, 101, 100, 101, 102, 100, 100, 99, 103, 
    116, 111, 119, 115, 116, 115, 127, 113, 54, 39, 52, 57, 70, 94, 123, 147, 160, 159, 145, 131, 119, 106, 99, 98, 100, 100, 101, 103, 100, 104, 
    120, 113, 122, 119, 119, 118, 114, 123, 88, 55, 68, 68, 62, 60, 66, 79, 101, 126, 146, 154, 156, 156, 144, 131, 118, 106, 99, 99, 98, 102, 
    124, 112, 120, 120, 118, 117, 110, 139, 108, 42, 53, 59, 57, 62, 61, 56, 57, 60, 68, 71, 90, 122, 146, 164, 165, 156, 142, 125, 109, 107, 
    130, 113, 117, 118, 118, 115, 118, 131, 78, 3, 0, 17, 46, 62, 68, 44, 19, 15, 35, 28, 7, 30, 69, 97, 100, 91, 99, 112, 111, 116, 
    126, 110, 113, 113, 115, 116, 127, 84, 38, 20, 0, 0, 0, 0, 9, 32, 38, 29, 9, 5, 3, 0, 0, 0, 23, 53, 65, 77, 89, 105, 
    126, 113, 116, 121, 122, 127, 133, 106, 98, 115, 92, 37, 28, 18, 37, 88, 113, 105, 46, 46, 71, 67, 43, 21, 59, 96, 100, 102, 103, 110, 
    156, 147, 150, 155, 155, 156, 155, 155, 155, 161, 155, 129, 127, 123, 121, 128, 126, 123, 102, 103, 109, 112, 104, 96, 99, 100, 98, 100, 102, 110, 
    96, 88, 87, 83, 79, 75, 72, 72, 68, 71, 70, 65, 63, 62, 70, 76, 72, 72, 77, 77, 75, 79, 84, 86, 82, 77, 73, 79, 85, 95, 
    72, 67, 63, 62, 59, 60, 66, 67, 66, 71, 67, 63, 63, 62, 67, 76, 77, 77, 79, 81, 82, 80, 81, 85, 87, 88, 89, 87, 85, 86, 
    94, 88, 90, 92, 85, 82, 82, 80, 82, 84, 82, 80, 75, 75, 72, 76, 75, 67, 67, 69, 68, 63, 60, 60, 62, 64, 65, 59, 57, 44, 
    62, 56, 60, 62, 60, 59, 57, 58, 59, 56, 53, 48, 47, 50, 51, 53, 53, 51, 49, 46, 46, 48, 49, 48, 47, 45, 44, 38, 22, 25, 
    54, 47, 50, 50, 50, 49, 48, 53, 54, 52, 49, 45, 44, 47, 50, 49, 52, 52, 48, 45, 43, 44, 48, 47, 44, 40, 31, 17, 30, 80, 
    51, 45, 45, 45, 44, 42, 43, 47, 47, 46, 37, 33, 35, 39, 40, 43, 43, 38, 35, 35, 40, 44, 44, 45, 44, 29, 18, 46, 87, 88, 
    51, 49, 49, 50, 49, 45, 47, 50, 49, 50, 51, 55, 55, 53, 55, 62, 60, 56, 54, 53, 51, 51, 48, 44, 32, 34, 69, 94, 77, 53, 
    
    -- channel=53
    0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 26, 18, 14, 18, 14, 15, 15, 14, 12, 9, 12, 8, 2, 8, 10, 9, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 18, 0, 4, 24, 20, 26, 23, 21, 18, 26, 27, 22, 21, 28, 22, 32, 18, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 55, 20, 16, 23, 2, 2, 15, 17, 19, 13, 14, 14, 2, 18, 10, 10, 9, 0, 9, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 39, 10, 24, 16, 7, 17, 19, 4, 3, 7, 29, 12, 17, 34, 14, 29, 3, 6, 27, 9, 2, 3, 1, 0, 
    0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 17, 0, 0, 0, 2, 1, 0, 7, 3, 4, 4, 0, 0, 6, 6, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 8, 0, 2, 0, 2, 4, 0, 1, 2, 1, 0, 8, 1, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 20, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 21, 31, 26, 23, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 37, 38, 22, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 10, 0, 0, 0, 0, 0, 5, 29, 27, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 17, 16, 0, 0, 0, 0, 18, 29, 24, 12, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 13, 0, 0, 0, 0, 3, 30, 38, 31, 19, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 11, 7, 6, 0, 0, 0, 5, 29, 41, 41, 32, 18, 12, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 30, 30, 5, 10, 0, 0, 0, 0, 16, 32, 40, 50, 45, 29, 21, 11, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 46, 31, 8, 15, 7, 7, 1, 0, 0, 0, 0, 13, 26, 37, 44, 45, 39, 28, 17, 8, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 30, 47, 0, 0, 0, 0, 9, 4, 0, 0, 0, 0, 0, 0, 0, 0, 16, 11, 7, 10, 10, 7, 2, 
    0, 0, 0, 0, 0, 0, 1, 30, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 2, 1, 1, 8, 32, 22, 0, 5, 13, 0, 0, 0, 0, 0, 4, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 27, 27, 29, 30, 32, 33, 32, 34, 42, 59, 41, 24, 16, 0, 4, 25, 43, 23, 3, 12, 25, 20, 0, 0, 5, 12, 16, 17, 14, 
    1, 6, 11, 9, 9, 8, 4, 6, 6, 2, 6, 6, 7, 12, 13, 11, 10, 8, 12, 16, 12, 12, 16, 21, 23, 17, 12, 13, 19, 24, 
    0, 3, 7, 4, 6, 5, 8, 11, 6, 9, 12, 7, 6, 0, 4, 11, 15, 19, 19, 18, 18, 21, 20, 22, 24, 25, 21, 25, 25, 26, 
    19, 20, 20, 21, 18, 18, 21, 18, 16, 18, 17, 17, 18, 17, 15, 15, 16, 13, 11, 14, 16, 12, 9, 9, 10, 10, 16, 17, 13, 3, 
    10, 5, 8, 11, 11, 12, 11, 5, 7, 6, 6, 7, 4, 5, 3, 5, 6, 4, 3, 3, 3, 2, 1, 1, 2, 4, 2, 3, 0, 0, 
    10, 1, 4, 3, 3, 6, 2, 0, 5, 4, 4, 0, 1, 1, 2, 0, 0, 6, 5, 1, 0, 0, 1, 4, 4, 3, 1, 0, 0, 0, 
    11, 0, 2, 2, 2, 2, 0, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 0, 26, 
    11, 3, 6, 2, 4, 3, 2, 4, 7, 12, 0, 0, 1, 2, 2, 1, 5, 2, 0, 0, 1, 3, 0, 5, 0, 0, 0, 0, 35, 19, 
    
    -- channel=54
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 11, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 16, 18, 19, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 17, 20, 19, 21, 27, 23, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 30, 28, 26, 22, 19, 18, 21, 29, 39, 38, 30, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 20, 31, 24, 17, 18, 14, 14, 17, 18, 23, 29, 36, 36, 35, 27, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 21, 12, 0, 0, 0, 0, 5, 0, 0, 13, 18, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 9, 8, 14, 17, 20, 21, 23, 24, 23, 17, 19, 18, 15, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 4, 5, 6, 10, 8, 11, 13, 14, 19, 21, 23, 23, 24, 25, 25, 25, 28, 27, 28, 23, 
    29, 29, 28, 29, 28, 27, 28, 31, 31, 31, 34, 33, 31, 30, 29, 27, 28, 27, 28, 31, 30, 29, 27, 26, 28, 29, 29, 26, 17, 1, 
    22, 22, 22, 22, 21, 21, 21, 23, 23, 26, 24, 22, 23, 24, 24, 22, 21, 23, 24, 24, 23, 23, 24, 24, 24, 22, 18, 6, 0, 0, 
    23, 22, 20, 26, 24, 22, 23, 25, 25, 26, 25, 23, 20, 22, 22, 23, 23, 24, 24, 24, 22, 23, 23, 24, 21, 14, 0, 0, 0, 18, 
    20, 21, 18, 19, 17, 18, 20, 20, 21, 20, 13, 5, 7, 9, 10, 11, 7, 7, 6, 10, 14, 22, 22, 20, 12, 0, 0, 0, 27, 29, 
    22, 26, 26, 25, 22, 21, 22, 23, 24, 21, 23, 19, 18, 19, 20, 23, 21, 19, 18, 21, 19, 23, 23, 11, 0, 0, 15, 30, 24, 22, 
    
    -- channel=55
    96, 94, 87, 82, 87, 86, 80, 83, 86, 90, 90, 96, 92, 94, 97, 94, 97, 96, 97, 98, 95, 95, 95, 98, 103, 102, 98, 96, 100, 87, 
    94, 92, 90, 84, 84, 57, 43, 49, 46, 56, 58, 57, 55, 57, 65, 59, 65, 66, 66, 67, 66, 60, 76, 83, 90, 91, 90, 93, 100, 87, 
    93, 90, 95, 91, 91, 48, 45, 48, 27, 29, 22, 21, 24, 27, 31, 20, 25, 29, 26, 28, 34, 21, 60, 71, 77, 91, 92, 94, 99, 85, 
    91, 90, 97, 91, 85, 49, 58, 55, 38, 54, 51, 41, 47, 45, 55, 50, 59, 66, 60, 63, 67, 60, 89, 88, 85, 94, 95, 95, 98, 83, 
    91, 90, 97, 92, 69, 27, 34, 28, 32, 49, 43, 27, 39, 32, 40, 38, 51, 50, 46, 52, 45, 55, 57, 59, 73, 85, 98, 95, 100, 82, 
    91, 90, 96, 88, 52, 21, 23, 22, 31, 33, 39, 25, 39, 28, 30, 26, 33, 29, 20, 34, 23, 51, 31, 46, 71, 75, 90, 92, 99, 80, 
    90, 89, 94, 85, 64, 55, 53, 57, 58, 53, 63, 55, 62, 58, 58, 55, 59, 58, 50, 61, 55, 73, 53, 70, 89, 86, 94, 95, 98, 81, 
    87, 88, 91, 85, 78, 72, 57, 65, 62, 61, 63, 62, 71, 69, 66, 61, 63, 62, 56, 62, 62, 77, 75, 82, 87, 89, 95, 96, 98, 81, 
    86, 91, 92, 88, 90, 83, 66, 74, 74, 74, 77, 74, 82, 80, 76, 73, 73, 74, 74, 81, 78, 91, 97, 86, 86, 91, 94, 92, 97, 82, 
    90, 97, 97, 89, 94, 90, 84, 94, 93, 94, 94, 94, 96, 92, 90, 87, 89, 93, 94, 97, 95, 99, 100, 89, 89, 92, 93, 91, 98, 83, 
    92, 91, 84, 64, 74, 85, 84, 94, 93, 93, 93, 91, 90, 89, 87, 86, 87, 89, 90, 95, 94, 93, 92, 89, 93, 96, 97, 97, 102, 84, 
    96, 83, 74, 56, 56, 62, 56, 66, 79, 86, 89, 88, 87, 87, 88, 88, 89, 91, 92, 93, 94, 92, 93, 96, 96, 96, 96, 95, 97, 80, 
    101, 93, 96, 90, 84, 72, 58, 55, 60, 69, 78, 86, 90, 91, 90, 90, 91, 90, 89, 89, 89, 88, 89, 90, 91, 91, 90, 90, 94, 79, 
    101, 98, 98, 93, 94, 92, 77, 69, 63, 63, 71, 81, 88, 89, 90, 89, 90, 89, 88, 90, 91, 91, 92, 93, 93, 93, 92, 92, 95, 80, 
    103, 101, 100, 97, 100, 102, 83, 63, 63, 55, 51, 59, 69, 78, 87, 90, 91, 90, 90, 92, 93, 92, 92, 93, 92, 92, 93, 92, 96, 80, 
    103, 103, 103, 99, 102, 101, 89, 58, 56, 59, 46, 50, 54, 58, 64, 72, 82, 86, 88, 90, 92, 91, 92, 92, 91, 91, 93, 92, 95, 80, 
    101, 103, 103, 99, 101, 101, 96, 54, 47, 60, 47, 54, 55, 53, 51, 49, 50, 56, 60, 72, 84, 86, 89, 90, 90, 90, 92, 91, 95, 78, 
    101, 103, 104, 100, 102, 103, 98, 44, 31, 49, 37, 48, 51, 53, 52, 52, 49, 42, 31, 34, 45, 51, 63, 77, 86, 92, 95, 93, 95, 78, 
    102, 102, 102, 100, 102, 101, 75, 34, 27, 41, 41, 46, 47, 49, 49, 51, 55, 53, 46, 43, 47, 39, 38, 48, 54, 63, 74, 81, 87, 75, 
    101, 100, 99, 98, 100, 94, 63, 54, 70, 63, 52, 52, 36, 53, 72, 80, 81, 62, 67, 65, 65, 58, 55, 81, 88, 89, 89, 84, 85, 70, 
    101, 98, 95, 97, 98, 95, 83, 99, 111, 92, 79, 91, 88, 104, 117, 108, 98, 82, 104, 107, 98, 92, 101, 122, 114, 102, 99, 95, 93, 77, 
    96, 89, 85, 87, 88, 85, 81, 85, 83, 71, 72, 89, 87, 94, 92, 78, 74, 73, 92, 88, 83, 83, 88, 95, 82, 75, 74, 72, 77, 68, 
    59, 44, 41, 41, 43, 43, 41, 39, 40, 35, 37, 42, 38, 43, 46, 43, 48, 48, 52, 48, 49, 51, 54, 53, 50, 51, 51, 50, 55, 49, 
    73, 61, 58, 60, 63, 65, 64, 65, 68, 65, 66, 65, 64, 61, 58, 49, 45, 46, 44, 44, 43, 42, 41, 39, 39, 37, 30, 27, 30, 30, 
    65, 50, 47, 45, 45, 43, 43, 43, 43, 42, 42, 39, 37, 33, 32, 27, 24, 25, 24, 22, 21, 21, 21, 19, 19, 17, 12, 10, 20, 35, 
    46, 30, 25, 24, 24, 25, 31, 33, 34, 34, 35, 33, 34, 33, 34, 35, 36, 39, 38, 38, 39, 41, 41, 42, 41, 40, 38, 44, 67, 84, 
    59, 45, 43, 44, 41, 44, 50, 50, 53, 53, 53, 49, 49, 49, 52, 53, 53, 54, 54, 55, 55, 54, 52, 52, 52, 54, 65, 86, 104, 101, 
    59, 44, 46, 48, 45, 49, 52, 50, 51, 51, 53, 50, 51, 54, 58, 58, 56, 56, 58, 58, 59, 57, 55, 53, 57, 73, 95, 104, 94, 79, 
    60, 46, 49, 52, 50, 53, 54, 52, 55, 60, 59, 57, 56, 60, 64, 63, 65, 64, 64, 59, 59, 57, 58, 67, 84, 102, 100, 85, 72, 71, 
    58, 45, 49, 49, 46, 46, 48, 48, 51, 57, 53, 50, 50, 54, 57, 55, 56, 55, 54, 49, 53, 56, 68, 90, 104, 97, 78, 63, 66, 69, 
    
    -- channel=56
    71, 24, 17, 6, 12, 48, 71, 71, 64, 60, 60, 69, 71, 69, 74, 71, 71, 73, 74, 76, 75, 73, 76, 76, 81, 85, 84, 82, 82, 102, 
    45, 0, 0, 0, 0, 57, 98, 121, 119, 93, 82, 85, 88, 84, 88, 89, 85, 84, 85, 83, 82, 88, 76, 62, 54, 54, 64, 67, 70, 93, 
    45, 1, 7, 1, 11, 56, 91, 165, 171, 153, 160, 154, 163, 164, 169, 166, 163, 163, 162, 152, 153, 158, 139, 119, 75, 57, 70, 74, 74, 97, 
    38, 0, 6, 0, 19, 62, 75, 151, 149, 142, 163, 155, 160, 160, 153, 152, 143, 143, 146, 130, 139, 144, 135, 138, 84, 54, 68, 68, 66, 89, 
    44, 3, 8, 0, 30, 91, 104, 163, 123, 122, 144, 136, 152, 166, 157, 145, 122, 129, 128, 119, 131, 125, 124, 129, 97, 66, 62, 64, 67, 88, 
    40, 1, 6, 7, 44, 101, 161, 206, 146, 135, 141, 141, 149, 172, 168, 159, 145, 152, 151, 159, 159, 140, 148, 140, 137, 107, 69, 61, 62, 81, 
    33, 0, 4, 0, 21, 68, 121, 161, 120, 102, 106, 114, 107, 120, 117, 115, 110, 122, 119, 135, 141, 129, 125, 106, 125, 105, 63, 52, 52, 73, 
    29, 0, 6, 0, 13, 44, 65, 80, 77, 68, 68, 79, 74, 79, 77, 76, 73, 79, 78, 93, 104, 92, 86, 64, 71, 71, 50, 42, 43, 64, 
    31, 0, 8, 1, 8, 18, 21, 28, 45, 47, 45, 46, 46, 48, 50, 50, 47, 44, 49, 60, 68, 68, 67, 50, 43, 46, 43, 38, 37, 60, 
    41, 0, 15, 1, 3, 5, 0, 0, 10, 9, 11, 10, 10, 14, 13, 14, 15, 16, 15, 25, 29, 32, 43, 41, 37, 40, 45, 43, 41, 62, 
    61, 13, 28, 20, 29, 35, 22, 5, 8, 9, 10, 13, 16, 19, 18, 15, 13, 17, 19, 24, 28, 29, 33, 37, 38, 41, 47, 46, 45, 67, 
    75, 21, 31, 30, 61, 89, 80, 52, 34, 24, 21, 23, 25, 27, 26, 26, 26, 28, 30, 33, 35, 36, 36, 38, 41, 43, 46, 46, 46, 70, 
    82, 13, 6, 7, 35, 86, 123, 124, 95, 61, 41, 35, 36, 36, 35, 36, 38, 39, 38, 39, 44, 42, 40, 40, 43, 44, 48, 48, 47, 71, 
    87, 22, 11, 0, 2, 15, 57, 102, 121, 112, 83, 62, 52, 47, 45, 48, 52, 54, 52, 52, 55, 52, 48, 43, 43, 43, 44, 41, 39, 59, 
    92, 38, 47, 43, 50, 32, 14, 31, 65, 106, 126, 118, 98, 78, 64, 57, 54, 53, 51, 51, 53, 51, 46, 42, 39, 36, 36, 34, 30, 49, 
    96, 47, 60, 53, 67, 76, 52, 19, 23, 73, 118, 146, 156, 139, 111, 87, 71, 62, 56, 51, 48, 46, 42, 41, 40, 38, 39, 35, 29, 46, 
    107, 63, 81, 71, 75, 84, 80, 42, 7, 54, 102, 118, 142, 162, 165, 151, 130, 104, 82, 62, 53, 46, 41, 42, 43, 41, 44, 41, 34, 49, 
    117, 76, 97, 85, 84, 84, 86, 64, 16, 54, 102, 107, 112, 118, 134, 154, 165, 163, 140, 113, 100, 89, 77, 71, 63, 52, 50, 44, 37, 51, 
    121, 76, 94, 84, 82, 81, 91, 63, 29, 62, 96, 105, 110, 108, 108, 110, 116, 124, 123, 124, 140, 153, 148, 138, 122, 97, 77, 60, 44, 50, 
    120, 72, 86, 83, 80, 80, 75, 49, 28, 33, 57, 75, 93, 97, 100, 94, 81, 72, 54, 61, 85, 114, 135, 148, 151, 131, 108, 88, 67, 63, 
    117, 65, 73, 79, 80, 75, 53, 31, 29, 5, 0, 8, 39, 59, 84, 72, 39, 18, 25, 41, 25, 26, 39, 73, 89, 70, 64, 72, 69, 67, 
    113, 64, 71, 81, 83, 80, 68, 51, 53, 41, 0, 0, 0, 14, 52, 66, 40, 0, 0, 22, 18, 0, 0, 11, 40, 41, 29, 32, 37, 47, 
    132, 87, 90, 102, 105, 107, 109, 108, 109, 103, 79, 59, 56, 53, 59, 59, 48, 31, 16, 20, 27, 23, 9, 3, 6, 9, 8, 12, 17, 33, 
    119, 76, 71, 75, 71, 72, 73, 73, 76, 75, 71, 67, 62, 59, 51, 35, 22, 19, 23, 21, 20, 21, 21, 14, 3, 0, 0, 4, 16, 42, 
    76, 40, 32, 32, 30, 36, 43, 50, 57, 55, 48, 40, 35, 34, 39, 42, 37, 40, 44, 43, 43, 45, 48, 49, 48, 47, 45, 48, 51, 74, 
    113, 86, 81, 78, 71, 73, 85, 96, 103, 104, 103, 97, 96, 95, 95, 98, 97, 99, 104, 104, 101, 98, 97, 98, 98, 99, 99, 92, 85, 111, 
    119, 102, 102, 105, 102, 100, 111, 121, 122, 116, 109, 101, 100, 105, 108, 113, 112, 108, 108, 110, 110, 110, 108, 106, 104, 102, 99, 97, 101, 118, 
    113, 99, 97, 101, 98, 100, 110, 115, 116, 112, 105, 101, 105, 113, 119, 123, 119, 114, 111, 112, 113, 115, 115, 112, 103, 88, 86, 100, 101, 113, 
    115, 101, 96, 100, 96, 98, 106, 109, 107, 102, 100, 94, 95, 104, 112, 114, 108, 105, 105, 107, 108, 113, 115, 108, 98, 95, 99, 94, 100, 132, 
    119, 109, 104, 103, 98, 98, 105, 110, 115, 115, 111, 105, 107, 115, 123, 123, 116, 111, 110, 108, 111, 120, 120, 116, 117, 109, 99, 100, 111, 134, 
    
    -- channel=57
    1, 5, 14, 12, 3, 0, 0, 0, 0, 2, 3, 1, 0, 0, 1, 3, 0, 0, 0, 1, 0, 0, 0, 1, 4, 3, 0, 0, 0, 3, 
    0, 5, 14, 19, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 3, 
    0, 6, 9, 12, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    1, 7, 7, 8, 4, 10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 
    1, 8, 7, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 8, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 7, 10, 3, 9, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 3, 
    0, 5, 7, 10, 28, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 8, 0, 0, 0, 3, 0, 4, 
    3, 3, 7, 9, 12, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 8, 0, 0, 1, 3, 0, 6, 
    7, 5, 10, 5, 4, 12, 18, 9, 14, 11, 14, 14, 12, 14, 10, 7, 8, 13, 12, 10, 12, 4, 0, 4, 0, 0, 0, 1, 0, 7, 
    6, 0, 0, 0, 0, 7, 23, 13, 14, 15, 12, 13, 11, 11, 11, 10, 10, 9, 12, 10, 12, 5, 0, 3, 2, 3, 2, 2, 0, 7, 
    4, 0, 0, 0, 0, 0, 0, 0, 5, 6, 3, 2, 1, 3, 2, 3, 3, 2, 3, 3, 3, 3, 2, 2, 3, 4, 2, 2, 0, 4, 
    4, 12, 16, 19, 0, 0, 0, 0, 0, 0, 3, 2, 2, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    5, 17, 24, 33, 40, 15, 0, 0, 0, 0, 0, 3, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    3, 1, 5, 11, 29, 42, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 0, 7, 
    3, 2, 3, 1, 2, 14, 33, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 2, 1, 7, 
    0, 0, 0, 0, 0, 0, 14, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 0, 1, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 5, 19, 1, 0, 0, 0, 0, 13, 23, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 23, 33, 43, 47, 19, 12, 22, 19, 33, 40, 32, 25, 23, 39, 33, 27, 19, 13, 19, 11, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 14, 7, 4, 29, 39, 28, 40, 18, 2, 8, 18, 39, 16, 21, 33, 39, 35, 6, 2, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 20, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 20, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 11, 0, 0, 0, 0, 0, 
    
    -- channel=58
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=59
    301, 334, 342, 320, 302, 292, 288, 288, 298, 312, 319, 320, 315, 311, 309, 308, 312, 313, 316, 320, 322, 320, 318, 320, 330, 350, 361, 366, 371, 345, 
    308, 340, 351, 331, 308, 292, 265, 241, 263, 288, 290, 299, 286, 279, 286, 290, 294, 293, 296, 303, 303, 298, 297, 305, 339, 364, 366, 371, 380, 354, 
    308, 338, 354, 354, 337, 287, 240, 225, 250, 258, 250, 258, 251, 246, 259, 258, 263, 268, 268, 273, 273, 262, 282, 307, 347, 373, 368, 373, 380, 353, 
    302, 334, 352, 356, 345, 269, 224, 218, 222, 222, 216, 222, 213, 208, 226, 228, 241, 248, 250, 251, 254, 237, 288, 331, 354, 370, 371, 375, 380, 353, 
    300, 330, 349, 352, 338, 270, 232, 212, 207, 214, 216, 209, 202, 196, 217, 227, 236, 246, 247, 241, 249, 239, 279, 317, 331, 355, 375, 378, 383, 355, 
    298, 327, 343, 345, 312, 233, 218, 210, 220, 237, 237, 216, 220, 213, 236, 244, 255, 260, 254, 252, 249, 260, 273, 289, 308, 340, 371, 377, 384, 354, 
    298, 325, 339, 337, 283, 210, 216, 221, 232, 234, 239, 224, 228, 224, 235, 235, 248, 248, 237, 241, 235, 265, 245, 257, 308, 342, 365, 371, 377, 350, 
    303, 324, 337, 331, 292, 268, 261, 253, 256, 248, 263, 259, 259, 257, 258, 256, 261, 264, 245, 247, 253, 280, 261, 280, 323, 346, 363, 368, 372, 346, 
    310, 328, 337, 336, 332, 329, 304, 287, 282, 283, 285, 280, 284, 287, 294, 300, 299, 294, 285, 286, 291, 307, 319, 339, 351, 358, 364, 367, 370, 343, 
    323, 336, 342, 346, 346, 334, 307, 298, 291, 289, 287, 286, 291, 296, 301, 303, 302, 299, 295, 297, 297, 312, 344, 358, 362, 363, 363, 363, 369, 342, 
    335, 351, 349, 334, 320, 312, 314, 323, 322, 317, 317, 319, 326, 330, 331, 327, 323, 323, 322, 325, 327, 335, 349, 355, 360, 362, 362, 365, 373, 345, 
    347, 355, 333, 292, 281, 289, 295, 309, 327, 344, 353, 353, 356, 360, 362, 360, 357, 357, 356, 355, 356, 358, 360, 363, 364, 366, 366, 368, 374, 347, 
    354, 338, 300, 257, 240, 249, 256, 270, 288, 310, 333, 351, 361, 367, 369, 367, 366, 364, 359, 357, 359, 360, 360, 362, 363, 366, 366, 368, 373, 346, 
    361, 354, 324, 286, 236, 198, 195, 210, 234, 266, 298, 329, 357, 371, 373, 372, 372, 368, 362, 358, 360, 362, 362, 361, 362, 363, 360, 361, 366, 339, 
    369, 385, 379, 367, 334, 269, 207, 173, 161, 188, 245, 290, 321, 346, 364, 370, 370, 366, 359, 356, 357, 359, 357, 357, 359, 358, 356, 359, 364, 336, 
    373, 389, 386, 385, 384, 365, 297, 210, 142, 118, 158, 217, 267, 298, 318, 334, 347, 355, 358, 357, 357, 360, 361, 362, 363, 362, 360, 361, 364, 336, 
    375, 393, 393, 391, 390, 390, 358, 261, 153, 86, 84, 115, 162, 217, 258, 281, 296, 307, 319, 327, 338, 353, 361, 363, 362, 361, 360, 360, 364, 337, 
    374, 394, 395, 392, 392, 387, 382, 298, 159, 75, 53, 58, 73, 102, 141, 184, 221, 246, 253, 258, 278, 304, 326, 339, 348, 355, 359, 360, 364, 336, 
    372, 390, 391, 388, 391, 389, 388, 278, 125, 60, 33, 39, 54, 61, 68, 82, 101, 127, 139, 160, 198, 238, 267, 281, 298, 314, 327, 340, 355, 332, 
    369, 385, 387, 387, 389, 391, 355, 228, 104, 58, 45, 35, 38, 46, 60, 91, 107, 94, 48, 42, 94, 136, 159, 186, 239, 294, 320, 332, 347, 329, 
    367, 379, 380, 384, 386, 379, 311, 237, 188, 139, 95, 70, 66, 94, 145, 185, 187, 147, 114, 106, 110, 107, 105, 150, 215, 262, 297, 326, 346, 330, 
    357, 370, 372, 373, 374, 365, 326, 301, 296, 259, 187, 154, 143, 178, 249, 291, 277, 213, 205, 223, 218, 190, 178, 226, 276, 295, 302, 310, 326, 314, 
    309, 317, 317, 314, 312, 308, 305, 302, 301, 289, 253, 234, 226, 236, 268, 291, 293, 270, 264, 267, 274, 269, 264, 272, 282, 289, 292, 293, 299, 282, 
    237, 239, 235, 230, 224, 221, 218, 212, 213, 210, 204, 201, 201, 210, 218, 219, 218, 218, 218, 219, 221, 224, 229, 227, 221, 216, 216, 215, 222, 209, 
    148, 145, 144, 138, 135, 132, 124, 120, 121, 113, 107, 105, 106, 116, 132, 138, 135, 130, 128, 128, 127, 129, 134, 136, 139, 140, 131, 124, 127, 119, 
    123, 122, 123, 117, 114, 111, 107, 107, 104, 99, 96, 92, 93, 92, 97, 96, 90, 88, 84, 80, 75, 75, 77, 80, 82, 81, 72, 65, 70, 96, 
    80, 78, 79, 76, 71, 62, 61, 62, 58, 52, 47, 44, 44, 44, 46, 48, 45, 38, 31, 28, 28, 29, 28, 27, 26, 27, 26, 36, 87, 133, 
    34, 29, 31, 30, 28, 25, 30, 30, 26, 21, 17, 19, 24, 26, 29, 36, 34, 27, 21, 21, 24, 26, 23, 20, 21, 25, 49, 106, 156, 137, 
    32, 25, 28, 29, 25, 27, 31, 29, 24, 20, 27, 32, 31, 31, 36, 41, 38, 35, 34, 34, 30, 26, 26, 27, 35, 74, 133, 160, 133, 89, 
    29, 20, 22, 21, 20, 23, 24, 21, 22, 28, 37, 41, 39, 41, 47, 47, 45, 42, 42, 37, 30, 28, 31, 47, 94, 149, 154, 112, 69, 47, 
    
    -- channel=60
    73, 83, 89, 87, 79, 70, 68, 70, 76, 76, 78, 79, 78, 77, 74, 76, 77, 78, 79, 79, 80, 80, 79, 79, 80, 82, 82, 83, 86, 71, 
    77, 85, 90, 85, 71, 56, 43, 42, 57, 65, 63, 64, 59, 57, 60, 62, 60, 62, 62, 63, 65, 61, 62, 75, 79, 83, 83, 86, 90, 74, 
    77, 87, 92, 93, 78, 48, 37, 37, 40, 40, 38, 43, 42, 38, 42, 45, 43, 47, 47, 47, 47, 46, 51, 72, 85, 88, 85, 86, 90, 74, 
    74, 86, 90, 93, 79, 47, 42, 43, 41, 43, 40, 38, 35, 35, 40, 45, 45, 49, 52, 49, 49, 48, 61, 82, 88, 89, 88, 88, 92, 75, 
    72, 85, 90, 91, 75, 37, 38, 42, 37, 40, 40, 35, 31, 33, 41, 48, 47, 53, 51, 47, 53, 48, 57, 70, 80, 87, 86, 84, 89, 75, 
    73, 85, 88, 87, 62, 21, 36, 40, 41, 45, 45, 39, 32, 34, 43, 48, 49, 47, 45, 43, 48, 49, 54, 55, 68, 84, 89, 92, 92, 75, 
    74, 86, 87, 85, 56, 22, 39, 45, 45, 46, 47, 42, 38, 41, 45, 48, 51, 47, 42, 43, 46, 50, 48, 56, 76, 85, 84, 88, 91, 76, 
    77, 86, 87, 84, 67, 56, 62, 61, 60, 54, 58, 58, 56, 54, 53, 58, 62, 58, 50, 51, 54, 61, 55, 61, 81, 91, 88, 91, 93, 76, 
    79, 87, 87, 87, 83, 81, 78, 73, 72, 72, 70, 73, 73, 72, 74, 77, 76, 72, 70, 67, 71, 78, 75, 79, 88, 92, 88, 89, 93, 75, 
    80, 87, 87, 90, 86, 82, 80, 79, 75, 74, 74, 74, 74, 75, 76, 80, 82, 79, 76, 72, 73, 79, 85, 86, 88, 88, 85, 87, 91, 75, 
    80, 90, 81, 78, 69, 69, 79, 83, 81, 78, 77, 78, 79, 81, 81, 81, 79, 79, 78, 76, 77, 79, 84, 87, 89, 88, 88, 90, 92, 76, 
    82, 92, 80, 70, 61, 49, 49, 62, 77, 87, 88, 87, 88, 90, 92, 91, 91, 91, 90, 88, 87, 89, 90, 90, 88, 87, 87, 86, 88, 73, 
    83, 90, 82, 74, 66, 60, 51, 47, 52, 63, 78, 87, 90, 92, 92, 90, 89, 88, 87, 85, 85, 86, 86, 86, 87, 88, 87, 88, 91, 75, 
    84, 88, 74, 62, 49, 45, 51, 48, 47, 50, 59, 73, 85, 90, 90, 89, 88, 87, 86, 86, 86, 89, 90, 90, 90, 90, 88, 90, 92, 76, 
    86, 94, 90, 89, 74, 52, 44, 41, 29, 31, 42, 48, 59, 75, 86, 90, 91, 88, 86, 84, 84, 85, 86, 86, 87, 88, 87, 89, 92, 76, 
    84, 92, 89, 92, 88, 79, 62, 51, 30, 11, 21, 35, 42, 45, 54, 68, 78, 86, 89, 88, 87, 89, 89, 89, 89, 89, 88, 89, 92, 77, 
    82, 90, 88, 90, 88, 87, 79, 63, 33, 0, 0, 8, 23, 36, 41, 41, 43, 52, 64, 72, 80, 88, 91, 91, 90, 89, 87, 88, 91, 76, 
    80, 89, 87, 90, 90, 87, 86, 70, 30, 0, 0, 0, 0, 4, 19, 31, 37, 38, 37, 37, 40, 51, 64, 73, 81, 87, 87, 89, 92, 77, 
    80, 88, 85, 89, 90, 87, 88, 59, 25, 3, 0, 0, 0, 0, 0, 0, 9, 21, 29, 33, 34, 35, 36, 35, 44, 55, 64, 77, 88, 76, 
    81, 88, 87, 91, 90, 90, 84, 53, 24, 19, 8, 0, 0, 0, 0, 15, 22, 13, 0, 1, 19, 24, 27, 31, 53, 71, 73, 74, 81, 74, 
    83, 87, 88, 91, 89, 87, 76, 62, 45, 34, 30, 23, 21, 24, 26, 33, 39, 37, 27, 18, 21, 27, 29, 33, 42, 55, 70, 78, 83, 78, 
    78, 82, 83, 83, 81, 78, 66, 56, 51, 45, 33, 26, 20, 28, 43, 54, 53, 41, 41, 42, 39, 33, 33, 44, 55, 61, 64, 66, 75, 72, 
    51, 55, 56, 56, 54, 52, 52, 51, 51, 50, 40, 32, 29, 35, 50, 67, 72, 64, 58, 60, 64, 62, 61, 64, 73, 79, 81, 77, 78, 68, 
    59, 61, 65, 65, 63, 62, 61, 60, 60, 60, 59, 60, 60, 62, 61, 63, 63, 62, 63, 63, 63, 63, 65, 65, 63, 62, 62, 58, 60, 48, 
    22, 23, 28, 27, 24, 20, 15, 12, 10, 9, 8, 7, 7, 12, 17, 19, 19, 16, 14, 14, 15, 15, 16, 16, 17, 18, 15, 14, 18, 7, 
    5, 4, 8, 8, 9, 7, 3, 2, 0, 0, 0, 1, 3, 3, 4, 4, 4, 2, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 4, 
    2, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 7, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 4, 0, 0, 0, 
    
    -- channel=61
    331, 396, 419, 413, 387, 354, 337, 341, 354, 377, 390, 390, 380, 375, 372, 377, 382, 380, 381, 386, 387, 386, 380, 384, 399, 421, 441, 446, 448, 413, 
    341, 402, 423, 428, 424, 375, 327, 307, 320, 359, 373, 374, 365, 361, 368, 373, 385, 385, 387, 394, 390, 381, 393, 408, 439, 455, 457, 456, 458, 419, 
    338, 391, 410, 426, 428, 390, 342, 291, 290, 301, 294, 296, 290, 291, 298, 308, 311, 310, 313, 320, 316, 306, 332, 370, 430, 450, 449, 450, 458, 422, 
    336, 387, 403, 419, 422, 390, 370, 338, 335, 326, 314, 316, 314, 312, 330, 346, 353, 357, 355, 362, 352, 350, 372, 394, 440, 456, 457, 459, 466, 431, 
    328, 382, 396, 413, 404, 353, 337, 306, 333, 334, 328, 327, 315, 308, 326, 347, 368, 371, 372, 373, 359, 369, 374, 388, 409, 433, 455, 457, 464, 431, 
    330, 379, 393, 406, 388, 336, 291, 269, 301, 311, 313, 305, 303, 297, 308, 312, 317, 324, 317, 311, 308, 332, 322, 333, 344, 391, 438, 446, 452, 422, 
    339, 383, 392, 409, 397, 367, 350, 332, 336, 344, 344, 338, 343, 345, 356, 355, 360, 359, 349, 345, 337, 358, 363, 373, 371, 400, 433, 440, 445, 415, 
    355, 389, 390, 406, 401, 396, 384, 361, 337, 340, 340, 331, 330, 333, 350, 360, 368, 360, 349, 345, 336, 358, 380, 415, 433, 430, 438, 443, 447, 412, 
    373, 404, 394, 406, 408, 406, 381, 354, 328, 323, 323, 320, 327, 336, 346, 349, 348, 343, 333, 335, 331, 345, 378, 418, 446, 439, 438, 439, 446, 410, 
    390, 425, 410, 415, 413, 410, 405, 397, 381, 381, 379, 383, 395, 403, 411, 410, 402, 393, 389, 388, 390, 399, 414, 427, 439, 437, 434, 434, 442, 411, 
    396, 420, 388, 358, 339, 358, 397, 431, 427, 422, 424, 428, 436, 442, 445, 443, 438, 429, 423, 421, 424, 430, 435, 434, 438, 440, 442, 445, 452, 420, 
    400, 412, 354, 287, 222, 211, 258, 337, 395, 427, 438, 440, 445, 451, 456, 456, 453, 448, 442, 438, 441, 444, 445, 442, 441, 442, 445, 447, 453, 419, 
    410, 441, 410, 363, 289, 202, 142, 156, 235, 328, 397, 434, 450, 458, 462, 462, 460, 455, 448, 441, 437, 438, 438, 437, 435, 435, 435, 436, 441, 408, 
    415, 456, 446, 441, 407, 346, 241, 150, 125, 180, 284, 379, 438, 463, 465, 458, 454, 448, 442, 436, 434, 435, 435, 436, 435, 435, 433, 432, 436, 404, 
    420, 470, 461, 461, 444, 430, 376, 253, 142, 95, 135, 222, 319, 398, 442, 455, 452, 444, 438, 435, 434, 436, 437, 439, 439, 440, 438, 437, 441, 408, 
    425, 476, 470, 478, 469, 454, 430, 331, 194, 84, 58, 86, 131, 210, 298, 369, 415, 435, 437, 434, 436, 437, 440, 440, 439, 438, 437, 437, 442, 411, 
    424, 473, 466, 476, 471, 464, 450, 359, 231, 96, 30, 45, 52, 70, 108, 163, 227, 292, 338, 377, 409, 436, 452, 449, 442, 436, 433, 432, 438, 410, 
    423, 470, 461, 470, 469, 467, 457, 351, 203, 56, 0, 1, 17, 40, 52, 56, 65, 81, 103, 143, 208, 288, 357, 397, 422, 436, 440, 441, 444, 414, 
    420, 468, 458, 466, 467, 468, 424, 310, 151, 8, 0, 0, 0, 16, 34, 43, 42, 30, 10, 0, 18, 61, 119, 177, 237, 304, 361, 403, 433, 417, 
    413, 463, 456, 460, 463, 458, 398, 297, 197, 114, 30, 0, 0, 4, 71, 135, 153, 99, 64, 44, 48, 34, 22, 69, 153, 246, 310, 354, 397, 395, 
    408, 460, 459, 461, 461, 460, 431, 393, 363, 335, 271, 190, 136, 162, 225, 306, 347, 292, 235, 213, 243, 229, 196, 208, 269, 346, 384, 393, 404, 390, 
    390, 437, 436, 430, 424, 417, 404, 404, 406, 386, 361, 333, 306, 323, 344, 361, 370, 355, 347, 332, 337, 343, 341, 345, 347, 353, 369, 377, 383, 365, 
    233, 262, 262, 246, 235, 225, 217, 211, 209, 197, 188, 187, 189, 213, 242, 255, 258, 252, 263, 267, 265, 268, 281, 294, 294, 289, 289, 289, 294, 280, 
    156, 175, 180, 171, 167, 161, 156, 151, 146, 141, 138, 134, 138, 149, 171, 189, 195, 192, 187, 189, 188, 190, 194, 201, 209, 214, 211, 202, 190, 173, 
    140, 152, 162, 158, 150, 137, 126, 116, 109, 102, 96, 95, 97, 101, 106, 105, 100, 88, 78, 76, 73, 70, 68, 71, 74, 76, 74, 64, 55, 54, 
    45, 46, 57, 57, 53, 43, 32, 24, 17, 7, 2, 1, 2, 4, 7, 7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 54, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 47, 62, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 60, 62, 21, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 22, 51, 47, 1, 0, 0, 
    
    -- channel=62
    110, 104, 90, 53, 48, 63, 73, 89, 99, 88, 72, 71, 67, 68, 75, 67, 67, 72, 75, 77, 73, 72, 74, 75, 81, 86, 79, 77, 84, 42, 
    117, 116, 109, 67, 39, 37, 62, 100, 111, 103, 86, 80, 73, 75, 86, 77, 69, 72, 71, 75, 73, 66, 80, 85, 83, 92, 93, 89, 94, 50, 
    113, 113, 114, 94, 70, 31, 47, 104, 114, 121, 133, 123, 114, 118, 130, 126, 120, 126, 123, 123, 122, 108, 132, 141, 106, 92, 94, 90, 94, 51, 
    114, 109, 113, 103, 88, 21, 18, 58, 47, 67, 85, 68, 62, 76, 88, 74, 70, 76, 70, 73, 79, 51, 96, 132, 104, 89, 90, 93, 97, 52, 
    112, 106, 109, 101, 86, 39, 77, 85, 35, 41, 48, 30, 36, 59, 69, 52, 42, 45, 34, 40, 51, 30, 70, 112, 117, 103, 88, 89, 96, 54, 
    110, 107, 107, 93, 72, 44, 105, 122, 86, 90, 91, 68, 73, 88, 107, 107, 111, 112, 98, 109, 110, 109, 110, 121, 154, 135, 102, 98, 106, 61, 
    102, 106, 107, 90, 50, 14, 41, 57, 67, 67, 69, 48, 45, 52, 65, 66, 77, 74, 59, 75, 71, 86, 57, 57, 121, 121, 97, 96, 107, 63, 
    93, 100, 110, 90, 53, 34, 28, 38, 60, 56, 67, 56, 54, 56, 61, 56, 50, 48, 37, 49, 53, 75, 46, 35, 75, 92, 91, 90, 99, 59, 
    82, 90, 105, 90, 81, 79, 62, 71, 85, 84, 92, 87, 87, 89, 94, 96, 91, 87, 78, 83, 87, 99, 107, 94, 82, 87, 93, 95, 99, 56, 
    77, 78, 93, 86, 95, 89, 55, 54, 59, 56, 60, 58, 60, 62, 64, 67, 66, 62, 55, 57, 57, 70, 105, 108, 93, 91, 95, 97, 100, 56, 
    85, 82, 96, 93, 113, 120, 80, 56, 55, 52, 56, 61, 66, 67, 63, 58, 56, 59, 57, 60, 62, 70, 89, 96, 93, 89, 87, 87, 95, 53, 
    91, 81, 91, 87, 120, 174, 172, 136, 109, 92, 89, 94, 98, 97, 94, 89, 87, 85, 84, 87, 90, 90, 87, 88, 90, 89, 87, 87, 97, 57, 
    92, 57, 33, 4, 14, 93, 173, 203, 186, 148, 115, 101, 98, 97, 93, 89, 86, 84, 83, 89, 95, 94, 91, 92, 95, 98, 99, 101, 106, 62, 
    98, 62, 33, 0, 0, 0, 0, 102, 184, 203, 171, 130, 104, 94, 93, 92, 93, 91, 88, 90, 97, 97, 96, 95, 95, 94, 95, 98, 104, 59, 
    103, 90, 91, 70, 25, 0, 0, 0, 53, 159, 200, 195, 164, 126, 102, 94, 94, 92, 87, 86, 89, 88, 87, 89, 89, 87, 86, 89, 98, 58, 
    104, 89, 91, 83, 81, 58, 0, 0, 0, 66, 140, 186, 212, 196, 160, 126, 104, 94, 89, 90, 94, 92, 91, 94, 94, 91, 90, 91, 98, 59, 
    106, 91, 96, 86, 85, 87, 55, 0, 0, 1, 54, 80, 138, 184, 202, 194, 175, 150, 127, 117, 114, 99, 89, 91, 92, 92, 93, 93, 100, 63, 
    104, 90, 99, 91, 89, 83, 77, 0, 0, 3, 47, 38, 50, 75, 114, 152, 180, 196, 192, 192, 194, 163, 127, 109, 98, 90, 87, 89, 98, 63, 
    105, 86, 95, 92, 90, 86, 80, 0, 0, 9, 56, 57, 50, 40, 34, 41, 62, 93, 121, 165, 216, 223, 200, 185, 166, 141, 122, 107, 102, 63, 
    112, 88, 94, 96, 94, 92, 60, 0, 0, 0, 0, 37, 55, 57, 43, 0, 0, 0, 0, 14, 59, 106, 140, 174, 177, 151, 142, 133, 120, 77, 
    116, 92, 92, 93, 94, 87, 18, 0, 0, 0, 0, 0, 0, 5, 30, 0, 0, 0, 0, 0, 0, 0, 0, 30, 66, 53, 68, 94, 105, 75, 
    121, 100, 100, 99, 102, 95, 52, 25, 33, 0, 0, 0, 0, 0, 55, 72, 29, 0, 0, 13, 0, 0, 0, 14, 73, 79, 82, 91, 100, 76, 
    167, 156, 154, 154, 155, 158, 161, 163, 170, 155, 112, 102, 108, 122, 149, 155, 146, 119, 110, 121, 128, 117, 105, 113, 128, 140, 147, 147, 143, 109, 
    148, 145, 139, 135, 131, 130, 127, 125, 129, 124, 121, 127, 132, 143, 145, 130, 124, 134, 137, 133, 136, 144, 149, 140, 130, 125, 127, 136, 147, 121, 
    58, 60, 54, 48, 44, 44, 40, 38, 41, 41, 41, 44, 52, 69, 89, 90, 83, 90, 98, 99, 99, 105, 114, 117, 119, 118, 111, 112, 123, 104, 
    82, 95, 93, 91, 88, 86, 85, 84, 79, 81, 84, 85, 88, 87, 93, 90, 77, 76, 83, 85, 82, 82, 83, 85, 88, 88, 78, 72, 73, 55, 
    60, 79, 76, 73, 65, 57, 57, 49, 40, 42, 46, 45, 44, 42, 41, 39, 28, 18, 19, 22, 24, 23, 21, 21, 23, 22, 15, 7, 11, 4, 
    9, 26, 23, 24, 19, 16, 21, 14, 8, 10, 15, 15, 12, 13, 14, 15, 12, 7, 6, 7, 8, 10, 10, 13, 14, 13, 3, 0, 16, 18, 
    10, 23, 20, 25, 18, 17, 20, 16, 11, 11, 13, 7, 3, 4, 8, 5, 0, 0, 0, 2, 5, 7, 7, 10, 9, 8, 13, 24, 31, 25, 
    4, 16, 14, 20, 16, 15, 15, 12, 10, 18, 18, 8, 3, 5, 13, 9, 3, 2, 2, 0, 3, 9, 7, 7, 12, 23, 32, 28, 20, 14, 
    
    -- channel=63
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=64
    41, 88, 68, 18, 23, 38, 34, 62, 113, 83, 11, 7, 47, 62, 20, 0, 21, 32, 15, 17, 61, 57, 0, 0, 108, 98, 29, 44, 36, 40, 
    33, 77, 44, 4, 31, 41, 31, 73, 114, 70, 16, 27, 61, 75, 16, 0, 35, 45, 11, 6, 61, 55, 0, 0, 109, 95, 7, 7, 25, 65, 
    24, 55, 29, 10, 42, 36, 29, 86, 116, 72, 40, 51, 60, 61, 11, 0, 28, 38, 10, 6, 63, 43, 0, 0, 80, 65, 0, 0, 31, 64, 
    23, 32, 38, 27, 45, 38, 36, 95, 117, 75, 48, 41, 34, 24, 6, 8, 30, 42, 40, 16, 48, 34, 0, 0, 44, 42, 0, 0, 18, 36, 
    52, 50, 36, 36, 37, 49, 54, 98, 110, 53, 15, 0, 0, 10, 36, 35, 18, 55, 81, 18, 12, 23, 0, 0, 22, 40, 0, 0, 11, 43, 
    78, 53, 18, 25, 26, 58, 72, 103, 86, 5, 0, 0, 0, 43, 82, 64, 3, 42, 101, 2, 0, 12, 0, 0, 13, 32, 0, 0, 37, 110, 
    75, 17, 0, 14, 40, 50, 67, 102, 48, 0, 0, 0, 27, 91, 100, 32, 0, 32, 59, 0, 0, 0, 0, 0, 0, 21, 0, 0, 85, 152, 
    63, 0, 0, 0, 59, 64, 47, 70, 5, 0, 0, 12, 71, 115, 48, 0, 0, 28, 1, 0, 0, 0, 0, 0, 0, 8, 0, 9, 120, 156, 
    61, 0, 0, 0, 42, 85, 65, 32, 0, 0, 0, 30, 98, 78, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 26, 140, 147, 
    72, 0, 0, 0, 12, 74, 81, 12, 0, 0, 0, 35, 59, 6, 0, 0, 0, 0, 0, 0, 7, 43, 0, 0, 0, 0, 0, 33, 142, 145, 
    90, 0, 0, 0, 0, 33, 54, 0, 0, 0, 0, 33, 36, 0, 0, 0, 0, 0, 0, 4, 22, 18, 0, 0, 13, 0, 0, 30, 137, 135, 
    86, 0, 0, 0, 0, 0, 4, 0, 0, 2, 0, 27, 31, 0, 0, 9, 10, 8, 5, 12, 16, 0, 0, 0, 15, 4, 0, 20, 123, 98, 
    59, 0, 0, 0, 0, 0, 0, 8, 20, 10, 12, 19, 8, 0, 8, 19, 20, 12, 9, 18, 3, 0, 0, 0, 10, 0, 0, 22, 105, 55, 
    55, 1, 0, 6, 0, 0, 0, 0, 30, 51, 21, 3, 2, 0, 0, 3, 12, 18, 12, 27, 1, 0, 0, 4, 24, 0, 0, 46, 105, 43, 
    50, 4, 0, 0, 0, 0, 0, 0, 0, 85, 51, 0, 0, 0, 0, 0, 2, 4, 0, 7, 8, 0, 0, 0, 25, 4, 0, 73, 121, 23, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 46, 58, 0, 0, 0, 0, 9, 1, 0, 0, 0, 0, 3, 0, 0, 16, 36, 7, 72, 117, 0, 
    0, 0, 0, 7, 13, 2, 3, 0, 0, 0, 17, 14, 0, 0, 0, 0, 0, 0, 0, 10, 2, 1, 0, 3, 45, 47, 42, 45, 73, 0, 
    0, 0, 4, 38, 38, 2, 0, 0, 14, 0, 0, 35, 9, 0, 0, 0, 0, 0, 0, 12, 3, 0, 6, 19, 59, 78, 56, 36, 20, 0, 
    0, 22, 34, 43, 46, 3, 0, 0, 8, 30, 0, 0, 2, 0, 0, 0, 0, 0, 4, 29, 2, 0, 14, 23, 62, 73, 36, 29, 0, 0, 
    40, 41, 20, 25, 47, 2, 0, 34, 0, 19, 29, 0, 0, 0, 0, 0, 0, 0, 6, 24, 6, 0, 19, 28, 52, 49, 23, 0, 0, 0, 
    71, 33, 0, 19, 47, 2, 0, 16, 3, 0, 16, 0, 0, 0, 0, 0, 0, 14, 18, 11, 8, 4, 12, 22, 33, 43, 10, 0, 0, 0, 
    41, 0, 0, 2, 32, 17, 0, 0, 7, 14, 0, 0, 0, 0, 0, 0, 0, 15, 21, 8, 0, 0, 5, 13, 25, 26, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 8, 0, 0, 15, 20, 0, 0, 0, 0, 0, 2, 0, 10, 22, 0, 0, 7, 10, 21, 33, 22, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 2, 18, 0, 0, 15, 0, 0, 23, 28, 23, 41, 52, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 10, 55, 48, 0, 0, 0, 0, 0, 23, 33, 22, 47, 93, 12, 0, 0, 12, 
    45, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 72, 60, 0, 0, 0, 0, 7, 15, 20, 35, 91, 94, 0, 0, 12, 30, 
    60, 87, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 22, 0, 0, 0, 2, 0, 20, 38, 65, 114, 68, 0, 0, 0, 0, 
    66, 92, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 30, 53, 89, 100, 28, 6, 0, 0, 0, 
    74, 64, 64, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 11, 0, 18, 20, 25, 48, 41, 52, 46, 0, 9, 0, 0, 0, 
    93, 43, 30, 66, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 19, 31, 48, 34, 17, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=65
    96, 104, 85, 62, 74, 108, 126, 127, 121, 88, 43, 68, 92, 96, 93, 87, 113, 134, 132, 136, 140, 131, 88, 96, 145, 122, 73, 102, 103, 92, 
    120, 119, 91, 69, 105, 132, 131, 129, 119, 73, 42, 82, 108, 107, 92, 91, 121, 131, 126, 130, 139, 126, 80, 100, 158, 123, 62, 85, 94, 105, 
    130, 125, 107, 91, 129, 137, 131, 130, 116, 61, 47, 83, 104, 100, 81, 91, 122, 116, 103, 116, 137, 123, 72, 105, 166, 126, 63, 92, 120, 135, 
    130, 120, 108, 115, 139, 132, 133, 129, 112, 56, 53, 77, 93, 95, 81, 102, 146, 143, 122, 125, 128, 120, 81, 106, 169, 145, 102, 138, 155, 147, 
    131, 140, 123, 121, 133, 125, 131, 125, 106, 52, 47, 69, 87, 98, 114, 127, 132, 127, 132, 119, 114, 119, 88, 113, 179, 181, 144, 154, 153, 146, 
    131, 131, 110, 121, 117, 115, 116, 111, 96, 46, 54, 91, 114, 129, 137, 125, 116, 115, 115, 89, 85, 128, 102, 124, 187, 195, 154, 151, 149, 166, 
    134, 111, 80, 109, 122, 126, 99, 91, 82, 47, 85, 132, 148, 154, 133, 92, 73, 123, 115, 57, 79, 141, 121, 140, 206, 197, 160, 160, 169, 174, 
    129, 102, 87, 134, 128, 130, 104, 78, 53, 52, 121, 155, 155, 145, 95, 46, 58, 112, 119, 81, 97, 144, 137, 145, 198, 201, 171, 175, 185, 161, 
    130, 102, 115, 178, 174, 130, 107, 100, 60, 75, 130, 138, 141, 122, 63, 58, 115, 133, 108, 118, 137, 162, 153, 145, 179, 191, 179, 185, 186, 144, 
    135, 100, 120, 186, 203, 166, 111, 100, 102, 125, 134, 122, 113, 70, 52, 101, 154, 150, 132, 142, 158, 168, 138, 135, 181, 191, 184, 190, 178, 117, 
    128, 95, 114, 183, 203, 196, 144, 88, 101, 130, 108, 91, 94, 73, 70, 110, 130, 127, 129, 122, 142, 146, 95, 110, 183, 196, 186, 182, 170, 108, 
    131, 91, 111, 174, 198, 205, 174, 97, 88, 93, 68, 59, 66, 86, 123, 133, 120, 106, 95, 85, 87, 93, 90, 133, 185, 186, 188, 187, 174, 109, 
    123, 80, 103, 149, 178, 191, 181, 136, 103, 75, 55, 62, 60, 46, 68, 97, 98, 88, 73, 72, 67, 63, 74, 114, 171, 169, 167, 182, 180, 107, 
    138, 105, 111, 142, 156, 176, 180, 148, 96, 84, 81, 57, 59, 61, 54, 52, 55, 60, 71, 82, 85, 81, 76, 88, 132, 160, 163, 188, 179, 110, 
    146, 122, 131, 153, 150, 163, 181, 149, 89, 60, 80, 67, 65, 74, 80, 70, 60, 54, 56, 66, 73, 95, 106, 102, 102, 132, 163, 182, 175, 113, 
    136, 115, 135, 151, 159, 157, 179, 148, 140, 116, 66, 48, 65, 63, 68, 88, 97, 82, 60, 64, 56, 59, 109, 131, 121, 111, 149, 180, 156, 79, 
    134, 122, 135, 154, 179, 171, 182, 151, 131, 151, 89, 42, 67, 77, 89, 79, 73, 91, 101, 106, 112, 92, 78, 102, 145, 146, 128, 167, 139, 74, 
    138, 141, 154, 150, 164, 156, 159, 153, 126, 134, 132, 90, 83, 88, 100, 100, 90, 81, 82, 87, 86, 97, 99, 99, 107, 142, 145, 153, 152, 98, 
    149, 155, 169, 165, 154, 133, 134, 148, 144, 109, 140, 137, 83, 82, 89, 93, 113, 106, 100, 112, 100, 89, 101, 103, 109, 121, 111, 118, 136, 138, 
    166, 171, 151, 142, 146, 122, 126, 145, 171, 135, 105, 135, 118, 95, 118, 118, 100, 112, 122, 111, 88, 85, 94, 99, 118, 116, 104, 118, 111, 150, 
    171, 152, 114, 119, 139, 120, 129, 142, 134, 162, 117, 77, 108, 120, 121, 134, 119, 111, 123, 119, 90, 91, 99, 94, 102, 118, 133, 137, 147, 182, 
    165, 107, 93, 147, 142, 129, 142, 154, 134, 141, 156, 86, 78, 121, 128, 123, 132, 130, 108, 102, 91, 81, 77, 84, 88, 109, 118, 140, 199, 220, 
    141, 95, 86, 129, 147, 137, 138, 161, 180, 146, 134, 129, 94, 102, 117, 125, 128, 134, 121, 92, 73, 89, 85, 88, 95, 107, 116, 153, 214, 207, 
    123, 111, 145, 170, 163, 157, 137, 146, 179, 166, 114, 111, 128, 99, 102, 123, 117, 116, 111, 94, 89, 89, 87, 94, 87, 102, 137, 172, 201, 194, 
    155, 178, 195, 198, 184, 166, 162, 163, 155, 149, 151, 127, 119, 109, 111, 127, 113, 111, 109, 87, 102, 109, 94, 87, 81, 96, 124, 153, 191, 189, 
    146, 154, 160, 180, 193, 188, 168, 176, 171, 139, 154, 179, 155, 135, 140, 131, 107, 94, 106, 103, 103, 120, 98, 71, 95, 123, 99, 130, 188, 178, 
    129, 115, 99, 141, 171, 191, 187, 167, 171, 172, 152, 149, 157, 155, 143, 109, 73, 77, 95, 113, 103, 92, 103, 104, 114, 120, 93, 129, 162, 143, 
    132, 119, 64, 78, 125, 157, 175, 186, 176, 174, 177, 159, 155, 164, 152, 131, 82, 70, 100, 103, 104, 114, 100, 107, 129, 98, 85, 134, 132, 109, 
    142, 126, 62, 42, 66, 132, 158, 186, 194, 179, 173, 176, 175, 167, 160, 163, 138, 102, 96, 105, 99, 119, 124, 117, 109, 84, 108, 116, 103, 163, 
    148, 122, 90, 76, 48, 84, 143, 172, 202, 210, 191, 177, 184, 175, 150, 130, 113, 117, 115, 127, 131, 139, 133, 125, 117, 102, 113, 92, 115, 187, 
    
    -- channel=66
    12, 30, 32, 15, 7, 40, 50, 48, 51, 50, 10, 7, 20, 29, 35, 12, 19, 33, 35, 29, 35, 50, 31, 0, 8, 60, 15, 20, 27, 18, 
    28, 32, 35, 8, 20, 53, 48, 45, 54, 41, 5, 16, 27, 38, 36, 8, 22, 37, 33, 24, 32, 54, 26, 0, 9, 61, 9, 7, 14, 28, 
    42, 21, 36, 10, 39, 55, 45, 42, 55, 30, 8, 25, 33, 36, 25, 6, 24, 36, 28, 24, 30, 52, 22, 0, 6, 49, 4, 11, 26, 48, 
    41, 16, 36, 21, 51, 49, 47, 40, 56, 25, 13, 22, 27, 22, 22, 24, 40, 43, 38, 37, 25, 46, 22, 0, 2, 47, 25, 34, 38, 43, 
    40, 40, 37, 32, 45, 42, 51, 34, 54, 19, 5, 5, 17, 22, 32, 45, 49, 34, 46, 48, 7, 34, 31, 0, 5, 56, 40, 42, 27, 38, 
    39, 61, 23, 28, 32, 35, 45, 28, 50, 8, 0, 6, 24, 31, 49, 57, 40, 18, 48, 40, 0, 30, 36, 2, 14, 60, 38, 41, 23, 62, 
    43, 55, 4, 21, 32, 36, 31, 22, 38, 0, 0, 27, 32, 44, 60, 38, 11, 15, 40, 17, 0, 28, 30, 18, 26, 61, 39, 45, 30, 79, 
    47, 44, 2, 27, 35, 44, 22, 15, 17, 0, 7, 30, 30, 54, 42, 0, 0, 28, 30, 5, 0, 20, 28, 25, 28, 60, 45, 47, 41, 87, 
    52, 44, 14, 42, 42, 51, 30, 18, 6, 0, 21, 20, 30, 44, 8, 0, 10, 35, 19, 9, 14, 30, 47, 11, 24, 58, 46, 51, 51, 83, 
    53, 46, 17, 49, 51, 49, 46, 30, 7, 20, 31, 4, 14, 9, 0, 0, 25, 29, 17, 17, 16, 43, 47, 0, 28, 58, 49, 56, 46, 69, 
    53, 43, 16, 51, 54, 49, 54, 24, 0, 22, 13, 0, 0, 0, 0, 7, 12, 9, 11, 7, 5, 18, 10, 0, 30, 59, 56, 54, 39, 64, 
    51, 37, 17, 51, 54, 51, 46, 9, 0, 0, 0, 0, 0, 0, 0, 6, 4, 1, 0, 0, 0, 0, 0, 0, 25, 61, 57, 43, 45, 58, 
    42, 30, 19, 40, 53, 45, 46, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 41, 44, 41, 52, 44, 
    48, 33, 26, 37, 53, 36, 48, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 37, 45, 57, 52, 
    51, 37, 35, 42, 45, 36, 44, 32, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 23, 47, 73, 55, 
    40, 30, 34, 35, 45, 43, 49, 47, 4, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 16, 41, 64, 34, 
    35, 23, 34, 32, 63, 46, 57, 43, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 28, 36, 45, 41, 
    39, 21, 42, 37, 65, 42, 49, 35, 31, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 37, 36, 40, 36, 
    42, 37, 60, 38, 54, 47, 28, 37, 33, 41, 20, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 18, 36, 36, 23, 
    48, 62, 45, 23, 46, 47, 20, 46, 46, 31, 43, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 23, 37, 19, 34, 
    57, 60, 7, 14, 41, 42, 30, 40, 43, 24, 38, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 38, 28, 26, 64, 
    55, 31, 0, 6, 25, 43, 43, 33, 38, 40, 36, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 19, 23, 58, 75, 
    35, 0, 0, 0, 7, 32, 41, 36, 49, 56, 36, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 34, 72, 62, 
    21, 1, 0, 6, 2, 12, 23, 32, 53, 51, 28, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 37, 67, 52, 
    44, 42, 32, 15, 6, 7, 13, 22, 39, 39, 28, 27, 15, 0, 0, 13, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 26, 57, 58, 
    37, 48, 35, 20, 16, 14, 11, 11, 19, 32, 38, 42, 32, 16, 22, 32, 21, 0, 0, 0, 0, 0, 0, 0, 0, 19, 33, 13, 59, 59, 
    21, 41, 31, 26, 15, 19, 8, 3, 8, 19, 27, 30, 26, 25, 20, 20, 15, 0, 0, 0, 0, 0, 0, 0, 10, 36, 8, 26, 57, 20, 
    24, 39, 21, 25, 3, 10, 12, 10, 5, 9, 17, 19, 19, 25, 18, 23, 18, 0, 0, 0, 0, 0, 0, 0, 25, 23, 2, 49, 9, 0, 
    29, 41, 6, 19, 4, 8, 14, 14, 10, 11, 13, 13, 15, 31, 24, 26, 24, 10, 0, 0, 0, 5, 11, 2, 15, 11, 17, 32, 0, 0, 
    42, 51, 0, 22, 15, 12, 12, 14, 25, 26, 21, 16, 17, 24, 5, 0, 0, 11, 3, 34, 29, 21, 11, 0, 11, 10, 14, 4, 2, 16, 
    
    -- channel=67
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=68
    60, 44, 33, 23, 33, 45, 43, 42, 45, 20, 19, 48, 57, 51, 51, 61, 80, 92, 90, 88, 75, 59, 52, 86, 99, 51, 62, 66, 38, 39, 
    68, 57, 32, 32, 59, 52, 43, 45, 43, 16, 26, 62, 71, 59, 50, 68, 69, 62, 58, 70, 77, 54, 47, 98, 112, 41, 31, 34, 33, 55, 
    70, 56, 30, 53, 72, 52, 47, 51, 39, 18, 41, 59, 66, 47, 25, 59, 77, 60, 54, 74, 84, 53, 49, 101, 113, 30, 28, 55, 66, 69, 
    67, 84, 56, 74, 71, 48, 55, 61, 36, 22, 36, 35, 37, 31, 27, 61, 80, 68, 65, 89, 89, 47, 54, 105, 112, 50, 55, 79, 85, 58, 
    63, 104, 81, 79, 57, 45, 52, 64, 37, 25, 17, 22, 32, 45, 57, 79, 87, 60, 54, 69, 75, 48, 63, 104, 118, 78, 68, 75, 76, 67, 
    65, 67, 63, 57, 57, 59, 41, 57, 37, 22, 19, 50, 67, 77, 87, 81, 71, 69, 48, 24, 63, 67, 59, 113, 138, 90, 77, 71, 80, 87, 
    62, 30, 42, 41, 47, 69, 49, 45, 18, 17, 55, 85, 85, 98, 83, 32, 15, 80, 65, 14, 63, 69, 61, 121, 149, 101, 89, 80, 99, 76, 
    53, 30, 62, 69, 50, 51, 66, 60, 11, 32, 80, 82, 94, 95, 42, 10, 32, 75, 55, 38, 82, 81, 102, 121, 139, 101, 92, 84, 104, 60, 
    48, 41, 79, 97, 81, 38, 49, 73, 47, 75, 99, 90, 85, 39, 3, 35, 91, 70, 56, 86, 101, 107, 122, 119, 125, 102, 90, 86, 96, 38, 
    50, 44, 84, 98, 107, 55, 30, 42, 54, 97, 113, 108, 81, 21, 7, 54, 80, 79, 94, 107, 116, 111, 68, 95, 122, 107, 92, 87, 85, 23, 
    58, 43, 84, 104, 110, 94, 45, 9, 52, 93, 93, 98, 86, 78, 98, 99, 88, 100, 111, 95, 111, 89, 53, 115, 125, 102, 105, 93, 86, 29, 
    42, 25, 71, 91, 105, 113, 74, 55, 95, 91, 84, 107, 86, 86, 114, 125, 122, 110, 99, 94, 94, 77, 79, 128, 124, 91, 91, 93, 95, 26, 
    45, 32, 65, 71, 99, 109, 99, 105, 111, 108, 112, 117, 98, 85, 92, 100, 100, 103, 106, 117, 104, 100, 87, 103, 126, 93, 79, 104, 92, 31, 
    65, 56, 75, 77, 76, 101, 108, 113, 80, 81, 114, 126, 114, 116, 113, 93, 84, 91, 101, 107, 109, 124, 104, 100, 99, 91, 91, 101, 89, 67, 
    61, 54, 73, 81, 55, 89, 101, 115, 120, 83, 76, 106, 109, 111, 110, 121, 127, 103, 90, 86, 75, 100, 135, 133, 84, 89, 98, 94, 80, 50, 
    60, 44, 65, 79, 81, 93, 104, 100, 152, 137, 43, 58, 104, 108, 111, 120, 119, 127, 127, 131, 112, 100, 114, 129, 142, 100, 97, 103, 52, 18, 
    66, 59, 62, 78, 97, 96, 106, 87, 110, 167, 87, 64, 106, 122, 129, 116, 104, 117, 119, 120, 126, 120, 103, 121, 133, 115, 118, 117, 59, 24, 
    64, 76, 82, 103, 78, 94, 84, 91, 70, 121, 156, 113, 91, 110, 105, 112, 129, 115, 109, 115, 120, 126, 115, 120, 93, 112, 84, 84, 90, 42, 
    66, 95, 101, 95, 62, 81, 68, 95, 105, 65, 135, 159, 107, 107, 103, 111, 124, 125, 126, 123, 108, 114, 116, 115, 112, 74, 47, 55, 59, 47, 
    79, 108, 76, 69, 65, 54, 74, 70, 104, 72, 61, 120, 128, 113, 121, 125, 107, 122, 145, 126, 109, 123, 125, 113, 117, 67, 74, 57, 26, 66, 
    92, 73, 67, 86, 68, 50, 87, 60, 44, 99, 64, 62, 112, 128, 132, 129, 121, 113, 124, 127, 117, 115, 121, 108, 101, 87, 80, 51, 69, 96, 
    90, 37, 47, 68, 63, 58, 77, 89, 53, 83, 104, 77, 95, 137, 140, 128, 139, 119, 114, 115, 110, 111, 120, 108, 111, 111, 66, 63, 105, 95, 
    64, 44, 77, 85, 81, 65, 60, 86, 105, 74, 74, 90, 115, 130, 142, 135, 131, 122, 111, 109, 111, 106, 116, 121, 123, 112, 90, 101, 100, 87, 
    84, 123, 167, 144, 113, 85, 74, 84, 99, 90, 61, 77, 118, 122, 139, 145, 140, 133, 112, 104, 123, 113, 121, 130, 110, 90, 108, 111, 87, 88, 
    97, 139, 182, 179, 156, 123, 97, 104, 83, 77, 102, 109, 128, 128, 143, 146, 144, 141, 124, 97, 138, 135, 116, 103, 104, 95, 85, 92, 81, 106, 
    76, 86, 133, 174, 183, 163, 130, 108, 94, 80, 99, 113, 115, 130, 115, 81, 90, 121, 125, 122, 122, 121, 120, 106, 112, 107, 54, 70, 94, 97, 
    73, 56, 71, 132, 163, 171, 161, 129, 111, 99, 91, 95, 99, 119, 100, 51, 46, 100, 129, 136, 121, 120, 113, 118, 119, 86, 29, 98, 103, 39, 
    81, 52, 30, 52, 120, 152, 167, 165, 134, 105, 98, 98, 97, 102, 110, 107, 88, 112, 130, 118, 123, 127, 115, 113, 92, 37, 59, 98, 76, 91, 
    88, 73, 46, 19, 65, 124, 160, 179, 176, 144, 115, 103, 103, 100, 104, 96, 97, 118, 125, 122, 143, 152, 127, 92, 45, 23, 64, 14, 63, 149, 
    102, 71, 65, 38, 32, 82, 134, 158, 176, 184, 161, 131, 117, 110, 111, 84, 65, 78, 102, 115, 116, 99, 80, 75, 53, 53, 58, 40, 97, 135, 
    
    -- channel=69
    0, 0, 11, 0, 0, 0, 0, 0, 3, 25, 0, 0, 0, 0, 9, 0, 0, 2, 10, 2, 0, 11, 3, 0, 0, 21, 0, 8, 5, 0, 
    0, 4, 11, 0, 0, 0, 0, 0, 11, 18, 0, 0, 0, 8, 10, 0, 0, 0, 2, 0, 0, 14, 0, 0, 0, 27, 0, 0, 0, 0, 
    1, 2, 5, 0, 0, 2, 0, 0, 18, 7, 0, 0, 8, 10, 0, 0, 0, 0, 0, 0, 1, 14, 0, 0, 8, 24, 0, 0, 0, 0, 
    13, 0, 4, 0, 6, 0, 0, 0, 19, 0, 0, 0, 2, 0, 0, 0, 2, 4, 0, 8, 9, 10, 0, 0, 6, 4, 0, 0, 0, 17, 
    0, 18, 13, 0, 2, 0, 4, 4, 23, 8, 0, 0, 0, 0, 0, 0, 8, 0, 0, 27, 5, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 24, 4, 0, 0, 0, 3, 3, 31, 12, 0, 0, 0, 0, 0, 26, 27, 0, 3, 12, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 
    2, 21, 0, 0, 0, 1, 0, 0, 31, 0, 0, 0, 0, 0, 32, 22, 0, 0, 21, 0, 0, 4, 0, 0, 1, 18, 0, 0, 0, 31, 
    8, 7, 0, 0, 0, 6, 6, 8, 5, 0, 0, 0, 0, 32, 48, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 49, 
    2, 0, 0, 0, 0, 0, 5, 28, 0, 0, 0, 0, 4, 42, 3, 0, 0, 7, 0, 0, 0, 0, 18, 0, 0, 6, 0, 0, 4, 48, 
    8, 1, 0, 0, 9, 0, 0, 14, 0, 0, 0, 8, 29, 4, 0, 0, 0, 0, 0, 0, 0, 7, 18, 0, 0, 3, 0, 0, 9, 34, 
    18, 3, 0, 0, 13, 1, 0, 0, 0, 0, 5, 8, 37, 6, 0, 0, 0, 0, 0, 0, 10, 33, 0, 0, 0, 7, 0, 0, 5, 27, 
    16, 0, 0, 0, 1, 18, 14, 0, 0, 2, 0, 0, 0, 0, 8, 15, 10, 4, 6, 0, 5, 0, 0, 0, 2, 2, 1, 0, 11, 38, 
    5, 0, 0, 0, 1, 4, 0, 0, 12, 5, 3, 15, 5, 0, 0, 1, 11, 13, 9, 9, 10, 0, 0, 0, 13, 13, 0, 0, 29, 29, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 13, 10, 1, 0, 0, 0, 0, 0, 8, 17, 14, 0, 0, 9, 4, 0, 0, 23, 24, 
    10, 0, 0, 0, 0, 0, 0, 26, 0, 0, 13, 9, 0, 5, 12, 2, 4, 0, 0, 0, 0, 5, 9, 9, 0, 0, 0, 0, 18, 37, 
    4, 0, 0, 0, 0, 0, 0, 7, 22, 1, 0, 0, 0, 0, 0, 5, 23, 12, 9, 8, 0, 0, 9, 20, 4, 5, 0, 2, 35, 11, 
    5, 0, 0, 0, 9, 0, 12, 0, 11, 42, 1, 0, 0, 4, 9, 2, 0, 0, 0, 8, 24, 4, 0, 0, 44, 15, 15, 28, 12, 0, 
    0, 0, 0, 0, 11, 0, 12, 0, 0, 25, 13, 0, 0, 0, 10, 3, 2, 3, 0, 0, 4, 9, 0, 1, 0, 18, 24, 20, 24, 0, 
    0, 0, 16, 15, 0, 7, 0, 4, 0, 0, 22, 32, 7, 0, 0, 0, 12, 2, 0, 9, 8, 0, 3, 13, 0, 25, 0, 0, 21, 0, 
    0, 17, 23, 0, 0, 4, 0, 0, 29, 0, 0, 24, 9, 0, 0, 0, 0, 0, 9, 19, 8, 1, 3, 9, 26, 14, 0, 7, 0, 0, 
    0, 41, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 11, 14, 1, 6, 6, 10, 9, 0, 20, 3, 0, 0, 
    23, 0, 0, 0, 0, 0, 3, 2, 0, 0, 14, 0, 0, 1, 7, 3, 11, 6, 0, 14, 6, 1, 5, 8, 3, 6, 6, 0, 0, 5, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 4, 7, 9, 6, 14, 7, 0, 1, 2, 7, 12, 21, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 17, 0, 0, 0, 1, 1, 19, 15, 6, 7, 13, 0, 0, 3, 14, 6, 3, 17, 3, 0, 0, 
    0, 11, 32, 27, 2, 0, 0, 0, 0, 1, 0, 0, 3, 0, 7, 31, 30, 16, 11, 0, 0, 11, 11, 13, 0, 1, 26, 0, 0, 0, 
    0, 5, 23, 22, 29, 7, 0, 0, 0, 0, 0, 4, 6, 0, 6, 15, 6, 0, 7, 0, 9, 14, 13, 0, 8, 32, 18, 0, 0, 17, 
    0, 0, 0, 18, 21, 24, 6, 0, 0, 0, 0, 0, 0, 6, 8, 0, 0, 0, 0, 25, 2, 0, 15, 7, 19, 58, 0, 0, 20, 0, 
    0, 4, 0, 0, 5, 9, 9, 2, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 5, 10, 4, 8, 6, 7, 37, 19, 0, 34, 20, 0, 
    5, 34, 0, 0, 0, 5, 7, 14, 10, 0, 0, 0, 0, 0, 0, 0, 0, 5, 13, 9, 7, 26, 32, 11, 5, 0, 0, 4, 0, 0, 
    9, 50, 0, 0, 0, 0, 9, 10, 15, 20, 4, 0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 24, 15, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=70
    13, 11, 12, 17, 16, 11, 15, 18, 24, 26, 33, 25, 26, 26, 23, 31, 25, 30, 32, 27, 19, 12, 15, 16, 12, 12, 42, 28, 10, 12, 
    5, 14, 4, 15, 14, 13, 13, 17, 21, 29, 39, 34, 41, 34, 27, 30, 17, 7, 11, 16, 17, 11, 13, 14, 10, 0, 11, 0, 0, 11, 
    0, 6, 0, 18, 15, 14, 13, 18, 19, 36, 46, 47, 40, 26, 12, 13, 16, 12, 12, 19, 24, 12, 11, 6, 0, 0, 0, 1, 6, 5, 
    8, 20, 16, 22, 19, 15, 14, 28, 22, 40, 39, 31, 11, 4, 7, 14, 16, 19, 24, 32, 39, 8, 3, 3, 0, 0, 0, 1, 3, 0, 
    25, 27, 46, 28, 16, 12, 13, 33, 27, 34, 20, 4, 0, 4, 14, 30, 37, 29, 16, 27, 34, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 20, 29, 12, 14, 16, 13, 29, 28, 27, 8, 2, 12, 24, 43, 52, 37, 33, 7, 5, 23, 7, 0, 0, 0, 0, 0, 0, 4, 11, 
    17, 8, 7, 0, 0, 8, 22, 18, 9, 15, 8, 12, 23, 39, 48, 34, 11, 6, 18, 2, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 
    4, 6, 7, 0, 0, 0, 21, 26, 2, 2, 1, 10, 30, 42, 30, 9, 7, 0, 0, 0, 0, 2, 12, 20, 0, 0, 0, 0, 12, 14, 
    7, 9, 15, 0, 0, 0, 1, 23, 25, 7, 8, 19, 16, 6, 0, 3, 9, 5, 0, 0, 8, 15, 25, 34, 0, 0, 0, 0, 10, 10, 
    5, 16, 18, 0, 0, 0, 0, 1, 17, 8, 16, 20, 1, 0, 0, 0, 0, 0, 12, 15, 23, 18, 0, 2, 0, 0, 0, 0, 5, 12, 
    16, 23, 25, 5, 0, 0, 0, 0, 0, 6, 8, 9, 1, 11, 13, 3, 0, 5, 14, 16, 11, 13, 0, 5, 1, 0, 1, 0, 4, 13, 
    4, 7, 17, 3, 1, 0, 0, 0, 0, 9, 4, 12, 14, 8, 12, 18, 20, 17, 3, 1, 0, 2, 4, 11, 13, 0, 0, 0, 1, 0, 
    0, 7, 8, 3, 0, 4, 0, 0, 6, 22, 21, 14, 7, 4, 0, 1, 5, 8, 14, 11, 3, 0, 0, 0, 6, 8, 0, 0, 0, 1, 
    7, 15, 14, 7, 0, 2, 0, 0, 0, 0, 13, 36, 16, 11, 7, 0, 0, 0, 5, 9, 5, 5, 0, 0, 0, 0, 0, 0, 14, 31, 
    8, 8, 7, 0, 0, 0, 0, 0, 3, 0, 0, 20, 15, 0, 0, 2, 7, 0, 0, 0, 0, 0, 2, 0, 0, 0, 6, 9, 10, 17, 
    2, 0, 0, 0, 0, 2, 3, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 2, 7, 4, 9, 1, 0, 0, 1, 4, 0, 14, 0, 0, 
    0, 0, 0, 1, 2, 21, 6, 14, 0, 0, 2, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 4, 1, 4, 0, 19, 30, 28, 15, 0, 
    0, 0, 2, 20, 11, 19, 12, 5, 5, 0, 24, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 13, 6, 28, 17, 21, 3, 
    0, 10, 16, 20, 13, 10, 20, 5, 30, 12, 0, 33, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 2, 0, 0, 0, 
    4, 13, 17, 6, 6, 5, 16, 9, 1, 30, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 2, 9, 3, 3, 4, 2, 0, 0, 0, 
    11, 3, 17, 11, 3, 6, 7, 5, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 1, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 8, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 11, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 13, 19, 22, 12, 0, 2, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 10, 1, 0, 0, 0, 0, 0, 6, 16, 18, 25, 30, 0, 5, 
    22, 26, 33, 12, 0, 0, 0, 0, 0, 0, 5, 14, 0, 14, 24, 34, 36, 16, 0, 0, 0, 4, 0, 0, 12, 27, 23, 30, 7, 20, 
    23, 24, 48, 50, 24, 3, 0, 0, 0, 2, 0, 7, 10, 14, 14, 6, 6, 12, 0, 0, 0, 0, 0, 13, 16, 29, 28, 18, 16, 20, 
    16, 24, 47, 58, 57, 14, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 21, 36, 24, 25, 19, 20, 0, 
    7, 14, 33, 30, 52, 47, 10, 0, 0, 0, 0, 0, 0, 0, 7, 11, 16, 9, 6, 0, 0, 2, 14, 22, 16, 18, 34, 13, 6, 0, 
    18, 22, 40, 21, 34, 55, 48, 11, 0, 0, 0, 0, 0, 0, 1, 0, 6, 25, 24, 21, 37, 38, 24, 6, 0, 0, 0, 0, 0, 3, 
    41, 37, 40, 21, 29, 44, 61, 50, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 25, 29, 27, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=71
    77, 70, 84, 95, 87, 100, 101, 80, 58, 78, 87, 89, 86, 80, 100, 100, 100, 107, 116, 109, 90, 101, 134, 105, 61, 105, 86, 89, 102, 80, 
    90, 74, 102, 99, 95, 108, 103, 74, 62, 79, 80, 83, 76, 74, 105, 104, 103, 111, 121, 111, 86, 106, 135, 106, 68, 117, 103, 104, 96, 71, 
    104, 82, 114, 98, 103, 107, 99, 65, 64, 69, 67, 74, 78, 83, 109, 106, 101, 106, 111, 107, 83, 113, 136, 116, 86, 128, 111, 105, 94, 94, 
    98, 82, 99, 96, 104, 95, 91, 55, 64, 66, 75, 87, 97, 101, 110, 105, 104, 99, 92, 106, 86, 115, 141, 123, 96, 129, 115, 120, 112, 115, 
    76, 84, 91, 98, 102, 82, 84, 49, 68, 80, 97, 110, 121, 109, 97, 99, 107, 80, 80, 115, 92, 116, 151, 129, 103, 132, 127, 139, 107, 95, 
    67, 106, 98, 105, 96, 73, 75, 46, 80, 102, 113, 132, 130, 98, 84, 88, 105, 72, 77, 124, 94, 122, 154, 138, 106, 134, 130, 136, 80, 68, 
    82, 130, 116, 112, 95, 83, 71, 54, 102, 116, 124, 147, 122, 92, 94, 108, 102, 81, 91, 119, 110, 139, 162, 147, 115, 131, 124, 123, 55, 60, 
    94, 138, 121, 121, 92, 92, 76, 69, 117, 122, 135, 138, 99, 92, 113, 119, 106, 111, 123, 126, 125, 139, 165, 151, 123, 134, 122, 110, 42, 60, 
    97, 133, 121, 126, 103, 91, 80, 89, 114, 115, 131, 111, 89, 111, 124, 121, 121, 142, 141, 141, 130, 127, 167, 145, 127, 137, 120, 102, 41, 66, 
    91, 125, 117, 131, 120, 94, 92, 117, 119, 116, 118, 88, 95, 123, 129, 133, 141, 149, 139, 140, 120, 132, 178, 145, 132, 140, 119, 100, 44, 65, 
    78, 115, 107, 129, 129, 111, 120, 140, 125, 124, 111, 71, 77, 98, 98, 115, 126, 126, 127, 116, 107, 125, 159, 133, 128, 140, 122, 96, 50, 73, 
    88, 116, 106, 123, 135, 124, 130, 124, 115, 111, 96, 68, 77, 88, 83, 90, 96, 102, 102, 89, 97, 105, 130, 124, 123, 143, 134, 102, 70, 96, 
    97, 112, 108, 110, 135, 128, 122, 102, 92, 84, 79, 75, 88, 89, 86, 84, 80, 80, 74, 67, 85, 85, 107, 104, 115, 135, 137, 105, 82, 100, 
    97, 109, 107, 105, 133, 129, 119, 117, 88, 69, 82, 76, 82, 86, 88, 86, 80, 77, 75, 64, 82, 83, 91, 91, 101, 128, 125, 94, 73, 95, 
    103, 115, 117, 120, 132, 132, 115, 121, 89, 49, 89, 85, 85, 90, 86, 81, 82, 87, 96, 86, 88, 85, 88, 86, 84, 113, 114, 79, 78, 119, 
    112, 118, 126, 115, 123, 117, 116, 110, 102, 65, 91, 91, 84, 83, 81, 82, 84, 83, 80, 77, 83, 80, 93, 75, 72, 87, 105, 79, 83, 124, 
    121, 118, 128, 102, 116, 105, 118, 108, 103, 93, 78, 75, 81, 70, 81, 85, 85, 91, 90, 83, 91, 84, 89, 71, 60, 66, 81, 85, 89, 129, 
    127, 103, 116, 87, 108, 108, 116, 119, 95, 102, 80, 64, 90, 85, 86, 85, 85, 91, 82, 77, 88, 84, 85, 76, 54, 67, 83, 92, 111, 135, 
    113, 89, 106, 92, 104, 117, 102, 112, 101, 86, 90, 75, 83, 92, 87, 81, 90, 90, 75, 77, 91, 85, 79, 78, 59, 85, 89, 106, 133, 138, 
    90, 100, 108, 100, 105, 122, 101, 103, 125, 95, 99, 103, 95, 91, 87, 89, 83, 83, 71, 71, 77, 77, 70, 76, 67, 83, 93, 120, 131, 133, 
    83, 112, 109, 100, 105, 120, 112, 115, 128, 117, 108, 117, 104, 96, 86, 92, 81, 78, 72, 78, 74, 80, 76, 79, 75, 82, 113, 125, 118, 133, 
    110, 141, 127, 126, 118, 123, 129, 120, 117, 113, 116, 115, 100, 98, 85, 87, 79, 76, 75, 85, 78, 82, 75, 80, 76, 96, 124, 119, 128, 147, 
    145, 153, 137, 139, 140, 144, 147, 121, 112, 119, 119, 120, 94, 97, 82, 85, 86, 76, 76, 94, 75, 81, 73, 78, 77, 100, 117, 111, 148, 154, 
    129, 126, 129, 148, 156, 163, 160, 129, 119, 133, 127, 115, 103, 89, 69, 74, 83, 74, 77, 95, 74, 68, 66, 80, 76, 85, 116, 119, 155, 140, 
    104, 114, 134, 145, 160, 166, 169, 154, 140, 135, 122, 104, 94, 73, 49, 64, 82, 75, 80, 82, 73, 68, 72, 79, 62, 60, 125, 126, 140, 129, 
    87, 102, 126, 134, 145, 167, 171, 171, 163, 150, 135, 124, 110, 91, 80, 88, 108, 87, 79, 82, 77, 73, 75, 61, 40, 71, 129, 118, 135, 127, 
    75, 83, 99, 128, 136, 161, 172, 170, 167, 170, 163, 154, 141, 130, 122, 116, 120, 96, 74, 81, 83, 69, 69, 46, 44, 98, 108, 124, 153, 135, 
    77, 90, 82, 117, 133, 151, 164, 168, 171, 178, 182, 181, 168, 159, 136, 116, 108, 89, 76, 84, 76, 64, 67, 53, 74, 106, 88, 140, 158, 120, 
    75, 105, 76, 102, 114, 140, 151, 158, 166, 173, 181, 186, 176, 181, 161, 131, 111, 95, 62, 65, 54, 59, 85, 89, 113, 123, 120, 169, 159, 116, 
    75, 118, 86, 97, 96, 116, 146, 150, 158, 164, 170, 173, 172, 187, 180, 150, 123, 115, 76, 80, 86, 105, 129, 120, 131, 129, 143, 157, 156, 139, 
    
    -- channel=72
    128, 97, 101, 132, 130, 116, 107, 99, 74, 78, 141, 154, 140, 128, 143, 185, 196, 195, 196, 187, 157, 127, 186, 220, 165, 135, 170, 154, 140, 134, 
    127, 105, 116, 155, 142, 118, 110, 96, 72, 95, 153, 158, 144, 128, 156, 191, 176, 170, 184, 184, 150, 128, 196, 232, 160, 118, 150, 143, 134, 118, 
    128, 128, 132, 164, 139, 118, 110, 94, 72, 107, 147, 149, 135, 122, 155, 182, 157, 144, 164, 176, 152, 133, 200, 232, 162, 120, 146, 149, 138, 107, 
    143, 143, 148, 159, 132, 116, 108, 97, 75, 107, 134, 140, 139, 132, 148, 170, 160, 149, 159, 172, 164, 149, 200, 233, 177, 135, 159, 165, 151, 128, 
    156, 162, 165, 156, 134, 111, 106, 101, 75, 108, 139, 154, 158, 160, 157, 152, 147, 144, 129, 165, 184, 156, 203, 239, 190, 150, 164, 166, 167, 143, 
    135, 145, 178, 156, 135, 109, 105, 103, 83, 137, 177, 193, 201, 187, 155, 150, 165, 135, 98, 150, 196, 170, 225, 250, 199, 153, 164, 163, 159, 122, 
    114, 126, 161, 144, 136, 118, 111, 102, 110, 183, 209, 225, 223, 174, 140, 150, 185, 151, 108, 152, 207, 204, 248, 269, 213, 162, 167, 161, 134, 74, 
    110, 134, 169, 133, 120, 124, 125, 107, 138, 203, 218, 227, 195, 145, 139, 169, 172, 162, 166, 183, 225, 233, 255, 271, 226, 176, 167, 155, 110, 50, 
    108, 150, 189, 157, 112, 105, 138, 141, 177, 211, 210, 194, 151, 129, 161, 199, 192, 190, 214, 226, 247, 236, 262, 281, 229, 178, 159, 138, 93, 53, 
    107, 153, 196, 172, 135, 93, 105, 165, 215, 219, 214, 186, 130, 129, 165, 199, 215, 230, 236, 246, 233, 209, 255, 283, 229, 181, 155, 130, 88, 57, 
    107, 155, 199, 178, 163, 112, 90, 161, 213, 215, 218, 206, 180, 178, 184, 196, 209, 230, 234, 242, 226, 208, 241, 267, 229, 189, 162, 141, 94, 59, 
    108, 150, 189, 184, 180, 155, 129, 168, 205, 227, 231, 220, 214, 235, 233, 221, 220, 221, 217, 211, 209, 220, 255, 271, 220, 187, 179, 157, 97, 70, 
    103, 138, 170, 173, 183, 188, 174, 191, 220, 239, 245, 243, 224, 227, 232, 231, 232, 228, 222, 208, 201, 204, 235, 262, 218, 193, 185, 163, 108, 98, 
    123, 147, 164, 155, 177, 198, 182, 182, 214, 235, 237, 251, 252, 241, 227, 222, 221, 229, 235, 228, 223, 212, 208, 212, 216, 204, 190, 164, 120, 128, 
    135, 158, 168, 154, 161, 188, 187, 192, 191, 185, 203, 245, 247, 252, 253, 238, 226, 225, 227, 217, 229, 237, 215, 192, 189, 200, 193, 146, 104, 146, 
    134, 157, 167, 169, 151, 176, 178, 211, 219, 162, 154, 213, 227, 232, 238, 247, 256, 245, 243, 227, 215, 228, 241, 228, 179, 187, 192, 135, 95, 149, 
    145, 153, 166, 173, 162, 179, 176, 195, 227, 200, 157, 180, 218, 234, 220, 224, 235, 246, 254, 255, 249, 230, 226, 229, 218, 183, 184, 154, 106, 145, 
    154, 166, 159, 163, 159, 174, 178, 184, 194, 223, 206, 179, 203, 224, 223, 227, 221, 224, 228, 220, 239, 245, 227, 212, 198, 170, 178, 173, 138, 148, 
    156, 157, 162, 170, 146, 166, 182, 186, 167, 196, 234, 205, 196, 208, 203, 214, 230, 231, 220, 207, 223, 239, 228, 212, 172, 139, 142, 136, 169, 176, 
    148, 142, 169, 171, 137, 159, 168, 178, 185, 159, 192, 233, 219, 217, 210, 197, 215, 229, 223, 207, 218, 230, 227, 214, 183, 143, 124, 118, 159, 181, 
    133, 154, 187, 174, 152, 155, 156, 141, 179, 170, 145, 200, 242, 229, 220, 214, 200, 204, 220, 213, 221, 235, 233, 222, 207, 174, 150, 152, 156, 168, 
    128, 159, 214, 197, 182, 176, 174, 153, 144, 177, 168, 185, 235, 248, 235, 223, 209, 191, 196, 215, 228, 226, 235, 237, 230, 201, 183, 181, 174, 179, 
    155, 183, 210, 214, 210, 199, 203, 196, 152, 148, 190, 208, 227, 252, 256, 230, 215, 196, 190, 204, 224, 223, 238, 249, 248, 231, 207, 194, 181, 186, 
    195, 233, 256, 248, 250, 233, 226, 215, 188, 159, 165, 203, 224, 250, 255, 232, 221, 202, 192, 216, 222, 212, 228, 242, 246, 231, 221, 208, 190, 200, 
    225, 265, 302, 298, 281, 275, 266, 238, 213, 214, 202, 196, 219, 246, 242, 229, 236, 225, 206, 223, 227, 215, 215, 228, 218, 191, 207, 224, 199, 195, 
    192, 227, 299, 318, 314, 294, 286, 276, 247, 234, 246, 245, 241, 234, 204, 197, 226, 244, 231, 212, 225, 225, 211, 217, 199, 156, 194, 220, 185, 195, 
    155, 164, 250, 306, 331, 325, 301, 283, 277, 266, 253, 265, 261, 236, 193, 159, 195, 235, 233, 226, 225, 223, 227, 216, 172, 159, 198, 185, 186, 200, 
    146, 129, 178, 256, 312, 332, 330, 300, 278, 280, 273, 275, 273, 260, 241, 199, 200, 230, 226, 225, 235, 216, 207, 197, 161, 170, 179, 196, 247, 221, 
    156, 134, 145, 181, 270, 321, 341, 331, 302, 275, 269, 278, 273, 269, 268, 250, 239, 235, 232, 224, 228, 215, 201, 175, 147, 154, 161, 212, 279, 266, 
    157, 169, 176, 153, 198, 282, 334, 350, 341, 312, 280, 270, 262, 264, 265, 243, 239, 247, 234, 208, 215, 208, 202, 176, 141, 147, 158, 200, 249, 247, 
    
    -- channel=73
    5, 0, 0, 4, 2, 0, 6, 0, 1, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 17, 0, 0, 0, 11, 0, 0, 
    5, 6, 0, 0, 2, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 1, 0, 0, 0, 19, 12, 0, 11, 17, 0, 0, 
    8, 14, 0, 0, 1, 0, 5, 2, 0, 0, 0, 0, 0, 3, 0, 5, 8, 0, 0, 0, 4, 0, 0, 25, 30, 0, 2, 7, 0, 6, 
    0, 7, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 10, 11, 0, 0, 2, 0, 0, 0, 13, 0, 0, 26, 28, 0, 0, 5, 14, 18, 
    0, 0, 0, 4, 0, 0, 0, 2, 0, 4, 13, 13, 5, 0, 0, 0, 4, 0, 0, 0, 22, 0, 0, 22, 18, 0, 0, 9, 8, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 17, 12, 6, 0, 0, 0, 0, 1, 11, 0, 0, 17, 0, 0, 9, 19, 0, 4, 2, 0, 0, 
    8, 4, 22, 5, 0, 0, 0, 0, 0, 9, 4, 1, 0, 0, 0, 2, 0, 11, 6, 0, 15, 6, 0, 0, 14, 0, 1, 0, 0, 0, 
    9, 0, 28, 20, 0, 0, 0, 14, 0, 2, 9, 0, 0, 0, 12, 15, 0, 7, 12, 0, 9, 0, 0, 0, 7, 0, 1, 0, 0, 0, 
    0, 0, 15, 24, 17, 0, 0, 9, 0, 0, 4, 0, 3, 7, 4, 0, 15, 7, 0, 0, 0, 0, 0, 3, 0, 0, 1, 0, 2, 0, 
    0, 0, 10, 9, 33, 3, 0, 0, 0, 0, 0, 8, 18, 17, 3, 3, 8, 0, 0, 0, 0, 0, 0, 9, 0, 0, 1, 0, 7, 0, 
    0, 0, 0, 2, 21, 29, 16, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 5, 0, 9, 0, 0, 3, 7, 7, 0, 
    0, 0, 0, 0, 4, 33, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 5, 6, 14, 0, 
    0, 0, 2, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 14, 0, 
    0, 0, 1, 0, 0, 4, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 15, 0, 1, 0, 4, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    4, 0, 1, 4, 0, 0, 0, 0, 11, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    9, 5, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 2, 0, 
    0, 1, 0, 0, 0, 0, 0, 4, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 4, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 23, 0, 0, 
    0, 0, 0, 2, 0, 0, 22, 5, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 0, 0, 
    15, 6, 14, 6, 0, 0, 5, 28, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 2, 
    29, 22, 20, 12, 1, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 8, 
    0, 0, 13, 15, 15, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 
    0, 0, 0, 8, 10, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 
    0, 0, 0, 0, 2, 6, 6, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 10, 7, 4, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 15, 
    9, 0, 0, 0, 0, 0, 0, 14, 13, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 24, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 12, 11, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 1, 0, 28, 0, 0, 10, 
    0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 8, 9, 9, 8, 25, 8, 0, 0, 0, 0, 0, 0, 10, 25, 10, 15, 28, 0, 3, 13, 
    
    -- channel=74
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=75
    69, 39, 0, 24, 59, 69, 76, 63, 0, 0, 5, 51, 66, 52, 60, 105, 136, 131, 132, 135, 111, 78, 121, 175, 118, 58, 42, 50, 71, 80, 
    96, 54, 37, 75, 87, 85, 88, 61, 0, 0, 22, 63, 63, 40, 61, 101, 120, 111, 121, 135, 102, 76, 134, 189, 115, 45, 41, 77, 105, 82, 
    113, 83, 86, 104, 98, 94, 96, 54, 0, 0, 8, 40, 32, 21, 72, 110, 108, 100, 117, 130, 94, 79, 142, 201, 134, 85, 92, 127, 127, 73, 
    133, 97, 107, 108, 97, 100, 95, 41, 0, 0, 0, 19, 35, 50, 95, 125, 124, 117, 117, 106, 82, 96, 156, 220, 186, 149, 147, 165, 143, 112, 
    136, 96, 92, 95, 98, 95, 84, 24, 0, 0, 1, 49, 85, 106, 115, 104, 96, 106, 84, 77, 87, 119, 172, 249, 237, 189, 173, 187, 182, 163, 
    82, 68, 79, 104, 100, 75, 68, 7, 0, 0, 73, 121, 145, 135, 84, 54, 79, 78, 39, 74, 106, 133, 203, 270, 256, 211, 191, 212, 198, 134, 
    41, 57, 92, 134, 124, 72, 49, 0, 0, 65, 139, 171, 172, 101, 14, 16, 101, 82, 30, 98, 131, 164, 234, 288, 264, 227, 213, 230, 165, 57, 
    53, 92, 143, 164, 141, 99, 46, 0, 40, 125, 173, 192, 137, 29, 0, 50, 115, 104, 95, 147, 170, 204, 230, 280, 263, 238, 226, 230, 126, 7, 
    76, 123, 191, 213, 158, 119, 74, 36, 96, 158, 180, 165, 80, 16, 54, 132, 140, 143, 169, 198, 220, 209, 207, 259, 257, 238, 231, 216, 93, 0, 
    79, 123, 196, 245, 195, 132, 81, 80, 150, 178, 177, 133, 58, 63, 137, 183, 190, 196, 204, 219, 205, 160, 201, 264, 258, 240, 233, 199, 73, 0, 
    61, 110, 186, 238, 234, 164, 101, 130, 170, 169, 166, 136, 109, 133, 169, 190, 198, 201, 195, 198, 161, 142, 204, 254, 259, 245, 221, 193, 72, 0, 
    58, 106, 168, 225, 246, 211, 176, 183, 169, 160, 157, 128, 135, 175, 191, 192, 178, 170, 170, 159, 145, 167, 216, 244, 240, 231, 226, 202, 77, 0, 
    70, 104, 149, 202, 230, 243, 239, 212, 176, 152, 146, 134, 129, 151, 165, 166, 163, 156, 160, 147, 148, 163, 204, 236, 212, 212, 235, 202, 98, 47, 
    100, 116, 149, 171, 216, 245, 240, 199, 189, 170, 139, 139, 159, 157, 149, 155, 158, 156, 160, 162, 167, 170, 199, 212, 211, 215, 231, 203, 114, 64, 
    113, 129, 157, 166, 215, 242, 239, 214, 181, 154, 132, 138, 172, 188, 197, 185, 162, 161, 166, 166, 189, 212, 210, 200, 214, 217, 216, 177, 79, 56, 
    112, 142, 171, 194, 208, 231, 228, 247, 220, 139, 136, 155, 171, 192, 207, 206, 207, 196, 195, 179, 177, 205, 233, 239, 194, 208, 203, 130, 57, 80, 
    138, 161, 197, 208, 199, 204, 200, 214, 243, 176, 170, 183, 186, 198, 193, 198, 217, 222, 227, 227, 207, 192, 222, 229, 205, 187, 163, 110, 67, 108, 
    180, 193, 203, 162, 171, 156, 182, 182, 219, 231, 198, 188, 199, 200, 220, 227, 209, 217, 223, 210, 207, 205, 212, 189, 184, 137, 130, 126, 82, 131, 
    208, 188, 173, 136, 139, 130, 172, 184, 159, 217, 212, 174, 200, 213, 231, 241, 240, 244, 237, 209, 207, 211, 206, 186, 134, 104, 102, 110, 137, 202, 
    197, 135, 141, 138, 114, 134, 150, 180, 154, 152, 193, 196, 216, 252, 255, 239, 253, 259, 230, 204, 204, 202, 193, 182, 135, 125, 96, 110, 193, 240, 
    142, 116, 139, 139, 120, 137, 132, 145, 190, 147, 147, 198, 239, 266, 270, 261, 247, 247, 229, 203, 195, 202, 189, 176, 160, 140, 129, 183, 223, 229, 
    105, 137, 185, 182, 154, 148, 159, 157, 192, 187, 152, 191, 251, 268, 269, 272, 246, 230, 207, 199, 197, 197, 189, 184, 163, 135, 172, 227, 229, 229, 
    156, 214, 242, 235, 193, 172, 195, 209, 177, 170, 188, 217, 243, 261, 264, 259, 246, 231, 205, 198, 207, 213, 203, 188, 161, 162, 189, 208, 223, 227, 
    233, 286, 296, 289, 256, 223, 219, 215, 184, 158, 193, 240, 245, 253, 249, 234, 225, 219, 210, 222, 222, 217, 193, 170, 159, 171, 171, 185, 228, 230, 
    244, 279, 302, 318, 303, 280, 262, 217, 197, 209, 214, 225, 235, 237, 210, 187, 192, 208, 212, 245, 232, 205, 180, 174, 147, 116, 133, 177, 229, 200, 
    170, 195, 239, 288, 312, 302, 289, 266, 230, 225, 236, 226, 226, 202, 157, 145, 170, 210, 233, 229, 228, 213, 182, 175, 131, 59, 113, 182, 190, 156, 
    109, 98, 142, 203, 272, 311, 309, 301, 274, 240, 226, 221, 218, 187, 144, 132, 174, 215, 230, 219, 220, 213, 198, 157, 80, 44, 133, 147, 143, 170, 
    95, 43, 47, 123, 197, 282, 325, 321, 303, 286, 262, 247, 239, 229, 207, 166, 175, 201, 205, 220, 228, 204, 171, 116, 51, 81, 110, 121, 192, 200, 
    99, 36, 5, 59, 136, 222, 296, 334, 329, 310, 300, 291, 269, 257, 243, 221, 194, 179, 185, 202, 193, 163, 135, 102, 89, 114, 93, 176, 269, 247, 
    74, 51, 35, 41, 75, 148, 231, 309, 345, 332, 321, 318, 295, 275, 253, 228, 201, 184, 166, 154, 140, 148, 170, 169, 163, 154, 158, 227, 280, 260, 
    
    -- channel=76
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 29, 13, 6, 7, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 30, 20, 9, 14, 19, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 14, 25, 22, 13, 21, 18, 0, 
    0, 0, 0, 3, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 24, 23, 20, 26, 10, 0, 
    0, 0, 7, 14, 9, 4, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 8, 22, 23, 25, 23, 5, 0, 
    0, 0, 9, 23, 15, 7, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 0, 0, 0, 0, 2, 0, 0, 10, 22, 23, 25, 19, 0, 0, 
    0, 0, 6, 17, 21, 8, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 3, 1, 0, 4, 0, 0, 0, 6, 27, 21, 13, 15, 0, 0, 
    0, 0, 6, 17, 21, 15, 0, 0, 0, 0, 0, 0, 2, 8, 8, 2, 0, 0, 0, 1, 0, 2, 2, 8, 24, 20, 15, 15, 0, 0, 
    0, 0, 1, 13, 15, 22, 13, 2, 0, 0, 0, 0, 0, 0, 4, 4, 5, 0, 0, 0, 0, 4, 13, 18, 15, 16, 17, 13, 0, 0, 
    0, 0, 0, 6, 14, 21, 17, 2, 15, 7, 0, 0, 0, 0, 0, 0, 2, 1, 1, 6, 0, 2, 15, 21, 24, 16, 23, 15, 0, 0, 
    0, 0, 1, 6, 19, 22, 18, 0, 0, 20, 0, 0, 3, 7, 4, 0, 0, 2, 4, 12, 17, 14, 10, 16, 27, 22, 24, 16, 0, 0, 
    0, 1, 4, 9, 10, 18, 14, 10, 0, 7, 13, 0, 0, 8, 14, 14, 9, 0, 0, 0, 0, 17, 24, 20, 7, 27, 21, 5, 0, 0, 
    0, 4, 13, 14, 9, 12, 8, 11, 12, 0, 13, 10, 2, 10, 7, 11, 19, 20, 20, 21, 9, 6, 17, 24, 18, 10, 5, 0, 0, 0, 
    8, 11, 5, 3, 6, 0, 6, 3, 17, 7, 0, 16, 17, 18, 23, 16, 11, 18, 18, 12, 10, 12, 13, 12, 20, 10, 8, 0, 0, 0, 
    15, 6, 3, 2, 0, 0, 4, 0, 0, 20, 0, 0, 16, 17, 23, 28, 22, 21, 27, 20, 14, 16, 15, 9, 8, 10, 1, 0, 2, 6, 
    15, 0, 2, 3, 0, 0, 1, 11, 0, 5, 13, 0, 12, 28, 28, 26, 32, 26, 19, 16, 12, 9, 11, 9, 6, 6, 0, 0, 17, 19, 
    2, 0, 0, 0, 0, 0, 0, 4, 12, 0, 0, 7, 15, 24, 34, 31, 29, 32, 23, 11, 11, 13, 11, 9, 8, 9, 3, 9, 12, 15, 
    0, 0, 13, 7, 1, 0, 0, 0, 11, 6, 0, 0, 19, 20, 28, 33, 28, 25, 18, 15, 12, 8, 8, 2, 0, 0, 12, 19, 16, 17, 
    0, 7, 12, 12, 3, 1, 6, 11, 2, 9, 8, 0, 14, 19, 25, 32, 31, 27, 18, 9, 18, 17, 9, 0, 0, 0, 3, 14, 13, 14, 
    0, 5, 12, 17, 14, 3, 0, 9, 4, 0, 12, 16, 11, 18, 19, 19, 16, 19, 21, 18, 17, 19, 9, 3, 7, 4, 0, 8, 10, 10, 
    9, 11, 11, 17, 15, 15, 7, 0, 1, 4, 1, 4, 5, 11, 10, 5, 2, 10, 18, 27, 16, 15, 13, 9, 0, 0, 0, 5, 7, 0, 
    5, 3, 0, 1, 11, 11, 16, 11, 0, 3, 9, 3, 3, 7, 12, 8, 0, 8, 20, 21, 24, 15, 5, 8, 0, 0, 0, 6, 0, 0, 
    0, 0, 0, 0, 2, 13, 14, 17, 14, 0, 0, 0, 0, 0, 0, 4, 1, 4, 17, 17, 15, 18, 14, 3, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 3, 12, 16, 24, 17, 6, 0, 0, 0, 0, 0, 0, 0, 12, 20, 18, 11, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 13, 18, 21, 24, 16, 8, 6, 6, 6, 0, 0, 3, 3, 0, 0, 0, 2, 0, 0, 0, 0, 2, 8, 
    0, 0, 0, 0, 0, 0, 0, 7, 14, 14, 20, 23, 19, 11, 5, 10, 11, 2, 1, 0, 2, 7, 10, 12, 4, 0, 0, 2, 16, 22, 
    
    -- channel=77
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 61, 22, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 75, 49, 0, 0, 4, 20, 0, 
    54, 9, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 0, 1, 0, 0, 34, 106, 101, 66, 24, 53, 48, 24, 
    37, 15, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 136, 148, 119, 58, 70, 72, 63, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 85, 160, 187, 151, 83, 102, 82, 57, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 39, 88, 172, 198, 179, 119, 137, 83, 14, 
    0, 0, 6, 56, 33, 2, 0, 0, 0, 0, 6, 21, 0, 0, 0, 0, 0, 0, 2, 22, 34, 65, 101, 158, 175, 183, 141, 149, 62, 0, 
    0, 0, 58, 129, 84, 16, 0, 0, 0, 9, 45, 16, 0, 0, 0, 0, 19, 27, 31, 74, 81, 68, 97, 132, 157, 174, 149, 139, 30, 0, 
    0, 8, 70, 149, 134, 56, 0, 0, 3, 46, 74, 46, 0, 0, 0, 13, 46, 55, 66, 96, 72, 33, 52, 94, 157, 169, 152, 133, 8, 0, 
    0, 0, 61, 152, 160, 106, 20, 0, 0, 46, 71, 61, 67, 72, 95, 98, 76, 68, 73, 75, 53, 33, 63, 105, 160, 162, 153, 131, 4, 0, 
    0, 0, 29, 126, 155, 150, 114, 68, 48, 71, 85, 75, 76, 94, 130, 135, 113, 93, 87, 73, 59, 48, 102, 132, 146, 137, 134, 120, 13, 0, 
    0, 0, 20, 88, 135, 155, 168, 145, 117, 99, 109, 105, 102, 84, 90, 99, 101, 108, 122, 125, 123, 100, 119, 121, 133, 129, 123, 113, 39, 0, 
    25, 15, 39, 73, 114, 138, 177, 154, 117, 99, 110, 114, 133, 133, 128, 113, 102, 107, 121, 133, 158, 165, 172, 135, 129, 119, 131, 110, 46, 8, 
    20, 14, 42, 74, 104, 127, 176, 200, 166, 104, 79, 84, 123, 150, 172, 177, 167, 142, 127, 115, 139, 176, 222, 211, 157, 130, 126, 83, 5, 0, 
    15, 14, 48, 91, 127, 140, 153, 198, 221, 160, 97, 68, 134, 167, 173, 188, 198, 199, 204, 193, 175, 167, 214, 247, 222, 167, 119, 61, 0, 0, 
    43, 44, 75, 88, 128, 118, 131, 146, 192, 206, 188, 136, 161, 197, 207, 194, 182, 194, 200, 204, 209, 193, 195, 202, 227, 172, 125, 58, 0, 0, 
    77, 92, 113, 82, 84, 62, 91, 105, 138, 194, 236, 215, 178, 177, 213, 222, 225, 219, 212, 200, 192, 193, 205, 185, 145, 106, 66, 25, 13, 34, 
    110, 99, 106, 53, 37, 29, 58, 97, 107, 141, 191, 228, 218, 204, 226, 234, 247, 254, 241, 220, 195, 183, 194, 180, 120, 60, 0, 0, 15, 77, 
    109, 80, 55, 14, 13, 16, 24, 63, 81, 82, 99, 161, 228, 252, 268, 263, 252, 263, 257, 231, 205, 195, 188, 171, 121, 77, 24, 24, 33, 98, 
    78, 46, 26, 27, 18, 17, 31, 36, 46, 69, 85, 107, 202, 272, 285, 289, 267, 255, 234, 221, 200, 192, 177, 162, 113, 87, 64, 84, 107, 125, 
    50, 19, 30, 52, 26, 24, 44, 74, 67, 72, 108, 143, 189, 271, 294, 291, 281, 259, 212, 201, 193, 192, 181, 168, 127, 91, 83, 107, 133, 117, 
    78, 111, 127, 128, 71, 34, 42, 85, 107, 71, 90, 162, 211, 257, 276, 284, 265, 248, 222, 201, 194, 208, 192, 171, 131, 105, 106, 114, 110, 88, 
    163, 233, 268, 235, 154, 93, 72, 72, 89, 92, 92, 159, 214, 253, 255, 266, 257, 241, 222, 230, 223, 230, 191, 152, 108, 82, 89, 85, 91, 81, 
    160, 220, 265, 277, 224, 166, 127, 92, 69, 94, 144, 189, 218, 233, 217, 209, 217, 230, 236, 243, 243, 238, 185, 142, 100, 49, 31, 35, 77, 57, 
    63, 86, 142, 214, 251, 218, 168, 127, 96, 84, 109, 156, 177, 166, 122, 94, 122, 185, 241, 247, 238, 224, 195, 153, 102, 21, 0, 0, 44, 27, 
    1, 0, 0, 82, 172, 223, 215, 174, 135, 111, 83, 89, 112, 112, 79, 44, 83, 156, 227, 254, 232, 207, 195, 145, 58, 0, 0, 0, 27, 0, 
    0, 0, 0, 0, 50, 164, 227, 236, 186, 135, 104, 87, 87, 98, 103, 107, 123, 161, 206, 223, 230, 213, 166, 83, 4, 0, 0, 17, 53, 59, 
    4, 0, 0, 0, 0, 80, 190, 251, 256, 205, 154, 123, 100, 96, 85, 98, 121, 145, 179, 209, 206, 186, 136, 44, 0, 0, 0, 7, 69, 137, 
    0, 0, 0, 0, 0, 0, 90, 192, 252, 265, 238, 193, 151, 136, 114, 89, 72, 84, 96, 120, 105, 95, 96, 78, 66, 49, 38, 76, 130, 129, 
    0, 0, 0, 0, 0, 0, 0, 78, 163, 215, 255, 255, 223, 207, 208, 200, 135, 69, 30, 38, 36, 76, 136, 164, 178, 149, 149, 170, 186, 155, 
    
    -- channel=78
    0, 0, 0, 2, 0, 0, 2, 0, 0, 0, 32, 12, 0, 0, 20, 34, 17, 17, 29, 14, 0, 0, 63, 33, 0, 0, 44, 4, 0, 8, 
    0, 0, 0, 14, 0, 0, 4, 0, 0, 0, 45, 34, 7, 0, 39, 36, 0, 0, 26, 17, 0, 0, 81, 40, 0, 0, 15, 0, 0, 0, 
    0, 0, 0, 12, 0, 0, 8, 0, 0, 11, 41, 40, 15, 0, 28, 31, 0, 0, 11, 15, 0, 0, 83, 42, 0, 0, 5, 4, 0, 0, 
    14, 0, 0, 9, 0, 13, 16, 0, 0, 6, 20, 15, 0, 0, 8, 29, 10, 0, 19, 32, 0, 0, 82, 53, 0, 0, 12, 17, 0, 0, 
    37, 23, 21, 9, 9, 10, 20, 0, 0, 0, 0, 0, 0, 0, 0, 23, 30, 5, 1, 52, 7, 0, 80, 78, 0, 0, 0, 14, 0, 0, 
    2, 24, 33, 5, 7, 0, 5, 0, 0, 3, 0, 0, 0, 0, 0, 40, 67, 0, 0, 45, 25, 0, 75, 92, 0, 0, 0, 22, 0, 0, 
    0, 2, 14, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 21, 61, 0, 0, 25, 10, 0, 50, 90, 1, 0, 9, 36, 0, 0, 
    0, 28, 28, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 3, 0, 0, 0, 9, 0, 0, 24, 72, 18, 1, 23, 31, 0, 0, 
    0, 68, 75, 0, 0, 0, 0, 0, 18, 18, 0, 0, 0, 0, 5, 20, 0, 0, 0, 4, 0, 0, 44, 67, 12, 13, 24, 9, 0, 0, 
    0, 83, 95, 38, 0, 0, 0, 26, 50, 19, 18, 0, 0, 0, 0, 0, 0, 0, 3, 16, 0, 0, 49, 59, 3, 23, 24, 0, 0, 0, 
    0, 88, 104, 60, 14, 0, 0, 0, 11, 0, 24, 7, 0, 17, 5, 0, 0, 0, 8, 26, 0, 0, 41, 37, 0, 31, 34, 0, 0, 0, 
    0, 67, 91, 71, 59, 0, 0, 0, 0, 0, 13, 0, 17, 70, 66, 37, 18, 9, 13, 5, 0, 0, 52, 46, 0, 19, 41, 0, 0, 0, 
    0, 30, 53, 53, 73, 43, 0, 0, 2, 16, 20, 0, 0, 7, 24, 31, 32, 31, 37, 17, 11, 3, 24, 40, 4, 8, 32, 0, 0, 0, 
    0, 31, 43, 25, 64, 67, 21, 0, 0, 11, 39, 34, 13, 1, 0, 0, 0, 16, 37, 38, 54, 39, 11, 0, 0, 27, 32, 0, 0, 19, 
    0, 33, 46, 10, 37, 53, 27, 15, 0, 0, 20, 70, 39, 25, 23, 8, 0, 0, 0, 0, 27, 72, 60, 0, 0, 16, 35, 0, 0, 36, 
    0, 10, 32, 24, 29, 47, 34, 74, 54, 0, 0, 42, 39, 25, 29, 31, 29, 15, 8, 0, 0, 36, 82, 67, 0, 2, 25, 0, 0, 39, 
    0, 0, 16, 30, 46, 59, 35, 56, 99, 17, 0, 0, 52, 51, 22, 16, 25, 38, 43, 35, 21, 7, 46, 74, 45, 29, 32, 0, 0, 32, 
    21, 12, 17, 6, 37, 50, 44, 25, 57, 108, 50, 0, 30, 51, 37, 33, 12, 12, 12, 9, 32, 30, 26, 21, 30, 29, 42, 26, 0, 7, 
    29, 24, 32, 4, 9, 41, 49, 37, 17, 84, 120, 43, 16, 28, 30, 32, 38, 41, 21, 4, 27, 33, 21, 16, 0, 0, 0, 9, 24, 37, 
    19, 15, 26, 0, 0, 40, 33, 35, 34, 9, 67, 107, 65, 42, 34, 19, 36, 55, 31, 11, 32, 37, 20, 20, 0, 0, 0, 0, 22, 38, 
    0, 16, 31, 0, 0, 34, 20, 0, 28, 0, 0, 71, 96, 54, 35, 36, 28, 35, 39, 32, 35, 36, 17, 6, 0, 0, 12, 31, 12, 6, 
    0, 1, 0, 0, 0, 7, 46, 0, 0, 22, 12, 39, 79, 66, 40, 49, 40, 17, 17, 32, 26, 22, 13, 0, 0, 0, 26, 52, 13, 1, 
    0, 0, 0, 0, 0, 0, 29, 43, 0, 9, 49, 61, 54, 64, 52, 44, 50, 25, 7, 33, 25, 17, 23, 8, 0, 2, 44, 31, 6, 1, 
    42, 73, 17, 0, 0, 0, 0, 6, 7, 10, 30, 50, 44, 55, 54, 50, 61, 35, 14, 48, 30, 8, 19, 13, 0, 21, 64, 32, 12, 9, 
    96, 134, 116, 35, 0, 0, 0, 0, 0, 32, 52, 45, 49, 58, 54, 76, 103, 71, 23, 50, 48, 13, 2, 10, 0, 0, 57, 50, 17, 10, 
    37, 91, 158, 128, 44, 0, 0, 0, 0, 0, 48, 51, 52, 36, 10, 37, 100, 95, 48, 37, 40, 19, 4, 15, 0, 0, 44, 47, 4, 0, 
    0, 6, 122, 164, 119, 51, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 43, 85, 59, 40, 32, 12, 21, 17, 0, 0, 47, 22, 0, 0, 
    0, 0, 14, 119, 141, 102, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 73, 57, 57, 48, 10, 7, 0, 0, 18, 31, 18, 31, 0, 
    0, 0, 0, 18, 117, 132, 106, 62, 0, 0, 0, 0, 0, 0, 0, 0, 29, 75, 69, 71, 77, 43, 6, 0, 0, 0, 0, 14, 68, 0, 
    0, 4, 0, 0, 40, 123, 135, 106, 72, 27, 0, 0, 0, 0, 0, 0, 0, 35, 57, 63, 68, 37, 11, 0, 0, 0, 0, 0, 24, 0, 
    
    -- channel=79
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=80
    56, 8, 0, 15, 33, 26, 22, 24, 35, 34, 34, 42, 45, 50, 36, 47, 80, 85, 67, 58, 63, 67, 69, 69, 61, 47, 40, 65, 80, 67, 
    16, 0, 11, 37, 32, 17, 23, 22, 25, 30, 29, 38, 42, 39, 36, 44, 82, 99, 76, 58, 59, 57, 57, 52, 43, 46, 56, 70, 69, 62, 
    2, 0, 23, 41, 24, 6, 18, 14, 15, 25, 20, 30, 40, 30, 27, 46, 72, 104, 84, 56, 56, 62, 59, 45, 45, 53, 63, 75, 60, 48, 
    19, 12, 19, 36, 14, 3, 12, 9, 15, 15, 16, 28, 39, 37, 22, 28, 50, 79, 82, 46, 38, 60, 62, 50, 50, 56, 62, 66, 53, 44, 
    36, 14, 2, 21, 12, 9, 9, 10, 8, 14, 16, 20, 33, 44, 22, 14, 29, 44, 57, 33, 18, 55, 64, 51, 60, 61, 57, 55, 50, 47, 
    47, 3, 0, 18, 13, 10, 7, 5, 4, 11, 16, 13, 25, 41, 25, 15, 19, 23, 31, 38, 29, 58, 73, 60, 72, 71, 55, 51, 52, 48, 
    46, 0, 4, 16, 13, 10, 0, 5, 8, 12, 17, 21, 30, 38, 34, 27, 20, 20, 25, 45, 39, 49, 75, 67, 68, 67, 50, 47, 52, 48, 
    22, 0, 8, 9, 10, 11, 5, 4, 7, 14, 19, 26, 36, 35, 37, 40, 37, 24, 20, 39, 23, 32, 81, 73, 57, 48, 46, 49, 52, 50, 
    22, 7, 0, 4, 7, 10, 9, 0, 2, 9, 21, 29, 30, 15, 17, 44, 52, 31, 19, 35, 24, 38, 97, 81, 51, 51, 57, 53, 52, 52, 
    20, 0, 14, 10, 0, 6, 1, 2, 6, 7, 6, 9, 23, 4, 0, 43, 61, 36, 24, 38, 37, 70, 111, 82, 47, 62, 63, 52, 51, 48, 
    0, 0, 23, 0, 0, 0, 5, 20, 22, 0, 0, 0, 26, 40, 34, 46, 67, 39, 18, 40, 55, 96, 120, 72, 51, 63, 62, 51, 49, 51, 
    0, 0, 1, 0, 0, 7, 18, 35, 17, 0, 0, 0, 36, 44, 70, 49, 36, 32, 10, 39, 74, 106, 109, 76, 62, 60, 61, 53, 53, 58, 
    0, 0, 0, 0, 6, 6, 16, 33, 0, 0, 0, 21, 24, 14, 33, 9, 0, 3, 6, 40, 82, 104, 101, 80, 59, 49, 57, 55, 62, 65, 
    27, 14, 0, 0, 11, 12, 7, 7, 0, 0, 0, 25, 3, 0, 0, 0, 0, 0, 0, 44, 78, 95, 94, 76, 54, 29, 43, 66, 70, 68, 
    71, 16, 0, 0, 13, 29, 8, 0, 0, 0, 0, 9, 2, 0, 0, 0, 0, 0, 1, 34, 73, 104, 101, 85, 49, 6, 16, 74, 89, 66, 
    59, 13, 0, 0, 9, 42, 16, 0, 0, 5, 0, 6, 21, 0, 0, 3, 7, 4, 12, 38, 100, 133, 116, 98, 36, 0, 2, 67, 111, 77, 
    54, 10, 0, 0, 0, 47, 45, 0, 0, 45, 0, 0, 47, 35, 38, 21, 28, 50, 56, 90, 134, 134, 114, 84, 27, 0, 0, 54, 121, 95, 
    66, 23, 0, 0, 0, 51, 95, 0, 0, 38, 0, 0, 72, 37, 24, 46, 55, 96, 104, 118, 123, 98, 91, 71, 23, 0, 0, 34, 125, 118, 
    69, 26, 0, 0, 0, 45, 138, 68, 0, 7, 0, 34, 83, 4, 0, 54, 94, 118, 103, 94, 86, 63, 86, 83, 30, 0, 0, 2, 123, 137, 
    56, 21, 0, 0, 0, 56, 164, 135, 42, 33, 47, 68, 90, 24, 6, 69, 114, 130, 97, 74, 74, 62, 89, 90, 41, 0, 0, 0, 108, 144, 
    54, 41, 0, 0, 18, 79, 152, 120, 64, 75, 81, 78, 82, 52, 48, 96, 119, 123, 106, 88, 93, 76, 73, 77, 45, 2, 0, 0, 89, 147, 
    58, 48, 11, 0, 26, 74, 99, 67, 56, 76, 68, 59, 53, 50, 77, 128, 127, 115, 108, 97, 104, 94, 75, 70, 53, 35, 0, 0, 64, 139, 
    55, 27, 26, 22, 12, 30, 37, 50, 67, 62, 41, 40, 43, 54, 108, 139, 117, 107, 103, 101, 108, 104, 89, 71, 50, 54, 34, 0, 26, 109, 
    41, 13, 33, 49, 19, 0, 0, 63, 55, 29, 46, 47, 50, 70, 98, 107, 97, 94, 97, 101, 109, 99, 89, 67, 40, 75, 76, 26, 16, 62, 
    26, 22, 34, 41, 33, 15, 0, 48, 50, 29, 63, 53, 39, 56, 72, 81, 81, 83, 84, 88, 93, 79, 72, 61, 53, 88, 78, 28, 45, 50, 
    42, 43, 23, 24, 40, 56, 25, 14, 66, 67, 62, 35, 16, 43, 72, 74, 66, 65, 63, 65, 70, 52, 44, 51, 61, 68, 42, 12, 52, 71, 
    58, 61, 20, 23, 57, 67, 37, 30, 59, 58, 41, 24, 17, 41, 68, 69, 48, 49, 54, 57, 53, 31, 29, 46, 50, 42, 36, 34, 64, 60, 
    62, 54, 16, 28, 60, 59, 32, 38, 60, 28, 24, 34, 29, 39, 58, 57, 44, 55, 60, 49, 40, 25, 28, 44, 42, 40, 52, 62, 60, 22, 
    40, 23, 14, 41, 47, 39, 26, 34, 35, 13, 31, 44, 43, 49, 51, 53, 52, 64, 57, 36, 36, 31, 28, 40, 43, 44, 59, 66, 33, 10, 
    13, 12, 40, 63, 47, 37, 32, 44, 33, 24, 40, 48, 57, 68, 56, 48, 51, 53, 46, 33, 35, 33, 26, 38, 48, 44, 52, 50, 31, 25, 
    
    -- channel=81
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    7, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 24, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 24, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    54, 17, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    55, 14, 3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 8, 0, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 27, 39, 31, 16, 18, 3, 0, 0, 0, 0, 14, 49, 19, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 5, 0, 0, 0, 0, 0, 5, 32, 47, 62, 57, 62, 66, 28, 0, 0, 0, 5, 26, 51, 20, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 0, 0, 8, 12, 16, 11, 3, 34, 73, 97, 74, 58, 84, 61, 29, 18, 20, 29, 35, 29, 1, 0, 0, 0, 0, 0, 0, 
    0, 1, 24, 16, 41, 46, 29, 31, 22, 11, 42, 78, 82, 59, 39, 20, 19, 31, 26, 47, 51, 41, 35, 13, 1, 0, 0, 0, 0, 0, 
    0, 0, 15, 27, 53, 49, 47, 37, 19, 24, 53, 56, 42, 33, 51, 42, 34, 57, 51, 57, 59, 45, 31, 13, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 48, 42, 47, 46, 38, 51, 64, 31, 2, 10, 49, 78, 85, 87, 81, 83, 65, 53, 34, 19, 5, 0, 0, 0, 6, 0, 
    0, 0, 0, 29, 55, 52, 49, 44, 54, 77, 67, 44, 29, 25, 51, 72, 75, 77, 81, 81, 74, 70, 45, 27, 6, 0, 1, 26, 23, 8, 
    0, 0, 0, 20, 54, 53, 45, 38, 54, 91, 73, 52, 47, 31, 35, 64, 53, 57, 67, 83, 99, 75, 36, 16, 0, 0, 7, 49, 54, 21, 
    0, 0, 0, 38, 64, 77, 67, 47, 61, 76, 30, 18, 46, 38, 13, 30, 44, 54, 65, 72, 67, 32, 2, 0, 0, 0, 6, 52, 78, 46, 
    0, 0, 0, 54, 85, 90, 77, 40, 58, 62, 20, 41, 62, 8, 0, 0, 0, 28, 33, 24, 8, 0, 0, 0, 0, 0, 9, 66, 94, 67, 
    0, 0, 0, 42, 90, 103, 103, 42, 23, 81, 74, 60, 41, 0, 0, 27, 9, 4, 10, 4, 0, 0, 0, 0, 0, 0, 6, 71, 118, 81, 
    0, 0, 0, 40, 82, 98, 105, 41, 0, 21, 69, 65, 32, 0, 0, 43, 53, 22, 3, 10, 24, 15, 5, 0, 0, 0, 6, 66, 123, 95, 
    0, 0, 0, 27, 70, 80, 62, 6, 0, 0, 0, 0, 0, 0, 0, 16, 42, 44, 26, 14, 19, 14, 9, 1, 0, 0, 0, 50, 102, 91, 
    0, 0, 0, 13, 53, 55, 20, 0, 0, 0, 0, 0, 0, 0, 0, 30, 30, 27, 30, 22, 24, 16, 8, 9, 0, 0, 0, 14, 67, 69, 
    0, 0, 0, 0, 32, 38, 8, 0, 0, 0, 0, 0, 0, 0, 5, 8, 0, 0, 0, 9, 22, 23, 7, 0, 0, 0, 0, 0, 38, 62, 
    0, 0, 0, 1, 1, 23, 52, 41, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 6, 2, 0, 0, 2, 0, 0, 3, 61, 
    0, 0, 0, 0, 0, 0, 25, 52, 35, 30, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 6, 3, 0, 3, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=82
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=83
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=84
    130, 81, 77, 115, 133, 130, 125, 133, 135, 122, 127, 131, 127, 116, 106, 108, 96, 79, 74, 79, 79, 77, 65, 66, 60, 59, 69, 93, 77, 68, 
    117, 112, 124, 131, 132, 126, 134, 137, 136, 131, 133, 124, 126, 123, 108, 116, 105, 85, 74, 78, 81, 83, 82, 73, 64, 70, 76, 91, 87, 75, 
    125, 145, 149, 143, 129, 128, 135, 130, 143, 138, 133, 134, 132, 131, 129, 127, 115, 80, 54, 64, 75, 79, 89, 92, 95, 92, 89, 87, 82, 78, 
    131, 145, 151, 140, 125, 138, 141, 138, 147, 140, 143, 149, 139, 133, 146, 137, 129, 95, 53, 52, 63, 67, 73, 80, 94, 99, 100, 88, 75, 82, 
    136, 134, 138, 135, 130, 140, 146, 146, 145, 144, 152, 152, 141, 128, 131, 147, 148, 131, 83, 59, 73, 87, 82, 83, 90, 99, 104, 97, 87, 89, 
    150, 119, 133, 143, 139, 145, 144, 144, 149, 150, 152, 152, 153, 138, 124, 142, 145, 142, 125, 95, 108, 119, 99, 95, 93, 96, 98, 97, 96, 93, 
    126, 105, 141, 143, 144, 145, 144, 152, 152, 160, 157, 156, 155, 151, 137, 137, 142, 149, 148, 129, 117, 113, 94, 91, 95, 83, 76, 87, 92, 94, 
    102, 127, 136, 134, 139, 139, 149, 159, 156, 155, 149, 150, 143, 143, 129, 121, 128, 144, 147, 145, 121, 121, 102, 89, 91, 79, 81, 91, 91, 95, 
    133, 135, 123, 137, 140, 145, 144, 146, 149, 153, 153, 150, 133, 126, 112, 106, 106, 123, 136, 148, 128, 136, 119, 97, 87, 89, 99, 98, 98, 94, 
    139, 116, 131, 152, 152, 151, 143, 143, 152, 166, 157, 125, 101, 111, 131, 124, 108, 108, 119, 129, 120, 131, 131, 91, 80, 88, 90, 90, 97, 94, 
    88, 113, 129, 117, 121, 135, 146, 147, 150, 154, 142, 122, 114, 110, 137, 160, 140, 110, 113, 112, 110, 116, 100, 59, 77, 88, 86, 87, 90, 93, 
    51, 131, 139, 120, 136, 147, 141, 147, 142, 132, 130, 150, 146, 116, 98, 103, 101, 83, 98, 105, 105, 106, 73, 54, 67, 80, 84, 84, 87, 93, 
    38, 137, 147, 146, 154, 149, 142, 138, 117, 116, 134, 161, 151, 136, 100, 52, 69, 78, 81, 99, 100, 88, 64, 49, 51, 67, 74, 76, 85, 88, 
    69, 118, 124, 146, 144, 138, 150, 137, 111, 130, 145, 135, 123, 129, 130, 86, 109, 113, 102, 116, 91, 74, 58, 45, 54, 69, 70, 66, 77, 82, 
    91, 78, 109, 146, 148, 135, 145, 141, 131, 142, 153, 142, 130, 140, 147, 132, 140, 134, 141, 123, 92, 86, 66, 63, 65, 70, 87, 72, 66, 76, 
    100, 73, 94, 135, 145, 127, 119, 140, 136, 153, 176, 172, 142, 140, 162, 164, 147, 143, 152, 143, 139, 109, 79, 65, 56, 73, 105, 99, 65, 64, 
    109, 98, 109, 131, 134, 130, 110, 136, 150, 156, 143, 141, 132, 147, 160, 160, 156, 144, 149, 156, 152, 101, 63, 40, 37, 73, 100, 113, 70, 51, 
    116, 115, 126, 139, 133, 133, 94, 113, 177, 133, 100, 140, 151, 135, 104, 87, 116, 122, 117, 111, 94, 55, 32, 31, 37, 71, 105, 114, 76, 44, 
    120, 90, 106, 139, 137, 137, 102, 71, 163, 152, 133, 162, 156, 116, 137, 105, 101, 97, 82, 66, 41, 36, 45, 42, 56, 77, 113, 121, 93, 37, 
    117, 92, 115, 139, 139, 143, 135, 48, 77, 132, 154, 169, 141, 110, 169, 165, 132, 93, 58, 58, 52, 64, 72, 47, 48, 71, 116, 139, 118, 48, 
    121, 113, 119, 136, 141, 136, 138, 50, 6, 46, 79, 106, 106, 90, 111, 138, 135, 99, 57, 57, 56, 64, 82, 60, 48, 66, 120, 150, 142, 71, 
    136, 115, 102, 128, 137, 128, 106, 43, 38, 44, 33, 35, 55, 52, 74, 101, 94, 84, 58, 48, 39, 36, 63, 74, 77, 72, 101, 146, 155, 84, 
    142, 118, 101, 115, 138, 127, 78, 63, 98, 80, 58, 54, 60, 71, 91, 67, 35, 34, 31, 30, 30, 21, 27, 56, 66, 66, 78, 132, 159, 107, 
    113, 114, 127, 116, 123, 133, 126, 117, 91, 70, 74, 93, 93, 95, 85, 52, 25, 15, 17, 20, 24, 19, 19, 28, 40, 71, 74, 92, 139, 142, 
    107, 121, 138, 117, 91, 111, 159, 154, 97, 119, 123, 115, 102, 92, 85, 72, 46, 33, 25, 18, 12, 12, 16, 8, 36, 78, 59, 52, 70, 114, 
    117, 126, 136, 130, 109, 103, 117, 149, 115, 120, 119, 101, 106, 115, 103, 94, 77, 61, 43, 38, 36, 28, 28, 25, 42, 56, 41, 56, 65, 78, 
    112, 118, 121, 131, 135, 126, 93, 119, 130, 107, 90, 82, 111, 128, 117, 100, 88, 80, 76, 77, 70, 60, 66, 70, 64, 60, 59, 77, 119, 80, 
    131, 106, 90, 122, 129, 118, 95, 95, 111, 89, 97, 100, 115, 126, 127, 105, 97, 103, 105, 96, 88, 89, 101, 99, 92, 89, 87, 93, 105, 76, 
    122, 96, 94, 124, 122, 109, 106, 116, 101, 94, 116, 114, 117, 125, 135, 122, 115, 113, 99, 99, 105, 108, 117, 114, 109, 105, 106, 98, 83, 88, 
    113, 108, 125, 127, 132, 132, 123, 126, 121, 128, 139, 128, 120, 115, 121, 124, 118, 107, 95, 104, 111, 113, 118, 122, 115, 117, 115, 96, 88, 99, 
    
    -- channel=85
    39, 12, 0, 0, 14, 22, 4, 5, 13, 11, 4, 18, 17, 11, 8, 6, 19, 17, 12, 8, 8, 9, 0, 2, 11, 4, 0, 8, 19, 8, 
    30, 0, 0, 1, 17, 11, 6, 19, 11, 11, 9, 7, 12, 15, 9, 7, 12, 15, 17, 11, 13, 13, 11, 11, 0, 0, 0, 11, 16, 10, 
    9, 2, 10, 12, 19, 1, 8, 14, 6, 15, 14, 8, 12, 15, 2, 12, 11, 10, 8, 4, 7, 8, 17, 15, 8, 10, 4, 10, 19, 9, 
    0, 14, 14, 20, 14, 3, 10, 5, 12, 13, 6, 14, 13, 12, 21, 14, 15, 5, 0, 0, 0, 0, 4, 9, 11, 14, 15, 13, 5, 2, 
    0, 23, 7, 11, 7, 4, 11, 12, 8, 6, 12, 17, 10, 9, 19, 14, 20, 16, 4, 1, 0, 0, 9, 0, 6, 13, 19, 17, 5, 6, 
    23, 24, 0, 15, 9, 6, 14, 7, 9, 8, 17, 13, 14, 14, 6, 7, 17, 21, 16, 0, 1, 10, 15, 10, 8, 15, 17, 12, 13, 10, 
    45, 0, 1, 17, 10, 16, 10, 5, 10, 15, 18, 10, 18, 20, 14, 10, 11, 11, 19, 6, 15, 8, 8, 9, 8, 14, 6, 3, 9, 8, 
    14, 0, 13, 8, 10, 7, 11, 12, 9, 14, 15, 6, 9, 14, 11, 1, 11, 17, 22, 18, 22, 0, 3, 8, 17, 10, 0, 4, 5, 9, 
    12, 20, 5, 6, 9, 3, 9, 10, 16, 13, 8, 9, 9, 11, 0, 0, 1, 14, 13, 15, 18, 7, 13, 23, 11, 5, 10, 14, 7, 12, 
    51, 8, 0, 21, 13, 16, 8, 2, 8, 14, 13, 2, 0, 8, 0, 0, 3, 7, 2, 11, 9, 9, 27, 37, 2, 5, 14, 12, 13, 11, 
    33, 0, 0, 14, 0, 1, 3, 0, 15, 21, 14, 0, 0, 6, 20, 35, 30, 17, 0, 1, 0, 1, 37, 23, 4, 11, 9, 8, 7, 9, 
    0, 0, 28, 0, 0, 1, 5, 7, 24, 9, 0, 0, 22, 0, 0, 33, 22, 7, 1, 0, 7, 21, 23, 3, 6, 12, 11, 10, 5, 9, 
    0, 0, 30, 0, 8, 18, 3, 12, 19, 0, 0, 9, 41, 31, 0, 0, 0, 0, 0, 0, 11, 17, 17, 8, 2, 4, 5, 3, 5, 12, 
    0, 18, 14, 0, 7, 15, 16, 22, 0, 0, 0, 10, 19, 14, 17, 0, 0, 4, 0, 0, 14, 7, 16, 3, 2, 5, 0, 0, 4, 11, 
    5, 17, 0, 0, 9, 6, 24, 18, 0, 0, 15, 8, 3, 0, 2, 0, 10, 10, 5, 20, 3, 12, 16, 7, 16, 9, 0, 0, 4, 11, 
    12, 0, 0, 0, 11, 5, 17, 10, 0, 0, 27, 19, 11, 8, 8, 19, 15, 14, 27, 23, 15, 36, 22, 23, 20, 0, 4, 0, 5, 11, 
    19, 9, 0, 0, 7, 0, 13, 14, 0, 9, 36, 12, 8, 10, 21, 32, 21, 20, 20, 24, 46, 51, 29, 16, 2, 0, 0, 5, 7, 8, 
    7, 22, 10, 0, 0, 0, 5, 20, 0, 38, 5, 0, 1, 36, 0, 0, 5, 18, 25, 26, 42, 35, 8, 5, 0, 0, 0, 1, 0, 15, 
    10, 18, 0, 0, 6, 13, 0, 21, 36, 35, 0, 0, 44, 52, 0, 0, 0, 18, 31, 23, 22, 2, 0, 7, 1, 0, 0, 0, 0, 18, 
    21, 5, 0, 0, 5, 19, 21, 11, 10, 32, 35, 33, 43, 20, 23, 39, 26, 22, 26, 13, 7, 2, 2, 7, 4, 2, 0, 2, 11, 22, 
    6, 10, 10, 0, 4, 16, 47, 35, 0, 0, 20, 38, 31, 10, 4, 35, 55, 31, 10, 1, 10, 21, 20, 14, 0, 0, 0, 7, 20, 31, 
    14, 20, 2, 1, 11, 16, 46, 26, 0, 0, 0, 0, 11, 9, 0, 12, 39, 34, 21, 6, 3, 8, 19, 15, 6, 0, 3, 8, 27, 30, 
    36, 21, 0, 5, 16, 28, 18, 0, 6, 26, 6, 0, 0, 0, 0, 24, 12, 10, 13, 10, 6, 1, 0, 7, 17, 0, 0, 15, 31, 22, 
    30, 13, 2, 7, 28, 31, 2, 0, 19, 0, 0, 1, 0, 4, 23, 16, 4, 0, 0, 0, 8, 10, 0, 9, 0, 0, 5, 9, 27, 35, 
    7, 0, 16, 9, 0, 4, 34, 38, 24, 0, 2, 18, 14, 8, 12, 9, 5, 0, 0, 0, 0, 0, 0, 0, 0, 2, 21, 0, 0, 35, 
    10, 12, 24, 17, 0, 0, 26, 21, 4, 20, 32, 29, 7, 5, 13, 18, 12, 5, 3, 0, 0, 0, 0, 0, 0, 13, 11, 0, 0, 3, 
    1, 17, 24, 8, 22, 20, 2, 12, 17, 25, 8, 3, 0, 17, 15, 21, 15, 7, 2, 8, 13, 5, 0, 0, 3, 0, 0, 0, 10, 21, 
    10, 24, 6, 0, 18, 30, 10, 0, 24, 28, 0, 1, 5, 15, 20, 19, 6, 4, 17, 19, 11, 2, 0, 10, 8, 3, 0, 0, 31, 24, 
    23, 21, 0, 6, 22, 13, 10, 7, 12, 0, 0, 16, 11, 16, 23, 17, 8, 15, 23, 11, 6, 6, 9, 7, 10, 8, 7, 20, 10, 0, 
    9, 0, 0, 20, 22, 17, 10, 17, 21, 8, 12, 16, 6, 11, 24, 19, 20, 17, 8, 6, 7, 8, 11, 9, 14, 10, 16, 13, 1, 0, 
    
    -- channel=86
    13, 16, 10, 23, 32, 32, 33, 31, 36, 32, 37, 39, 43, 44, 39, 40, 32, 35, 39, 41, 36, 31, 31, 26, 24, 22, 26, 30, 30, 30, 
    10, 15, 18, 26, 31, 35, 30, 29, 34, 30, 34, 35, 33, 38, 36, 37, 45, 41, 44, 46, 40, 36, 33, 26, 23, 22, 26, 29, 36, 31, 
    19, 20, 29, 30, 31, 34, 26, 26, 31, 30, 28, 32, 36, 37, 44, 38, 38, 35, 29, 38, 40, 38, 36, 40, 38, 31, 32, 30, 28, 30, 
    18, 18, 35, 24, 26, 32, 29, 30, 28, 29, 33, 34, 38, 39, 40, 44, 31, 30, 19, 17, 25, 22, 21, 29, 31, 34, 33, 30, 26, 26, 
    14, 19, 28, 19, 23, 27, 30, 30, 26, 28, 30, 34, 33, 33, 32, 40, 41, 35, 22, 7, 15, 26, 24, 33, 34, 37, 39, 36, 31, 27, 
    15, 28, 20, 23, 27, 28, 27, 25, 25, 29, 27, 33, 33, 35, 32, 34, 36, 33, 30, 29, 28, 43, 35, 36, 41, 40, 43, 39, 33, 31, 
    14, 20, 21, 28, 29, 27, 27, 30, 28, 31, 37, 38, 33, 39, 40, 38, 39, 42, 37, 38, 22, 29, 25, 31, 39, 34, 28, 28, 30, 29, 
    18, 22, 24, 21, 22, 27, 28, 36, 33, 27, 25, 29, 28, 29, 29, 27, 30, 40, 40, 36, 24, 29, 24, 26, 34, 31, 30, 28, 31, 29, 
    33, 34, 18, 17, 24, 25, 26, 23, 23, 27, 29, 25, 18, 8, 9, 5, 15, 27, 39, 38, 32, 33, 36, 32, 44, 37, 39, 38, 36, 30, 
    49, 42, 21, 32, 37, 24, 22, 26, 29, 38, 26, 3, 0, 0, 12, 10, 11, 20, 29, 26, 31, 39, 48, 46, 43, 37, 36, 36, 35, 33, 
    44, 36, 7, 3, 0, 5, 18, 27, 25, 29, 13, 0, 0, 3, 21, 41, 48, 28, 27, 20, 21, 36, 34, 37, 39, 44, 42, 37, 36, 32, 
    28, 29, 12, 10, 3, 8, 14, 17, 20, 19, 8, 11, 7, 14, 11, 0, 17, 5, 4, 15, 13, 29, 35, 39, 38, 42, 41, 38, 36, 36, 
    14, 26, 34, 23, 6, 8, 16, 7, 1, 4, 7, 15, 17, 12, 0, 0, 0, 0, 0, 0, 10, 23, 26, 31, 29, 33, 34, 33, 36, 35, 
    26, 27, 30, 16, 4, 4, 12, 9, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 8, 18, 27, 28, 30, 27, 18, 25, 36, 
    23, 17, 23, 19, 9, 14, 12, 16, 2, 0, 0, 2, 3, 12, 7, 0, 0, 0, 0, 0, 0, 8, 31, 39, 38, 30, 21, 17, 11, 32, 
    25, 15, 7, 8, 3, 7, 3, 14, 11, 2, 20, 25, 10, 13, 25, 23, 17, 11, 15, 23, 35, 41, 53, 49, 40, 37, 21, 21, 12, 22, 
    22, 19, 18, 3, 0, 5, 10, 17, 38, 5, 10, 5, 5, 28, 50, 39, 49, 39, 48, 63, 66, 63, 52, 38, 33, 29, 22, 8, 10, 15, 
    31, 28, 28, 9, 0, 0, 7, 13, 52, 6, 0, 13, 19, 12, 19, 0, 20, 44, 48, 55, 46, 40, 33, 25, 33, 25, 22, 2, 0, 6, 
    25, 14, 11, 6, 0, 0, 18, 21, 55, 59, 29, 30, 25, 17, 29, 15, 11, 33, 42, 39, 21, 23, 33, 32, 40, 33, 19, 2, 0, 0, 
    15, 15, 21, 18, 2, 3, 32, 42, 48, 65, 73, 66, 54, 47, 53, 52, 45, 42, 36, 45, 42, 41, 44, 34, 28, 26, 26, 10, 0, 0, 
    20, 21, 25, 25, 14, 15, 27, 33, 28, 24, 43, 52, 56, 48, 46, 44, 55, 63, 50, 49, 50, 46, 51, 43, 32, 29, 33, 30, 10, 3, 
    24, 23, 20, 20, 19, 14, 8, 8, 12, 23, 23, 15, 13, 20, 33, 50, 61, 64, 60, 53, 50, 45, 49, 57, 52, 47, 33, 40, 27, 10, 
    29, 29, 18, 13, 21, 9, 0, 3, 17, 31, 19, 21, 18, 30, 38, 37, 37, 39, 42, 45, 46, 46, 45, 46, 47, 43, 38, 47, 44, 24, 
    21, 19, 26, 25, 18, 21, 20, 12, 0, 8, 3, 18, 33, 28, 22, 25, 22, 26, 30, 37, 39, 41, 45, 35, 37, 46, 47, 52, 47, 44, 
    25, 26, 21, 20, 12, 17, 27, 37, 12, 30, 44, 27, 24, 15, 15, 23, 21, 22, 22, 22, 21, 23, 27, 23, 31, 44, 36, 31, 24, 20, 
    26, 25, 29, 26, 18, 25, 17, 36, 37, 19, 37, 27, 24, 21, 23, 23, 26, 19, 13, 15, 18, 16, 15, 15, 18, 19, 17, 16, 30, 19, 
    24, 23, 30, 32, 24, 32, 32, 25, 35, 31, 22, 13, 21, 22, 27, 22, 20, 18, 21, 25, 22, 18, 19, 16, 16, 17, 21, 28, 39, 34, 
    39, 21, 16, 18, 25, 20, 19, 23, 8, 12, 20, 20, 24, 23, 26, 24, 25, 31, 31, 31, 24, 23, 24, 20, 20, 23, 28, 33, 25, 17, 
    23, 11, 12, 11, 19, 19, 16, 19, 14, 12, 14, 21, 29, 31, 35, 40, 36, 33, 26, 26, 29, 27, 25, 24, 20, 24, 26, 25, 24, 24, 
    18, 15, 21, 25, 34, 40, 32, 26, 26, 36, 33, 32, 33, 34, 35, 43, 36, 29, 24, 24, 27, 24, 23, 24, 22, 24, 25, 20, 19, 21, 
    
    -- channel=87
    73, 78, 69, 49, 49, 48, 44, 49, 45, 50, 43, 41, 39, 39, 48, 38, 33, 34, 37, 30, 30, 32, 35, 38, 41, 39, 35, 22, 28, 31, 
    83, 75, 64, 54, 58, 52, 46, 55, 48, 52, 49, 45, 42, 44, 41, 36, 26, 29, 37, 30, 28, 30, 31, 37, 36, 33, 28, 24, 31, 33, 
    75, 69, 63, 58, 64, 56, 53, 59, 52, 55, 53, 46, 43, 45, 40, 37, 36, 35, 44, 37, 30, 25, 26, 28, 24, 27, 25, 26, 36, 33, 
    66, 75, 65, 64, 68, 58, 57, 60, 56, 57, 54, 50, 46, 45, 47, 43, 46, 44, 47, 50, 40, 29, 33, 28, 24, 25, 27, 31, 37, 34, 
    63, 82, 68, 69, 67, 60, 63, 62, 64, 58, 59, 57, 51, 48, 54, 47, 52, 50, 49, 52, 42, 23, 29, 24, 17, 21, 26, 29, 33, 33, 
    70, 80, 68, 67, 64, 62, 66, 64, 66, 57, 59, 56, 49, 46, 56, 53, 58, 52, 48, 39, 39, 23, 29, 26, 15, 21, 27, 27, 30, 32, 
    78, 76, 65, 66, 65, 63, 66, 61, 62, 53, 56, 49, 46, 42, 49, 49, 51, 46, 48, 39, 55, 41, 41, 36, 25, 31, 34, 32, 31, 32, 
    74, 67, 68, 68, 67, 62, 65, 62, 63, 58, 59, 53, 50, 52, 53, 49, 46, 44, 45, 38, 62, 47, 41, 44, 35, 35, 31, 32, 30, 32, 
    64, 64, 68, 67, 65, 65, 71, 71, 66, 61, 61, 62, 62, 71, 63, 52, 47, 46, 43, 38, 57, 44, 34, 48, 35, 29, 28, 32, 30, 33, 
    67, 56, 53, 62, 63, 67, 73, 65, 63, 70, 87, 88, 74, 78, 63, 50, 49, 55, 46, 41, 47, 28, 30, 48, 36, 30, 33, 35, 32, 32, 
    85, 54, 70, 85, 79, 78, 73, 62, 71, 91, 107, 89, 66, 56, 43, 41, 38, 58, 52, 42, 41, 26, 35, 47, 33, 30, 33, 35, 32, 30, 
    81, 49, 77, 79, 73, 75, 70, 61, 83, 99, 100, 74, 63, 61, 48, 71, 62, 70, 67, 43, 37, 25, 32, 36, 32, 34, 34, 36, 29, 27, 
    56, 51, 77, 72, 70, 77, 68, 70, 97, 93, 78, 64, 69, 73, 68, 91, 76, 85, 74, 51, 43, 29, 35, 35, 38, 41, 36, 38, 27, 26, 
    33, 56, 78, 70, 71, 72, 72, 79, 98, 89, 80, 73, 83, 84, 75, 85, 75, 84, 73, 59, 50, 37, 38, 33, 41, 51, 42, 38, 31, 28, 
    27, 60, 69, 61, 64, 60, 75, 86, 96, 85, 84, 68, 74, 80, 71, 75, 74, 81, 73, 68, 45, 35, 29, 28, 46, 56, 51, 34, 34, 34, 
    31, 58, 66, 65, 70, 56, 80, 95, 77, 67, 75, 60, 65, 66, 59, 64, 63, 65, 57, 45, 18, 22, 21, 27, 52, 56, 54, 33, 31, 37, 
    24, 52, 62, 66, 74, 48, 67, 99, 55, 68, 91, 63, 44, 52, 36, 56, 41, 37, 33, 17, 10, 24, 24, 37, 54, 62, 60, 43, 29, 41, 
    14, 48, 63, 71, 78, 53, 45, 97, 55, 73, 91, 47, 34, 76, 56, 61, 39, 25, 30, 22, 30, 36, 27, 38, 48, 63, 68, 55, 27, 42, 
    22, 56, 71, 74, 75, 52, 17, 65, 48, 52, 62, 36, 32, 70, 40, 33, 21, 17, 33, 29, 36, 32, 13, 26, 39, 62, 74, 68, 27, 46, 
    26, 46, 62, 67, 64, 41, 3, 44, 35, 30, 34, 23, 19, 38, 14, 5, 8, 10, 29, 22, 22, 24, 11, 28, 40, 63, 75, 70, 28, 42, 
    21, 35, 54, 60, 54, 34, 18, 51, 39, 33, 35, 28, 20, 31, 14, 4, 14, 14, 26, 24, 22, 27, 20, 27, 36, 48, 67, 64, 30, 37, 
    23, 33, 45, 55, 50, 45, 48, 51, 32, 32, 39, 39, 39, 32, 9, 6, 21, 22, 28, 29, 24, 28, 25, 22, 30, 33, 56, 60, 34, 31, 
    28, 34, 32, 46, 59, 66, 65, 37, 32, 28, 31, 24, 25, 16, 7, 21, 36, 32, 33, 28, 25, 29, 30, 34, 39, 24, 40, 50, 41, 32, 
    36, 30, 23, 32, 55, 65, 60, 40, 68, 47, 31, 24, 21, 16, 20, 28, 34, 29, 29, 24, 23, 30, 31, 42, 39, 13, 30, 38, 41, 36, 
    34, 27, 31, 38, 49, 49, 61, 41, 59, 37, 21, 32, 30, 24, 25, 27, 31, 29, 35, 32, 32, 40, 39, 43, 32, 19, 41, 52, 36, 42, 
    25, 26, 37, 32, 37, 34, 58, 52, 42, 46, 36, 43, 29, 21, 19, 27, 33, 34, 39, 35, 35, 45, 42, 41, 37, 37, 48, 48, 22, 38, 
    18, 26, 39, 23, 23, 27, 47, 36, 33, 48, 38, 43, 28, 21, 18, 29, 35, 31, 28, 27, 31, 42, 35, 35, 38, 40, 37, 30, 19, 43, 
    12, 33, 36, 23, 25, 31, 45, 33, 37, 49, 28, 31, 26, 24, 19, 27, 27, 18, 20, 23, 28, 37, 32, 32, 37, 36, 29, 30, 38, 51, 
    29, 41, 28, 23, 27, 30, 34, 30, 41, 41, 24, 28, 24, 21, 22, 21, 24, 20, 25, 27, 27, 34, 34, 30, 35, 32, 28, 33, 44, 38, 
    35, 34, 18, 17, 20, 21, 25, 22, 34, 28, 21, 27, 24, 23, 28, 25, 29, 27, 30, 30, 30, 36, 37, 29, 31, 30, 31, 37, 41, 32, 
    
    -- channel=88
    280, 283, 297, 321, 328, 329, 334, 338, 345, 341, 347, 343, 328, 309, 298, 278, 237, 204, 196, 199, 197, 196, 192, 191, 196, 201, 208, 198, 177, 173, 
    305, 323, 332, 339, 338, 343, 342, 346, 357, 349, 353, 352, 348, 333, 326, 305, 266, 224, 202, 201, 200, 203, 195, 192, 198, 205, 215, 209, 194, 190, 
    327, 341, 345, 339, 343, 353, 351, 359, 365, 360, 366, 362, 359, 355, 348, 336, 294, 234, 198, 196, 202, 214, 214, 218, 221, 221, 218, 212, 210, 206, 
    330, 333, 348, 342, 349, 365, 363, 366, 373, 371, 377, 376, 371, 368, 371, 360, 322, 252, 199, 196, 208, 214, 216, 233, 237, 237, 229, 215, 217, 218, 
    304, 314, 342, 336, 352, 370, 372, 373, 374, 381, 386, 389, 374, 364, 381, 382, 354, 297, 236, 229, 239, 232, 220, 229, 235, 239, 238, 228, 221, 224, 
    280, 313, 334, 340, 354, 363, 374, 376, 377, 382, 389, 397, 376, 360, 369, 380, 370, 345, 299, 283, 287, 276, 250, 242, 233, 233, 241, 239, 231, 231, 
    279, 312, 328, 346, 357, 365, 372, 376, 383, 391, 393, 398, 378, 364, 357, 360, 357, 359, 349, 328, 318, 307, 265, 246, 228, 224, 235, 235, 234, 234, 
    274, 302, 325, 342, 356, 369, 378, 383, 384, 395, 390, 377, 354, 346, 339, 333, 335, 348, 357, 340, 322, 303, 258, 232, 227, 222, 225, 228, 232, 232, 
    270, 306, 322, 335, 356, 365, 375, 388, 391, 394, 370, 341, 307, 299, 298, 287, 295, 323, 343, 334, 327, 306, 250, 219, 229, 231, 231, 232, 230, 232, 
    278, 321, 320, 335, 360, 369, 370, 384, 389, 393, 349, 304, 261, 256, 266, 256, 262, 290, 312, 308, 306, 289, 229, 210, 221, 226, 231, 234, 234, 232, 
    276, 318, 304, 333, 355, 356, 360, 366, 365, 377, 336, 282, 225, 239, 266, 246, 249, 261, 272, 267, 261, 237, 199, 192, 203, 216, 222, 228, 231, 233, 
    266, 307, 298, 322, 326, 331, 340, 334, 332, 353, 331, 290, 237, 220, 233, 236, 245, 244, 249, 242, 222, 196, 161, 165, 187, 212, 220, 227, 226, 227, 
    251, 295, 320, 335, 320, 314, 311, 299, 309, 328, 317, 303, 281, 252, 201, 188, 216, 210, 230, 222, 196, 177, 145, 147, 168, 200, 217, 222, 218, 217, 
    224, 272, 317, 326, 308, 309, 302, 289, 299, 311, 300, 304, 312, 301, 248, 207, 216, 221, 222, 207, 189, 161, 138, 139, 159, 196, 213, 212, 203, 204, 
    224, 252, 300, 314, 298, 295, 300, 302, 302, 308, 300, 301, 313, 318, 293, 257, 254, 254, 243, 219, 191, 156, 142, 140, 164, 212, 216, 199, 185, 190, 
    230, 244, 288, 304, 293, 283, 287, 309, 317, 300, 306, 314, 312, 326, 315, 287, 279, 278, 274, 247, 202, 160, 146, 144, 176, 226, 237, 197, 164, 175, 
    258, 253, 277, 288, 280, 261, 262, 301, 308, 277, 310, 321, 296, 299, 324, 308, 294, 277, 272, 254, 205, 161, 145, 138, 179, 230, 249, 209, 151, 147, 
    269, 273, 294, 280, 262, 241, 234, 279, 287, 255, 291, 303, 266, 270, 295, 288, 283, 251, 228, 204, 171, 151, 138, 132, 176, 233, 252, 212, 141, 120, 
    261, 272, 299, 283, 254, 223, 187, 232, 277, 256, 276, 287, 253, 267, 275, 237, 238, 211, 176, 152, 134, 141, 140, 141, 184, 238, 269, 223, 133, 102, 
    262, 261, 285, 283, 257, 228, 163, 160, 242, 265, 259, 256, 244, 278, 314, 263, 217, 187, 162, 147, 134, 148, 152, 149, 196, 245, 278, 245, 146, 95, 
    269, 266, 287, 286, 259, 231, 168, 133, 162, 198, 217, 221, 217, 244, 293, 274, 223, 178, 154, 154, 149, 159, 163, 157, 187, 239, 279, 269, 182, 117, 
    266, 262, 279, 281, 259, 220, 187, 176, 150, 137, 155, 179, 193, 216, 226, 208, 194, 165, 136, 127, 123, 138, 165, 172, 187, 225, 270, 283, 218, 146, 
    272, 266, 268, 273, 257, 231, 222, 223, 209, 194, 180, 184, 201, 209, 187, 155, 136, 127, 115, 105, 92, 97, 130, 159, 188, 212, 240, 284, 250, 172, 
    287, 292, 271, 265, 274, 268, 254, 241, 240, 245, 231, 226, 230, 227, 190, 145, 114, 102, 99, 95, 89, 87, 100, 132, 172, 187, 198, 259, 265, 202, 
    282, 292, 283, 261, 267, 297, 296, 271, 257, 256, 241, 244, 248, 236, 206, 172, 141, 122, 110, 102, 95, 99, 109, 134, 164, 172, 176, 212, 247, 229, 
    285, 282, 282, 274, 250, 262, 296, 287, 260, 262, 256, 252, 258, 250, 236, 213, 186, 163, 149, 136, 128, 135, 147, 152, 166, 176, 180, 196, 191, 202, 
    266, 257, 279, 290, 267, 246, 258, 283, 240, 229, 249, 258, 274, 271, 254, 238, 224, 205, 190, 189, 190, 199, 203, 195, 195, 202, 215, 230, 204, 189, 
    252, 238, 270, 280, 268, 261, 253, 255, 245, 245, 253, 261, 282, 282, 266, 254, 250, 236, 226, 235, 241, 253, 255, 247, 241, 242, 244, 238, 235, 225, 
    269, 256, 267, 270, 266, 264, 267, 255, 244, 264, 277, 281, 293, 288, 278, 273, 266, 255, 251, 262, 269, 280, 281, 273, 264, 262, 252, 239, 239, 250, 
    283, 283, 279, 269, 269, 272, 277, 280, 272, 284, 287, 287, 288, 279, 278, 280, 273, 263, 256, 269, 280, 287, 291, 282, 272, 268, 260, 249, 252, 263, 
    
    -- channel=89
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=90
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=91
    71, 67, 92, 99, 87, 82, 92, 94, 83, 82, 76, 69, 53, 45, 56, 57, 37, 9, 0, 3, 7, 2, 5, 0, 3, 16, 38, 26, 12, 1, 
    125, 131, 130, 112, 95, 101, 102, 102, 97, 90, 76, 75, 62, 48, 58, 51, 29, 2, 0, 0, 7, 9, 3, 2, 15, 27, 40, 30, 13, 12, 
    164, 159, 143, 110, 99, 107, 105, 115, 107, 102, 96, 84, 71, 64, 60, 57, 29, 0, 0, 0, 8, 19, 19, 24, 33, 37, 33, 23, 17, 21, 
    173, 160, 144, 120, 116, 116, 116, 124, 120, 120, 116, 100, 88, 84, 66, 69, 48, 13, 0, 0, 9, 19, 21, 32, 40, 42, 31, 21, 30, 35, 
    160, 144, 145, 132, 128, 130, 130, 133, 134, 135, 124, 110, 98, 88, 87, 90, 84, 50, 24, 24, 33, 25, 17, 19, 31, 34, 30, 30, 36, 41, 
    135, 143, 153, 141, 135, 131, 137, 146, 144, 136, 130, 122, 105, 89, 94, 101, 111, 97, 70, 67, 62, 43, 34, 23, 22, 19, 25, 36, 41, 48, 
    134, 153, 149, 147, 139, 136, 144, 150, 152, 134, 132, 128, 118, 99, 93, 99, 109, 110, 101, 86, 77, 66, 50, 28, 8, 8, 26, 37, 44, 50, 
    144, 137, 143, 147, 142, 147, 150, 147, 145, 137, 141, 128, 120, 105, 104, 107, 105, 99, 104, 89, 90, 84, 62, 30, 11, 19, 30, 36, 44, 46, 
    119, 124, 149, 147, 148, 143, 147, 151, 151, 145, 146, 131, 124, 120, 125, 116, 98, 89, 103, 101, 118, 111, 71, 26, 25, 36, 35, 39, 41, 46, 
    79, 132, 150, 140, 145, 148, 152, 156, 158, 151, 156, 164, 169, 167, 155, 134, 100, 84, 98, 105, 121, 110, 47, 15, 25, 30, 31, 37, 39, 46, 
    67, 135, 140, 151, 171, 176, 172, 162, 150, 158, 192, 211, 193, 192, 174, 124, 89, 86, 95, 106, 106, 71, 19, 10, 12, 14, 19, 24, 37, 45, 
    78, 132, 142, 171, 188, 186, 184, 154, 139, 179, 243, 238, 186, 154, 138, 113, 101, 114, 118, 117, 94, 36, 0, 0, 1, 10, 15, 21, 32, 36, 
    95, 130, 171, 207, 210, 195, 179, 149, 159, 209, 247, 213, 169, 136, 100, 114, 130, 140, 155, 136, 89, 34, 0, 0, 0, 3, 16, 23, 25, 26, 
    67, 96, 167, 207, 210, 203, 176, 160, 197, 227, 220, 191, 175, 182, 165, 185, 186, 188, 189, 144, 99, 41, 0, 0, 0, 5, 28, 36, 20, 15, 
    43, 79, 150, 199, 199, 191, 177, 187, 229, 248, 222, 190, 184, 206, 223, 235, 229, 231, 207, 171, 127, 53, 10, 0, 0, 31, 53, 52, 27, 8, 
    39, 76, 151, 199, 197, 179, 177, 198, 255, 253, 219, 197, 201, 217, 219, 213, 219, 222, 209, 186, 114, 39, 0, 0, 0, 53, 90, 71, 35, 10, 
    66, 85, 144, 196, 206, 173, 165, 190, 235, 210, 201, 210, 201, 175, 171, 174, 173, 175, 165, 135, 53, 0, 0, 0, 0, 60, 120, 99, 47, 8, 
    79, 95, 152, 206, 224, 180, 158, 174, 170, 171, 202, 202, 154, 116, 128, 157, 133, 102, 75, 37, 0, 0, 0, 0, 0, 66, 129, 131, 70, 8, 
    64, 96, 167, 220, 234, 186, 119, 127, 122, 153, 197, 179, 112, 112, 106, 114, 83, 29, 0, 0, 0, 0, 0, 0, 0, 69, 151, 169, 92, 15, 
    74, 97, 156, 217, 235, 191, 66, 30, 75, 119, 138, 112, 81, 122, 130, 103, 46, 0, 0, 0, 0, 0, 0, 0, 0, 75, 168, 200, 116, 25, 
    99, 101, 147, 199, 208, 164, 28, 0, 0, 37, 56, 43, 25, 56, 99, 85, 25, 0, 0, 0, 0, 0, 0, 0, 0, 73, 157, 206, 136, 39, 
    92, 86, 133, 171, 170, 117, 28, 0, 0, 0, 0, 0, 0, 24, 41, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 126, 177, 132, 50, 
    78, 81, 120, 149, 138, 106, 90, 71, 9, 0, 0, 0, 6, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 78, 126, 114, 51, 
    85, 102, 105, 120, 133, 139, 135, 95, 57, 52, 52, 32, 33, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 75, 102, 54, 
    88, 106, 101, 100, 133, 165, 149, 114, 112, 80, 58, 43, 49, 45, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 93, 81, 
    97, 99, 100, 104, 108, 114, 139, 129, 130, 98, 63, 59, 73, 68, 51, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 46, 55, 
    95, 84, 102, 122, 106, 66, 93, 114, 79, 54, 58, 81, 91, 84, 64, 41, 33, 31, 20, 3, 0, 2, 13, 8, 2, 4, 26, 60, 19, 14, 
    66, 60, 100, 110, 93, 68, 75, 91, 68, 69, 70, 80, 89, 88, 68, 57, 59, 52, 32, 25, 31, 47, 54, 51, 45, 44, 47, 47, 26, 42, 
    65, 76, 101, 95, 80, 76, 87, 76, 74, 95, 92, 89, 89, 86, 72, 66, 62, 46, 40, 43, 55, 70, 75, 77, 72, 68, 51, 32, 43, 74, 
    86, 113, 111, 97, 80, 79, 96, 99, 97, 100, 90, 85, 82, 76, 66, 59, 53, 46, 50, 58, 71, 81, 91, 90, 86, 74, 58, 55, 68, 85, 
    
    -- channel=92
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 12, 7, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 12, 1, 8, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 3, 14, 2, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 6, 2, 0, 0, 0, 6, 8, 2, 0, 2, 2, 5, 4, 6, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 1, 0, 0, 7, 13, 0, 0, 0, 2, 14, 17, 15, 14, 11, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 6, 6, 0, 0, 16, 8, 0, 0, 2, 4, 5, 6, 11, 9, 6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 7, 2, 0, 0, 12, 8, 5, 11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 16, 10, 11, 0, 0, 1, 0, 2, 0, 0, 6, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 1, 0, 
    0, 0, 1, 19, 19, 9, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 9, 0, 
    0, 0, 0, 18, 18, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 11, 0, 
    0, 0, 0, 12, 14, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 11, 0, 
    0, 0, 0, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=93
    113, 87, 103, 91, 84, 89, 97, 103, 84, 81, 65, 53, 42, 34, 36, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 11, 5, 0, 
    151, 142, 136, 102, 88, 86, 98, 107, 95, 99, 86, 76, 63, 57, 52, 41, 0, 0, 0, 0, 0, 0, 5, 20, 30, 37, 24, 7, 3, 1, 
    154, 146, 129, 108, 99, 100, 112, 115, 113, 116, 107, 98, 81, 71, 74, 62, 28, 0, 0, 0, 0, 0, 0, 12, 33, 44, 32, 13, 4, 11, 
    141, 135, 114, 113, 112, 110, 123, 128, 124, 126, 119, 106, 87, 72, 73, 80, 75, 37, 0, 0, 0, 11, 13, 10, 25, 34, 31, 28, 25, 30, 
    142, 129, 114, 135, 126, 118, 128, 131, 139, 133, 127, 117, 108, 86, 73, 76, 97, 89, 75, 58, 52, 45, 36, 20, 17, 16, 17, 27, 38, 43, 
    136, 110, 127, 137, 130, 131, 136, 141, 150, 143, 137, 127, 125, 106, 92, 85, 102, 108, 110, 88, 70, 40, 29, 10, 0, 0, 0, 15, 33, 43, 
    123, 112, 127, 127, 129, 130, 141, 147, 147, 137, 137, 127, 122, 101, 90, 79, 93, 103, 115, 100, 94, 56, 40, 7, 0, 2, 9, 24, 34, 42, 
    123, 119, 125, 135, 139, 130, 131, 134, 148, 145, 143, 135, 127, 114, 104, 89, 78, 82, 103, 105, 119, 92, 59, 18, 0, 15, 28, 35, 35, 42, 
    98, 101, 135, 151, 147, 144, 141, 141, 149, 147, 144, 139, 144, 160, 162, 141, 96, 72, 83, 98, 111, 86, 41, 7, 0, 2, 9, 19, 30, 42, 
    32, 74, 124, 128, 135, 151, 159, 147, 140, 134, 161, 183, 186, 189, 186, 171, 121, 86, 83, 97, 93, 43, 0, 0, 0, 0, 0, 2, 17, 37, 
    3, 94, 165, 161, 169, 181, 171, 143, 128, 130, 189, 227, 224, 162, 101, 93, 71, 80, 92, 106, 89, 27, 0, 0, 0, 0, 0, 0, 11, 28, 
    4, 99, 186, 200, 218, 207, 176, 138, 134, 152, 210, 222, 205, 167, 100, 80, 68, 103, 118, 113, 85, 12, 0, 0, 0, 0, 0, 0, 1, 15, 
    18, 78, 151, 196, 215, 208, 186, 167, 172, 195, 218, 187, 167, 174, 181, 197, 175, 199, 179, 144, 93, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 55, 125, 196, 219, 197, 184, 191, 221, 242, 251, 210, 191, 204, 230, 264, 253, 250, 231, 191, 118, 44, 0, 0, 0, 0, 15, 16, 0, 0, 
    46, 59, 119, 187, 213, 182, 166, 189, 245, 263, 267, 238, 224, 226, 241, 262, 247, 247, 243, 219, 145, 58, 0, 0, 0, 1, 65, 58, 12, 0, 
    84, 104, 144, 195, 221, 179, 160, 183, 216, 228, 218, 209, 220, 200, 193, 207, 204, 204, 186, 161, 86, 0, 0, 0, 0, 2, 84, 88, 34, 0, 
    97, 122, 166, 214, 239, 187, 139, 157, 175, 206, 188, 196, 190, 149, 90, 112, 108, 103, 68, 16, 0, 0, 0, 0, 0, 15, 98, 115, 53, 0, 
    91, 100, 144, 222, 261, 211, 109, 102, 119, 200, 214, 202, 175, 155, 124, 130, 67, 16, 0, 0, 0, 0, 0, 0, 0, 30, 122, 158, 84, 0, 
    109, 111, 150, 218, 260, 223, 90, 9, 0, 105, 173, 153, 123, 139, 168, 189, 93, 0, 0, 0, 0, 0, 0, 0, 0, 33, 134, 202, 132, 23, 
    128, 129, 156, 201, 229, 185, 51, 0, 0, 0, 0, 23, 29, 61, 78, 107, 69, 0, 0, 0, 0, 0, 0, 0, 0, 25, 133, 211, 159, 53, 
    140, 125, 133, 171, 187, 132, 27, 0, 0, 0, 0, 0, 0, 2, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 98, 173, 154, 61, 
    139, 123, 128, 149, 153, 125, 70, 24, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 115, 132, 66, 
    116, 129, 141, 136, 140, 156, 152, 100, 49, 15, 33, 41, 39, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 92, 86, 
    116, 129, 143, 122, 108, 139, 184, 155, 124, 88, 89, 74, 67, 47, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 65, 
    129, 137, 144, 142, 126, 96, 122, 121, 125, 93, 77, 82, 90, 94, 67, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    112, 116, 133, 144, 152, 102, 79, 86, 95, 64, 36, 74, 104, 123, 92, 51, 26, 15, 4, 0, 0, 0, 0, 0, 0, 0, 0, 25, 31, 24, 
    105, 97, 107, 122, 126, 92, 83, 58, 68, 78, 67, 100, 111, 125, 107, 80, 61, 58, 53, 35, 27, 39, 48, 51, 39, 31, 30, 25, 19, 42, 
    95, 109, 115, 129, 123, 100, 108, 99, 87, 97, 109, 124, 114, 121, 112, 99, 79, 65, 60, 54, 64, 79, 88, 88, 82, 72, 54, 38, 24, 62, 
    108, 141, 150, 148, 134, 130, 132, 128, 136, 141, 134, 126, 100, 90, 85, 82, 77, 62, 60, 67, 82, 94, 106, 110, 108, 91, 72, 53, 58, 85, 
    140, 163, 146, 117, 100, 108, 125, 112, 117, 115, 120, 115, 88, 62, 47, 50, 67, 70, 79, 84, 92, 105, 116, 120, 116, 104, 92, 89, 92, 97, 
    
    -- channel=94
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 10, 7, 0, 0, 17, 23, 10, 0, 0, 0, 6, 15, 31, 7, 0, 0, 
    0, 0, 0, 0, 1, 21, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 34, 21, 8, 0, 0, 0, 2, 16, 11, 5, 6, 
    6, 4, 0, 0, 0, 10, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 31, 27, 24, 26, 17, 7, 1, 0, 10, 10, 
    12, 16, 0, 0, 0, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 12, 1, 17, 38, 33, 21, 2, 0, 8, 17, 
    0, 14, 5, 0, 0, 6, 0, 3, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 19, 24, 24, 18, 5, 7, 13, 
    0, 25, 12, 0, 0, 2, 3, 5, 0, 0, 0, 0, 0, 0, 0, 11, 3, 0, 0, 0, 4, 0, 0, 16, 17, 22, 33, 27, 18, 20, 
    0, 33, 15, 4, 3, 5, 9, 4, 4, 0, 0, 5, 0, 0, 0, 11, 17, 11, 0, 0, 0, 0, 0, 4, 5, 6, 22, 22, 20, 22, 
    4, 23, 15, 5, 0, 6, 17, 11, 2, 0, 6, 0, 0, 0, 0, 5, 22, 27, 19, 0, 0, 0, 0, 0, 2, 2, 8, 12, 15, 19, 
    24, 29, 16, 2, 0, 0, 6, 8, 0, 0, 5, 0, 0, 0, 0, 0, 0, 28, 40, 10, 15, 0, 0, 0, 22, 23, 20, 22, 18, 18, 
    57, 53, 22, 24, 14, 0, 0, 0, 4, 8, 8, 0, 0, 18, 4, 0, 0, 11, 37, 20, 28, 18, 0, 7, 32, 21, 22, 29, 24, 22, 
    90, 50, 0, 18, 11, 0, 2, 0, 3, 15, 19, 0, 0, 40, 66, 22, 0, 10, 27, 13, 14, 0, 0, 21, 31, 12, 13, 23, 27, 27, 
    112, 45, 0, 5, 0, 0, 1, 0, 0, 28, 50, 25, 0, 10, 31, 43, 19, 10, 27, 8, 0, 0, 0, 18, 33, 21, 16, 23, 26, 26, 
    101, 76, 57, 45, 13, 8, 0, 0, 8, 37, 42, 24, 12, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 6, 17, 15, 10, 18, 23, 25, 
    49, 77, 93, 50, 12, 21, 10, 0, 17, 28, 0, 0, 9, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 13, 0, 0, 9, 20, 
    0, 59, 99, 56, 10, 16, 33, 34, 35, 23, 0, 0, 0, 46, 40, 32, 30, 34, 9, 0, 0, 0, 0, 7, 25, 37, 0, 0, 0, 19, 
    0, 36, 86, 59, 14, 0, 33, 70, 54, 35, 48, 21, 9, 53, 64, 51, 50, 56, 46, 24, 0, 0, 6, 18, 50, 68, 31, 0, 0, 13, 
    0, 31, 69, 46, 11, 0, 17, 98, 62, 16, 68, 46, 9, 49, 74, 77, 71, 68, 83, 71, 18, 1, 3, 11, 55, 76, 57, 0, 0, 0, 
    12, 55, 91, 58, 19, 0, 0, 121, 73, 0, 42, 36, 0, 19, 18, 27, 53, 50, 60, 42, 7, 0, 0, 0, 42, 74, 64, 0, 0, 0, 
    0, 40, 97, 76, 31, 0, 0, 100, 146, 58, 62, 37, 0, 34, 0, 0, 0, 0, 11, 0, 0, 0, 0, 4, 49, 85, 80, 2, 0, 0, 
    0, 21, 82, 86, 49, 0, 0, 23, 171, 156, 118, 67, 30, 109, 106, 10, 0, 0, 3, 15, 13, 21, 0, 0, 46, 95, 107, 37, 0, 0, 
    1, 28, 84, 89, 48, 4, 0, 0, 44, 88, 106, 88, 54, 89, 113, 62, 8, 0, 5, 33, 36, 46, 14, 0, 24, 89, 128, 82, 0, 0, 
    3, 19, 67, 77, 34, 0, 0, 0, 0, 0, 0, 20, 17, 31, 35, 24, 33, 17, 8, 16, 17, 42, 50, 33, 32, 69, 124, 113, 0, 0, 
    17, 26, 36, 53, 34, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 11, 12, 14, 4, 13, 42, 48, 50, 44, 90, 127, 29, 0, 
    24, 45, 24, 28, 50, 34, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 2, 0, 0, 7, 26, 52, 25, 51, 122, 90, 0, 
    19, 41, 24, 2, 34, 82, 61, 0, 0, 0, 0, 11, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 39, 8, 16, 64, 80, 46, 
    30, 32, 36, 10, 0, 23, 82, 48, 6, 19, 18, 27, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 6, 31, 
    24, 30, 65, 48, 6, 0, 41, 60, 0, 0, 8, 31, 46, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 0, 
    13, 13, 57, 41, 12, 0, 13, 25, 1, 11, 3, 12, 34, 25, 0, 0, 7, 9, 7, 2, 0, 6, 1, 0, 0, 0, 0, 16, 13, 11, 
    10, 8, 27, 14, 2, 3, 14, 0, 0, 20, 10, 9, 26, 31, 20, 10, 13, 9, 14, 17, 10, 16, 14, 1, 0, 2, 0, 0, 11, 38, 
    14, 21, 18, 19, 32, 32, 33, 19, 19, 31, 17, 12, 13, 20, 36, 28, 12, 1, 7, 19, 16, 18, 24, 9, 6, 8, 0, 0, 15, 35, 
    
    -- channel=95
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=96
    16, 36, 43, 32, 39, 52, 51, 54, 67, 73, 72, 65, 65, 77, 84, 79, 79, 77, 90, 88, 86, 81, 90, 98, 121, 120, 79, 77, 93, 93, 
    42, 55, 56, 52, 60, 73, 74, 76, 84, 88, 86, 79, 77, 86, 91, 87, 89, 90, 85, 82, 83, 86, 96, 112, 134, 110, 62, 68, 93, 95, 
    58, 62, 64, 69, 82, 87, 89, 89, 92, 95, 93, 86, 85, 91, 92, 89, 90, 87, 85, 80, 73, 89, 106, 115, 117, 84, 54, 65, 95, 97, 
    67, 72, 84, 92, 96, 96, 99, 96, 95, 96, 94, 89, 89, 90, 90, 86, 86, 84, 82, 62, 54, 84, 114, 109, 94, 64, 46, 67, 92, 99, 
    84, 96, 104, 103, 97, 99, 101, 96, 92, 90, 90, 87, 88, 84, 82, 80, 80, 80, 73, 48, 57, 108, 105, 92, 82, 48, 47, 71, 92, 102, 
    99, 103, 100, 95, 94, 97, 97, 90, 86, 83, 85, 83, 83, 78, 76, 74, 72, 74, 67, 58, 102, 136, 86, 65, 70, 50, 68, 83, 97, 100, 
    93, 95, 90, 89, 89, 91, 90, 85, 82, 80, 81, 74, 72, 67, 68, 68, 63, 65, 68, 90, 135, 133, 61, 42, 61, 75, 87, 91, 96, 97, 
    88, 91, 88, 90, 88, 88, 89, 84, 80, 72, 70, 60, 59, 60, 65, 69, 65, 67, 80, 107, 127, 103, 46, 39, 76, 88, 91, 91, 93, 96, 
    87, 92, 90, 91, 90, 88, 90, 86, 79, 66, 67, 55, 55, 59, 54, 43, 28, 18, 61, 90, 90, 87, 52, 53, 89, 94, 92, 93, 93, 96, 
    87, 92, 91, 91, 90, 89, 92, 86, 81, 69, 61, 33, 12, 14, 0, 0, 0, 0, 15, 37, 37, 108, 99, 71, 73, 87, 95, 95, 94, 97, 
    87, 92, 91, 90, 91, 89, 91, 85, 71, 50, 28, 0, 0, 0, 2, 3, 18, 32, 44, 0, 0, 114, 158, 105, 62, 46, 99, 103, 96, 98, 
    88, 91, 90, 88, 93, 91, 90, 72, 51, 34, 18, 8, 45, 91, 96, 89, 108, 117, 43, 0, 0, 83, 180, 144, 72, 38, 86, 117, 99, 99, 
    88, 90, 90, 89, 98, 96, 80, 59, 46, 61, 70, 66, 97, 140, 133, 92, 103, 97, 0, 0, 0, 23, 143, 180, 103, 60, 85, 115, 101, 97, 
    87, 88, 92, 88, 87, 89, 69, 62, 72, 98, 71, 53, 95, 123, 109, 62, 40, 5, 0, 0, 0, 0, 95, 171, 137, 87, 91, 76, 74, 95, 
    88, 89, 93, 86, 61, 57, 70, 67, 101, 77, 43, 48, 79, 53, 18, 0, 0, 0, 0, 0, 0, 6, 117, 154, 131, 121, 75, 10, 10, 94, 
    90, 90, 94, 93, 66, 54, 71, 76, 86, 92, 61, 77, 32, 0, 0, 0, 0, 0, 0, 0, 0, 85, 180, 136, 93, 115, 34, 0, 0, 109, 
    93, 89, 72, 91, 92, 76, 66, 70, 111, 117, 71, 84, 0, 0, 0, 0, 0, 0, 0, 0, 12, 153, 170, 70, 46, 42, 0, 0, 0, 116, 
    94, 53, 12, 64, 117, 87, 56, 91, 136, 108, 60, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 90, 90, 19, 0, 0, 0, 0, 5, 116, 
    68, 0, 0, 56, 150, 106, 62, 109, 135, 106, 64, 39, 0, 0, 0, 0, 0, 0, 23, 14, 0, 0, 24, 0, 0, 0, 1, 14, 45, 138, 
    35, 0, 0, 85, 153, 111, 78, 120, 136, 100, 70, 44, 0, 0, 0, 0, 0, 85, 135, 101, 27, 0, 0, 0, 4, 9, 17, 54, 111, 163, 
    31, 0, 36, 69, 121, 116, 99, 135, 122, 69, 38, 15, 0, 0, 0, 0, 67, 175, 160, 93, 68, 0, 0, 0, 32, 38, 61, 115, 167, 142, 
    52, 91, 96, 10, 74, 125, 118, 132, 100, 37, 0, 0, 0, 0, 0, 0, 137, 194, 105, 78, 90, 47, 0, 0, 40, 56, 106, 166, 147, 87, 
    78, 106, 68, 0, 42, 132, 135, 110, 72, 18, 5, 0, 0, 0, 0, 24, 175, 155, 71, 91, 101, 85, 4, 0, 10, 72, 151, 159, 96, 66, 
    91, 80, 55, 0, 33, 140, 135, 83, 36, 5, 18, 0, 0, 0, 0, 48, 176, 124, 53, 80, 96, 111, 48, 0, 0, 105, 174, 134, 82, 76, 
    91, 69, 61, 3, 27, 127, 112, 37, 0, 0, 0, 0, 0, 0, 0, 44, 163, 115, 30, 53, 98, 115, 85, 0, 12, 134, 172, 121, 90, 87, 
    87, 60, 57, 14, 33, 104, 87, 22, 0, 0, 0, 0, 0, 3, 7, 59, 161, 115, 34, 41, 99, 127, 114, 55, 57, 141, 152, 113, 98, 89, 
    87, 71, 61, 49, 68, 120, 102, 70, 63, 65, 77, 79, 78, 85, 87, 109, 156, 93, 36, 71, 100, 134, 126, 98, 99, 132, 122, 104, 99, 86, 
    83, 89, 96, 90, 106, 121, 110, 101, 98, 98, 103, 103, 105, 110, 112, 117, 132, 79, 33, 66, 96, 117, 137, 113, 107, 111, 105, 99, 92, 80, 
    82, 94, 99, 93, 84, 74, 87, 98, 87, 83, 85, 86, 88, 92, 97, 99, 104, 82, 63, 69, 98, 138, 133, 109, 103, 103, 100, 94, 83, 76, 
    78, 76, 62, 50, 43, 47, 85, 97, 75, 66, 67, 69, 73, 76, 81, 86, 92, 89, 74, 78, 114, 130, 109, 98, 98, 99, 95, 88, 79, 78, 
    
    -- channel=97
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 27, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 47, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 109, 78, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 95, 23, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 59, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 71, 52, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 82, 89, 87, 56, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 32, 40, 59, 91, 134, 190, 191, 143, 129, 89, 49, 40, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 90, 168, 189, 192, 201, 218, 229, 210, 222, 235, 146, 58, 34, 27, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 108, 159, 182, 158, 127, 102, 105, 93, 98, 204, 282, 213, 101, 42, 26, 46, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 79, 79, 101, 110, 64, 31, 37, 52, 43, 96, 213, 281, 262, 169, 54, 28, 45, 42, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 54, 80, 39, 44, 89, 101, 67, 49, 60, 77, 82, 164, 257, 270, 279, 218, 71, 20, 28, 28, 9, 0, 
    0, 0, 0, 0, 0, 0, 37, 69, 89, 74, 64, 82, 111, 84, 68, 70, 73, 113, 182, 249, 262, 262, 250, 176, 72, 26, 24, 29, 48, 34, 
    0, 0, 0, 0, 5, 74, 121, 111, 117, 110, 88, 98, 113, 90, 137, 208, 240, 268, 286, 280, 261, 260, 203, 64, 18, 44, 28, 49, 111, 119, 
    0, 0, 0, 0, 64, 80, 87, 104, 126, 95, 61, 70, 68, 87, 223, 303, 300, 292, 282, 272, 270, 230, 122, 31, 34, 66, 81, 119, 169, 169, 
    0, 0, 0, 76, 136, 113, 87, 96, 97, 54, 47, 72, 81, 114, 241, 290, 273, 260, 265, 266, 265, 238, 165, 111, 121, 159, 188, 196, 182, 177, 
    0, 0, 50, 189, 207, 134, 78, 87, 76, 39, 40, 78, 113, 151, 247, 274, 255, 264, 267, 246, 246, 265, 248, 219, 222, 232, 220, 202, 188, 161, 
    0, 0, 163, 261, 219, 153, 86, 88, 68, 37, 43, 69, 94, 156, 252, 264, 254, 275, 222, 146, 118, 167, 229, 252, 257, 243, 225, 210, 181, 120, 
    0, 19, 177, 221, 200, 166, 100, 77, 47, 38, 54, 84, 99, 158, 255, 255, 264, 249, 125, 57, 53, 59, 130, 217, 256, 239, 209, 190, 132, 38, 
    0, 30, 93, 103, 154, 168, 108, 77, 46, 45, 83, 145, 159, 196, 253, 254, 266, 194, 68, 67, 83, 62, 65, 144, 206, 202, 192, 144, 48, 0, 
    0, 20, 72, 93, 146, 181, 116, 66, 53, 65, 109, 154, 155, 212, 268, 270, 264, 165, 67, 70, 65, 61, 54, 91, 166, 200, 181, 94, 7, 0, 
    0, 14, 83, 114, 151, 186, 132, 80, 81, 107, 139, 150, 169, 239, 272, 268, 250, 155, 78, 89, 90, 79, 49, 63, 135, 198, 161, 62, 4, 0, 
    0, 4, 68, 109, 147, 183, 129, 82, 94, 125, 153, 157, 175, 221, 232, 236, 224, 144, 79, 106, 102, 83, 54, 47, 100, 159, 118, 41, 8, 2, 
    0, 0, 51, 89, 131, 165, 137, 109, 137, 176, 212, 227, 231, 239, 242, 244, 225, 137, 67, 109, 144, 117, 82, 46, 65, 107, 77, 27, 13, 12, 
    0, 0, 40, 91, 122, 139, 118, 109, 118, 127, 139, 147, 152, 156, 152, 147, 142, 100, 71, 86, 97, 90, 57, 38, 32, 39, 29, 21, 21, 18, 
    0, 0, 35, 72, 96, 88, 68, 62, 60, 57, 60, 58, 58, 55, 52, 47, 44, 33, 53, 97, 84, 80, 66, 31, 22, 21, 21, 22, 25, 23, 
    0, 28, 63, 84, 91, 90, 96, 97, 85, 88, 89, 83, 77, 69, 64, 56, 50, 43, 44, 73, 108, 104, 60, 29, 26, 28, 28, 28, 29, 32, 
    
    -- channel=98
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 35, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 14, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 12, 16, 23, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 48, 72, 20, 25, 50, 6, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 52, 75, 76, 76, 89, 108, 83, 35, 52, 55, 27, 24, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 44, 77, 78, 55, 29, 50, 60, 22, 37, 75, 53, 48, 31, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 2, 14, 46, 35, 19, 0, 19, 9, 1, 65, 89, 59, 72, 40, 13, 16, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 21, 48, 21, 6, 0, 0, 0, 40, 88, 80, 79, 98, 30, 3, 15, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 12, 32, 20, 15, 50, 29, 0, 0, 0, 12, 46, 81, 77, 76, 105, 82, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 31, 31, 43, 61, 41, 34, 66, 11, 4, 59, 75, 89, 93, 89, 74, 85, 83, 20, 0, 0, 0, 0, 18, 0, 
    0, 0, 0, 0, 0, 39, 40, 34, 58, 47, 33, 23, 58, 15, 53, 109, 110, 102, 90, 87, 76, 63, 40, 0, 0, 0, 16, 35, 52, 21, 
    0, 0, 0, 0, 56, 68, 45, 28, 53, 30, 28, 29, 65, 30, 73, 110, 101, 85, 94, 107, 98, 70, 52, 28, 26, 52, 66, 67, 56, 42, 
    0, 0, 0, 42, 90, 81, 39, 28, 49, 24, 29, 43, 73, 39, 82, 106, 87, 94, 134, 127, 111, 98, 83, 78, 80, 89, 84, 69, 65, 67, 
    0, 0, 41, 105, 86, 90, 39, 39, 41, 23, 24, 34, 61, 38, 88, 101, 77, 124, 124, 70, 64, 86, 79, 88, 103, 104, 86, 79, 84, 56, 
    0, 0, 90, 90, 61, 88, 43, 43, 30, 25, 15, 36, 66, 45, 90, 89, 79, 131, 60, 20, 32, 55, 63, 73, 104, 98, 78, 88, 65, 10, 
    0, 0, 50, 52, 39, 83, 55, 42, 26, 31, 32, 75, 76, 52, 93, 83, 89, 115, 29, 29, 31, 36, 55, 48, 74, 77, 78, 76, 19, 0, 
    0, 0, 28, 57, 39, 81, 65, 40, 28, 36, 47, 79, 58, 66, 106, 87, 96, 100, 24, 25, 28, 30, 47, 39, 50, 74, 86, 55, 0, 0, 
    0, 0, 28, 66, 48, 83, 78, 45, 36, 42, 51, 67, 57, 83, 103, 81, 90, 94, 34, 28, 34, 32, 36, 40, 37, 74, 87, 41, 0, 0, 
    0, 0, 15, 55, 50, 75, 74, 41, 42, 52, 60, 72, 72, 88, 95, 84, 90, 96, 35, 30, 37, 44, 34, 41, 31, 67, 70, 27, 1, 0, 
    0, 0, 0, 43, 51, 78, 79, 64, 79, 93, 103, 109, 109, 113, 115, 105, 94, 90, 32, 45, 57, 52, 36, 38, 31, 49, 40, 16, 7, 3, 
    0, 0, 0, 42, 60, 75, 67, 61, 69, 72, 75, 77, 79, 80, 79, 72, 62, 58, 23, 39, 37, 28, 34, 26, 18, 20, 16, 12, 12, 9, 
    0, 0, 1, 33, 47, 41, 29, 36, 39, 36, 36, 34, 33, 32, 30, 26, 22, 28, 26, 33, 35, 39, 38, 18, 12, 12, 12, 11, 12, 8, 
    0, 0, 11, 31, 42, 41, 46, 63, 54, 48, 50, 46, 42, 37, 32, 28, 23, 26, 33, 39, 46, 47, 28, 15, 14, 14, 15, 14, 13, 10, 
    
    -- channel=99
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=100
    186, 202, 208, 212, 224, 230, 229, 228, 223, 211, 199, 193, 193, 193, 182, 169, 160, 153, 159, 133, 137, 119, 112, 89, 68, 73, 72, 80, 88, 90, 
    222, 223, 211, 201, 210, 216, 207, 205, 199, 187, 177, 171, 171, 172, 163, 152, 146, 143, 122, 119, 127, 112, 95, 90, 76, 37, 40, 71, 91, 94, 
    211, 205, 191, 186, 191, 191, 180, 175, 171, 164, 155, 150, 150, 150, 144, 137, 130, 129, 121, 116, 111, 88, 75, 84, 57, 25, 31, 70, 94, 94, 
    182, 185, 185, 185, 172, 166, 157, 152, 150, 145, 137, 132, 134, 134, 131, 127, 120, 119, 123, 113, 83, 71, 73, 56, 43, 40, 45, 77, 95, 94, 
    169, 169, 163, 154, 143, 143, 138, 134, 132, 130, 124, 121, 122, 123, 124, 122, 119, 117, 120, 102, 85, 96, 83, 53, 51, 51, 72, 98, 110, 103, 
    144, 136, 129, 123, 123, 125, 123, 121, 121, 121, 120, 120, 120, 118, 119, 119, 120, 116, 109, 93, 102, 88, 67, 73, 68, 71, 101, 115, 118, 103, 
    113, 112, 112, 114, 115, 116, 113, 115, 117, 119, 120, 119, 118, 116, 116, 114, 119, 120, 109, 101, 94, 47, 31, 68, 80, 97, 108, 111, 113, 103, 
    104, 107, 110, 114, 114, 117, 114, 116, 118, 121, 116, 109, 119, 125, 131, 128, 132, 130, 111, 102, 66, 7, 5, 51, 89, 108, 109, 106, 110, 103, 
    105, 109, 112, 116, 115, 118, 117, 118, 119, 120, 118, 122, 131, 126, 127, 111, 94, 73, 41, 43, 21, 0, 17, 60, 85, 100, 105, 103, 105, 101, 
    107, 111, 112, 115, 114, 117, 117, 118, 117, 118, 127, 115, 88, 59, 56, 57, 65, 78, 88, 67, 12, 0, 6, 65, 98, 84, 83, 94, 100, 99, 
    112, 114, 113, 116, 113, 116, 116, 115, 114, 105, 90, 65, 79, 97, 120, 143, 159, 177, 202, 149, 87, 33, 0, 26, 69, 83, 76, 78, 91, 94, 
    113, 117, 115, 118, 112, 115, 117, 112, 97, 76, 85, 108, 132, 139, 150, 157, 138, 131, 134, 98, 119, 110, 4, 0, 9, 66, 81, 75, 82, 89, 
    115, 117, 115, 118, 114, 113, 115, 95, 79, 99, 121, 111, 95, 74, 55, 58, 55, 45, 18, 13, 105, 140, 58, 0, 0, 20, 74, 70, 70, 80, 
    117, 119, 115, 116, 116, 93, 80, 68, 96, 105, 73, 50, 57, 42, 14, 9, 31, 3, 0, 13, 104, 121, 104, 36, 0, 0, 36, 44, 37, 41, 
    116, 119, 114, 108, 105, 83, 62, 78, 70, 47, 46, 58, 69, 40, 0, 0, 0, 0, 0, 79, 103, 94, 143, 131, 42, 11, 22, 21, 9, 15, 
    113, 118, 113, 96, 88, 105, 98, 81, 42, 47, 58, 79, 91, 47, 6, 5, 38, 68, 112, 122, 102, 126, 161, 104, 67, 32, 0, 0, 31, 51, 
    112, 116, 110, 75, 48, 67, 72, 51, 70, 47, 41, 46, 36, 40, 89, 117, 136, 148, 142, 122, 119, 120, 62, 10, 37, 7, 0, 7, 80, 96, 
    114, 112, 80, 41, 25, 31, 37, 47, 54, 31, 29, 29, 0, 49, 127, 131, 128, 118, 114, 126, 152, 96, 0, 0, 4, 22, 31, 65, 85, 113, 
    116, 92, 48, 71, 42, 13, 19, 41, 27, 20, 17, 45, 25, 71, 112, 110, 99, 90, 123, 167, 197, 168, 74, 26, 41, 62, 73, 79, 76, 122, 
    105, 71, 113, 151, 61, 7, 11, 43, 26, 13, 7, 22, 17, 72, 102, 100, 85, 108, 139, 123, 124, 177, 153, 94, 79, 82, 89, 85, 102, 125, 
    79, 87, 178, 168, 79, 15, 14, 38, 15, 13, 0, 0, 0, 63, 99, 89, 91, 127, 82, 22, 15, 71, 139, 133, 106, 96, 84, 96, 115, 73, 
    77, 105, 90, 77, 71, 14, 25, 29, 8, 5, 3, 19, 19, 71, 87, 77, 108, 86, 17, 17, 21, 2, 75, 125, 102, 67, 68, 91, 60, 19, 
    94, 94, 9, 21, 67, 23, 25, 16, 4, 0, 17, 51, 39, 76, 95, 97, 113, 35, 14, 17, 16, 0, 25, 96, 86, 55, 73, 52, 19, 21, 
    90, 72, 25, 22, 69, 41, 21, 11, 7, 0, 20, 23, 35, 100, 108, 113, 92, 18, 29, 15, 10, 10, 0, 61, 88, 82, 70, 28, 23, 41, 
    71, 58, 41, 21, 66, 43, 3, 0, 0, 0, 4, 0, 33, 85, 84, 95, 66, 12, 33, 30, 7, 1, 0, 28, 88, 96, 57, 19, 25, 38, 
    59, 56, 39, 19, 60, 57, 20, 11, 34, 69, 93, 89, 114, 130, 131, 148, 111, 31, 25, 53, 52, 39, 13, 12, 75, 93, 44, 12, 18, 27, 
    53, 47, 51, 42, 72, 83, 53, 53, 71, 96, 117, 123, 129, 134, 132, 145, 125, 52, 33, 44, 60, 26, 12, 5, 43, 48, 18, 10, 14, 20, 
    54, 41, 47, 39, 59, 45, 13, 11, 18, 24, 29, 33, 39, 42, 42, 48, 51, 18, 53, 52, 32, 18, 24, 10, 16, 13, 8, 10, 11, 13, 
    61, 54, 35, 13, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 31, 53, 49, 58, 25, 8, 8, 7, 7, 8, 11, 12, 
    57, 52, 26, 0, 0, 0, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 26, 17, 4, 5, 5, 3, 5, 7, 8, 14, 
    
    -- channel=101
    20, 22, 27, 27, 27, 31, 34, 32, 35, 35, 32, 31, 30, 32, 32, 28, 20, 2, 39, 47, 23, 27, 33, 11, 0, 19, 22, 16, 20, 18, 
    30, 30, 31, 25, 27, 34, 34, 33, 36, 34, 31, 29, 27, 30, 31, 27, 25, 25, 24, 25, 23, 16, 19, 4, 14, 24, 12, 12, 20, 19, 
    31, 27, 28, 19, 29, 33, 33, 32, 32, 30, 29, 27, 25, 30, 28, 25, 24, 27, 20, 19, 20, 6, 0, 9, 28, 15, 2, 6, 16, 16, 
    28, 23, 27, 32, 37, 31, 31, 30, 29, 28, 27, 25, 25, 27, 25, 24, 22, 22, 21, 28, 16, 0, 0, 10, 10, 7, 0, 7, 13, 15, 
    23, 29, 36, 39, 34, 27, 28, 26, 27, 26, 24, 22, 25, 26, 22, 23, 23, 19, 24, 30, 0, 4, 32, 6, 5, 6, 0, 13, 16, 26, 
    31, 35, 36, 27, 25, 25, 28, 24, 23, 23, 22, 23, 23, 24, 21, 19, 17, 15, 21, 0, 0, 29, 45, 20, 23, 6, 11, 20, 25, 29, 
    24, 25, 25, 22, 23, 23, 24, 21, 22, 21, 23, 25, 15, 11, 12, 16, 15, 16, 15, 0, 6, 32, 14, 10, 15, 15, 21, 26, 25, 22, 
    19, 21, 21, 21, 23, 22, 23, 21, 22, 21, 21, 20, 10, 14, 15, 20, 17, 17, 11, 1, 20, 15, 0, 0, 6, 15, 18, 21, 21, 19, 
    20, 22, 23, 21, 23, 23, 24, 22, 24, 26, 18, 13, 8, 14, 11, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 11, 19, 19, 19, 
    22, 22, 23, 22, 22, 22, 24, 23, 23, 20, 12, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 16, 16, 6, 4, 15, 18, 20, 
    23, 22, 23, 22, 23, 23, 22, 23, 18, 11, 12, 6, 0, 0, 0, 0, 7, 19, 62, 73, 0, 0, 0, 0, 39, 12, 2, 7, 14, 19, 
    23, 21, 23, 21, 24, 24, 21, 23, 23, 8, 0, 0, 0, 13, 30, 39, 37, 42, 79, 57, 0, 7, 0, 0, 0, 20, 10, 13, 9, 15, 
    22, 21, 24, 23, 21, 23, 24, 30, 0, 0, 0, 19, 9, 20, 33, 36, 15, 19, 22, 0, 0, 32, 10, 0, 0, 0, 16, 31, 16, 12, 
    23, 21, 24, 24, 20, 12, 16, 0, 0, 10, 29, 9, 5, 21, 7, 3, 0, 4, 0, 0, 0, 21, 22, 8, 0, 0, 8, 23, 3, 0, 
    24, 22, 25, 26, 30, 0, 0, 0, 12, 19, 6, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 23, 83, 29, 0, 9, 12, 0, 0, 
    24, 23, 27, 20, 18, 7, 1, 22, 0, 7, 8, 5, 39, 34, 0, 0, 0, 0, 0, 0, 0, 0, 53, 106, 34, 21, 12, 0, 0, 0, 
    24, 24, 24, 0, 0, 1, 32, 3, 0, 25, 5, 0, 46, 0, 0, 0, 0, 0, 10, 2, 0, 7, 68, 17, 2, 5, 0, 0, 0, 0, 
    28, 29, 15, 0, 0, 0, 1, 0, 30, 26, 14, 0, 0, 0, 0, 4, 8, 11, 3, 0, 13, 28, 5, 0, 0, 0, 0, 0, 0, 11, 
    34, 39, 0, 0, 0, 3, 0, 0, 23, 16, 8, 4, 0, 0, 0, 7, 5, 0, 0, 38, 72, 58, 16, 0, 0, 0, 0, 0, 0, 20, 
    50, 5, 0, 5, 29, 9, 0, 0, 30, 7, 0, 0, 0, 0, 0, 6, 0, 0, 26, 53, 58, 73, 47, 0, 0, 0, 1, 2, 0, 56, 
    31, 0, 9, 78, 32, 17, 0, 13, 27, 5, 0, 0, 0, 0, 0, 1, 0, 20, 77, 14, 0, 22, 34, 20, 7, 11, 10, 0, 46, 74, 
    0, 0, 46, 50, 10, 17, 0, 23, 12, 11, 0, 0, 0, 0, 0, 0, 0, 86, 46, 0, 0, 0, 0, 7, 22, 14, 0, 35, 67, 27, 
    3, 20, 10, 0, 0, 4, 12, 22, 3, 0, 0, 0, 0, 0, 0, 0, 21, 69, 0, 0, 9, 0, 0, 2, 14, 0, 7, 58, 30, 0, 
    19, 22, 0, 0, 0, 14, 22, 15, 0, 0, 0, 2, 0, 0, 2, 0, 38, 46, 0, 0, 0, 0, 0, 0, 0, 0, 40, 45, 7, 0, 
    14, 5, 3, 0, 0, 12, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 31, 0, 0, 0, 0, 0, 0, 0, 23, 54, 29, 2, 5, 
    9, 4, 3, 0, 0, 25, 28, 0, 0, 0, 6, 0, 0, 13, 19, 22, 41, 39, 3, 4, 2, 14, 0, 0, 0, 40, 53, 17, 3, 5, 
    4, 10, 1, 1, 0, 38, 34, 2, 2, 14, 33, 42, 39, 42, 46, 65, 80, 60, 0, 0, 15, 28, 8, 0, 0, 38, 32, 6, 2, 4, 
    2, 0, 0, 0, 5, 25, 9, 0, 0, 0, 4, 7, 10, 16, 16, 26, 45, 41, 0, 0, 18, 0, 13, 5, 3, 11, 6, 3, 1, 0, 
    6, 2, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 2, 18, 29, 7, 1, 1, 0, 0, 0, 0, 
    6, 11, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 27, 14, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=102
    80, 88, 88, 92, 97, 100, 101, 104, 102, 100, 95, 93, 93, 92, 90, 87, 87, 91, 77, 66, 80, 69, 58, 58, 51, 46, 54, 58, 60, 63, 
    97, 99, 93, 88, 88, 98, 98, 96, 95, 92, 88, 85, 86, 85, 84, 81, 80, 78, 73, 65, 71, 70, 61, 57, 52, 43, 39, 51, 58, 65, 
    86, 86, 80, 82, 84, 92, 90, 87, 85, 84, 81, 78, 79, 79, 78, 75, 75, 71, 71, 67, 53, 43, 43, 54, 49, 38, 39, 44, 55, 61, 
    75, 79, 86, 88, 85, 85, 82, 81, 80, 78, 74, 72, 72, 73, 73, 69, 70, 66, 65, 58, 33, 13, 23, 38, 37, 38, 40, 37, 51, 55, 
    88, 84, 83, 80, 75, 78, 75, 76, 74, 72, 69, 67, 67, 67, 69, 66, 66, 65, 62, 50, 41, 27, 32, 39, 30, 40, 39, 50, 65, 60, 
    81, 75, 72, 71, 68, 71, 68, 69, 69, 68, 66, 64, 65, 63, 64, 60, 61, 58, 51, 51, 51, 42, 42, 51, 45, 49, 54, 64, 71, 65, 
    69, 67, 66, 68, 66, 66, 64, 65, 66, 67, 65, 58, 53, 51, 52, 48, 51, 53, 50, 56, 49, 38, 37, 48, 54, 59, 64, 63, 66, 67, 
    63, 65, 66, 67, 65, 67, 64, 64, 65, 63, 57, 46, 43, 45, 55, 57, 57, 58, 51, 48, 32, 13, 14, 32, 46, 61, 69, 64, 65, 67, 
    62, 65, 65, 67, 65, 66, 66, 65, 63, 59, 56, 52, 56, 44, 39, 25, 0, 0, 0, 0, 0, 0, 8, 31, 35, 47, 63, 64, 64, 65, 
    63, 64, 64, 66, 64, 65, 66, 65, 63, 60, 56, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 49, 44, 35, 56, 64, 64, 
    64, 65, 63, 65, 65, 63, 65, 64, 58, 41, 8, 0, 0, 0, 0, 21, 35, 45, 39, 10, 0, 0, 0, 11, 40, 47, 35, 35, 59, 62, 
    65, 65, 63, 65, 65, 61, 66, 57, 37, 10, 9, 30, 42, 42, 62, 74, 74, 61, 38, 5, 0, 0, 0, 0, 29, 36, 42, 34, 53, 62, 
    64, 65, 63, 63, 65, 63, 62, 42, 31, 38, 50, 44, 31, 25, 31, 36, 48, 25, 0, 0, 0, 0, 0, 0, 0, 36, 42, 43, 46, 56, 
    64, 66, 64, 62, 56, 44, 25, 32, 37, 43, 22, 16, 10, 13, 22, 15, 12, 0, 0, 0, 0, 0, 0, 0, 0, 21, 33, 30, 21, 17, 
    63, 65, 63, 56, 38, 28, 8, 19, 14, 2, 16, 22, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 37, 18, 27, 9, 0, 0, 
    63, 62, 60, 54, 41, 44, 37, 14, 14, 16, 37, 42, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 36, 42, 20, 0, 0, 0, 0, 
    64, 61, 51, 37, 14, 20, 20, 25, 25, 36, 35, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    65, 44, 11, 0, 0, 7, 23, 30, 20, 37, 32, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    56, 12, 0, 0, 0, 0, 12, 25, 24, 40, 37, 32, 9, 0, 0, 0, 0, 0, 0, 11, 16, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    40, 15, 0, 0, 0, 0, 11, 28, 35, 43, 38, 21, 0, 0, 0, 0, 0, 0, 27, 57, 45, 32, 10, 0, 0, 0, 0, 0, 13, 40, 
    47, 55, 38, 38, 8, 0, 15, 24, 35, 30, 13, 0, 0, 0, 0, 0, 0, 0, 28, 27, 28, 20, 29, 5, 0, 0, 0, 13, 43, 46, 
    65, 63, 22, 7, 2, 0, 10, 29, 33, 15, 4, 0, 0, 0, 0, 0, 0, 0, 22, 22, 37, 34, 22, 26, 0, 0, 0, 18, 37, 35, 
    65, 44, 11, 0, 0, 0, 2, 22, 23, 6, 3, 0, 0, 0, 0, 0, 0, 0, 22, 10, 11, 29, 27, 24, 0, 0, 0, 17, 34, 36, 
    59, 42, 20, 0, 1, 0, 1, 19, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 6, 4, 20, 25, 24, 18, 0, 4, 28, 44, 48, 
    53, 43, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 1, 0, 0, 18, 26, 40, 25, 22, 38, 46, 47, 
    48, 41, 21, 0, 0, 0, 0, 0, 0, 2, 1, 4, 3, 3, 5, 10, 12, 2, 12, 7, 21, 18, 36, 38, 57, 55, 45, 41, 42, 44, 
    45, 36, 36, 32, 36, 39, 48, 56, 60, 63, 64, 65, 67, 67, 66, 61, 58, 40, 37, 10, 13, 18, 20, 46, 53, 48, 44, 44, 43, 40, 
    39, 38, 34, 41, 44, 40, 32, 29, 34, 37, 36, 37, 39, 40, 42, 43, 41, 36, 41, 34, 5, 15, 31, 46, 45, 44, 43, 43, 41, 36, 
    37, 35, 25, 10, 0, 0, 0, 0, 11, 13, 10, 10, 13, 16, 20, 22, 26, 34, 32, 38, 47, 43, 43, 42, 41, 41, 40, 40, 36, 35, 
    28, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 14, 19, 18, 16, 17, 28, 35, 33, 31, 32, 33, 31, 31, 
    
    -- channel=103
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 10, 3, 16, 21, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 7, 14, 27, 21, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 10, 13, 11, 18, 22, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 26, 21, 23, 23, 21, 20, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 16, 17, 33, 26, 25, 23, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 21, 6, 23, 35, 17, 15, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 11, 12, 12, 31, 35, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 10, 16, 32, 45, 41, 12, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 3, 12, 17, 36, 58, 75, 56, 63, 59, 44, 44, 18, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 48, 69, 84, 93, 99, 102, 95, 69, 98, 86, 41, 46, 20, 25, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 44, 76, 70, 59, 52, 44, 36, 30, 40, 107, 88, 35, 45, 29, 44, 28, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 29, 37, 42, 23, 16, 18, 21, 12, 18, 71, 124, 98, 54, 41, 39, 46, 36, 3, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 12, 12, 23, 36, 26, 24, 27, 37, 20, 47, 116, 126, 100, 82, 43, 40, 48, 33, 10, 7, 1, 0, 
    0, 0, 0, 0, 0, 0, 14, 10, 14, 22, 44, 43, 24, 32, 34, 55, 62, 110, 148, 123, 104, 96, 39, 37, 38, 33, 24, 38, 29, 9, 
    0, 0, 0, 0, 11, 15, 24, 32, 31, 49, 50, 36, 44, 85, 103, 134, 143, 156, 140, 113, 109, 65, 10, 24, 11, 15, 45, 77, 61, 14, 
    0, 0, 0, 0, 16, 21, 32, 42, 33, 39, 42, 29, 82, 127, 125, 134, 125, 117, 105, 109, 76, 16, 0, 21, 7, 19, 75, 100, 73, 4, 
    0, 0, 0, 7, 34, 44, 49, 37, 21, 37, 53, 44, 119, 131, 101, 102, 101, 104, 107, 111, 70, 26, 41, 53, 41, 63, 92, 89, 69, 0, 
    0, 9, 49, 31, 41, 47, 45, 18, 22, 35, 54, 52, 124, 114, 89, 101, 108, 110, 105, 105, 86, 66, 81, 85, 77, 78, 79, 73, 67, 0, 
    0, 64, 77, 43, 41, 49, 43, 10, 25, 26, 41, 45, 112, 97, 90, 104, 104, 73, 51, 53, 68, 70, 82, 93, 88, 84, 79, 73, 46, 0, 
    27, 63, 54, 39, 38, 52, 31, 7, 24, 30, 46, 57, 121, 94, 91, 106, 71, 21, 18, 30, 52, 75, 77, 85, 82, 79, 70, 43, 14, 4, 
    19, 7, 27, 47, 29, 52, 23, 15, 31, 54, 71, 83, 129, 96, 96, 99, 27, 14, 35, 44, 44, 74, 78, 60, 63, 66, 43, 14, 5, 23, 
    0, 0, 49, 80, 34, 45, 20, 24, 40, 69, 69, 76, 119, 94, 106, 85, 9, 39, 40, 31, 30, 52, 77, 58, 63, 59, 22, 12, 26, 35, 
    0, 8, 58, 85, 35, 36, 26, 39, 54, 74, 60, 87, 118, 95, 102, 63, 11, 60, 42, 37, 36, 37, 68, 66, 62, 40, 11, 25, 32, 28, 
    1, 21, 47, 82, 35, 28, 34, 50, 68, 78, 67, 103, 106, 85, 96, 55, 23, 67, 47, 39, 36, 26, 56, 71, 50, 18, 11, 27, 22, 20, 
    6, 24, 41, 79, 46, 38, 63, 84, 101, 107, 100, 121, 111, 100, 108, 65, 30, 67, 60, 50, 40, 33, 40, 66, 34, 6, 16, 24, 20, 23, 
    5, 26, 34, 69, 43, 36, 56, 63, 65, 59, 49, 59, 54, 54, 56, 30, 9, 57, 48, 39, 16, 18, 21, 43, 17, 3, 18, 23, 22, 27, 
    5, 17, 19, 34, 15, 10, 24, 22, 22, 19, 15, 19, 18, 18, 17, 6, 0, 49, 39, 34, 31, 21, 23, 31, 19, 18, 26, 24, 24, 29, 
    9, 11, 14, 25, 21, 31, 37, 36, 37, 35, 34, 33, 32, 29, 26, 22, 17, 45, 38, 35, 30, 17, 18, 26, 24, 25, 28, 29, 32, 35, 
    10, 15, 30, 47, 62, 66, 51, 48, 49, 48, 48, 46, 43, 39, 35, 34, 31, 41, 35, 26, 12, 5, 23, 29, 29, 29, 31, 35, 40, 39, 
    23, 36, 58, 71, 76, 66, 47, 54, 59, 59, 61, 59, 59, 57, 53, 50, 45, 48, 50, 40, 26, 30, 36, 36, 36, 35, 37, 40, 43, 38, 
    
    -- channel=104
    605, 624, 632, 651, 669, 678, 680, 670, 646, 617, 591, 579, 575, 558, 532, 511, 474, 440, 418, 379, 385, 374, 308, 260, 179, 151, 187, 234, 270, 287, 
    660, 650, 630, 628, 625, 623, 611, 594, 570, 544, 519, 510, 508, 497, 476, 458, 428, 398, 382, 372, 368, 348, 293, 222, 129, 110, 170, 241, 284, 298, 
    622, 600, 575, 560, 551, 547, 529, 510, 491, 470, 450, 444, 445, 439, 424, 411, 391, 380, 368, 350, 329, 296, 244, 184, 119, 116, 180, 250, 292, 299, 
    538, 516, 499, 489, 478, 474, 457, 444, 431, 415, 400, 396, 398, 399, 391, 382, 371, 373, 362, 327, 284, 209, 167, 158, 139, 163, 218, 270, 297, 292, 
    453, 435, 427, 425, 415, 410, 401, 396, 390, 380, 370, 368, 373, 379, 379, 374, 367, 370, 353, 316, 247, 142, 108, 134, 164, 216, 260, 296, 306, 295, 
    391, 378, 373, 372, 371, 369, 366, 368, 370, 368, 361, 360, 366, 372, 375, 372, 370, 370, 348, 299, 206, 107, 118, 160, 205, 262, 300, 321, 323, 309, 
    342, 342, 346, 349, 349, 348, 349, 356, 361, 367, 363, 358, 364, 369, 375, 375, 373, 367, 332, 261, 150, 75, 128, 206, 258, 306, 327, 331, 327, 318, 
    323, 332, 341, 345, 347, 346, 348, 354, 359, 365, 365, 363, 363, 361, 368, 368, 360, 350, 300, 209, 107, 58, 127, 220, 287, 325, 334, 328, 322, 313, 
    322, 334, 344, 347, 349, 350, 349, 352, 355, 362, 358, 346, 342, 328, 330, 323, 302, 278, 223, 132, 71, 48, 108, 197, 257, 295, 313, 317, 312, 302, 
    328, 337, 343, 347, 348, 349, 350, 351, 351, 349, 325, 295, 273, 242, 238, 233, 209, 182, 111, 45, 31, 25, 83, 165, 191, 230, 265, 293, 300, 292, 
    340, 342, 343, 346, 345, 346, 348, 343, 325, 303, 273, 240, 205, 164, 165, 175, 174, 169, 119, 68, 39, 0, 21, 117, 157, 171, 201, 246, 280, 281, 
    348, 345, 343, 345, 343, 343, 339, 318, 295, 261, 218, 186, 169, 143, 149, 167, 166, 150, 132, 146, 107, 0, 0, 32, 107, 148, 152, 183, 241, 265, 
    350, 347, 343, 343, 338, 332, 313, 294, 264, 213, 179, 158, 121, 79, 87, 108, 105, 72, 87, 134, 110, 24, 0, 0, 43, 116, 127, 136, 193, 237, 
    348, 347, 344, 337, 313, 297, 270, 250, 195, 158, 137, 122, 78, 32, 36, 70, 74, 49, 80, 93, 66, 45, 0, 0, 3, 66, 92, 98, 140, 194, 
    344, 345, 337, 319, 284, 241, 199, 163, 133, 107, 114, 113, 70, 28, 24, 37, 58, 57, 65, 66, 57, 68, 35, 0, 23, 42, 63, 82, 96, 126, 
    340, 339, 322, 288, 250, 196, 130, 110, 76, 76, 115, 114, 71, 64, 49, 27, 48, 64, 69, 68, 79, 65, 52, 81, 77, 44, 61, 88, 77, 77, 
    334, 326, 291, 238, 172, 137, 99, 81, 54, 59, 88, 84, 86, 131, 105, 79, 92, 93, 86, 80, 66, 37, 36, 76, 86, 47, 52, 78, 80, 68, 
    324, 293, 253, 167, 65, 48, 58, 60, 42, 51, 64, 49, 64, 139, 114, 77, 75, 79, 82, 83, 52, 0, 0, 35, 54, 37, 37, 62, 87, 77, 
    301, 271, 215, 84, 0, 1, 37, 44, 28, 55, 72, 58, 61, 111, 75, 43, 49, 64, 76, 101, 101, 41, 0, 7, 26, 31, 39, 54, 82, 78, 
    286, 275, 172, 42, 0, 0, 30, 37, 33, 55, 59, 59, 73, 99, 53, 35, 56, 46, 53, 113, 155, 132, 67, 21, 18, 25, 39, 62, 68, 75, 
    281, 257, 145, 53, 0, 0, 24, 34, 41, 45, 35, 21, 52, 85, 45, 45, 48, 3, 26, 61, 96, 142, 131, 64, 18, 25, 55, 54, 58, 88, 
    259, 187, 104, 73, 20, 0, 15, 28, 41, 48, 40, 6, 28, 69, 38, 46, 16, 0, 30, 39, 37, 83, 131, 96, 30, 25, 34, 34, 61, 98, 
    234, 133, 45, 49, 30, 0, 6, 28, 39, 46, 44, 24, 55, 64, 35, 36, 0, 0, 40, 43, 42, 46, 94, 103, 44, 13, 4, 22, 74, 113, 
    210, 128, 44, 40, 38, 0, 0, 26, 35, 28, 18, 24, 67, 64, 44, 34, 0, 0, 40, 26, 22, 30, 67, 109, 78, 14, 0, 36, 97, 130, 
    184, 127, 54, 38, 30, 0, 0, 9, 17, 5, 0, 8, 52, 51, 41, 24, 0, 0, 42, 25, 10, 8, 44, 102, 105, 31, 4, 50, 99, 124, 
    166, 121, 65, 41, 37, 0, 0, 15, 28, 30, 18, 25, 53, 55, 54, 34, 0, 0, 57, 42, 13, 4, 32, 86, 108, 48, 27, 57, 85, 103, 
    161, 135, 89, 65, 58, 29, 28, 56, 72, 90, 95, 99, 102, 101, 100, 87, 37, 23, 63, 59, 34, 29, 34, 64, 88, 65, 52, 61, 73, 87, 
    160, 133, 103, 76, 58, 42, 42, 48, 52, 60, 63, 69, 72, 72, 72, 77, 65, 73, 77, 43, 38, 25, 32, 55, 66, 61, 62, 67, 69, 79, 
    151, 114, 70, 37, 17, 9, 1, 0, 5, 9, 8, 14, 20, 25, 27, 37, 44, 64, 91, 70, 42, 33, 43, 59, 61, 59, 63, 67, 71, 79, 
    130, 94, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 13, 21, 29, 42, 50, 41, 33, 46, 54, 55, 53, 55, 60, 67, 74, 
    
    -- channel=105
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 8, 7, 10, 12, 19, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 56, 18, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 50, 57, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 58, 34, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 43, 16, 1, 9, 29, 42, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 58, 49, 70, 45, 1, 9, 6, 0, 0, 0, 0, 0, 0, 26, 30, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 66, 78, 46, 30, 3, 3, 5, 0, 0, 0, 0, 0, 0, 9, 20, 30, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 23, 22, 0, 0, 0, 4, 0, 0, 0, 0, 0, 25, 27, 4, 0, 13, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 7, 0, 0, 0, 0, 0, 38, 51, 19, 17, 23, 14, 0, 0, 0, 7, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 11, 10, 1, 3, 0, 0, 0, 4, 51, 38, 15, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 10, 3, 0, 0, 0, 0, 0, 0, 26, 9, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 12, 0, 0, 0, 0, 8, 22, 15, 0, 20, 11, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 27, 0, 0, 0, 0, 11, 19, 15, 0, 28, 14, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 33, 0, 0, 0, 6, 0, 0, 11, 8, 21, 5, 0, 12, 0, 0, 0, 0, 0, 0, 10, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 27, 0, 0, 4, 14, 3, 13, 7, 0, 9, 0, 10, 12, 0, 15, 4, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 26, 17, 10, 22, 32, 36, 42, 7, 3, 13, 4, 22, 8, 0, 13, 20, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 16, 4, 3, 0, 0, 4, 0, 0, 0, 0, 1, 6, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 18, 22, 12, 3, 7, 11, 10, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 27, 26, 21, 17, 11, 17, 20, 20, 20, 18, 16, 14, 10, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=106
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=107
    0, 0, 0, 4, 12, 11, 11, 10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 1, 0, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 35, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 51, 18, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 13, 8, 13, 33, 58, 89, 58, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 54, 89, 108, 135, 168, 195, 170, 128, 109, 75, 21, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 108, 159, 190, 209, 232, 260, 274, 216, 205, 207, 125, 50, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 107, 172, 213, 217, 199, 182, 180, 163, 153, 267, 322, 196, 79, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 45, 87, 105, 134, 128, 83, 40, 16, 3, 0, 66, 278, 375, 284, 137, 15, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 32, 55, 44, 46, 68, 41, 0, 0, 0, 0, 0, 165, 329, 386, 360, 220, 54, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 39, 44, 43, 30, 35, 56, 25, 0, 0, 54, 103, 197, 322, 377, 398, 402, 254, 55, 0, 0, 0, 0, 16, 9, 
    0, 0, 0, 0, 16, 40, 58, 58, 55, 32, 43, 50, 23, 73, 167, 237, 296, 364, 397, 406, 414, 335, 146, 34, 0, 0, 0, 74, 123, 59, 
    0, 0, 0, 0, 43, 60, 67, 84, 34, 6, 11, 18, 77, 233, 358, 409, 426, 426, 419, 421, 377, 222, 57, 4, 0, 1, 87, 188, 207, 103, 
    0, 0, 11, 69, 51, 28, 44, 44, 0, 0, 0, 0, 120, 306, 401, 416, 402, 405, 415, 412, 326, 187, 91, 68, 101, 142, 197, 236, 249, 129, 
    0, 0, 162, 169, 82, 26, 24, 0, 0, 0, 0, 1, 132, 294, 367, 368, 370, 391, 375, 345, 305, 239, 203, 213, 238, 256, 259, 252, 244, 106, 
    0, 137, 267, 207, 101, 31, 17, 0, 0, 0, 0, 15, 153, 291, 349, 354, 373, 325, 225, 201, 249, 263, 279, 308, 308, 287, 261, 244, 172, 23, 
    34, 192, 226, 178, 103, 45, 7, 0, 0, 0, 0, 35, 184, 298, 341, 358, 330, 165, 43, 34, 98, 192, 260, 302, 295, 263, 243, 173, 42, 0, 
    34, 79, 116, 145, 106, 65, 0, 0, 0, 0, 28, 84, 201, 304, 347, 358, 234, 50, 0, 0, 0, 71, 177, 238, 247, 231, 176, 48, 0, 0, 
    0, 0, 33, 113, 108, 67, 0, 0, 0, 16, 91, 132, 245, 330, 358, 329, 154, 25, 0, 0, 0, 0, 87, 159, 204, 197, 84, 0, 0, 0, 
    0, 0, 29, 113, 118, 61, 0, 0, 0, 54, 101, 163, 279, 337, 355, 293, 131, 32, 0, 0, 0, 0, 29, 118, 184, 149, 21, 0, 0, 0, 
    0, 0, 33, 114, 118, 60, 0, 0, 56, 120, 153, 229, 306, 335, 347, 278, 133, 45, 22, 30, 16, 0, 0, 82, 140, 85, 0, 0, 0, 0, 
    0, 0, 26, 105, 120, 64, 25, 55, 121, 174, 196, 239, 273, 291, 297, 229, 97, 33, 53, 62, 28, 0, 0, 29, 59, 0, 0, 0, 0, 0, 
    0, 0, 17, 76, 89, 45, 31, 57, 106, 146, 165, 181, 191, 195, 194, 143, 37, 2, 42, 74, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 26, 11, 0, 0, 0, 0, 8, 17, 26, 30, 28, 25, 9, 0, 0, 5, 20, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 34, 41, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=108
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 12, 16, 25, 31, 35, 17, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 7, 7, 12, 24, 29, 21, 25, 40, 29, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 30, 33, 25, 22, 34, 32, 26, 52, 65, 44, 21, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 26, 32, 20, 1, 0, 0, 0, 4, 59, 83, 66, 42, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 2, 0, 0, 0, 0, 0, 34, 70, 90, 85, 54, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 1, 17, 28, 43, 66, 84, 95, 95, 48, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 24, 33, 45, 64, 82, 92, 95, 69, 23, 0, 0, 0, 0, 3, 6, 0, 
    0, 0, 0, 0, 7, 4, 5, 8, 0, 0, 0, 0, 0, 28, 63, 80, 88, 92, 96, 97, 93, 62, 11, 0, 0, 0, 16, 29, 28, 5, 
    0, 0, 0, 25, 13, 0, 0, 1, 0, 0, 0, 0, 7, 55, 91, 101, 97, 98, 95, 89, 73, 51, 23, 9, 19, 26, 36, 46, 47, 12, 
    0, 0, 34, 47, 27, 0, 0, 0, 0, 0, 0, 0, 6, 58, 88, 91, 89, 90, 72, 53, 41, 37, 44, 48, 55, 60, 57, 52, 47, 2, 
    0, 16, 47, 53, 33, 0, 0, 0, 0, 0, 0, 0, 18, 60, 83, 84, 90, 71, 42, 39, 41, 34, 55, 75, 75, 63, 52, 47, 21, 0, 
    0, 38, 33, 36, 28, 0, 0, 0, 0, 0, 0, 8, 32, 63, 81, 84, 81, 35, 10, 6, 18, 27, 41, 67, 68, 59, 51, 25, 0, 0, 
    0, 30, 33, 32, 29, 8, 0, 0, 0, 0, 0, 3, 31, 70, 84, 87, 61, 6, 0, 0, 0, 3, 21, 50, 64, 58, 37, 0, 0, 0, 
    0, 0, 6, 15, 23, 11, 0, 0, 0, 0, 11, 20, 49, 74, 82, 78, 40, 0, 0, 0, 0, 0, 0, 23, 48, 48, 13, 0, 0, 0, 
    0, 0, 0, 14, 24, 9, 0, 0, 0, 5, 21, 32, 56, 73, 81, 72, 35, 0, 0, 0, 0, 0, 0, 6, 34, 31, 0, 0, 0, 0, 
    0, 0, 3, 19, 25, 15, 0, 0, 10, 29, 42, 58, 72, 83, 87, 73, 38, 0, 0, 1, 1, 0, 0, 0, 18, 12, 0, 0, 0, 0, 
    0, 0, 4, 18, 23, 7, 0, 0, 6, 13, 19, 30, 41, 47, 49, 37, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 4, 0, 0, 0, 5, 16, 22, 26, 29, 30, 31, 17, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=109
    68, 53, 44, 38, 35, 28, 20, 13, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 34, 34, 24, 20, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 36, 38, 23, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 21, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 31, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 15, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 23, 15, 17, 11, 10, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 27, 36, 48, 35, 26, 18, 17, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 11, 30, 35, 58, 73, 103, 150, 193, 175, 125, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 87, 151, 220, 258, 287, 331, 357, 343, 320, 234, 113, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 103, 174, 224, 252, 241, 221, 207, 181, 184, 281, 338, 278, 76, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 34, 79, 117, 143, 120, 74, 18, 0, 0, 0, 11, 181, 351, 377, 189, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 13, 40, 55, 45, 38, 17, 0, 0, 0, 0, 0, 44, 232, 396, 431, 299, 92, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 22, 21, 31, 4, 9, 17, 0, 0, 0, 0, 0, 80, 225, 368, 454, 451, 341, 189, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 20, 57, 73, 64, 15, 2, 9, 17, 27, 58, 110, 198, 264, 359, 443, 478, 481, 405, 254, 116, 0, 0, 0, 0, 66, 59, 
    0, 0, 0, 0, 0, 11, 51, 44, 10, 0, 0, 0, 27, 168, 336, 461, 490, 514, 512, 502, 439, 300, 108, 0, 0, 0, 4, 100, 207, 156, 
    0, 0, 15, 9, 5, 0, 0, 0, 0, 0, 0, 0, 40, 218, 412, 492, 476, 476, 482, 497, 445, 281, 104, 31, 48, 116, 177, 230, 272, 184, 
    0, 37, 119, 129, 82, 0, 0, 0, 0, 0, 0, 0, 102, 251, 393, 439, 431, 439, 453, 470, 457, 388, 298, 225, 223, 264, 290, 283, 263, 155, 
    11, 135, 260, 278, 148, 6, 0, 0, 0, 0, 0, 0, 103, 252, 383, 419, 414, 375, 310, 252, 276, 349, 395, 377, 349, 333, 309, 280, 210, 80, 
    39, 163, 293, 283, 150, 38, 0, 0, 0, 0, 0, 0, 93, 245, 379, 412, 359, 248, 101, 0, 8, 142, 296, 390, 369, 321, 277, 202, 95, 0, 
    23, 64, 121, 133, 103, 55, 0, 0, 0, 0, 0, 27, 169, 272, 379, 392, 276, 131, 0, 0, 0, 0, 127, 268, 309, 264, 178, 79, 0, 0, 
    0, 0, 0, 44, 75, 59, 0, 0, 0, 0, 0, 103, 236, 318, 409, 378, 216, 56, 0, 0, 0, 0, 17, 143, 238, 210, 103, 0, 0, 0, 
    0, 0, 0, 64, 80, 67, 0, 0, 0, 0, 25, 127, 244, 348, 420, 349, 178, 41, 0, 0, 0, 0, 0, 63, 187, 181, 51, 0, 0, 0, 
    0, 0, 0, 74, 78, 54, 0, 0, 0, 33, 86, 167, 258, 342, 385, 310, 158, 41, 0, 0, 0, 0, 0, 3, 108, 114, 0, 0, 0, 0, 
    0, 0, 0, 64, 85, 72, 13, 0, 81, 183, 248, 304, 339, 373, 391, 319, 172, 53, 0, 38, 24, 0, 0, 0, 2, 7, 0, 0, 0, 0, 
    0, 0, 0, 59, 66, 59, 26, 19, 77, 142, 190, 229, 237, 245, 250, 208, 106, 33, 0, 22, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 24, 50, 64, 53, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=110
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 43, 15, 5, 0, 0, 5, 9, 9, 11, 17, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 13, 0, 1, 25, 13, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    11, 13, 11, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 37, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    16, 11, 4, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 38, 16, 35, 6, 0, 8, 11, 4, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 34, 0, 0, 43, 33, 9, 11, 6, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 1, 0, 0, 5, 19, 1, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 2, 0, 0, 5, 8, 1, 4, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 2, 0, 2, 13, 28, 21, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 5, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 4, 15, 19, 6, 17, 6, 0, 20, 53, 97, 130, 78, 45, 0, 0, 0, 39, 65, 22, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 8, 18, 20, 38, 89, 117, 130, 164, 181, 183, 187, 200, 232, 99, 0, 0, 0, 72, 90, 7, 0, 0, 0, 
    0, 0, 0, 3, 0, 1, 7, 23, 41, 57, 92, 121, 93, 62, 80, 96, 65, 44, 130, 221, 142, 0, 0, 0, 0, 96, 56, 4, 0, 0, 
    0, 0, 0, 8, 0, 0, 9, 43, 46, 37, 50, 60, 10, 0, 0, 20, 0, 0, 74, 140, 112, 49, 0, 0, 0, 31, 51, 27, 0, 0, 
    3, 2, 0, 11, 8, 0, 3, 19, 2, 1, 32, 36, 0, 0, 0, 0, 0, 0, 47, 81, 86, 83, 0, 0, 0, 0, 20, 32, 0, 0, 
    5, 7, 6, 21, 54, 46, 28, 9, 0, 13, 65, 54, 28, 19, 0, 0, 0, 31, 64, 75, 84, 55, 12, 45, 17, 0, 6, 55, 2, 0, 
    6, 11, 14, 6, 34, 72, 66, 53, 10, 25, 65, 46, 100, 172, 106, 76, 107, 116, 102, 94, 50, 0, 0, 27, 18, 0, 0, 69, 51, 0, 
    11, 16, 14, 0, 0, 22, 74, 47, 2, 20, 47, 19, 126, 233, 159, 114, 120, 119, 113, 108, 15, 0, 0, 0, 0, 0, 24, 63, 76, 0, 
    20, 46, 33, 0, 0, 0, 60, 11, 0, 24, 70, 68, 157, 206, 124, 89, 99, 110, 133, 175, 147, 11, 0, 0, 16, 41, 51, 54, 65, 0, 
    54, 137, 100, 0, 0, 0, 37, 0, 0, 21, 59, 89, 186, 194, 104, 87, 102, 92, 122, 202, 267, 230, 116, 48, 45, 58, 63, 60, 44, 0, 
    113, 205, 173, 82, 0, 0, 13, 0, 0, 15, 18, 30, 149, 172, 95, 94, 67, 9, 36, 78, 151, 262, 253, 139, 76, 76, 78, 56, 20, 6, 
    117, 122, 140, 153, 10, 0, 0, 0, 0, 36, 45, 32, 124, 138, 81, 78, 0, 0, 7, 10, 18, 144, 254, 194, 88, 64, 43, 3, 0, 9, 
    72, 13, 45, 129, 29, 0, 0, 0, 8, 63, 88, 88, 150, 124, 81, 47, 0, 0, 20, 9, 0, 44, 178, 192, 92, 31, 0, 0, 0, 12, 
    53, 27, 37, 117, 51, 0, 0, 2, 25, 55, 52, 90, 162, 129, 102, 30, 0, 0, 18, 0, 0, 0, 108, 192, 130, 13, 0, 0, 18, 26, 
    49, 57, 56, 114, 61, 0, 0, 6, 29, 25, 0, 54, 117, 99, 88, 8, 0, 0, 47, 0, 0, 0, 43, 170, 151, 16, 0, 4, 27, 28, 
    38, 56, 58, 101, 69, 0, 0, 42, 80, 91, 73, 97, 124, 122, 126, 54, 0, 0, 78, 43, 0, 0, 7, 120, 134, 28, 0, 10, 20, 23, 
    25, 56, 66, 100, 95, 45, 69, 122, 167, 198, 202, 206, 208, 203, 204, 149, 35, 45, 90, 72, 24, 0, 0, 59, 79, 26, 4, 9, 15, 25, 
    11, 38, 57, 84, 74, 46, 54, 70, 87, 99, 104, 111, 115, 113, 113, 100, 53, 85, 89, 40, 4, 0, 0, 8, 15, 4, 3, 6, 9, 19, 
    15, 8, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 95, 73, 34, 0, 0, 0, 0, 0, 0, 2, 6, 13, 
    25, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 62, 26, 0, 0, 0, 0, 0, 0, 0, 8, 10, 
    
    -- channel=111
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=112
    40, 45, 46, 39, 34, 39, 41, 38, 29, 20, 23, 36, 43, 45, 50, 56, 59, 57, 60, 67, 69, 74, 78, 80, 81, 79, 76, 80, 82, 78, 
    41, 45, 49, 39, 36, 59, 47, 28, 26, 18, 8, 19, 35, 40, 43, 54, 61, 59, 63, 70, 67, 70, 71, 68, 67, 64, 60, 63, 65, 62, 
    42, 43, 49, 39, 39, 75, 49, 11, 27, 28, 13, 11, 23, 29, 34, 51, 57, 54, 55, 59, 54, 52, 50, 48, 46, 44, 46, 52, 56, 60, 
    44, 42, 49, 46, 48, 69, 44, 19, 38, 36, 22, 15, 17, 20, 21, 32, 37, 33, 35, 34, 35, 31, 34, 38, 38, 40, 48, 55, 62, 68, 
    47, 44, 48, 58, 70, 69, 40, 37, 37, 28, 21, 16, 14, 12, 9, 13, 8, 7, 20, 26, 27, 27, 34, 45, 46, 49, 58, 66, 71, 74, 
    47, 45, 49, 67, 90, 83, 44, 32, 32, 24, 22, 21, 16, 3, 0, 9, 4, 0, 14, 25, 25, 29, 40, 53, 56, 59, 64, 66, 68, 69, 
    45, 41, 41, 51, 75, 83, 44, 27, 26, 16, 17, 18, 10, 4, 2, 8, 12, 7, 8, 12, 12, 24, 45, 48, 49, 55, 57, 57, 57, 57, 
    29, 18, 10, 4, 35, 83, 60, 26, 18, 0, 0, 1, 0, 10, 10, 6, 8, 8, 5, 0, 1, 11, 30, 35, 36, 45, 47, 46, 45, 44, 
    0, 0, 0, 0, 36, 111, 70, 30, 27, 0, 0, 0, 0, 17, 16, 3, 5, 6, 3, 0, 0, 0, 13, 24, 25, 34, 37, 36, 36, 38, 
    0, 0, 0, 0, 61, 136, 65, 28, 41, 4, 0, 0, 0, 16, 20, 4, 4, 8, 2, 0, 0, 0, 7, 15, 13, 22, 31, 35, 39, 44, 
    0, 0, 0, 0, 59, 134, 69, 17, 29, 0, 0, 0, 9, 7, 15, 3, 3, 11, 7, 3, 9, 6, 0, 9, 8, 16, 32, 40, 46, 54, 
    0, 0, 0, 0, 39, 109, 94, 26, 12, 0, 0, 0, 12, 5, 8, 0, 0, 15, 12, 6, 14, 14, 0, 0, 14, 17, 33, 47, 58, 68, 
    2, 5, 6, 2, 13, 61, 89, 58, 34, 22, 1, 2, 15, 11, 2, 0, 0, 11, 12, 8, 16, 16, 0, 0, 23, 24, 37, 60, 71, 75, 
    4, 3, 0, 0, 0, 19, 40, 53, 70, 63, 12, 5, 21, 11, 0, 0, 0, 0, 10, 11, 15, 15, 0, 0, 24, 37, 42, 59, 66, 62, 
    0, 0, 0, 0, 0, 21, 7, 18, 64, 63, 0, 0, 22, 12, 0, 0, 0, 0, 8, 14, 15, 11, 9, 0, 16, 38, 36, 44, 47, 48, 
    0, 0, 0, 0, 0, 35, 0, 0, 26, 20, 8, 0, 16, 23, 1, 0, 0, 0, 8, 13, 11, 7, 13, 3, 7, 28, 23, 29, 51, 67, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 31, 14, 0, 30, 15, 0, 0, 0, 3, 6, 5, 5, 13, 8, 1, 23, 31, 47, 78, 93, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 40, 41, 0, 28, 23, 0, 0, 0, 0, 0, 0, 5, 13, 11, 5, 30, 57, 72, 91, 90, 
    0, 0, 0, 0, 0, 0, 20, 24, 0, 0, 34, 57, 0, 9, 22, 0, 0, 0, 0, 0, 0, 5, 14, 14, 13, 39, 72, 77, 81, 80, 
    0, 0, 0, 20, 39, 0, 32, 39, 0, 0, 35, 42, 0, 4, 15, 0, 0, 0, 0, 0, 1, 12, 20, 20, 19, 32, 62, 75, 74, 78, 
    0, 0, 0, 64, 87, 18, 32, 29, 6, 13, 31, 22, 13, 29, 18, 0, 0, 0, 0, 2, 11, 15, 18, 23, 25, 22, 43, 74, 77, 74, 
    0, 0, 8, 75, 69, 8, 23, 47, 38, 34, 24, 9, 17, 57, 48, 13, 12, 11, 6, 7, 9, 7, 14, 28, 33, 24, 29, 66, 84, 74, 
    16, 35, 44, 53, 37, 21, 35, 62, 67, 46, 24, 0, 3, 46, 66, 34, 16, 13, 0, 0, 0, 0, 15, 41, 45, 32, 26, 50, 78, 78, 
    47, 41, 35, 34, 37, 39, 39, 41, 49, 53, 28, 0, 0, 37, 56, 30, 8, 1, 0, 0, 0, 3, 8, 33, 51, 40, 35, 36, 59, 81, 
    35, 33, 35, 38, 36, 29, 23, 29, 42, 49, 44, 23, 19, 30, 39, 30, 8, 0, 0, 0, 0, 10, 10, 19, 40, 49, 44, 36, 41, 74, 
    40, 39, 33, 25, 23, 27, 37, 50, 57, 51, 53, 59, 41, 22, 28, 32, 16, 5, 0, 0, 0, 20, 14, 14, 34, 50, 53, 46, 39, 59, 
    37, 30, 26, 28, 39, 53, 64, 71, 62, 38, 42, 61, 42, 26, 35, 45, 33, 26, 20, 7, 13, 20, 18, 19, 39, 57, 60, 55, 50, 52, 
    34, 39, 47, 55, 64, 73, 75, 72, 52, 28, 38, 56, 42, 36, 55, 61, 54, 48, 47, 37, 26, 23, 25, 35, 56, 67, 62, 61, 63, 59, 
    58, 68, 74, 71, 69, 72, 71, 70, 52, 31, 40, 50, 48, 58, 68, 67, 65, 56, 57, 55, 44, 42, 47, 55, 67, 72, 66, 66, 73, 71, 
    81, 84, 76, 68, 66, 69, 72, 73, 56, 34, 46, 47, 56, 74, 69, 71, 70, 59, 62, 68, 60, 60, 66, 66, 70, 76, 75, 72, 76, 79, 
    
    -- channel=113
    118, 118, 113, 107, 104, 107, 114, 106, 100, 101, 97, 95, 98, 100, 100, 97, 92, 88, 85, 86, 83, 81, 77, 72, 65, 58, 52, 52, 52, 45, 
    120, 120, 115, 108, 102, 105, 113, 99, 92, 90, 90, 88, 86, 88, 89, 88, 88, 83, 81, 80, 72, 68, 65, 60, 56, 50, 45, 44, 42, 36, 
    118, 117, 112, 104, 98, 105, 101, 81, 80, 75, 75, 84, 82, 73, 70, 75, 80, 76, 75, 69, 61, 57, 52, 48, 44, 39, 38, 42, 44, 42, 
    118, 116, 112, 103, 100, 104, 78, 63, 81, 77, 65, 71, 80, 72, 61, 59, 62, 65, 69, 64, 53, 48, 46, 48, 50, 51, 55, 57, 56, 53, 
    114, 114, 111, 102, 97, 95, 69, 58, 75, 63, 49, 43, 47, 49, 47, 51, 51, 51, 61, 68, 67, 63, 64, 67, 68, 67, 69, 67, 64, 59, 
    107, 107, 106, 99, 87, 78, 71, 65, 61, 53, 44, 38, 33, 25, 18, 24, 42, 61, 78, 87, 90, 84, 80, 76, 73, 76, 79, 71, 58, 47, 
    102, 100, 98, 96, 81, 58, 46, 51, 62, 53, 46, 43, 33, 21, 20, 20, 27, 53, 82, 89, 85, 80, 80, 78, 68, 68, 65, 54, 41, 29, 
    96, 96, 97, 95, 78, 58, 35, 35, 52, 46, 38, 36, 31, 28, 28, 28, 27, 29, 49, 68, 75, 80, 73, 62, 55, 53, 48, 39, 31, 22, 
    93, 94, 97, 99, 102, 109, 64, 33, 49, 51, 54, 58, 56, 53, 43, 28, 29, 32, 32, 39, 52, 62, 65, 56, 45, 42, 34, 25, 19, 14, 
    100, 110, 124, 138, 156, 154, 83, 36, 51, 55, 66, 80, 90, 82, 64, 42, 33, 33, 30, 26, 34, 51, 62, 61, 42, 30, 24, 23, 26, 28, 
    137, 149, 162, 171, 184, 155, 78, 43, 53, 44, 54, 78, 98, 100, 78, 55, 44, 40, 30, 25, 27, 41, 52, 49, 40, 30, 30, 34, 38, 41, 
    161, 164, 169, 175, 185, 155, 77, 47, 54, 47, 51, 79, 88, 85, 78, 62, 52, 52, 40, 31, 34, 39, 43, 39, 33, 33, 38, 46, 52, 57, 
    167, 168, 168, 166, 167, 155, 90, 47, 62, 73, 71, 84, 89, 71, 65, 61, 63, 71, 59, 44, 43, 42, 37, 44, 44, 42, 50, 63, 71, 69, 
    165, 162, 157, 152, 150, 149, 113, 47, 40, 69, 77, 77, 90, 74, 55, 56, 69, 85, 74, 59, 51, 43, 36, 48, 59, 57, 60, 69, 69, 61, 
    152, 148, 146, 144, 143, 145, 139, 95, 66, 46, 37, 43, 53, 50, 44, 56, 75, 92, 88, 71, 57, 46, 39, 47, 61, 62, 57, 59, 53, 37, 
    144, 141, 139, 142, 150, 152, 149, 133, 128, 80, 20, 43, 52, 49, 50, 63, 89, 106, 102, 85, 64, 52, 47, 48, 58, 64, 48, 34, 26, 21, 
    142, 145, 151, 157, 165, 155, 127, 124, 124, 117, 84, 85, 72, 62, 55, 66, 88, 105, 104, 89, 70, 59, 57, 53, 57, 62, 47, 30, 24, 19, 
    154, 156, 160, 164, 172, 180, 150, 145, 170, 155, 119, 107, 79, 85, 73, 70, 88, 103, 104, 92, 78, 69, 66, 60, 57, 58, 46, 28, 18, 3, 
    163, 169, 180, 201, 229, 241, 228, 179, 162, 166, 153, 124, 79, 92, 81, 72, 86, 100, 101, 93, 82, 76, 70, 63, 56, 53, 37, 7, 0, 0, 
    202, 222, 241, 256, 265, 246, 253, 216, 149, 142, 160, 141, 75, 80, 83, 68, 78, 92, 91, 84, 80, 78, 73, 64, 53, 41, 19, 0, 0, 0, 
    259, 264, 263, 266, 239, 189, 202, 196, 137, 121, 132, 122, 84, 79, 81, 65, 73, 85, 84, 78, 75, 75, 72, 61, 44, 27, 10, 0, 0, 0, 
    271, 270, 269, 268, 206, 122, 113, 117, 111, 108, 100, 89, 79, 74, 75, 69, 73, 84, 82, 79, 78, 71, 60, 46, 26, 10, 9, 5, 0, 0, 
    270, 270, 268, 252, 188, 123, 119, 109, 92, 87, 72, 64, 66, 66, 50, 54, 76, 85, 82, 77, 74, 72, 65, 50, 28, 2, 1, 12, 2, 0, 
    260, 237, 202, 169, 149, 137, 136, 124, 84, 57, 54, 46, 53, 77, 67, 39, 44, 59, 63, 71, 85, 94, 81, 51, 18, 0, 0, 10, 10, 0, 
    172, 150, 141, 136, 133, 120, 102, 92, 89, 62, 32, 27, 45, 76, 79, 62, 58, 67, 73, 83, 99, 106, 91, 70, 27, 0, 0, 0, 13, 10, 
    120, 122, 122, 112, 97, 85, 81, 79, 83, 77, 55, 45, 57, 64, 65, 63, 60, 69, 77, 92, 116, 121, 99, 78, 52, 13, 0, 0, 1, 19, 
    104, 94, 83, 79, 79, 75, 67, 56, 47, 38, 37, 33, 27, 30, 47, 48, 41, 47, 60, 84, 115, 119, 96, 74, 51, 22, 0, 0, 0, 9, 
    76, 69, 67, 66, 63, 53, 38, 17, 0, 0, 13, 34, 23, 9, 15, 15, 12, 19, 30, 44, 69, 79, 67, 51, 34, 12, 0, 0, 0, 0, 
    64, 57, 50, 39, 27, 12, 0, 0, 0, 0, 8, 27, 18, 9, 0, 0, 0, 0, 0, 2, 9, 20, 25, 22, 11, 0, 0, 0, 0, 0, 
    51, 36, 17, 0, 0, 0, 0, 0, 0, 0, 0, 17, 11, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=114
    36, 35, 36, 32, 29, 26, 30, 24, 15, 6, 5, 9, 17, 24, 26, 26, 25, 24, 20, 24, 25, 24, 25, 23, 22, 19, 16, 12, 15, 11, 
    37, 36, 36, 33, 25, 23, 36, 17, 3, 0, 0, 0, 2, 9, 12, 18, 23, 22, 17, 19, 17, 15, 16, 12, 12, 8, 4, 1, 2, 0, 
    36, 35, 33, 32, 21, 24, 36, 0, 0, 0, 0, 0, 0, 0, 0, 6, 18, 16, 13, 10, 6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 36, 33, 33, 22, 22, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 35, 32, 31, 22, 19, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 2, 0, 
    32, 32, 30, 27, 24, 20, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 3, 0, 0, 2, 3, 4, 8, 4, 0, 0, 
    27, 28, 25, 24, 15, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    22, 21, 16, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 7, 5, 5, 0, 14, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 10, 15, 21, 13, 40, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 26, 30, 35, 27, 41, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 34, 36, 39, 33, 30, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    41, 39, 39, 37, 33, 21, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 37, 34, 30, 24, 14, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    34, 30, 25, 20, 15, 18, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 20, 18, 18, 18, 20, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 21, 21, 17, 11, 0, 14, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 14, 10, 6, 9, 3, 13, 19, 0, 19, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 12, 16, 23, 48, 41, 28, 50, 20, 17, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 42, 44, 45, 83, 64, 44, 61, 25, 7, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    58, 59, 53, 53, 89, 50, 31, 36, 9, 2, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    65, 70, 73, 70, 66, 13, 0, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    86, 93, 92, 72, 46, 17, 9, 12, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    89, 74, 60, 47, 40, 34, 24, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 39, 40, 37, 32, 20, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 29, 25, 16, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=115
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=116
    60, 60, 56, 60, 60, 61, 68, 72, 75, 88, 88, 76, 67, 69, 67, 58, 52, 50, 50, 52, 49, 45, 42, 40, 37, 33, 30, 30, 24, 20, 
    58, 60, 55, 57, 58, 60, 74, 75, 69, 82, 96, 91, 78, 71, 72, 68, 62, 53, 53, 53, 50, 47, 41, 36, 31, 26, 24, 26, 24, 24, 
    59, 59, 56, 53, 61, 65, 56, 65, 82, 89, 102, 113, 108, 92, 86, 77, 66, 55, 52, 46, 43, 39, 34, 34, 35, 35, 36, 39, 39, 40, 
    60, 61, 60, 53, 65, 71, 39, 66, 94, 92, 93, 103, 111, 110, 107, 97, 72, 52, 43, 44, 45, 47, 49, 52, 54, 56, 55, 58, 60, 59, 
    58, 60, 62, 55, 61, 72, 62, 75, 85, 89, 92, 94, 106, 110, 106, 106, 91, 78, 63, 63, 67, 71, 72, 72, 69, 70, 70, 70, 68, 65, 
    57, 56, 59, 58, 55, 51, 60, 73, 84, 94, 97, 102, 105, 106, 107, 107, 103, 111, 105, 89, 81, 80, 89, 88, 74, 67, 66, 64, 61, 59, 
    57, 55, 55, 56, 37, 12, 32, 69, 84, 88, 83, 85, 86, 92, 109, 116, 109, 110, 117, 107, 98, 98, 96, 87, 73, 63, 61, 62, 64, 62, 
    51, 46, 43, 41, 30, 27, 40, 67, 81, 87, 84, 80, 80, 86, 99, 117, 116, 110, 112, 113, 113, 114, 99, 85, 78, 71, 68, 67, 66, 66, 
    42, 43, 49, 55, 69, 76, 56, 65, 75, 92, 102, 98, 98, 99, 98, 111, 117, 116, 113, 116, 119, 122, 118, 101, 91, 81, 76, 76, 76, 78, 
    62, 74, 83, 90, 108, 82, 54, 69, 69, 75, 95, 100, 114, 118, 104, 110, 115, 114, 115, 118, 118, 120, 125, 114, 106, 96, 91, 90, 89, 87, 
    93, 98, 103, 108, 125, 68, 39, 70, 70, 55, 78, 94, 103, 115, 108, 110, 111, 106, 111, 118, 116, 114, 120, 111, 107, 110, 103, 97, 92, 90, 
    104, 107, 109, 109, 123, 77, 25, 62, 86, 75, 89, 109, 96, 106, 112, 109, 110, 106, 105, 112, 118, 111, 116, 111, 105, 112, 107, 99, 93, 89, 
    106, 107, 104, 102, 107, 95, 31, 27, 57, 91, 114, 128, 121, 115, 115, 106, 110, 104, 99, 106, 116, 112, 109, 119, 108, 108, 109, 99, 90, 83, 
    98, 99, 97, 94, 93, 104, 81, 32, 27, 59, 86, 97, 106, 104, 109, 106, 109, 103, 98, 102, 112, 112, 104, 119, 112, 99, 104, 98, 83, 68, 
    91, 90, 90, 90, 95, 107, 125, 100, 73, 33, 30, 67, 85, 91, 105, 114, 119, 114, 108, 107, 110, 110, 105, 111, 114, 94, 92, 82, 68, 63, 
    90, 94, 98, 104, 104, 85, 89, 115, 90, 54, 42, 86, 93, 82, 98, 114, 123, 118, 113, 109, 106, 107, 107, 103, 113, 97, 87, 81, 77, 84, 
    97, 99, 98, 93, 88, 69, 38, 104, 124, 107, 79, 91, 108, 97, 100, 112, 117, 114, 112, 108, 105, 105, 109, 102, 110, 102, 92, 101, 100, 94, 
    85, 82, 84, 93, 112, 131, 73, 96, 155, 139, 122, 81, 119, 121, 104, 113, 113, 111, 111, 109, 108, 106, 109, 103, 106, 107, 97, 101, 90, 73, 
    86, 102, 117, 131, 159, 195, 170, 119, 153, 142, 164, 99, 112, 129, 115, 111, 111, 110, 110, 111, 111, 111, 112, 108, 106, 110, 87, 77, 70, 63, 
    130, 141, 145, 141, 154, 184, 211, 157, 136, 134, 170, 122, 110, 136, 126, 113, 111, 112, 112, 112, 114, 120, 118, 113, 108, 106, 77, 61, 67, 67, 
    151, 150, 155, 161, 120, 109, 130, 115, 114, 133, 148, 130, 115, 125, 123, 117, 116, 118, 119, 120, 121, 118, 109, 103, 97, 98, 88, 67, 67, 71, 
    155, 166, 188, 197, 108, 74, 83, 78, 96, 115, 122, 122, 113, 88, 77, 106, 124, 125, 124, 120, 110, 102, 104, 104, 100, 96, 100, 86, 70, 70, 
    185, 177, 162, 143, 96, 92, 108, 89, 65, 70, 91, 99, 97, 83, 57, 68, 88, 97, 102, 102, 97, 101, 106, 100, 98, 92, 102, 106, 79, 66, 
    145, 121, 103, 99, 102, 98, 98, 88, 62, 47, 51, 61, 83, 106, 79, 60, 76, 86, 93, 96, 91, 96, 108, 107, 89, 87, 96, 109, 96, 71, 
    93, 94, 94, 90, 84, 78, 77, 88, 96, 83, 66, 70, 100, 109, 93, 73, 82, 94, 99, 104, 101, 97, 108, 120, 106, 95, 88, 97, 107, 90, 
    87, 85, 78, 73, 73, 82, 90, 100, 109, 106, 84, 74, 85, 93, 96, 86, 87, 96, 99, 117, 125, 112, 107, 115, 118, 104, 97, 91, 103, 105, 
    72, 70, 71, 81, 92, 102, 105, 103, 93, 83, 84, 75, 72, 77, 94, 98, 93, 96, 93, 110, 127, 119, 107, 101, 108, 108, 102, 91, 92, 102, 
    68, 77, 88, 98, 103, 99, 91, 84, 78, 77, 88, 87, 75, 81, 97, 95, 88, 91, 85, 86, 102, 108, 106, 105, 105, 99, 92, 91, 87, 89, 
    87, 94, 96, 93, 88, 79, 73, 73, 75, 84, 94, 93, 81, 94, 94, 87, 84, 83, 80, 78, 85, 93, 100, 104, 97, 83, 82, 89, 87, 80, 
    91, 85, 79, 75, 76, 79, 76, 75, 74, 85, 94, 93, 90, 90, 85, 89, 85, 83, 86, 83, 79, 80, 84, 87, 85, 79, 78, 83, 85, 77, 
    
    -- channel=117
    0, 0, 0, 0, 0, 0, 3, 5, 5, 7, 3, 0, 0, 3, 6, 3, 1, 3, 0, 2, 5, 4, 6, 6, 4, 3, 1, 0, 2, 0, 
    0, 0, 0, 2, 0, 0, 13, 11, 0, 3, 7, 0, 0, 1, 1, 3, 5, 4, 1, 6, 4, 3, 4, 1, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 2, 0, 0, 22, 2, 0, 2, 7, 12, 10, 3, 0, 0, 5, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 2, 0, 0, 0, 11, 7, 0, 5, 8, 0, 6, 13, 13, 9, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 
    1, 2, 2, 0, 3, 22, 6, 0, 9, 6, 0, 0, 0, 5, 7, 8, 7, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 4, 7, 8, 
    0, 0, 1, 0, 0, 14, 19, 8, 4, 1, 1, 0, 4, 3, 0, 0, 3, 4, 1, 2, 3, 0, 0, 5, 5, 4, 7, 8, 8, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 14, 6, 0, 5, 9, 5, 3, 7, 7, 7, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 5, 7, 9, 4, 2, 0, 2, 4, 3, 4, 4, 
    0, 0, 0, 0, 0, 1, 19, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 4, 1, 0, 4, 5, 3, 1, 0, 
    0, 0, 0, 0, 0, 28, 25, 0, 0, 0, 0, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 1, 4, 6, 6, 4, 2, 1, 2, 2, 
    0, 0, 0, 0, 4, 21, 16, 0, 0, 0, 0, 0, 0, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 6, 5, 5, 5, 
    0, 0, 0, 1, 19, 14, 6, 0, 12, 0, 0, 0, 0, 0, 2, 4, 0, 0, 0, 0, 0, 0, 3, 0, 0, 2, 6, 5, 5, 7, 
    1, 2, 4, 2, 14, 15, 0, 0, 0, 7, 7, 12, 5, 4, 3, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 4, 8, 10, 13, 
    3, 3, 3, 1, 1, 18, 8, 0, 0, 0, 11, 1, 7, 10, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 3, 5, 10, 14, 13, 
    0, 0, 0, 0, 0, 7, 37, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 7, 8, 5, 
    0, 0, 0, 0, 0, 0, 15, 5, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 3, 3, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 8, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 9, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 25, 0, 13, 0, 9, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 25, 26, 
    0, 0, 0, 0, 0, 36, 12, 2, 11, 25, 4, 20, 7, 8, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 14, 15, 11, 
    0, 0, 0, 0, 22, 42, 52, 48, 15, 0, 32, 36, 2, 2, 14, 1, 0, 0, 0, 0, 0, 3, 5, 1, 0, 4, 5, 5, 4, 6, 
    0, 0, 0, 0, 28, 7, 24, 38, 6, 4, 30, 27, 0, 2, 20, 8, 0, 0, 0, 0, 0, 5, 0, 0, 0, 6, 4, 0, 4, 8, 
    1, 6, 16, 49, 51, 0, 0, 0, 1, 17, 17, 9, 0, 0, 12, 9, 9, 7, 3, 3, 7, 1, 0, 0, 0, 6, 10, 3, 6, 8, 
    17, 23, 39, 60, 33, 2, 0, 0, 2, 3, 2, 4, 2, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 5, 5, 8, 12, 8, 5, 
    42, 38, 26, 14, 9, 8, 21, 21, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 18, 13, 3, 
    20, 10, 6, 8, 14, 11, 5, 10, 16, 6, 0, 0, 0, 15, 10, 1, 0, 0, 0, 0, 0, 0, 4, 11, 0, 0, 0, 11, 16, 8, 
    4, 7, 13, 9, 2, 0, 2, 6, 19, 27, 6, 0, 11, 13, 5, 2, 0, 0, 0, 0, 1, 6, 1, 6, 8, 5, 3, 5, 13, 17, 
    8, 5, 1, 0, 3, 7, 14, 18, 24, 23, 9, 1, 0, 0, 2, 11, 6, 0, 0, 4, 16, 16, 7, 1, 2, 10, 14, 7, 8, 19, 
    0, 0, 2, 9, 14, 19, 22, 21, 17, 3, 2, 11, 8, 0, 1, 12, 8, 5, 0, 2, 10, 16, 11, 4, 7, 18, 16, 9, 6, 11, 
    5, 10, 17, 19, 20, 18, 14, 9, 9, 2, 4, 14, 3, 1, 16, 11, 9, 9, 5, 1, 1, 4, 9, 14, 17, 17, 12, 10, 9, 8, 
    19, 21, 21, 17, 13, 10, 11, 8, 8, 2, 5, 13, 1, 13, 14, 11, 14, 9, 6, 7, 5, 0, 7, 13, 12, 11, 10, 10, 11, 8, 
    
    -- channel=118
    7, 9, 9, 11, 12, 10, 11, 18, 18, 22, 27, 19, 16, 18, 18, 16, 16, 18, 22, 24, 27, 27, 28, 31, 31, 31, 29, 27, 24, 22, 
    7, 8, 9, 8, 13, 16, 17, 28, 19, 20, 30, 30, 23, 20, 24, 26, 23, 23, 24, 26, 29, 29, 26, 23, 19, 16, 12, 12, 12, 13, 
    8, 8, 9, 8, 16, 21, 13, 26, 29, 38, 45, 48, 47, 40, 36, 33, 25, 24, 19, 18, 15, 11, 9, 8, 8, 9, 8, 9, 11, 14, 
    11, 11, 12, 12, 18, 21, 19, 28, 40, 47, 51, 51, 53, 56, 54, 47, 27, 11, 0, 1, 3, 3, 7, 8, 10, 12, 11, 15, 20, 25, 
    14, 14, 15, 16, 23, 32, 44, 41, 38, 46, 50, 54, 57, 59, 56, 49, 38, 21, 6, 2, 8, 11, 12, 12, 16, 19, 21, 24, 28, 31, 
    16, 15, 15, 19, 26, 32, 40, 49, 48, 55, 58, 60, 59, 57, 59, 57, 50, 44, 34, 19, 11, 12, 18, 24, 22, 18, 18, 21, 24, 26, 
    15, 14, 11, 6, 1, 0, 16, 47, 49, 50, 45, 39, 42, 45, 51, 62, 58, 51, 46, 37, 28, 28, 24, 21, 20, 15, 15, 19, 24, 25, 
    2, 0, 0, 0, 0, 0, 13, 44, 45, 45, 38, 26, 27, 33, 40, 52, 58, 59, 54, 49, 44, 37, 31, 21, 19, 17, 17, 18, 17, 18, 
    0, 0, 0, 0, 0, 0, 23, 44, 45, 49, 48, 32, 29, 29, 35, 49, 55, 58, 60, 57, 55, 50, 45, 35, 24, 15, 12, 15, 17, 20, 
    0, 0, 0, 0, 0, 0, 17, 45, 42, 39, 41, 35, 32, 41, 37, 45, 52, 51, 56, 60, 59, 56, 55, 44, 33, 23, 17, 18, 19, 20, 
    0, 0, 0, 0, 0, 0, 0, 36, 36, 23, 21, 29, 25, 35, 41, 41, 45, 42, 47, 55, 59, 56, 56, 48, 33, 30, 23, 18, 18, 21, 
    0, 0, 0, 0, 0, 0, 0, 22, 45, 35, 27, 30, 30, 30, 42, 41, 41, 35, 39, 48, 55, 56, 54, 52, 35, 30, 28, 21, 23, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 19, 42, 57, 54, 50, 47, 48, 43, 37, 30, 31, 41, 50, 55, 55, 54, 44, 34, 36, 29, 28, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 41, 44, 33, 40, 44, 40, 32, 24, 26, 34, 45, 53, 57, 53, 52, 38, 39, 37, 30, 23, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 8, 17, 27, 39, 41, 39, 30, 30, 35, 43, 51, 55, 51, 53, 41, 33, 28, 17, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 12, 28, 43, 39, 34, 31, 33, 40, 45, 52, 50, 50, 41, 29, 30, 28, 39, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 16, 24, 42, 39, 32, 30, 31, 36, 41, 48, 50, 48, 46, 39, 48, 52, 52, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 28, 24, 39, 40, 33, 30, 31, 33, 37, 43, 49, 48, 52, 49, 53, 50, 43, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 16, 10, 14, 31, 31, 38, 39, 33, 30, 31, 33, 37, 44, 51, 52, 53, 45, 39, 42, 41, 
    0, 0, 0, 0, 0, 23, 39, 32, 25, 29, 33, 35, 32, 37, 42, 43, 38, 33, 32, 33, 37, 44, 51, 55, 54, 49, 39, 29, 35, 42, 
    0, 0, 0, 0, 0, 8, 13, 17, 39, 51, 52, 50, 49, 46, 51, 55, 45, 41, 41, 43, 44, 44, 44, 45, 47, 43, 39, 30, 29, 41, 
    0, 0, 0, 0, 0, 0, 0, 11, 38, 56, 59, 57, 50, 37, 28, 54, 66, 58, 55, 45, 34, 31, 36, 44, 51, 47, 39, 35, 28, 35, 
    8, 15, 6, 0, 0, 0, 11, 21, 18, 28, 51, 52, 41, 29, 21, 27, 42, 43, 40, 34, 26, 26, 32, 37, 42, 50, 43, 40, 33, 28, 
    12, 4, 1, 6, 12, 13, 5, 1, 2, 2, 13, 27, 35, 31, 29, 27, 33, 37, 33, 27, 16, 13, 26, 37, 34, 40, 46, 40, 39, 30, 
    8, 15, 18, 15, 6, 3, 4, 7, 12, 22, 26, 36, 49, 45, 37, 31, 35, 41, 34, 28, 18, 16, 27, 37, 45, 41, 44, 41, 41, 39, 
    21, 17, 10, 7, 8, 14, 23, 35, 40, 40, 37, 29, 34, 44, 45, 39, 41, 46, 43, 44, 39, 32, 36, 42, 45, 47, 49, 49, 45, 43, 
    11, 11, 13, 19, 29, 39, 47, 51, 46, 37, 30, 27, 28, 36, 40, 48, 53, 56, 55, 54, 53, 46, 41, 42, 46, 51, 53, 54, 48, 44, 
    14, 22, 32, 42, 49, 50, 47, 46, 42, 41, 35, 29, 30, 39, 43, 51, 52, 54, 55, 52, 51, 52, 50, 53, 56, 53, 52, 53, 51, 48, 
    36, 46, 50, 50, 48, 44, 42, 45, 44, 46, 41, 34, 37, 40, 47, 50, 50, 50, 48, 48, 52, 55, 56, 57, 57, 52, 52, 53, 53, 51, 
    52, 50, 47, 47, 46, 50, 49, 47, 45, 48, 43, 35, 42, 39, 47, 53, 52, 52, 52, 50, 49, 51, 49, 49, 52, 52, 52, 53, 54, 52, 
    
    -- channel=119
    75, 72, 72, 72, 72, 63, 64, 67, 79, 91, 95, 88, 78, 70, 65, 65, 63, 64, 59, 57, 55, 50, 49, 48, 47, 47, 47, 45, 48, 48, 
    75, 73, 72, 76, 70, 54, 70, 75, 85, 99, 105, 98, 91, 85, 76, 67, 61, 60, 56, 57, 57, 53, 55, 57, 58, 58, 57, 54, 54, 52, 
    74, 74, 70, 75, 66, 53, 80, 79, 84, 96, 103, 103, 100, 99, 92, 77, 71, 64, 64, 65, 69, 67, 68, 66, 66, 63, 59, 54, 53, 50, 
    73, 73, 69, 72, 64, 60, 80, 77, 86, 101, 110, 113, 112, 112, 109, 97, 93, 82, 78, 77, 76, 74, 70, 68, 67, 62, 56, 50, 47, 43, 
    71, 72, 68, 63, 53, 55, 71, 77, 97, 110, 116, 119, 122, 127, 126, 116, 107, 91, 81, 78, 76, 75, 69, 65, 63, 56, 50, 47, 44, 43, 
    71, 73, 68, 57, 47, 53, 72, 83, 103, 116, 118, 120, 126, 132, 131, 120, 111, 97, 84, 84, 83, 78, 70, 63, 60, 54, 52, 51, 49, 47, 
    73, 77, 75, 73, 63, 60, 81, 91, 118, 133, 132, 132, 135, 131, 129, 123, 119, 112, 101, 94, 91, 85, 77, 72, 61, 52, 51, 52, 52, 52, 
    86, 93, 98, 101, 74, 57, 83, 96, 124, 140, 134, 138, 136, 129, 130, 128, 129, 124, 118, 112, 109, 105, 95, 83, 65, 54, 54, 57, 59, 58, 
    103, 106, 107, 108, 62, 55, 86, 94, 116, 134, 124, 132, 132, 125, 132, 134, 135, 134, 131, 127, 127, 122, 109, 95, 76, 61, 60, 60, 60, 57, 
    102, 101, 102, 104, 57, 60, 92, 92, 108, 132, 125, 125, 130, 124, 133, 139, 139, 138, 140, 138, 137, 135, 122, 107, 85, 65, 60, 59, 59, 57, 
    98, 96, 97, 99, 66, 59, 91, 93, 108, 132, 133, 127, 134, 134, 135, 144, 138, 136, 138, 139, 138, 140, 135, 115, 95, 72, 61, 59, 56, 53, 
    93, 90, 91, 93, 77, 59, 74, 84, 97, 117, 128, 128, 134, 138, 136, 144, 134, 130, 133, 134, 133, 138, 143, 122, 101, 80, 62, 56, 51, 46, 
    89, 87, 88, 91, 87, 72, 72, 81, 81, 91, 107, 112, 121, 133, 136, 144, 135, 131, 132, 132, 130, 136, 144, 127, 103, 88, 64, 53, 49, 46, 
    91, 90, 92, 95, 92, 83, 83, 79, 67, 82, 107, 108, 119, 133, 138, 146, 141, 138, 134, 133, 132, 138, 141, 133, 107, 94, 70, 57, 54, 54, 
    99, 99, 100, 98, 87, 77, 89, 76, 74, 92, 114, 106, 109, 124, 131, 142, 142, 139, 134, 134, 136, 141, 139, 140, 116, 103, 88, 71, 62, 53, 
    105, 102, 102, 103, 99, 87, 124, 111, 97, 108, 92, 102, 97, 112, 128, 138, 144, 141, 136, 138, 140, 143, 139, 143, 126, 112, 100, 73, 50, 34, 
    109, 114, 123, 131, 135, 113, 131, 133, 101, 115, 79, 107, 92, 100, 124, 139, 146, 144, 140, 142, 143, 144, 141, 144, 134, 112, 93, 57, 34, 28, 
    133, 139, 141, 135, 133, 117, 109, 129, 108, 125, 71, 104, 93, 94, 124, 141, 148, 145, 144, 145, 145, 145, 144, 145, 136, 106, 81, 50, 33, 31, 
    139, 135, 126, 99, 102, 97, 79, 111, 112, 122, 74, 99, 104, 101, 126, 143, 147, 147, 146, 145, 144, 141, 143, 143, 134, 104, 75, 49, 31, 28, 
    126, 126, 115, 68, 80, 81, 68, 104, 114, 114, 87, 105, 114, 109, 127, 139, 144, 145, 145, 139, 134, 134, 137, 139, 129, 105, 71, 46, 31, 26, 
    125, 121, 102, 59, 90, 104, 97, 118, 113, 107, 105, 121, 120, 109, 120, 124, 135, 138, 137, 130, 128, 134, 139, 137, 122, 102, 68, 43, 36, 30, 
    105, 89, 73, 60, 96, 109, 101, 105, 108, 109, 122, 136, 128, 102, 102, 105, 115, 127, 132, 130, 132, 136, 132, 122, 106, 90, 67, 44, 40, 36, 
    74, 73, 77, 78, 86, 82, 81, 87, 99, 114, 129, 140, 121, 91, 88, 103, 118, 132, 141, 138, 134, 133, 126, 111, 97, 79, 64, 50, 44, 41, 
    81, 83, 80, 72, 68, 70, 78, 85, 94, 106, 125, 128, 109, 87, 86, 102, 114, 132, 146, 144, 135, 132, 127, 110, 93, 77, 61, 56, 48, 42, 
    77, 73, 73, 72, 74, 74, 75, 69, 68, 73, 80, 88, 90, 96, 97, 107, 117, 131, 148, 144, 131, 129, 128, 117, 96, 78, 62, 57, 53, 43, 
    70, 73, 78, 78, 75, 67, 60, 51, 52, 59, 59, 67, 85, 99, 98, 105, 117, 124, 135, 130, 120, 125, 131, 127, 103, 81, 60, 53, 54, 48, 
    75, 73, 71, 66, 60, 54, 48, 43, 52, 61, 56, 61, 80, 84, 84, 87, 97, 102, 107, 109, 109, 121, 129, 126, 101, 78, 57, 47, 48, 49, 
    68, 59, 52, 49, 49, 48, 46, 42, 51, 56, 54, 60, 73, 65, 64, 64, 71, 76, 79, 87, 93, 102, 103, 98, 82, 67, 51, 40, 39, 43, 
    47, 41, 40, 43, 45, 44, 42, 37, 45, 49, 49, 59, 62, 54, 51, 45, 49, 55, 57, 63, 71, 71, 70, 66, 59, 51, 42, 34, 32, 36, 
    36, 34, 37, 36, 35, 33, 35, 34, 43, 47, 44, 58, 51, 48, 43, 33, 37, 42, 42, 46, 53, 49, 47, 46, 41, 36, 34, 32, 30, 32, 
    
    -- channel=120
    107, 104, 107, 112, 116, 117, 115, 136, 178, 204, 205, 186, 162, 143, 126, 114, 107, 109, 113, 108, 106, 98, 94, 93, 90, 89, 89, 87, 82, 82, 
    107, 105, 107, 113, 121, 121, 127, 163, 198, 228, 242, 224, 204, 191, 173, 146, 121, 116, 119, 119, 119, 112, 108, 107, 102, 99, 97, 94, 91, 92, 
    106, 104, 105, 114, 123, 117, 139, 191, 217, 249, 280, 278, 262, 248, 229, 193, 151, 130, 124, 126, 129, 124, 122, 121, 116, 112, 108, 107, 107, 109, 
    109, 108, 108, 115, 125, 119, 148, 206, 240, 270, 299, 319, 323, 317, 296, 249, 189, 150, 132, 132, 138, 140, 141, 140, 137, 135, 129, 127, 127, 127, 
    113, 113, 112, 115, 125, 134, 162, 217, 257, 288, 310, 330, 345, 357, 353, 314, 251, 195, 159, 152, 156, 164, 165, 157, 149, 143, 136, 137, 141, 141, 
    116, 117, 118, 111, 112, 140, 189, 236, 274, 305, 323, 335, 351, 368, 372, 358, 323, 271, 218, 190, 187, 195, 187, 168, 152, 141, 136, 140, 147, 152, 
    119, 118, 116, 104, 99, 124, 186, 255, 286, 308, 317, 325, 340, 362, 376, 375, 363, 337, 291, 252, 235, 229, 214, 184, 157, 140, 140, 151, 160, 166, 
    118, 118, 115, 109, 107, 109, 174, 258, 289, 302, 298, 298, 314, 334, 361, 385, 383, 368, 348, 323, 306, 285, 250, 209, 178, 158, 162, 174, 184, 192, 
    117, 118, 121, 128, 129, 115, 174, 254, 280, 298, 296, 295, 302, 315, 341, 378, 393, 387, 383, 379, 368, 344, 301, 247, 213, 193, 195, 202, 204, 208, 
    129, 134, 141, 151, 137, 116, 171, 240, 258, 287, 301, 308, 307, 314, 332, 364, 382, 387, 397, 402, 400, 381, 346, 292, 252, 228, 220, 220, 217, 214, 
    148, 152, 155, 158, 128, 98, 150, 221, 234, 265, 294, 305, 311, 324, 331, 347, 359, 362, 383, 398, 399, 385, 361, 323, 286, 258, 236, 223, 212, 201, 
    152, 153, 153, 155, 131, 90, 124, 199, 228, 250, 285, 299, 305, 328, 337, 340, 339, 332, 352, 377, 385, 380, 370, 338, 299, 271, 239, 211, 194, 180, 
    148, 148, 147, 149, 141, 103, 97, 162, 224, 249, 284, 309, 313, 331, 346, 342, 331, 315, 327, 355, 372, 374, 376, 351, 305, 270, 236, 199, 175, 162, 
    147, 147, 146, 150, 154, 139, 106, 121, 165, 207, 259, 298, 313, 334, 350, 346, 332, 308, 313, 338, 361, 372, 377, 359, 313, 269, 234, 193, 166, 157, 
    150, 151, 154, 159, 166, 172, 167, 155, 127, 151, 212, 253, 280, 317, 348, 353, 336, 312, 310, 330, 354, 370, 370, 357, 318, 267, 233, 202, 177, 174, 
    162, 163, 164, 165, 163, 170, 194, 213, 173, 147, 188, 221, 254, 292, 335, 355, 342, 319, 313, 325, 347, 365, 364, 354, 326, 276, 242, 218, 199, 198, 
    164, 166, 163, 160, 149, 133, 171, 222, 211, 186, 198, 212, 256, 276, 321, 347, 338, 318, 312, 323, 340, 356, 358, 352, 333, 294, 258, 236, 214, 209, 
    154, 155, 154, 152, 149, 130, 143, 215, 248, 226, 210, 203, 264, 286, 316, 344, 335, 317, 313, 321, 336, 350, 356, 352, 337, 299, 257, 233, 212, 202, 
    144, 148, 155, 167, 179, 195, 176, 199, 266, 275, 238, 215, 284, 311, 323, 343, 337, 321, 319, 326, 337, 348, 354, 353, 333, 291, 242, 216, 202, 197, 
    149, 156, 165, 168, 187, 251, 247, 232, 279, 302, 285, 263, 305, 327, 327, 340, 341, 330, 326, 331, 341, 351, 356, 351, 326, 282, 230, 205, 199, 197, 
    159, 159, 162, 136, 146, 229, 259, 261, 288, 311, 320, 315, 315, 312, 311, 330, 340, 336, 333, 330, 333, 345, 349, 341, 316, 281, 237, 208, 201, 202, 
    165, 166, 163, 131, 124, 175, 202, 229, 270, 308, 333, 332, 297, 266, 268, 303, 331, 335, 333, 325, 321, 328, 331, 323, 303, 284, 256, 220, 207, 209, 
    167, 165, 163, 148, 135, 156, 166, 174, 218, 266, 304, 310, 279, 219, 208, 259, 303, 318, 322, 310, 301, 302, 312, 312, 297, 287, 271, 239, 214, 211, 
    167, 156, 145, 140, 139, 151, 163, 158, 163, 197, 241, 274, 275, 236, 206, 228, 270, 296, 304, 296, 286, 287, 300, 298, 293, 286, 279, 260, 230, 211, 
    149, 145, 142, 144, 147, 154, 163, 174, 170, 168, 197, 237, 266, 262, 247, 249, 276, 299, 303, 294, 275, 275, 307, 314, 296, 283, 276, 272, 253, 220, 
    148, 150, 153, 158, 164, 176, 188, 198, 201, 199, 201, 223, 254, 269, 266, 266, 285, 303, 305, 301, 282, 278, 305, 326, 314, 288, 274, 271, 267, 236, 
    154, 158, 168, 182, 197, 207, 212, 216, 217, 222, 215, 207, 228, 263, 269, 272, 283, 290, 292, 299, 293, 287, 299, 314, 308, 287, 275, 268, 265, 249, 
    161, 173, 189, 205, 216, 221, 222, 223, 225, 235, 232, 217, 227, 248, 256, 268, 273, 272, 268, 277, 286, 289, 290, 292, 286, 273, 268, 263, 255, 248, 
    179, 190, 203, 217, 224, 224, 221, 225, 233, 245, 241, 232, 241, 248, 252, 257, 257, 258, 253, 254, 266, 277, 277, 274, 267, 259, 260, 257, 245, 237, 
    189, 198, 208, 220, 225, 226, 223, 225, 233, 248, 249, 241, 243, 243, 250, 254, 256, 257, 252, 245, 248, 252, 253, 254, 253, 248, 249, 246, 236, 223, 
    
    -- channel=121
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 7, 13, 23, 15, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 14, 14, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 4, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 22, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 17, 30, 23, 0, 3, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 19, 18, 12, 15, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=122
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=123
    102, 96, 92, 90, 99, 107, 103, 100, 110, 111, 109, 104, 94, 79, 67, 60, 54, 50, 46, 36, 26, 16, 4, 0, 0, 0, 0, 0, 0, 0, 
    102, 95, 90, 88, 98, 99, 82, 85, 104, 114, 114, 108, 97, 85, 73, 60, 47, 44, 38, 29, 18, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    98, 93, 86, 88, 92, 70, 66, 86, 96, 103, 114, 110, 97, 87, 75, 61, 43, 37, 32, 28, 23, 16, 16, 15, 15, 17, 21, 21, 19, 17, 
    95, 93, 84, 88, 81, 47, 64, 83, 82, 83, 94, 104, 102, 91, 76, 59, 49, 49, 53, 51, 52, 50, 53, 54, 54, 56, 56, 50, 41, 31, 
    88, 88, 80, 79, 68, 40, 45, 61, 67, 66, 69, 80, 82, 81, 86, 79, 75, 78, 89, 91, 91, 90, 90, 83, 78, 74, 66, 54, 41, 26, 
    79, 81, 76, 62, 38, 23, 29, 46, 57, 61, 64, 63, 65, 73, 85, 97, 107, 110, 112, 114, 116, 118, 103, 83, 77, 71, 60, 46, 31, 18, 
    73, 75, 73, 53, 25, 16, 23, 37, 52, 60, 67, 66, 73, 86, 91, 93, 103, 119, 119, 118, 120, 116, 100, 80, 69, 61, 51, 39, 27, 18, 
    79, 89, 97, 97, 84, 41, 19, 30, 51, 66, 76, 83, 94, 98, 98, 94, 94, 104, 112, 116, 121, 113, 100, 86, 73, 61, 52, 45, 41, 37, 
    120, 142, 162, 184, 164, 72, 25, 34, 61, 82, 100, 117, 125, 113, 102, 99, 100, 98, 102, 108, 117, 119, 109, 98, 83, 73, 67, 62, 61, 59, 
    188, 210, 231, 250, 193, 89, 34, 34, 58, 87, 115, 146, 147, 123, 111, 106, 104, 103, 100, 103, 113, 121, 118, 108, 94, 88, 86, 84, 81, 77, 
    240, 252, 262, 266, 186, 91, 43, 36, 50, 87, 121, 148, 154, 131, 117, 112, 110, 107, 102, 101, 106, 110, 110, 113, 109, 101, 100, 98, 91, 83, 
    252, 254, 254, 254, 189, 97, 59, 48, 57, 96, 134, 142, 147, 132, 118, 118, 118, 110, 105, 105, 101, 101, 105, 111, 113, 108, 105, 102, 91, 76, 
    241, 238, 235, 233, 204, 120, 72, 66, 85, 101, 125, 138, 132, 120, 114, 127, 128, 121, 115, 111, 101, 95, 109, 112, 113, 109, 103, 95, 77, 56, 
    223, 221, 220, 223, 222, 174, 102, 80, 80, 70, 87, 121, 123, 115, 116, 134, 144, 140, 129, 119, 103, 93, 108, 113, 108, 104, 90, 71, 53, 39, 
    213, 218, 226, 236, 240, 219, 166, 127, 72, 50, 79, 104, 112, 112, 121, 145, 159, 157, 142, 123, 105, 97, 102, 110, 100, 91, 74, 60, 51, 45, 
    225, 233, 243, 250, 241, 227, 218, 199, 162, 116, 123, 120, 119, 125, 129, 152, 166, 166, 149, 128, 113, 106, 100, 108, 99, 87, 75, 69, 60, 44, 
    242, 253, 269, 285, 284, 252, 269, 260, 241, 206, 182, 157, 140, 135, 131, 145, 161, 164, 151, 135, 123, 117, 105, 107, 104, 97, 89, 68, 38, 8, 
    280, 305, 337, 367, 377, 327, 322, 322, 279, 260, 203, 182, 155, 143, 138, 142, 157, 161, 154, 145, 136, 128, 113, 108, 108, 94, 70, 33, 0, 0, 
    361, 390, 421, 443, 436, 392, 329, 305, 270, 286, 209, 175, 160, 148, 138, 143, 155, 159, 157, 154, 148, 136, 119, 107, 101, 72, 36, 0, 0, 0, 
    438, 455, 465, 438, 385, 355, 285, 241, 233, 260, 196, 153, 153, 142, 134, 142, 153, 157, 157, 156, 152, 133, 115, 100, 87, 56, 24, 0, 0, 0, 
    471, 474, 456, 353, 266, 245, 222, 201, 192, 190, 155, 133, 139, 128, 119, 132, 148, 154, 153, 146, 134, 121, 110, 96, 81, 61, 32, 13, 0, 0, 
    466, 449, 396, 262, 190, 174, 166, 160, 138, 120, 109, 110, 109, 103, 101, 106, 124, 133, 133, 128, 124, 123, 112, 91, 68, 62, 49, 27, 5, 0, 
    385, 345, 299, 230, 195, 177, 144, 111, 91, 78, 76, 91, 101, 74, 60, 72, 95, 110, 119, 126, 134, 134, 121, 95, 62, 56, 57, 37, 18, 0, 
    268, 235, 209, 188, 168, 156, 138, 103, 74, 62, 70, 98, 117, 81, 47, 51, 71, 95, 118, 142, 157, 154, 129, 91, 64, 50, 53, 47, 30, 14, 
    176, 164, 152, 143, 135, 129, 129, 121, 93, 63, 64, 86, 95, 90, 77, 75, 84, 105, 135, 165, 173, 164, 144, 106, 69, 45, 43, 51, 44, 24, 
    126, 123, 121, 120, 123, 122, 119, 110, 91, 67, 60, 66, 72, 83, 84, 81, 87, 107, 143, 173, 171, 156, 141, 123, 85, 54, 30, 39, 49, 29, 
    101, 102, 109, 114, 112, 98, 77, 53, 41, 48, 47, 41, 47, 71, 75, 63, 67, 81, 112, 139, 140, 131, 123, 117, 88, 51, 21, 20, 36, 32, 
    96, 96, 92, 82, 67, 47, 25, 7, 9, 36, 53, 44, 48, 53, 43, 33, 35, 38, 53, 75, 88, 94, 94, 86, 58, 27, 8, 3, 13, 23, 
    77, 61, 42, 28, 17, 4, 0, 0, 3, 33, 51, 48, 55, 35, 15, 3, 0, 4, 11, 21, 34, 49, 52, 40, 18, 1, 0, 0, 0, 3, 
    27, 8, 0, 0, 0, 0, 0, 0, 0, 24, 42, 46, 42, 20, 2, 0, 0, 0, 0, 0, 0, 6, 6, 1, 0, 0, 0, 0, 0, 0, 
    
    -- channel=124
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 9, 12, 13, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 21, 26, 30, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 34, 36, 38, 24, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    34, 35, 35, 37, 23, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 32, 33, 33, 25, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 28, 28, 29, 27, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 26, 28, 29, 28, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 25, 28, 32, 34, 35, 17, 12, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 34, 42, 51, 51, 47, 38, 13, 16, 9, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 55, 62, 67, 63, 52, 56, 37, 17, 15, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    65, 69, 78, 84, 70, 56, 45, 32, 13, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    83, 91, 96, 92, 61, 41, 21, 8, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    97, 98, 91, 70, 43, 29, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    90, 82, 66, 39, 23, 8, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    64, 62, 55, 36, 19, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 38, 27, 17, 12, 11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 9, 7, 7, 6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=125
    36, 29, 23, 23, 34, 38, 40, 26, 11, 9, 15, 17, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    34, 28, 20, 22, 25, 9, 6, 0, 0, 0, 0, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 28, 20, 21, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    20, 20, 14, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 24, 25, 29, 28, 26, 26, 25, 24, 13, 0, 0, 
    7, 6, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 53, 58, 53, 53, 47, 39, 29, 21, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 52, 52, 45, 36, 27, 20, 13, 3, 0, 0, 0, 
    0, 3, 12, 23, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 22, 25, 18, 19, 22, 22, 8, 0, 0, 0, 
    37, 62, 92, 125, 104, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 23, 30, 35, 26, 16, 10, 8, 
    134, 167, 196, 220, 162, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 38, 52, 52, 44, 40, 34, 
    217, 236, 248, 256, 176, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 58, 71, 64, 56, 45, 
    245, 250, 249, 244, 183, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 49, 73, 73, 61, 43, 
    236, 235, 229, 221, 189, 107, 3, 0, 0, 0, 1, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 34, 57, 63, 46, 20, 
    209, 209, 209, 208, 201, 165, 95, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 24, 30, 13, 0, 
    188, 195, 206, 217, 219, 204, 184, 123, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    194, 211, 227, 236, 223, 185, 173, 159, 130, 52, 11, 8, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 3, 
    213, 231, 248, 265, 262, 210, 201, 196, 208, 184, 113, 92, 56, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    248, 279, 320, 363, 395, 360, 301, 263, 258, 265, 168, 140, 77, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    352, 401, 447, 481, 504, 483, 401, 305, 233, 267, 191, 155, 74, 47, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    481, 513, 527, 491, 454, 406, 341, 270, 176, 190, 157, 124, 51, 22, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    546, 555, 537, 428, 311, 199, 149, 134, 93, 95, 64, 41, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    547, 542, 500, 371, 236, 110, 52, 32, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    477, 424, 357, 264, 196, 133, 83, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    306, 253, 209, 170, 153, 124, 88, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    155, 136, 125, 114, 103, 91, 78, 66, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    85, 77, 76, 74, 75, 77, 79, 68, 46, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 45, 27, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 46, 53, 61, 67, 60, 43, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 42, 46, 39, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    34, 23, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=126
    22, 18, 19, 27, 37, 39, 32, 24, 19, 10, 0, 0, 7, 18, 17, 11, 9, 12, 10, 9, 13, 10, 7, 5, 4, 5, 7, 0, 0, 0, 
    23, 18, 16, 25, 35, 30, 33, 26, 4, 5, 3, 0, 0, 0, 9, 14, 15, 17, 9, 4, 8, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 18, 11, 23, 30, 3, 23, 30, 0, 0, 16, 3, 0, 0, 0, 0, 12, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 24, 14, 23, 25, 0, 9, 25, 0, 0, 2, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 3, 4, 6, 
    26, 28, 19, 19, 23, 10, 16, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 13, 19, 16, 15, 13, 11, 
    20, 24, 21, 10, 5, 20, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 28, 19, 9, 6, 8, 9, 13, 23, 23, 16, 9, 3, 0, 
    16, 16, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 26, 16, 8, 1, 1, 13, 17, 9, 4, 0, 0, 0, 
    6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 8, 0, 0, 1, 11, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    6, 16, 24, 33, 0, 0, 0, 0, 0, 11, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 12, 5, 0, 0, 0, 0, 
    40, 46, 50, 52, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 22, 10, 7, 7, 7, 
    54, 55, 56, 57, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 29, 22, 15, 14, 15, 
    61, 58, 54, 52, 17, 0, 0, 0, 31, 32, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 34, 23, 18, 15, 
    54, 51, 47, 42, 29, 0, 0, 0, 0, 16, 49, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 32, 22, 11, 4, 
    40, 38, 37, 37, 31, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 7, 0, 0, 
    33, 35, 39, 38, 14, 0, 40, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 10, 
    36, 36, 35, 23, 0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 19, 14, 11, 
    23, 18, 20, 23, 12, 0, 0, 32, 25, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 22, 10, 0, 
    20, 32, 50, 67, 97, 71, 0, 4, 53, 60, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    63, 78, 79, 55, 101, 160, 64, 15, 50, 75, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    89, 92, 75, 0, 9, 92, 54, 20, 34, 41, 11, 0, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    101, 116, 102, 0, 0, 0, 0, 0, 3, 7, 0, 0, 0, 0, 13, 28, 6, 0, 0, 0, 0, 0, 0, 0, 0, 9, 1, 0, 0, 0, 
    125, 124, 106, 46, 16, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 5, 0, 0, 0, 0, 0, 0, 0, 0, 15, 25, 0, 0, 0, 
    104, 79, 64, 59, 54, 48, 23, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 12, 0, 0, 
    57, 53, 51, 47, 40, 29, 24, 11, 0, 0, 0, 6, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 27, 2, 0, 
    45, 43, 34, 24, 20, 23, 31, 38, 35, 19, 2, 3, 14, 6, 0, 0, 0, 0, 22, 35, 0, 0, 0, 0, 0, 0, 0, 20, 25, 0, 
    24, 22, 24, 26, 27, 28, 31, 28, 30, 32, 0, 0, 0, 7, 0, 0, 0, 2, 31, 54, 27, 0, 0, 0, 0, 0, 0, 10, 25, 11, 
    16, 25, 32, 33, 29, 20, 15, 9, 16, 30, 7, 0, 0, 0, 0, 0, 0, 3, 11, 29, 29, 9, 0, 0, 0, 0, 2, 7, 14, 23, 
    28, 31, 30, 24, 13, 0, 0, 0, 19, 36, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 19, 14, 3, 0, 0, 3, 8, 6, 15, 
    31, 21, 14, 10, 5, 0, 0, 0, 15, 35, 18, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 5, 4, 0, 0, 0, 7, 3, 2, 
    
    -- channel=127
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=128
    98, 81, 0, 0, 0, 6, 10, 10, 9, 0, 0, 0, 0, 0, 0, 0, 18, 73, 90, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    97, 92, 0, 0, 0, 19, 8, 0, 2, 12, 0, 0, 0, 0, 0, 0, 0, 49, 95, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    96, 97, 28, 0, 0, 28, 0, 0, 0, 15, 10, 0, 0, 0, 0, 0, 0, 47, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    95, 98, 53, 0, 0, 26, 0, 0, 0, 11, 36, 22, 13, 0, 0, 0, 12, 44, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    95, 97, 72, 0, 0, 1, 0, 0, 0, 2, 52, 57, 36, 15, 8, 13, 36, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    97, 92, 50, 0, 0, 0, 0, 0, 0, 0, 35, 55, 37, 16, 33, 35, 35, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    71, 52, 0, 0, 0, 0, 23, 0, 0, 0, 2, 21, 19, 16, 42, 37, 21, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 9, 44, 0, 0, 0, 0, 0, 3, 24, 52, 31, 18, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 46, 0, 0, 0, 0, 0, 4, 38, 60, 42, 16, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 21, 31, 0, 0, 0, 0, 0, 21, 55, 61, 25, 13, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 9, 0, 0, 0, 0, 0, 34, 58, 40, 0, 6, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 1, 26, 37, 6, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 14, 0, 0, 0, 2, 6, 0, 0, 27, 39, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 19, 39, 0, 0, 4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 53, 0, 0, 0, 0, 0, 0, 2, 4, 10, 14, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 27, 0, 5, 3, 0, 0, 39, 25, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 50, 0, 0, 12, 0, 0, 38, 31, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 43, 3, 0, 0, 0, 0, 25, 16, 18, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 12, 0, 0, 0, 27, 14, 2, 15, 0, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 24, 32, 3, 0, 0, 0, 0, 19, 18, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 3, 27, 41, 10, 0, 0, 0, 0, 13, 24, 16, 12, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 17, 53, 35, 0, 0, 0, 0, 0, 14, 16, 16, 29, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 29, 54, 12, 0, 0, 3, 0, 0, 12, 15, 20, 31, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 54, 15, 0, 0, 0, 0, 0, 4, 38, 43, 1, 0, 1, 10, 0, 0, 14, 19, 23, 21, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 26, 94, 20, 0, 0, 0, 0, 0, 18, 38, 36, 5, 0, 12, 12, 4, 16, 21, 16, 12, 16, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 22, 66, 0, 0, 0, 5, 2, 9, 25, 44, 39, 5, 0, 17, 17, 18, 35, 29, 5, 0, 8, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 14, 0, 0, 7, 12, 10, 22, 32, 53, 36, 0, 2, 19, 15, 26, 41, 24, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 23, 13, 15, 28, 45, 58, 23, 0, 11, 14, 12, 28, 36, 18, 0, 0, 2, 20, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 3, 31, 36, 22, 19, 38, 58, 49, 11, 7, 18, 7, 11, 25, 28, 10, 3, 6, 11, 17, 
    0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 29, 67, 67, 41, 29, 42, 54, 34, 9, 22, 16, 3, 12, 25, 22, 17, 20, 14, 5, 7, 
    
    -- channel=129
    37, 21, 0, 0, 46, 64, 75, 83, 77, 73, 63, 56, 58, 62, 70, 81, 87, 85, 72, 68, 56, 43, 72, 75, 63, 64, 65, 65, 63, 58, 
    37, 26, 0, 0, 49, 82, 94, 107, 108, 100, 94, 89, 88, 89, 92, 105, 115, 111, 85, 52, 33, 59, 105, 100, 87, 85, 83, 80, 75, 69, 
    37, 33, 3, 0, 41, 83, 94, 112, 134, 132, 113, 108, 104, 99, 98, 106, 117, 133, 125, 70, 32, 86, 133, 125, 115, 108, 99, 93, 88, 81, 
    35, 37, 13, 0, 30, 72, 80, 110, 150, 164, 142, 121, 123, 123, 118, 120, 124, 135, 124, 86, 73, 131, 162, 151, 139, 131, 122, 118, 117, 110, 
    34, 34, 21, 0, 22, 65, 74, 106, 158, 187, 172, 134, 114, 107, 115, 130, 132, 137, 123, 95, 114, 169, 184, 179, 176, 168, 162, 156, 148, 141, 
    39, 34, 26, 2, 25, 77, 87, 105, 151, 198, 191, 145, 108, 88, 92, 114, 120, 119, 114, 115, 142, 175, 169, 172, 188, 188, 188, 193, 182, 175, 
    30, 35, 28, 8, 33, 95, 125, 127, 149, 192, 194, 158, 111, 90, 98, 95, 95, 96, 95, 127, 173, 188, 170, 177, 193, 194, 198, 202, 193, 189, 
    62, 27, 11, 33, 98, 150, 149, 130, 146, 184, 190, 178, 146, 122, 118, 101, 81, 93, 96, 127, 179, 184, 171, 199, 218, 217, 225, 206, 185, 189, 
    150, 116, 83, 113, 156, 161, 148, 111, 120, 171, 191, 186, 174, 160, 140, 119, 106, 108, 111, 125, 166, 174, 171, 205, 219, 214, 210, 183, 162, 180, 
    165, 158, 154, 161, 166, 167, 151, 106, 112, 160, 180, 178, 178, 171, 154, 118, 102, 118, 114, 124, 158, 176, 190, 214, 221, 222, 206, 175, 157, 163, 
    170, 163, 160, 166, 174, 172, 142, 110, 131, 164, 177, 176, 173, 166, 144, 115, 108, 123, 114, 128, 154, 166, 193, 225, 233, 231, 214, 182, 164, 160, 
    173, 171, 164, 160, 173, 164, 130, 124, 152, 179, 181, 177, 172, 150, 118, 106, 128, 137, 123, 139, 156, 156, 183, 223, 235, 232, 219, 191, 171, 161, 
    171, 169, 160, 146, 152, 142, 126, 140, 154, 175, 178, 166, 168, 160, 128, 110, 148, 161, 143, 154, 162, 159, 177, 217, 232, 233, 226, 208, 185, 167, 
    176, 166, 152, 137, 127, 104, 113, 156, 151, 140, 136, 148, 164, 153, 139, 148, 161, 162, 158, 153, 147, 151, 174, 200, 220, 229, 232, 232, 204, 178, 
    182, 172, 151, 136, 114, 76, 101, 165, 176, 173, 162, 178, 193, 160, 113, 130, 151, 145, 145, 146, 151, 152, 171, 189, 199, 215, 230, 242, 214, 192, 
    183, 174, 155, 139, 118, 77, 107, 177, 192, 194, 193, 185, 176, 170, 146, 128, 134, 137, 130, 135, 154, 146, 140, 170, 192, 202, 219, 219, 198, 200, 
    190, 172, 150, 134, 129, 97, 105, 177, 199, 179, 174, 182, 174, 166, 171, 132, 97, 121, 128, 108, 128, 132, 82, 68, 127, 179, 203, 194, 173, 189, 
    198, 173, 142, 128, 136, 138, 134, 171, 201, 197, 203, 206, 185, 176, 177, 134, 88, 110, 121, 101, 129, 137, 90, 56, 60, 103, 140, 145, 148, 177, 
    203, 183, 153, 143, 155, 167, 166, 168, 190, 202, 214, 226, 212, 197, 187, 157, 106, 98, 112, 108, 125, 120, 94, 95, 78, 75, 101, 108, 107, 142, 
    203, 193, 175, 169, 175, 177, 184, 179, 172, 177, 192, 199, 196, 205, 190, 168, 142, 103, 104, 130, 127, 99, 89, 100, 90, 93, 113, 114, 101, 101, 
    206, 200, 186, 174, 176, 179, 175, 178, 178, 173, 180, 171, 163, 183, 185, 186, 189, 147, 122, 136, 113, 88, 91, 105, 107, 119, 126, 109, 98, 97, 
    205, 204, 194, 175, 166, 182, 180, 175, 185, 190, 180, 147, 137, 161, 165, 171, 181, 162, 142, 120, 89, 89, 106, 116, 121, 130, 117, 100, 100, 105, 
    201, 203, 198, 174, 160, 185, 199, 192, 186, 183, 171, 135, 130, 152, 156, 155, 157, 153, 138, 99, 72, 95, 118, 119, 120, 128, 115, 105, 100, 90, 
    199, 196, 199, 175, 159, 184, 204, 205, 193, 179, 155, 130, 139, 158, 156, 152, 155, 149, 125, 88, 79, 106, 120, 114, 124, 134, 119, 111, 103, 85, 
    197, 191, 191, 176, 162, 182, 201, 199, 187, 165, 119, 96, 136, 160, 149, 145, 150, 140, 114, 89, 89, 109, 114, 103, 117, 129, 118, 105, 97, 96, 
    195, 187, 180, 170, 165, 178, 198, 196, 183, 141, 62, 52, 125, 153, 138, 132, 132, 121, 108, 85, 86, 105, 107, 103, 108, 109, 103, 96, 96, 95, 
    192, 181, 172, 161, 155, 170, 199, 203, 189, 145, 69, 61, 121, 141, 121, 117, 117, 109, 97, 76, 85, 101, 99, 97, 100, 86, 77, 89, 101, 100, 
    188, 175, 163, 155, 151, 159, 195, 210, 192, 162, 127, 123, 135, 120, 105, 102, 97, 98, 80, 63, 83, 94, 90, 91, 92, 78, 72, 82, 99, 109, 
    182, 167, 158, 151, 146, 153, 189, 209, 194, 172, 160, 153, 128, 100, 90, 93, 94, 88, 63, 65, 87, 90, 90, 95, 89, 76, 73, 85, 100, 109, 
    170, 151, 152, 149, 136, 139, 175, 199, 191, 176, 161, 147, 121, 96, 86, 89, 89, 73, 59, 72, 84, 79, 87, 96, 88, 78, 80, 91, 95, 97, 
    
    -- channel=130
    18, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 13, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 14, 12, 0, 0, 0, 0, 0, 8, 7, 3, 0, 0, 0, 0, 0, 0, 0, 6, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 14, 14, 0, 0, 0, 0, 0, 17, 18, 23, 13, 5, 1, 0, 0, 0, 0, 8, 7, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    12, 13, 14, 0, 0, 0, 0, 0, 17, 27, 35, 27, 15, 8, 0, 3, 3, 12, 9, 1, 0, 16, 19, 9, 6, 5, 0, 0, 0, 0, 
    5, 8, 15, 0, 0, 0, 0, 5, 15, 35, 38, 28, 14, 0, 0, 13, 6, 15, 9, 0, 0, 27, 18, 7, 15, 15, 10, 17, 14, 8, 
    0, 0, 0, 0, 0, 0, 2, 21, 19, 36, 32, 22, 10, 0, 0, 13, 0, 7, 9, 0, 11, 36, 15, 6, 21, 17, 22, 35, 24, 17, 
    0, 0, 0, 0, 0, 0, 14, 30, 19, 31, 33, 27, 14, 7, 7, 15, 1, 6, 14, 7, 14, 31, 11, 18, 31, 25, 34, 36, 20, 15, 
    0, 0, 0, 0, 4, 0, 15, 21, 8, 27, 37, 31, 22, 21, 22, 28, 9, 14, 22, 8, 13, 18, 6, 21, 24, 16, 25, 19, 11, 13, 
    6, 10, 7, 6, 5, 2, 18, 6, 1, 24, 32, 28, 27, 30, 33, 27, 8, 17, 24, 8, 16, 18, 9, 23, 24, 16, 19, 11, 5, 9, 
    6, 9, 12, 7, 7, 8, 12, 0, 5, 26, 35, 31, 31, 31, 32, 18, 4, 22, 22, 9, 20, 20, 9, 26, 30, 22, 17, 12, 3, 7, 
    7, 10, 13, 1, 6, 8, 0, 3, 18, 36, 47, 35, 26, 28, 21, 6, 5, 31, 19, 20, 28, 17, 6, 25, 32, 26, 18, 12, 8, 5, 
    5, 7, 9, 0, 4, 4, 0, 10, 24, 36, 40, 23, 24, 33, 25, 6, 17, 39, 26, 31, 29, 14, 5, 21, 29, 29, 20, 13, 20, 4, 
    8, 6, 7, 0, 0, 0, 0, 8, 13, 16, 18, 18, 31, 40, 33, 10, 20, 34, 30, 18, 20, 15, 5, 14, 23, 27, 22, 25, 32, 9, 
    12, 11, 11, 0, 0, 0, 0, 9, 24, 29, 31, 39, 40, 32, 19, 15, 10, 16, 27, 8, 17, 18, 16, 16, 19, 23, 23, 38, 31, 12, 
    14, 18, 16, 0, 0, 0, 0, 11, 38, 41, 30, 37, 40, 29, 18, 32, 4, 0, 24, 6, 4, 15, 23, 14, 12, 18, 25, 38, 20, 9, 
    12, 23, 18, 3, 0, 0, 0, 13, 33, 30, 20, 32, 37, 29, 22, 28, 2, 0, 16, 0, 0, 0, 0, 0, 0, 10, 19, 25, 8, 2, 
    13, 20, 14, 0, 0, 0, 2, 21, 34, 37, 33, 38, 39, 32, 28, 17, 7, 0, 3, 0, 0, 3, 0, 0, 0, 0, 0, 5, 0, 2, 
    15, 16, 18, 7, 12, 12, 10, 25, 33, 37, 41, 49, 43, 39, 37, 13, 4, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 1, 
    18, 18, 26, 21, 22, 21, 18, 20, 21, 21, 33, 48, 35, 37, 36, 12, 6, 3, 0, 1, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 18, 28, 32, 21, 19, 19, 14, 14, 15, 28, 36, 18, 28, 31, 25, 22, 12, 0, 12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 19, 25, 38, 19, 17, 21, 17, 16, 19, 21, 17, 4, 13, 20, 20, 21, 9, 5, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 18, 20, 38, 19, 22, 29, 26, 19, 19, 18, 4, 0, 7, 11, 10, 10, 5, 8, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    22, 17, 16, 31, 20, 25, 36, 35, 22, 26, 29, 0, 0, 9, 9, 5, 7, 7, 3, 0, 0, 0, 3, 3, 0, 3, 0, 0, 0, 0, 
    20, 15, 14, 22, 22, 25, 34, 34, 21, 29, 22, 0, 0, 10, 7, 1, 5, 4, 0, 0, 0, 0, 2, 0, 0, 7, 1, 0, 0, 0, 
    19, 12, 10, 16, 23, 22, 30, 30, 19, 16, 0, 0, 0, 10, 2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 4, 0, 0, 0, 0, 
    18, 10, 5, 9, 22, 20, 28, 32, 24, 8, 0, 0, 0, 5, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 10, 1, 6, 22, 19, 29, 34, 31, 16, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 11, 0, 3, 25, 22, 29, 36, 33, 21, 8, 6, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 9, 0, 0, 27, 26, 24, 33, 31, 20, 13, 18, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=131
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=132
    18, 9, 32, 114, 141, 142, 138, 120, 106, 123, 139, 139, 136, 134, 133, 133, 123, 85, 43, 65, 76, 96, 131, 139, 144, 144, 147, 150, 149, 148, 
    18, 13, 17, 97, 146, 149, 141, 114, 94, 94, 118, 132, 128, 121, 121, 127, 129, 114, 74, 50, 52, 104, 135, 142, 150, 152, 153, 154, 152, 151, 
    17, 18, 9, 74, 143, 146, 135, 114, 99, 84, 90, 119, 135, 138, 136, 133, 136, 138, 107, 56, 58, 119, 139, 141, 144, 145, 147, 150, 151, 151, 
    17, 18, 6, 52, 134, 139, 120, 120, 110, 98, 80, 99, 124, 140, 150, 148, 148, 145, 112, 61, 77, 136, 155, 154, 148, 145, 143, 141, 142, 140, 
    21, 22, 12, 35, 112, 118, 98, 112, 115, 116, 95, 81, 94, 104, 118, 140, 143, 134, 113, 73, 89, 127, 145, 147, 143, 140, 139, 140, 140, 139, 
    4, 22, 27, 11, 55, 95, 106, 115, 122, 128, 109, 73, 62, 65, 84, 103, 111, 99, 99, 98, 115, 126, 138, 131, 129, 126, 128, 143, 149, 148, 
    0, 0, 0, 0, 61, 121, 123, 124, 135, 129, 119, 95, 63, 65, 79, 68, 80, 75, 81, 117, 136, 130, 136, 142, 141, 142, 150, 156, 160, 155, 
    64, 33, 13, 55, 116, 133, 119, 109, 122, 124, 129, 121, 97, 92, 87, 76, 84, 78, 82, 115, 139, 122, 130, 154, 148, 149, 158, 146, 152, 163, 
    128, 98, 90, 120, 129, 135, 125, 90, 97, 113, 122, 121, 120, 114, 104, 86, 81, 84, 85, 106, 133, 131, 147, 155, 150, 154, 150, 136, 139, 159, 
    138, 123, 127, 133, 137, 146, 122, 88, 96, 106, 113, 116, 123, 123, 114, 79, 75, 78, 78, 98, 118, 138, 163, 159, 157, 166, 146, 137, 139, 148, 
    145, 135, 133, 140, 151, 155, 112, 98, 117, 120, 122, 130, 121, 106, 88, 71, 70, 74, 70, 94, 109, 126, 158, 163, 161, 166, 148, 131, 137, 142, 
    148, 145, 139, 141, 157, 164, 118, 104, 125, 136, 135, 129, 113, 102, 77, 64, 82, 83, 75, 100, 115, 118, 151, 164, 165, 166, 154, 127, 130, 137, 
    148, 147, 141, 139, 146, 154, 134, 110, 101, 98, 90, 93, 98, 94, 98, 94, 102, 90, 100, 102, 97, 118, 151, 162, 166, 169, 163, 142, 133, 131, 
    150, 149, 140, 146, 126, 123, 144, 118, 103, 90, 80, 109, 116, 82, 73, 108, 114, 93, 113, 105, 96, 126, 167, 177, 168, 166, 166, 169, 143, 134, 
    145, 151, 145, 159, 122, 97, 148, 130, 119, 121, 113, 114, 119, 96, 59, 110, 139, 106, 104, 129, 122, 118, 177, 214, 198, 172, 172, 177, 152, 150, 
    140, 144, 144, 158, 132, 77, 127, 141, 123, 110, 101, 92, 98, 102, 92, 93, 133, 129, 101, 130, 121, 103, 110, 154, 191, 196, 196, 176, 160, 163, 
    143, 129, 126, 132, 132, 88, 108, 141, 135, 113, 116, 102, 83, 93, 109, 67, 100, 145, 109, 110, 130, 127, 83, 77, 125, 166, 175, 158, 166, 181, 
    152, 125, 112, 113, 125, 120, 107, 125, 143, 142, 149, 140, 114, 102, 110, 78, 64, 129, 110, 94, 136, 139, 118, 92, 94, 115, 126, 122, 144, 185, 
    154, 132, 116, 126, 130, 133, 133, 123, 127, 133, 140, 153, 144, 128, 117, 96, 54, 91, 101, 108, 137, 126, 127, 118, 91, 98, 117, 117, 123, 144, 
    153, 140, 121, 136, 138, 128, 139, 131, 118, 115, 124, 135, 143, 145, 128, 129, 109, 88, 109, 132, 132, 108, 115, 114, 98, 112, 128, 122, 112, 109, 
    155, 147, 125, 132, 141, 129, 124, 129, 127, 129, 126, 108, 125, 134, 126, 138, 144, 112, 126, 134, 119, 100, 109, 113, 114, 119, 120, 107, 108, 118, 
    153, 154, 133, 123, 135, 138, 129, 128, 133, 143, 130, 100, 111, 122, 121, 126, 131, 124, 132, 116, 100, 105, 113, 118, 119, 115, 109, 100, 107, 112, 
    149, 156, 146, 120, 130, 141, 140, 138, 141, 145, 150, 129, 119, 127, 128, 127, 126, 133, 126, 95, 97, 115, 120, 119, 125, 122, 109, 114, 108, 93, 
    146, 152, 156, 126, 131, 141, 138, 138, 142, 146, 156, 147, 134, 134, 135, 138, 138, 138, 114, 98, 109, 120, 117, 109, 131, 131, 122, 119, 103, 99, 
    146, 149, 154, 136, 141, 147, 135, 129, 139, 129, 101, 118, 137, 139, 140, 140, 141, 131, 113, 105, 111, 118, 114, 107, 121, 129, 129, 110, 104, 102, 
    146, 148, 148, 140, 142, 149, 138, 128, 144, 114, 54, 82, 134, 143, 137, 139, 137, 122, 116, 104, 110, 115, 109, 107, 110, 109, 110, 113, 110, 98, 
    148, 150, 144, 136, 138, 145, 139, 133, 139, 115, 74, 106, 141, 136, 130, 129, 120, 118, 108, 95, 106, 111, 100, 104, 100, 94, 97, 108, 110, 108, 
    152, 153, 141, 130, 134, 142, 140, 138, 130, 120, 116, 135, 132, 125, 123, 118, 112, 116, 92, 91, 108, 109, 102, 102, 97, 91, 89, 99, 115, 119, 
    150, 148, 143, 125, 121, 141, 141, 137, 130, 123, 124, 131, 133, 129, 128, 119, 109, 102, 78, 94, 104, 103, 102, 106, 97, 84, 90, 107, 118, 114, 
    139, 140, 152, 137, 115, 133, 140, 137, 133, 131, 135, 135, 126, 122, 129, 119, 109, 85, 79, 99, 99, 98, 104, 107, 96, 97, 109, 110, 103, 101, 
    
    -- channel=133
    3, 0, 0, 0, 0, 4, 5, 3, 0, 3, 6, 3, 0, 2, 4, 2, 0, 0, 0, 7, 17, 0, 0, 2, 0, 1, 0, 1, 3, 5, 
    4, 0, 0, 0, 0, 12, 15, 9, 0, 0, 1, 1, 1, 0, 0, 0, 11, 6, 0, 10, 0, 0, 0, 0, 0, 1, 1, 2, 3, 3, 
    3, 1, 0, 0, 0, 17, 20, 3, 0, 0, 0, 2, 9, 7, 0, 0, 0, 14, 31, 19, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 
    2, 3, 0, 0, 0, 16, 15, 0, 0, 0, 0, 0, 10, 21, 17, 9, 8, 22, 31, 5, 0, 0, 5, 1, 0, 0, 0, 0, 0, 0, 
    4, 4, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 9, 6, 14, 19, 35, 27, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 
    0, 2, 1, 0, 0, 0, 0, 0, 0, 4, 10, 0, 0, 0, 0, 11, 13, 20, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 
    0, 0, 0, 0, 0, 0, 3, 4, 0, 12, 16, 6, 0, 0, 0, 2, 0, 1, 0, 0, 0, 13, 0, 0, 0, 0, 0, 13, 11, 1, 
    0, 0, 0, 0, 0, 0, 3, 10, 1, 5, 11, 16, 0, 0, 5, 3, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 7, 18, 10, 0, 
    14, 3, 0, 0, 0, 0, 14, 5, 0, 0, 5, 7, 5, 8, 5, 18, 0, 0, 0, 0, 5, 2, 0, 0, 0, 0, 9, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 29, 0, 0, 0, 0, 0, 4, 15, 29, 14, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 6, 2, 0, 0, 
    2, 0, 0, 0, 0, 13, 19, 0, 0, 0, 1, 0, 6, 14, 24, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 1, 0, 0, 7, 29, 7, 0, 0, 8, 16, 18, 12, 14, 6, 0, 0, 4, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 2, 0, 8, 37, 0, 0, 0, 0, 10, 0, 0, 20, 12, 0, 0, 8, 0, 0, 2, 0, 0, 0, 0, 1, 4, 0, 0, 0, 
    1, 0, 1, 0, 9, 25, 0, 9, 0, 0, 0, 0, 0, 0, 6, 0, 3, 2, 7, 0, 0, 0, 0, 0, 0, 1, 0, 5, 12, 0, 
    2, 3, 5, 2, 10, 13, 0, 2, 1, 0, 0, 2, 21, 9, 0, 0, 15, 0, 10, 0, 0, 0, 21, 31, 18, 1, 0, 23, 13, 0, 
    0, 3, 7, 15, 10, 0, 0, 0, 0, 2, 0, 0, 3, 7, 0, 10, 20, 0, 0, 3, 0, 0, 3, 30, 32, 18, 15, 30, 9, 0, 
    0, 0, 1, 7, 15, 0, 0, 2, 12, 0, 0, 0, 0, 0, 1, 3, 2, 2, 16, 2, 0, 15, 0, 0, 0, 14, 29, 30, 10, 0, 
    1, 1, 0, 0, 0, 0, 0, 0, 7, 6, 9, 7, 0, 0, 7, 0, 0, 0, 15, 0, 0, 39, 18, 0, 0, 0, 0, 5, 3, 14, 
    5, 3, 0, 0, 0, 6, 0, 0, 0, 0, 4, 23, 17, 0, 15, 1, 0, 0, 0, 0, 4, 27, 10, 11, 0, 0, 0, 0, 0, 5, 
    1, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 16, 13, 16, 21, 10, 0, 0, 0, 1, 24, 15, 0, 9, 0, 0, 1, 14, 0, 0, 
    1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 9, 0, 4, 5, 6, 20, 3, 0, 24, 29, 0, 0, 0, 0, 0, 13, 12, 2, 0, 
    2, 1, 0, 3, 0, 0, 0, 0, 0, 0, 11, 1, 0, 0, 0, 0, 10, 3, 10, 32, 9, 0, 0, 2, 0, 2, 10, 0, 0, 11, 
    0, 4, 1, 4, 0, 0, 1, 0, 0, 9, 27, 14, 0, 0, 1, 0, 0, 2, 28, 20, 0, 0, 3, 11, 0, 8, 6, 0, 10, 10, 
    0, 1, 8, 6, 0, 0, 0, 3, 0, 7, 48, 28, 0, 1, 4, 4, 4, 18, 26, 6, 0, 0, 8, 4, 2, 16, 7, 16, 13, 1, 
    0, 0, 10, 6, 0, 0, 0, 0, 0, 13, 41, 8, 0, 6, 8, 5, 13, 23, 15, 10, 0, 3, 9, 0, 3, 18, 21, 11, 0, 1, 
    0, 0, 4, 5, 1, 0, 0, 0, 3, 22, 5, 0, 0, 13, 12, 9, 18, 16, 20, 12, 0, 2, 11, 0, 3, 17, 18, 5, 6, 5, 
    3, 2, 5, 4, 0, 0, 0, 0, 17, 28, 0, 0, 0, 18, 8, 11, 15, 10, 25, 4, 0, 7, 5, 0, 11, 8, 1, 4, 4, 2, 
    9, 8, 4, 3, 2, 0, 0, 2, 12, 13, 0, 0, 11, 14, 9, 9, 7, 18, 23, 0, 0, 9, 3, 1, 7, 7, 0, 0, 0, 5, 
    15, 13, 2, 0, 1, 0, 0, 5, 6, 0, 0, 10, 20, 20, 10, 11, 9, 25, 5, 0, 6, 7, 2, 3, 11, 2, 0, 0, 6, 10, 
    19, 10, 9, 3, 0, 0, 0, 5, 9, 5, 0, 15, 29, 25, 23, 18, 17, 19, 0, 0, 8, 3, 0, 11, 10, 0, 0, 9, 7, 5, 
    
    -- channel=134
    34, 34, 27, 33, 18, 2, 3, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    34, 35, 28, 33, 28, 9, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    34, 34, 30, 30, 37, 17, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    34, 32, 31, 28, 40, 24, 7, 0, 0, 0, 0, 0, 8, 14, 15, 9, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    34, 36, 35, 25, 28, 11, 0, 0, 0, 0, 0, 0, 0, 9, 12, 15, 22, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 29, 28, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 10, 31, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 15, 29, 18, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 4, 18, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 6, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 12, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 4, 6, 0, 0, 3, 1, 7, 9, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 7, 13, 7, 3, 1, 6, 6, 6, 6, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 4, 13, 11, 14, 4, 2, 0, 2, 2, 5, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 11, 15, 13, 13, 5, 6, 3, 0, 0, 2, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 5, 16, 18, 13, 13, 10, 13, 9, 7, 5, 2, 0, 0, 0, 0, 5, 7, 2, 
    4, 9, 7, 11, 7, 6, 0, 0, 0, 0, 0, 7, 23, 34, 35, 29, 18, 10, 10, 9, 9, 6, 3, 0, 2, 7, 13, 9, 1, 0, 
    
    -- channel=135
    26, 31, 77, 74, 71, 82, 85, 85, 83, 90, 92, 89, 90, 95, 98, 98, 87, 66, 59, 70, 100, 90, 90, 96, 94, 95, 97, 96, 93, 91, 
    27, 26, 70, 78, 62, 77, 88, 88, 85, 87, 98, 95, 97, 104, 104, 103, 89, 59, 47, 82, 111, 94, 99, 101, 98, 99, 101, 100, 97, 95, 
    27, 25, 59, 80, 55, 71, 92, 88, 86, 83, 91, 87, 84, 92, 96, 96, 83, 57, 55, 100, 115, 103, 112, 112, 110, 107, 106, 103, 97, 95, 
    27, 26, 46, 76, 55, 69, 92, 90, 87, 76, 77, 73, 66, 77, 80, 80, 71, 64, 74, 114, 111, 107, 116, 118, 116, 117, 115, 112, 110, 107, 
    26, 24, 36, 78, 74, 82, 98, 98, 88, 73, 66, 63, 65, 70, 67, 70, 60, 71, 94, 117, 111, 118, 127, 126, 123, 124, 123, 120, 120, 120, 
    36, 30, 57, 103, 104, 96, 98, 102, 86, 77, 73, 71, 78, 73, 60, 69, 61, 75, 102, 108, 98, 120, 133, 127, 128, 127, 119, 121, 124, 127, 
    75, 82, 110, 121, 107, 87, 88, 101, 84, 81, 83, 83, 84, 74, 64, 73, 67, 75, 97, 97, 90, 122, 131, 116, 113, 107, 98, 112, 126, 131, 
    98, 110, 127, 116, 106, 89, 87, 103, 88, 82, 84, 86, 81, 71, 59, 71, 62, 69, 91, 94, 98, 131, 133, 121, 117, 106, 105, 119, 131, 136, 
    113, 122, 124, 117, 114, 88, 92, 108, 93, 87, 89, 87, 76, 63, 57, 69, 66, 67, 90, 91, 104, 134, 135, 133, 130, 117, 122, 132, 137, 142, 
    120, 122, 124, 123, 114, 91, 105, 113, 96, 91, 92, 81, 67, 55, 60, 76, 67, 71, 92, 89, 104, 134, 137, 140, 136, 129, 132, 139, 139, 142, 
    120, 116, 121, 119, 111, 100, 109, 107, 91, 83, 83, 76, 66, 64, 77, 88, 71, 82, 92, 87, 103, 133, 139, 143, 143, 141, 140, 145, 144, 147, 
    124, 118, 123, 108, 104, 108, 99, 95, 79, 71, 79, 75, 69, 74, 89, 89, 73, 88, 86, 82, 103, 128, 136, 141, 145, 147, 146, 143, 152, 158, 
    130, 122, 127, 95, 91, 115, 91, 100, 95, 94, 104, 90, 70, 70, 88, 76, 70, 91, 89, 89, 108, 129, 132, 140, 144, 149, 144, 135, 155, 161, 
    132, 124, 125, 85, 78, 117, 88, 103, 104, 98, 95, 84, 72, 73, 88, 82, 73, 89, 102, 92, 99, 116, 125, 132, 143, 146, 134, 129, 152, 154, 
    129, 121, 116, 81, 63, 105, 87, 94, 96, 95, 86, 83, 84, 78, 65, 77, 78, 76, 101, 88, 79, 81, 96, 111, 126, 135, 123, 132, 152, 148, 
    123, 119, 111, 88, 66, 93, 93, 94, 103, 112, 100, 94, 93, 81, 52, 73, 89, 67, 96, 97, 81, 76, 86, 102, 108, 106, 106, 132, 152, 147, 
    124, 123, 120, 102, 80, 86, 92, 100, 107, 115, 105, 99, 102, 87, 61, 71, 94, 64, 92, 101, 73, 77, 85, 91, 101, 97, 96, 122, 138, 138, 
    131, 130, 132, 113, 94, 92, 93, 101, 104, 104, 98, 98, 97, 87, 79, 74, 92, 81, 94, 94, 67, 79, 75, 77, 95, 96, 93, 106, 114, 121, 
    137, 131, 133, 116, 100, 98, 98, 104, 109, 104, 92, 97, 93, 88, 98, 92, 94, 100, 91, 77, 64, 82, 75, 81, 95, 88, 78, 87, 93, 104, 
    140, 129, 128, 121, 109, 103, 107, 112, 115, 101, 88, 99, 90, 88, 100, 91, 86, 97, 75, 66, 72, 86, 84, 88, 87, 75, 69, 80, 84, 86, 
    140, 127, 120, 125, 116, 109, 114, 114, 114, 96, 88, 105, 95, 92, 97, 89, 84, 84, 60, 70, 83, 88, 85, 88, 80, 72, 75, 77, 71, 65, 
    138, 128, 115, 129, 120, 110, 113, 112, 107, 96, 93, 107, 101, 97, 98, 92, 88, 73, 62, 82, 92, 85, 83, 91, 80, 77, 81, 73, 68, 68, 
    137, 131, 116, 132, 123, 108, 107, 104, 91, 76, 84, 94, 94, 97, 97, 91, 83, 67, 69, 89, 89, 78, 80, 90, 77, 76, 76, 71, 72, 74, 
    136, 132, 122, 133, 127, 110, 104, 100, 69, 48, 72, 83, 86, 94, 93, 84, 75, 67, 72, 86, 81, 76, 79, 84, 71, 71, 71, 73, 72, 68, 
    135, 131, 126, 133, 132, 116, 107, 100, 63, 45, 80, 82, 78, 88, 88, 78, 72, 67, 69, 82, 78, 73, 78, 73, 63, 67, 72, 76, 74, 73, 
    133, 130, 129, 132, 139, 126, 111, 101, 74, 67, 91, 78, 73, 82, 81, 73, 69, 60, 68, 79, 74, 71, 76, 66, 61, 68, 76, 78, 76, 78, 
    129, 127, 127, 131, 144, 132, 114, 103, 92, 86, 85, 67, 69, 80, 77, 71, 67, 56, 75, 78, 73, 73, 76, 65, 63, 71, 77, 80, 78, 73, 
    123, 125, 122, 125, 143, 132, 111, 102, 101, 94, 84, 71, 75, 80, 72, 67, 58, 58, 79, 72, 71, 74, 74, 65, 68, 75, 79, 77, 73, 69, 
    120, 126, 122, 118, 137, 129, 104, 100, 105, 99, 83, 70, 66, 68, 64, 59, 54, 68, 77, 68, 72, 76, 71, 69, 74, 77, 73, 71, 72, 73, 
    116, 119, 118, 107, 123, 124, 97, 93, 98, 87, 66, 54, 52, 56, 56, 52, 57, 72, 71, 66, 75, 75, 69, 71, 69, 67, 65, 74, 78, 77, 
    
    -- channel=136
    56, 82, 178, 283, 302, 289, 259, 228, 239, 272, 294, 296, 293, 291, 287, 260, 212, 158, 137, 152, 197, 249, 266, 287, 306, 311, 316, 319, 317, 319, 
    57, 71, 153, 273, 308, 283, 241, 193, 176, 205, 246, 261, 259, 260, 262, 250, 217, 156, 106, 127, 205, 252, 259, 280, 297, 305, 313, 317, 316, 317, 
    58, 63, 126, 247, 302, 276, 233, 179, 139, 142, 186, 222, 232, 238, 247, 246, 233, 188, 134, 140, 213, 244, 249, 266, 278, 286, 296, 301, 300, 302, 
    59, 58, 102, 214, 289, 273, 239, 186, 134, 113, 131, 178, 214, 235, 250, 246, 232, 192, 155, 166, 220, 238, 247, 255, 257, 258, 266, 271, 271, 274, 
    63, 60, 84, 176, 263, 263, 233, 196, 150, 109, 100, 130, 168, 207, 233, 228, 216, 189, 165, 173, 204, 221, 240, 242, 230, 229, 234, 235, 238, 241, 
    76, 76, 82, 156, 242, 246, 217, 194, 161, 117, 94, 97, 126, 161, 179, 184, 182, 170, 176, 181, 185, 191, 216, 215, 196, 201, 211, 216, 229, 233, 
    80, 87, 114, 169, 215, 229, 215, 196, 171, 131, 113, 97, 108, 131, 132, 141, 151, 150, 175, 195, 191, 192, 221, 206, 184, 197, 204, 219, 242, 243, 
    114, 112, 154, 194, 220, 226, 204, 195, 185, 148, 136, 127, 122, 124, 124, 120, 138, 140, 162, 194, 196, 206, 236, 220, 205, 220, 224, 241, 267, 262, 
    203, 185, 200, 221, 230, 222, 187, 183, 180, 153, 147, 150, 146, 135, 122, 128, 140, 138, 154, 187, 204, 224, 244, 233, 225, 234, 242, 259, 283, 289, 
    231, 224, 227, 233, 237, 221, 192, 186, 171, 147, 144, 151, 150, 140, 124, 123, 133, 127, 144, 174, 203, 240, 258, 241, 238, 245, 251, 268, 288, 303, 
    242, 231, 235, 248, 246, 223, 202, 199, 177, 151, 145, 145, 142, 131, 124, 126, 122, 112, 134, 158, 183, 233, 262, 246, 239, 247, 250, 267, 289, 302, 
    260, 248, 245, 262, 258, 236, 216, 202, 188, 163, 149, 152, 134, 113, 116, 129, 116, 110, 133, 144, 170, 222, 256, 250, 241, 242, 237, 246, 267, 284, 
    267, 258, 252, 258, 251, 253, 230, 180, 167, 153, 148, 147, 129, 118, 124, 136, 126, 127, 137, 142, 174, 219, 256, 255, 249, 244, 236, 226, 239, 267, 
    267, 258, 252, 242, 225, 250, 243, 174, 143, 130, 134, 132, 109, 102, 139, 157, 146, 149, 157, 158, 173, 227, 264, 267, 258, 252, 246, 224, 233, 261, 
    265, 257, 249, 228, 198, 225, 244, 185, 158, 143, 140, 141, 121, 96, 122, 163, 178, 171, 182, 190, 188, 235, 284, 293, 278, 263, 254, 240, 251, 266, 
    259, 254, 249, 227, 182, 197, 230, 186, 150, 148, 142, 123, 125, 124, 116, 160, 215, 199, 187, 212, 200, 199, 262, 315, 310, 285, 263, 258, 279, 281, 
    247, 238, 235, 224, 185, 170, 203, 192, 156, 142, 132, 113, 112, 123, 115, 140, 215, 222, 187, 216, 209, 175, 196, 251, 292, 292, 276, 274, 298, 295, 
    245, 226, 220, 216, 192, 172, 184, 196, 185, 174, 159, 129, 113, 116, 109, 120, 187, 219, 198, 217, 218, 205, 207, 199, 225, 251, 249, 262, 299, 306, 
    249, 228, 218, 214, 197, 188, 185, 190, 194, 194, 185, 167, 148, 127, 120, 120, 144, 191, 207, 204, 207, 220, 232, 205, 203, 219, 218, 224, 258, 292, 
    248, 231, 220, 218, 201, 193, 198, 190, 184, 188, 178, 181, 188, 161, 151, 148, 134, 170, 209, 201, 199, 217, 223, 206, 203, 207, 205, 209, 221, 244, 
    248, 231, 213, 212, 207, 187, 192, 198, 191, 182, 167, 180, 200, 184, 180, 183, 169, 178, 201, 199, 208, 213, 210, 202, 200, 197, 195, 205, 209, 211, 
    250, 238, 214, 207, 214, 189, 178, 186, 194, 186, 166, 176, 199, 189, 183, 187, 187, 192, 189, 198, 219, 214, 201, 198, 199, 186, 189, 197, 196, 197, 
    253, 252, 225, 212, 220, 197, 179, 178, 187, 189, 178, 188, 201, 194, 191, 190, 191, 189, 184, 199, 221, 215, 200, 203, 201, 185, 192, 190, 185, 187, 
    252, 263, 245, 228, 228, 201, 179, 179, 187, 182, 195, 223, 217, 204, 208, 209, 200, 191, 188, 202, 221, 212, 198, 207, 209, 196, 194, 195, 192, 189, 
    253, 268, 267, 255, 244, 212, 178, 177, 173, 157, 189, 243, 232, 212, 221, 223, 211, 199, 193, 207, 221, 209, 196, 202, 205, 201, 201, 199, 194, 190, 
    254, 269, 275, 274, 263, 228, 186, 175, 159, 130, 164, 232, 230, 219, 230, 227, 215, 206, 195, 210, 218, 204, 197, 196, 190, 199, 209, 205, 194, 186, 
    255, 268, 277, 278, 266, 238, 191, 174, 165, 147, 167, 209, 221, 222, 228, 224, 216, 203, 196, 215, 211, 199, 195, 192, 182, 187, 204, 212, 203, 194, 
    256, 266, 276, 274, 263, 240, 190, 170, 174, 178, 189, 205, 212, 221, 224, 214, 206, 193, 198, 213, 204, 198, 194, 188, 179, 187, 202, 209, 207, 199, 
    256, 269, 274, 266, 255, 238, 190, 168, 174, 185, 199, 202, 207, 220, 221, 208, 194, 186, 201, 206, 199, 202, 200, 187, 182, 190, 200, 203, 206, 199, 
    253, 274, 280, 262, 241, 236, 197, 172, 180, 186, 188, 189, 206, 221, 223, 205, 182, 184, 195, 195, 194, 202, 198, 191, 191, 193, 196, 199, 202, 198, 
    
    -- channel=137
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 19, 0, 0, 0, 0, 4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 2, 20, 6, 0, 0, 0, 0, 0, 1, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 18, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 2, 0, 8, 3, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=138
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=139
    0, 0, 47, 145, 213, 221, 206, 197, 206, 214, 211, 214, 214, 217, 222, 218, 185, 134, 104, 78, 133, 223, 257, 261, 258, 257, 259, 256, 250, 244, 
    0, 0, 27, 137, 212, 221, 206, 208, 213, 225, 225, 226, 231, 240, 253, 257, 236, 171, 94, 74, 170, 261, 291, 290, 284, 280, 278, 275, 268, 261, 
    0, 0, 3, 115, 189, 203, 203, 224, 233, 234, 236, 235, 237, 247, 260, 275, 270, 207, 116, 113, 220, 297, 319, 316, 307, 300, 296, 291, 282, 273, 
    0, 0, 0, 86, 155, 179, 206, 239, 265, 258, 242, 227, 225, 236, 252, 265, 255, 199, 144, 182, 277, 326, 338, 334, 328, 320, 317, 314, 305, 296, 
    0, 0, 0, 52, 129, 177, 219, 258, 296, 283, 235, 195, 174, 192, 221, 226, 213, 182, 168, 237, 310, 340, 351, 356, 354, 350, 349, 344, 334, 324, 
    0, 0, 0, 49, 169, 222, 235, 266, 307, 298, 240, 185, 154, 163, 173, 171, 162, 169, 203, 275, 317, 329, 344, 369, 375, 380, 386, 372, 362, 361, 
    14, 0, 12, 137, 238, 258, 249, 262, 292, 305, 271, 214, 189, 177, 148, 143, 139, 160, 227, 296, 321, 333, 365, 387, 394, 397, 381, 363, 363, 382, 
    111, 87, 155, 246, 289, 275, 236, 241, 277, 308, 302, 270, 244, 211, 168, 142, 140, 163, 221, 289, 310, 346, 397, 410, 415, 407, 364, 345, 359, 384, 
    252, 235, 272, 305, 317, 276, 208, 216, 268, 304, 312, 307, 280, 236, 178, 153, 156, 168, 211, 275, 308, 357, 405, 421, 421, 394, 348, 327, 348, 382, 
    313, 311, 319, 331, 331, 274, 213, 226, 270, 300, 310, 309, 279, 225, 159, 150, 162, 170, 208, 263, 312, 367, 412, 434, 433, 397, 354, 326, 333, 368, 
    327, 321, 328, 339, 329, 269, 241, 259, 284, 300, 304, 285, 252, 200, 161, 165, 182, 181, 217, 259, 297, 362, 419, 443, 442, 412, 369, 339, 328, 345, 
    338, 325, 325, 334, 315, 264, 260, 278, 286, 278, 271, 263, 235, 185, 175, 209, 213, 207, 237, 258, 279, 351, 415, 442, 443, 425, 386, 356, 332, 331, 
    341, 325, 319, 312, 282, 258, 264, 268, 264, 253, 259, 269, 247, 211, 201, 236, 239, 239, 243, 257, 291, 350, 408, 439, 446, 439, 414, 377, 348, 353, 
    341, 322, 318, 280, 240, 251, 271, 281, 263, 253, 274, 271, 236, 216, 239, 251, 247, 255, 248, 264, 298, 345, 389, 422, 442, 451, 442, 390, 370, 390, 
    344, 319, 311, 260, 213, 247, 281, 316, 313, 292, 291, 286, 249, 214, 241, 243, 233, 248, 262, 268, 284, 325, 344, 366, 405, 442, 438, 393, 389, 409, 
    340, 310, 296, 259, 208, 253, 297, 323, 324, 315, 304, 289, 274, 255, 228, 226, 228, 231, 250, 255, 263, 252, 269, 311, 356, 393, 384, 370, 392, 416, 
    329, 293, 277, 270, 237, 261, 307, 326, 327, 333, 324, 305, 297, 283, 218, 203, 221, 211, 222, 251, 249, 188, 173, 225, 284, 321, 324, 335, 371, 401, 
    330, 291, 279, 291, 289, 288, 315, 339, 350, 362, 357, 334, 318, 301, 237, 194, 219, 203, 220, 268, 253, 204, 167, 166, 199, 242, 264, 291, 336, 368, 
    350, 314, 307, 313, 321, 323, 316, 329, 345, 358, 366, 351, 336, 315, 275, 227, 230, 223, 243, 260, 226, 208, 195, 178, 194, 226, 231, 234, 266, 315, 
    368, 338, 331, 326, 328, 339, 327, 320, 330, 339, 331, 324, 328, 321, 313, 285, 253, 255, 262, 234, 191, 196, 204, 207, 228, 238, 220, 204, 212, 249, 
    377, 349, 331, 323, 326, 335, 342, 341, 345, 328, 295, 293, 304, 317, 331, 327, 291, 279, 247, 197, 175, 201, 220, 233, 243, 235, 208, 200, 200, 195, 
    382, 355, 325, 317, 332, 345, 353, 360, 365, 330, 283, 280, 291, 306, 314, 316, 305, 277, 211, 172, 188, 217, 231, 240, 246, 229, 207, 200, 186, 160, 
    380, 362, 322, 315, 338, 361, 368, 367, 360, 326, 276, 273, 296, 307, 306, 303, 296, 251, 184, 173, 202, 225, 228, 240, 246, 231, 218, 191, 165, 153, 
    373, 363, 323, 317, 338, 360, 370, 366, 345, 289, 242, 263, 302, 312, 308, 300, 280, 226, 182, 181, 207, 218, 217, 239, 242, 230, 211, 188, 176, 166, 
    365, 355, 325, 317, 332, 351, 360, 355, 305, 215, 196, 252, 297, 303, 292, 282, 253, 211, 178, 180, 201, 206, 201, 217, 219, 205, 188, 189, 183, 170, 
    358, 341, 317, 308, 326, 347, 357, 349, 271, 173, 185, 258, 284, 276, 266, 247, 221, 192, 159, 168, 190, 191, 190, 189, 178, 171, 177, 185, 183, 176, 
    348, 326, 303, 291, 312, 345, 363, 350, 288, 220, 232, 262, 258, 244, 232, 215, 197, 161, 137, 161, 180, 176, 180, 169, 150, 145, 165, 189, 201, 197, 
    330, 308, 290, 277, 295, 335, 360, 349, 316, 288, 282, 263, 237, 218, 205, 189, 169, 125, 126, 156, 168, 168, 172, 162, 142, 140, 165, 195, 204, 196, 
    302, 292, 278, 263, 280, 314, 345, 346, 326, 312, 295, 254, 207, 188, 179, 167, 139, 107, 131, 151, 159, 166, 175, 160, 144, 154, 174, 185, 187, 181, 
    268, 274, 266, 242, 252, 284, 322, 335, 326, 309, 272, 212, 164, 149, 143, 138, 110, 110, 135, 141, 148, 165, 172, 162, 159, 162, 160, 164, 176, 182, 
    
    -- channel=140
    0, 0, 0, 0, 1, 11, 14, 15, 12, 4, 0, 4, 4, 7, 11, 14, 17, 19, 12, 0, 0, 10, 15, 15, 14, 14, 12, 11, 10, 8, 
    0, 0, 0, 0, 1, 14, 20, 29, 26, 23, 13, 14, 17, 20, 24, 26, 24, 17, 4, 0, 1, 22, 27, 25, 22, 21, 19, 17, 16, 14, 
    0, 0, 0, 0, 0, 11, 19, 35, 38, 36, 27, 17, 14, 16, 22, 27, 29, 23, 5, 0, 12, 30, 37, 36, 32, 30, 27, 24, 22, 19, 
    0, 0, 0, 0, 0, 5, 20, 37, 49, 48, 39, 25, 18, 15, 18, 23, 24, 17, 10, 13, 28, 35, 37, 38, 38, 36, 36, 37, 35, 33, 
    0, 0, 0, 0, 0, 5, 24, 40, 57, 55, 44, 28, 15, 16, 21, 18, 20, 15, 13, 32, 47, 48, 50, 52, 52, 51, 50, 47, 44, 42, 
    0, 0, 0, 0, 2, 14, 23, 39, 57, 58, 47, 33, 18, 16, 19, 15, 15, 16, 19, 38, 48, 46, 53, 65, 68, 70, 67, 56, 51, 52, 
    0, 0, 0, 0, 12, 21, 27, 32, 48, 58, 50, 35, 27, 22, 16, 14, 11, 15, 25, 42, 49, 48, 56, 63, 68, 68, 60, 51, 49, 58, 
    0, 0, 0, 17, 28, 31, 28, 31, 44, 55, 53, 43, 37, 30, 20, 6, 8, 14, 25, 42, 45, 52, 65, 68, 73, 71, 54, 44, 43, 50, 
    21, 14, 23, 35, 38, 31, 19, 27, 44, 56, 57, 54, 45, 36, 22, 15, 15, 18, 24, 39, 39, 47, 63, 69, 68, 62, 45, 34, 38, 45, 
    41, 40, 40, 42, 41, 30, 19, 26, 44, 55, 56, 55, 46, 34, 18, 15, 20, 21, 26, 38, 42, 48, 63, 69, 67, 58, 44, 30, 30, 37, 
    40, 41, 41, 41, 39, 28, 26, 31, 42, 50, 50, 47, 43, 34, 22, 20, 28, 24, 32, 40, 41, 51, 66, 72, 71, 63, 49, 36, 29, 31, 
    39, 38, 37, 41, 32, 21, 33, 39, 42, 41, 41, 43, 37, 25, 25, 33, 33, 29, 37, 38, 35, 50, 66, 72, 72, 67, 56, 47, 33, 31, 
    39, 37, 35, 38, 27, 17, 36, 44, 50, 50, 48, 51, 46, 31, 19, 35, 40, 34, 35, 44, 43, 47, 62, 71, 73, 70, 64, 57, 43, 41, 
    38, 36, 34, 32, 25, 19, 39, 46, 41, 41, 44, 41, 42, 44, 39, 35, 42, 40, 30, 40, 42, 40, 48, 63, 72, 73, 71, 58, 50, 53, 
    40, 32, 31, 25, 23, 23, 40, 57, 52, 44, 50, 52, 41, 34, 39, 24, 26, 37, 29, 31, 39, 39, 26, 34, 55, 69, 69, 56, 51, 57, 
    42, 31, 28, 24, 23, 39, 48, 60, 63, 63, 62, 58, 51, 42, 35, 26, 17, 28, 29, 30, 40, 35, 34, 31, 35, 47, 49, 46, 48, 58, 
    42, 32, 28, 31, 28, 42, 55, 55, 56, 59, 60, 63, 60, 53, 36, 26, 13, 17, 23, 25, 27, 11, 12, 26, 31, 38, 39, 35, 38, 50, 
    40, 32, 29, 37, 39, 44, 58, 57, 56, 60, 61, 60, 61, 58, 38, 27, 23, 13, 25, 33, 26, 9, 1, 6, 14, 26, 32, 33, 34, 36, 
    45, 36, 34, 40, 47, 48, 51, 57, 60, 63, 67, 60, 60, 59, 49, 37, 35, 24, 29, 30, 20, 11, 11, 11, 15, 20, 21, 20, 27, 35, 
    50, 45, 44, 43, 48, 55, 52, 50, 55, 60, 57, 52, 54, 54, 51, 41, 33, 32, 31, 23, 12, 13, 16, 19, 23, 23, 20, 16, 18, 25, 
    52, 49, 47, 43, 46, 55, 58, 55, 55, 54, 48, 45, 46, 52, 57, 53, 41, 37, 28, 13, 8, 15, 21, 24, 29, 28, 21, 17, 14, 10, 
    52, 48, 47, 41, 47, 56, 60, 62, 64, 55, 43, 43, 44, 47, 53, 55, 47, 38, 20, 9, 11, 19, 24, 26, 32, 28, 21, 18, 14, 8, 
    51, 46, 42, 40, 47, 61, 64, 63, 62, 51, 31, 37, 44, 43, 47, 46, 43, 31, 14, 7, 12, 20, 23, 24, 28, 26, 22, 13, 10, 7, 
    49, 44, 36, 37, 45, 61, 67, 64, 60, 41, 20, 32, 45, 43, 42, 42, 37, 25, 12, 6, 14, 20, 22, 26, 25, 23, 19, 14, 10, 5, 
    46, 41, 33, 31, 39, 56, 64, 62, 54, 33, 20, 33, 44, 40, 36, 36, 29, 20, 10, 7, 14, 17, 16, 22, 21, 15, 12, 14, 13, 12, 
    43, 36, 28, 26, 35, 50, 59, 59, 42, 20, 21, 38, 39, 32, 29, 25, 20, 15, 2, 4, 11, 13, 14, 15, 13, 10, 8, 10, 13, 12, 
    40, 33, 25, 21, 31, 49, 59, 60, 43, 21, 23, 32, 31, 24, 21, 19, 15, 6, 0, 4, 9, 11, 12, 11, 6, 2, 6, 12, 15, 14, 
    34, 27, 22, 19, 27, 45, 60, 61, 50, 37, 35, 34, 26, 17, 15, 12, 8, 0, 0, 2, 5, 6, 9, 8, 3, 1, 6, 12, 14, 15, 
    27, 23, 18, 19, 26, 37, 56, 61, 52, 47, 43, 28, 11, 5, 6, 8, 3, 0, 0, 1, 4, 6, 10, 6, 4, 5, 7, 9, 11, 13, 
    17, 15, 9, 11, 21, 27, 47, 57, 51, 44, 34, 18, 3, 0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 6, 5, 2, 3, 6, 11, 12, 
    
    -- channel=141
    0, 0, 0, 73, 191, 227, 212, 209, 199, 190, 196, 210, 217, 217, 223, 242, 243, 187, 96, 46, 113, 219, 297, 306, 295, 291, 286, 281, 277, 268, 
    0, 0, 0, 44, 155, 210, 211, 230, 245, 222, 209, 219, 245, 257, 264, 277, 278, 237, 154, 108, 164, 266, 333, 328, 315, 307, 301, 297, 294, 288, 
    0, 0, 0, 13, 109, 178, 203, 251, 298, 278, 237, 210, 225, 253, 273, 291, 284, 236, 168, 164, 227, 317, 365, 358, 346, 335, 326, 318, 312, 303, 
    0, 0, 0, 0, 65, 150, 194, 260, 332, 328, 270, 195, 160, 177, 206, 238, 235, 211, 182, 213, 262, 324, 353, 364, 366, 366, 363, 358, 350, 338, 
    0, 0, 0, 0, 58, 163, 222, 276, 343, 359, 296, 200, 137, 125, 134, 159, 154, 163, 197, 269, 312, 337, 346, 367, 385, 391, 392, 393, 388, 383, 
    0, 0, 0, 26, 139, 223, 251, 284, 337, 371, 333, 258, 191, 153, 128, 121, 110, 142, 205, 295, 341, 362, 378, 415, 444, 440, 421, 405, 392, 402, 
    93, 37, 63, 160, 255, 260, 229, 246, 300, 362, 361, 329, 280, 227, 177, 146, 130, 155, 215, 289, 333, 368, 395, 446, 472, 448, 406, 370, 365, 399, 
    254, 226, 235, 282, 309, 267, 215, 210, 255, 335, 359, 351, 327, 277, 200, 168, 143, 164, 215, 272, 326, 380, 414, 457, 470, 427, 367, 320, 321, 375, 
    297, 297, 311, 325, 325, 272, 223, 217, 261, 327, 350, 348, 323, 269, 200, 157, 143, 160, 205, 253, 312, 379, 428, 465, 468, 420, 352, 299, 292, 336, 
    325, 320, 323, 335, 332, 279, 240, 248, 298, 344, 355, 337, 295, 226, 170, 160, 160, 175, 210, 249, 299, 359, 415, 467, 467, 421, 355, 297, 273, 295, 
    332, 326, 323, 323, 318, 285, 261, 267, 302, 328, 331, 315, 276, 217, 179, 192, 204, 222, 235, 263, 300, 349, 405, 461, 469, 436, 378, 316, 272, 274, 
    327, 315, 316, 294, 281, 274, 268, 271, 254, 253, 270, 270, 262, 240, 232, 249, 256, 261, 255, 270, 294, 347, 408, 454, 469, 458, 424, 363, 311, 299, 
    326, 309, 313, 277, 248, 252, 272, 314, 282, 267, 281, 293, 273, 231, 240, 267, 276, 268, 267, 281, 301, 355, 409, 452, 466, 472, 458, 410, 366, 344, 
    324, 307, 317, 285, 245, 253, 281, 352, 342, 329, 321, 315, 296, 264, 245, 261, 275, 264, 268, 284, 310, 326, 372, 427, 460, 473, 458, 426, 396, 386, 
    313, 288, 299, 290, 257, 268, 289, 362, 354, 339, 323, 304, 292, 292, 260, 243, 243, 248, 255, 257, 272, 234, 228, 290, 383, 442, 430, 402, 392, 402, 
    304, 263, 258, 279, 287, 299, 308, 364, 386, 377, 357, 343, 316, 300, 260, 213, 200, 218, 250, 245, 259, 226, 147, 140, 226, 314, 338, 344, 366, 401, 
    313, 265, 252, 283, 321, 346, 338, 358, 393, 423, 427, 410, 379, 340, 277, 211, 184, 180, 236, 248, 256, 246, 187, 146, 153, 197, 229, 261, 307, 369, 
    331, 294, 288, 312, 353, 373, 361, 351, 360, 390, 410, 423, 417, 378, 326, 256, 208, 187, 235, 261, 243, 227, 193, 186, 183, 193, 214, 221, 232, 284, 
    350, 318, 313, 328, 357, 368, 364, 355, 347, 352, 355, 370, 383, 389, 376, 337, 298, 257, 250, 261, 219, 199, 190, 208, 224, 233, 229, 215, 200, 212, 
    367, 338, 319, 321, 348, 365, 361, 365, 373, 357, 327, 315, 322, 353, 371, 368, 353, 318, 260, 228, 191, 188, 207, 235, 252, 247, 221, 200, 191, 189, 
    374, 350, 321, 315, 339, 381, 390, 386, 391, 373, 326, 297, 297, 327, 346, 346, 338, 313, 239, 187, 169, 199, 230, 253, 261, 245, 217, 190, 174, 155, 
    371, 354, 320, 314, 333, 391, 420, 420, 406, 381, 343, 321, 315, 332, 345, 340, 328, 283, 214, 168, 173, 213, 239, 261, 264, 258, 229, 196, 170, 138, 
    361, 346, 316, 315, 331, 385, 417, 421, 397, 350, 321, 318, 334, 346, 345, 341, 319, 265, 199, 173, 188, 213, 226, 245, 258, 263, 231, 201, 175, 155, 
    352, 329, 302, 304, 326, 375, 403, 402, 349, 273, 237, 259, 322, 341, 329, 316, 291, 239, 187, 176, 185, 202, 209, 218, 225, 229, 212, 190, 172, 159, 
    343, 313, 279, 274, 306, 359, 398, 393, 331, 238, 201, 226, 297, 317, 294, 275, 249, 204, 168, 161, 171, 184, 191, 187, 179, 174, 175, 183, 184, 171, 
    334, 297, 260, 241, 273, 337, 391, 393, 344, 286, 271, 264, 286, 274, 246, 227, 204, 160, 137, 136, 155, 169, 170, 160, 149, 133, 144, 176, 196, 196, 
    320, 282, 241, 216, 248, 316, 384, 391, 358, 330, 326, 300, 265, 233, 211, 193, 165, 122, 112, 117, 150, 162, 164, 150, 133, 124, 139, 172, 199, 202, 
    288, 261, 227, 197, 222, 291, 370, 387, 364, 340, 325, 285, 238, 207, 186, 172, 133, 95, 94, 110, 141, 152, 161, 150, 137, 130, 146, 172, 186, 181, 
    241, 231, 219, 188, 197, 255, 344, 379, 366, 345, 301, 241, 183, 154, 150, 141, 107, 86, 90, 111, 131, 145, 156, 157, 149, 146, 152, 159, 163, 169, 
    182, 178, 184, 161, 163, 208, 297, 354, 345, 314, 254, 172, 93, 66, 75, 88, 88, 85, 94, 107, 122, 139, 153, 153, 142, 137, 133, 142, 160, 175, 
    
    -- channel=142
    6, 30, 133, 134, 38, 9, 24, 21, 18, 25, 26, 14, 7, 13, 18, 2, 0, 0, 0, 39, 96, 82, 20, 10, 11, 8, 11, 10, 8, 9, 
    8, 15, 115, 158, 67, 21, 43, 39, 11, 16, 40, 36, 15, 14, 22, 25, 0, 0, 0, 7, 109, 82, 22, 20, 21, 18, 19, 17, 14, 13, 
    11, 9, 88, 159, 84, 25, 64, 70, 21, 0, 27, 56, 47, 40, 34, 38, 36, 0, 0, 9, 102, 68, 21, 19, 19, 19, 22, 22, 20, 18, 
    10, 7, 61, 147, 94, 25, 79, 103, 56, 0, 4, 60, 88, 95, 84, 66, 50, 10, 0, 36, 98, 72, 42, 28, 21, 19, 19, 18, 17, 17, 
    10, 10, 40, 126, 96, 14, 56, 113, 92, 17, 0, 16, 61, 95, 103, 90, 68, 40, 26, 57, 71, 65, 68, 55, 40, 37, 30, 19, 15, 12, 
    0, 6, 20, 84, 73, 0, 24, 106, 110, 41, 0, 0, 0, 41, 54, 71, 63, 58, 83, 88, 44, 42, 67, 55, 40, 44, 42, 39, 43, 38, 
    0, 0, 0, 47, 44, 0, 22, 112, 126, 67, 4, 0, 0, 0, 0, 25, 38, 49, 112, 125, 56, 50, 86, 65, 49, 54, 45, 57, 74, 68, 
    0, 0, 0, 45, 37, 0, 6, 106, 140, 94, 51, 12, 0, 0, 0, 13, 35, 46, 105, 130, 63, 58, 99, 79, 65, 56, 33, 54, 90, 91, 
    0, 0, 22, 43, 27, 0, 0, 71, 120, 96, 74, 58, 31, 8, 1, 31, 51, 50, 95, 119, 75, 73, 83, 64, 48, 15, 0, 26, 76, 102, 
    15, 26, 48, 47, 27, 0, 0, 56, 85, 72, 68, 62, 44, 26, 13, 37, 43, 39, 86, 106, 89, 103, 92, 62, 44, 1, 0, 3, 47, 89, 
    27, 30, 52, 59, 32, 0, 0, 64, 82, 70, 72, 59, 30, 11, 21, 43, 28, 21, 73, 87, 79, 110, 108, 70, 47, 8, 0, 0, 23, 58, 
    34, 33, 49, 57, 41, 15, 18, 60, 94, 92, 91, 70, 22, 0, 18, 45, 20, 19, 63, 73, 75, 106, 105, 75, 54, 24, 0, 0, 0, 25, 
    26, 28, 42, 36, 35, 68, 41, 20, 48, 56, 71, 62, 22, 22, 59, 66, 24, 37, 62, 57, 75, 105, 98, 74, 64, 49, 8, 0, 0, 23, 
    22, 25, 42, 11, 2, 97, 71, 2, 0, 5, 42, 51, 14, 17, 85, 90, 31, 38, 63, 52, 60, 108, 112, 81, 68, 68, 45, 0, 8, 42, 
    23, 34, 56, 13, 0, 97, 109, 39, 33, 42, 55, 61, 38, 4, 44, 90, 58, 24, 72, 83, 56, 104, 156, 147, 104, 82, 57, 27, 43, 51, 
    10, 34, 70, 45, 0, 71, 123, 66, 37, 47, 35, 30, 53, 43, 11, 66, 99, 29, 55, 93, 40, 26, 115, 190, 177, 126, 68, 57, 76, 56, 
    0, 6, 56, 65, 11, 34, 95, 81, 40, 38, 22, 0, 27, 44, 0, 10, 101, 52, 30, 82, 29, 0, 0, 89, 162, 148, 89, 88, 112, 79, 
    0, 0, 29, 61, 42, 32, 57, 84, 90, 90, 69, 31, 23, 24, 0, 0, 52, 62, 39, 73, 41, 0, 0, 0, 61, 88, 60, 79, 130, 125, 
    0, 0, 29, 63, 57, 52, 42, 56, 87, 103, 105, 93, 70, 35, 5, 0, 0, 33, 50, 49, 30, 41, 34, 0, 23, 44, 26, 40, 93, 131, 
    15, 0, 35, 74, 65, 60, 49, 38, 46, 58, 68, 104, 108, 67, 54, 12, 0, 9, 49, 34, 25, 44, 41, 22, 34, 42, 29, 30, 46, 77, 
    32, 6, 20, 72, 77, 49, 46, 48, 45, 28, 19, 72, 99, 81, 91, 79, 23, 21, 27, 26, 37, 44, 41, 45, 45, 32, 22, 32, 41, 45, 
    45, 17, 2, 60, 96, 61, 45, 54, 56, 26, 1, 38, 65, 61, 70, 73, 51, 28, 1, 19, 53, 49, 45, 57, 42, 14, 14, 25, 30, 28, 
    47, 30, 0, 44, 103, 88, 66, 63, 56, 41, 38, 51, 51, 47, 54, 53, 43, 14, 0, 22, 58, 51, 47, 69, 51, 14, 19, 15, 7, 8, 
    41, 36, 2, 35, 94, 94, 79, 76, 58, 51, 97, 113, 65, 47, 59, 59, 41, 8, 0, 36, 61, 46, 46, 79, 69, 38, 30, 21, 15, 17, 
    34, 31, 11, 37, 88, 90, 68, 62, 28, 3, 96, 145, 76, 46, 62, 61, 40, 17, 16, 47, 60, 40, 43, 68, 68, 59, 44, 32, 23, 18, 
    28, 21, 10, 34, 88, 97, 63, 44, 0, 0, 38, 109, 66, 46, 59, 54, 39, 25, 25, 56, 57, 36, 44, 50, 44, 54, 60, 45, 19, 4, 
    27, 18, 3, 21, 85, 108, 73, 39, 0, 0, 17, 57, 42, 44, 50, 41, 35, 19, 30, 60, 49, 30, 37, 30, 19, 36, 59, 56, 35, 20, 
    32, 25, 0, 8, 82, 120, 84, 43, 23, 24, 40, 33, 25, 38, 39, 28, 25, 8, 35, 56, 41, 35, 32, 17, 10, 27, 48, 56, 49, 35, 
    39, 40, 2, 0, 76, 135, 99, 53, 39, 40, 35, 24, 29, 49, 46, 28, 12, 9, 43, 46, 40, 44, 35, 15, 8, 25, 42, 52, 50, 34, 
    43, 59, 22, 0, 56, 143, 119, 66, 52, 47, 29, 22, 44, 73, 70, 40, 8, 19, 40, 33, 38, 47, 36, 20, 22, 34, 42, 46, 43, 30, 
    
    -- channel=143
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=144
    0, 0, 0, 0, 0, 7, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 26, 29, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 55, 75, 30, 48, 38, 30, 58, 34, 25, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 82, 119, 58, 68, 60, 53, 74, 58, 59, 69, 45, 49, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 64, 129, 61, 33, 30, 34, 46, 32, 38, 50, 51, 56, 49, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 42, 126, 51, 0, 0, 0, 17, 22, 21, 35, 33, 39, 35, 15, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 37, 129, 46, 0, 0, 0, 12, 47, 40, 37, 30, 26, 33, 8, 2, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 57, 135, 35, 0, 38, 10, 29, 72, 50, 34, 27, 19, 35, 9, 6, 25, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 0, 26, 35, 94, 123, 35, 10, 54, 27, 42, 68, 51, 38, 32, 27, 41, 21, 1, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 44, 63, 88, 115, 60, 31, 57, 52, 59, 62, 55, 51, 48, 50, 59, 37, 17, 26, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 39, 23, 71, 129, 94, 49, 42, 50, 62, 66, 65, 64, 66, 67, 55, 41, 40, 33, 26, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 43, 15, 77, 116, 92, 39, 28, 38, 46, 74, 81, 68, 60, 48, 23, 25, 51, 41, 16, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 35, 47, 30, 61, 76, 58, 37, 50, 58, 52, 77, 95, 79, 59, 47, 35, 49, 81, 70, 37, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 43, 63, 37, 12, 12, 44, 66, 70, 86, 94, 84, 85, 94, 87, 74, 74, 79, 92, 105, 90, 72, 57, 42, 34, 35, 2, 0, 0, 0, 
    0, 90, 98, 29, 0, 0, 63, 115, 73, 85, 88, 85, 74, 75, 94, 96, 93, 100, 92, 93, 99, 88, 86, 70, 50, 45, 21, 0, 0, 0, 
    9, 94, 96, 6, 0, 26, 116, 111, 53, 47, 29, 46, 51, 60, 95, 94, 69, 72, 41, 26, 78, 82, 69, 55, 11, 7, 8, 0, 0, 0, 
    1, 84, 89, 0, 0, 106, 146, 58, 26, 42, 28, 36, 39, 51, 61, 31, 5, 10, 0, 0, 31, 38, 12, 0, 0, 4, 18, 0, 0, 0, 
    2, 95, 105, 0, 15, 147, 135, 34, 27, 78, 83, 74, 52, 52, 24, 0, 21, 36, 4, 12, 49, 36, 28, 0, 0, 66, 72, 30, 0, 0, 
    0, 97, 128, 35, 37, 137, 113, 58, 57, 88, 100, 87, 71, 71, 6, 2, 81, 75, 47, 55, 73, 66, 62, 31, 35, 115, 105, 30, 0, 0, 
    0, 87, 137, 75, 55, 101, 101, 95, 85, 73, 79, 80, 68, 67, 53, 49, 71, 75, 69, 75, 82, 63, 58, 55, 66, 90, 71, 28, 0, 0, 
    0, 86, 127, 69, 70, 78, 92, 110, 97, 79, 63, 46, 25, 67, 107, 62, 24, 51, 73, 62, 66, 31, 5, 87, 87, 23, 25, 48, 0, 0, 
    0, 98, 145, 56, 53, 75, 68, 103, 107, 92, 70, 41, 18, 67, 145, 74, 0, 2, 52, 28, 33, 0, 0, 90, 125, 21, 26, 80, 0, 0, 
    8, 116, 167, 77, 29, 33, 46, 98, 121, 102, 85, 77, 60, 94, 139, 77, 0, 15, 58, 24, 30, 19, 19, 133, 147, 58, 74, 86, 0, 0, 
    17, 101, 152, 73, 23, 0, 37, 111, 122, 108, 102, 96, 87, 101, 104, 85, 48, 3, 0, 0, 3, 2, 73, 158, 119, 79, 78, 52, 0, 0, 
    12, 47, 80, 60, 25, 0, 54, 110, 98, 108, 113, 103, 97, 94, 87, 93, 64, 0, 0, 0, 0, 0, 84, 161, 121, 81, 60, 30, 0, 0, 
    0, 5, 33, 61, 64, 12, 60, 98, 78, 101, 123, 111, 95, 91, 78, 70, 44, 0, 0, 6, 22, 20, 116, 179, 128, 76, 41, 25, 0, 0, 
    0, 10, 38, 63, 76, 31, 65, 96, 70, 98, 124, 107, 87, 82, 73, 59, 43, 19, 29, 43, 27, 23, 129, 177, 116, 69, 39, 29, 0, 0, 
    15, 35, 42, 46, 66, 64, 85, 88, 72, 95, 111, 103, 84, 79, 75, 70, 67, 61, 56, 43, 27, 28, 115, 172, 109, 67, 49, 30, 0, 0, 
    32, 34, 34, 37, 68, 100, 101, 72, 74, 93, 97, 94, 83, 76, 77, 76, 69, 63, 60, 51, 44, 44, 97, 148, 114, 68, 49, 11, 0, 0, 
    22, 17, 20, 25, 58, 123, 113, 69, 76, 85, 82, 77, 73, 68, 71, 71, 59, 50, 53, 50, 47, 47, 77, 113, 104, 62, 25, 0, 0, 0, 
    
    -- channel=145
    225, 218, 208, 211, 220, 216, 204, 186, 180, 166, 164, 166, 168, 166, 158, 171, 188, 218, 234, 230, 221, 223, 229, 230, 217, 192, 185, 202, 199, 178, 
    235, 234, 232, 225, 228, 231, 213, 184, 197, 205, 193, 205, 214, 216, 226, 236, 242, 248, 247, 245, 234, 224, 224, 233, 228, 213, 206, 214, 204, 184, 
    248, 246, 246, 245, 250, 257, 230, 188, 200, 216, 212, 222, 224, 225, 247, 250, 248, 250, 236, 234, 234, 218, 211, 227, 231, 229, 225, 211, 200, 201, 
    262, 261, 260, 258, 261, 269, 253, 209, 211, 219, 219, 232, 216, 217, 232, 228, 239, 247, 234, 230, 210, 204, 207, 221, 226, 225, 216, 198, 194, 215, 
    261, 260, 260, 261, 265, 258, 226, 187, 188, 199, 196, 213, 202, 197, 203, 194, 206, 209, 195, 206, 202, 187, 209, 222, 214, 220, 208, 188, 187, 208, 
    261, 261, 259, 263, 264, 260, 239, 181, 159, 185, 194, 205, 217, 227, 228, 217, 206, 203, 188, 166, 191, 214, 213, 227, 219, 208, 199, 176, 168, 187, 
    261, 259, 260, 264, 252, 253, 265, 207, 170, 209, 221, 231, 243, 261, 272, 265, 254, 242, 240, 213, 179, 211, 225, 230, 229, 206, 188, 173, 148, 161, 
    259, 258, 263, 264, 240, 248, 263, 208, 181, 251, 271, 288, 289, 269, 262, 258, 256, 257, 251, 261, 238, 190, 186, 219, 225, 212, 206, 201, 174, 151, 
    256, 257, 262, 265, 255, 262, 263, 199, 188, 235, 227, 252, 276, 251, 245, 248, 246, 258, 248, 254, 257, 214, 192, 205, 215, 227, 236, 207, 170, 153, 
    247, 253, 260, 269, 257, 250, 235, 190, 191, 226, 219, 231, 249, 241, 239, 243, 243, 254, 249, 248, 263, 234, 214, 228, 242, 252, 255, 230, 199, 204, 
    234, 247, 257, 266, 219, 191, 199, 179, 178, 207, 215, 213, 221, 223, 220, 221, 227, 229, 223, 232, 248, 234, 214, 211, 230, 249, 261, 260, 260, 260, 
    211, 231, 249, 243, 211, 209, 205, 161, 148, 169, 202, 203, 202, 211, 209, 205, 204, 200, 195, 201, 206, 206, 194, 169, 190, 236, 255, 253, 259, 261, 
    191, 220, 233, 205, 182, 201, 205, 164, 135, 156, 194, 215, 215, 198, 183, 179, 177, 178, 185, 190, 171, 160, 166, 176, 216, 251, 263, 253, 251, 260, 
    175, 194, 202, 167, 140, 145, 164, 183, 187, 206, 200, 197, 212, 205, 179, 172, 182, 201, 220, 223, 188, 158, 163, 175, 196, 210, 224, 240, 249, 258, 
    171, 185, 185, 153, 132, 117, 150, 190, 195, 194, 188, 177, 183, 180, 165, 158, 150, 150, 154, 147, 146, 143, 134, 146, 163, 185, 191, 186, 224, 256, 
    186, 200, 166, 104, 101, 136, 211, 198, 160, 158, 130, 105, 110, 109, 121, 117, 110, 114, 120, 105, 108, 121, 117, 130, 139, 149, 164, 155, 192, 242, 
    175, 181, 154, 85, 83, 150, 213, 175, 130, 141, 145, 151, 149, 134, 140, 99, 71, 70, 67, 76, 99, 82, 65, 68, 75, 127, 160, 150, 175, 226, 
    199, 209, 187, 116, 113, 162, 155, 112, 120, 144, 159, 185, 194, 178, 166, 125, 125, 143, 140, 154, 200, 172, 130, 135, 130, 173, 199, 189, 185, 212, 
    213, 212, 183, 116, 127, 167, 118, 74, 119, 152, 145, 130, 140, 164, 166, 155, 202, 224, 218, 225, 231, 225, 218, 214, 218, 225, 204, 171, 147, 176, 
    213, 218, 190, 113, 124, 153, 112, 84, 107, 122, 122, 104, 107, 105, 121, 171, 201, 165, 151, 168, 175, 168, 157, 153, 178, 202, 158, 125, 129, 162, 
    214, 226, 206, 108, 84, 122, 110, 96, 89, 88, 116, 113, 111, 104, 122, 129, 148, 162, 173, 170, 164, 163, 148, 152, 182, 167, 139, 129, 127, 154, 
    216, 228, 212, 136, 88, 100, 114, 103, 86, 66, 79, 94, 112, 119, 124, 96, 86, 103, 125, 116, 113, 114, 109, 130, 125, 104, 133, 158, 136, 145, 
    227, 235, 208, 127, 122, 116, 105, 119, 100, 74, 63, 78, 116, 159, 164, 87, 66, 128, 159, 142, 142, 142, 147, 208, 168, 91, 137, 183, 137, 137, 
    240, 243, 203, 111, 101, 138, 132, 153, 125, 85, 70, 66, 70, 99, 116, 75, 70, 132, 169, 170, 182, 182, 173, 224, 173, 84, 96, 109, 95, 141, 
    232, 237, 194, 111, 81, 108, 160, 192, 139, 95, 77, 63, 54, 55, 58, 63, 72, 75, 89, 126, 148, 160, 165, 151, 100, 79, 82, 84, 94, 151, 
    220, 224, 211, 165, 136, 139, 162, 184, 139, 113, 86, 65, 56, 57, 58, 62, 56, 57, 126, 216, 240, 230, 229, 204, 103, 67, 75, 90, 117, 162, 
    211, 218, 233, 234, 197, 160, 165, 173, 138, 131, 109, 71, 50, 50, 53, 60, 61, 64, 129, 208, 222, 216, 217, 196, 95, 52, 65, 100, 132, 167, 
    217, 230, 233, 223, 195, 160, 170, 169, 135, 135, 114, 77, 57, 57, 61, 70, 92, 112, 127, 143, 151, 171, 187, 158, 83, 54, 67, 105, 131, 166, 
    238, 237, 224, 210, 200, 178, 163, 143, 126, 127, 111, 83, 69, 69, 74, 78, 84, 93, 107, 121, 137, 160, 185, 153, 79, 58, 71, 103, 124, 177, 
    233, 227, 225, 217, 206, 184, 158, 119, 118, 117, 104, 92, 81, 78, 84, 87, 88, 92, 101, 112, 124, 137, 154, 147, 93, 65, 78, 97, 124, 192, 
    
    -- channel=146
    42, 36, 39, 41, 37, 40, 49, 35, 35, 35, 28, 26, 26, 27, 19, 25, 32, 39, 44, 42, 43, 43, 42, 37, 39, 26, 22, 22, 41, 26, 
    47, 46, 46, 44, 40, 48, 65, 49, 50, 65, 56, 56, 67, 57, 58, 68, 57, 59, 49, 48, 50, 49, 40, 39, 39, 29, 31, 34, 36, 26, 
    55, 54, 54, 53, 49, 54, 89, 76, 72, 100, 80, 91, 99, 82, 96, 97, 75, 84, 59, 50, 54, 48, 32, 38, 41, 34, 35, 35, 25, 30, 
    62, 61, 61, 59, 59, 64, 110, 103, 98, 122, 102, 116, 115, 102, 116, 111, 102, 109, 78, 56, 46, 40, 29, 39, 35, 30, 33, 31, 23, 34, 
    62, 62, 62, 60, 65, 61, 96, 107, 94, 110, 101, 111, 110, 103, 110, 110, 110, 110, 92, 69, 42, 33, 32, 42, 33, 33, 29, 30, 24, 27, 
    62, 62, 60, 63, 75, 59, 85, 115, 79, 90, 84, 95, 111, 117, 124, 121, 116, 114, 104, 84, 55, 44, 41, 39, 38, 35, 22, 23, 21, 23, 
    62, 61, 58, 68, 78, 58, 103, 136, 81, 97, 98, 96, 126, 143, 145, 143, 132, 131, 126, 101, 86, 66, 39, 43, 47, 28, 14, 16, 22, 23, 
    61, 60, 59, 68, 75, 68, 123, 135, 86, 124, 133, 112, 143, 151, 142, 143, 132, 131, 141, 121, 108, 82, 37, 39, 39, 28, 29, 37, 29, 18, 
    60, 59, 59, 67, 94, 96, 128, 127, 89, 127, 133, 115, 142, 144, 137, 139, 132, 130, 143, 127, 119, 103, 52, 37, 43, 42, 43, 40, 18, 10, 
    54, 57, 57, 70, 107, 92, 116, 119, 100, 127, 130, 125, 136, 137, 138, 137, 136, 137, 142, 133, 131, 120, 89, 68, 60, 52, 53, 45, 34, 34, 
    48, 52, 55, 68, 82, 65, 106, 117, 108, 110, 122, 120, 122, 124, 128, 128, 131, 131, 123, 120, 123, 115, 106, 76, 52, 51, 64, 61, 61, 61, 
    41, 47, 57, 70, 65, 58, 110, 109, 90, 85, 110, 115, 120, 124, 123, 123, 120, 114, 97, 101, 108, 95, 85, 54, 42, 55, 67, 61, 61, 61, 
    39, 41, 59, 58, 52, 50, 90, 80, 83, 92, 115, 119, 119, 124, 113, 106, 101, 101, 97, 104, 98, 79, 78, 72, 73, 77, 80, 64, 58, 62, 
    23, 29, 59, 46, 42, 25, 46, 81, 112, 113, 120, 121, 123, 122, 108, 106, 111, 120, 123, 116, 100, 83, 83, 82, 87, 90, 97, 75, 52, 61, 
    20, 34, 67, 46, 26, 0, 30, 100, 119, 116, 112, 101, 102, 93, 84, 91, 89, 91, 98, 87, 79, 80, 80, 90, 100, 91, 96, 80, 45, 56, 
    31, 26, 60, 35, 9, 3, 68, 110, 93, 74, 59, 42, 60, 51, 60, 73, 58, 52, 63, 40, 45, 67, 58, 71, 67, 67, 83, 72, 44, 48, 
    28, 19, 63, 31, 3, 18, 99, 95, 69, 60, 62, 59, 83, 58, 70, 44, 12, 11, 26, 6, 23, 39, 10, 22, 26, 48, 76, 75, 64, 42, 
    45, 41, 82, 46, 9, 36, 91, 59, 56, 69, 85, 85, 93, 77, 88, 36, 37, 59, 67, 60, 73, 70, 49, 63, 49, 72, 103, 97, 83, 35, 
    48, 40, 80, 58, 24, 47, 67, 43, 65, 74, 77, 73, 81, 77, 85, 58, 96, 111, 100, 98, 108, 107, 101, 103, 77, 99, 113, 86, 72, 27, 
    48, 38, 83, 62, 36, 46, 55, 46, 64, 59, 66, 64, 63, 54, 72, 73, 89, 86, 82, 89, 92, 92, 78, 79, 84, 97, 90, 64, 66, 25, 
    51, 39, 83, 55, 31, 40, 51, 46, 54, 47, 65, 57, 60, 40, 66, 80, 75, 69, 82, 88, 78, 86, 61, 56, 93, 79, 56, 60, 81, 27, 
    58, 46, 91, 61, 29, 49, 45, 38, 44, 35, 47, 42, 58, 37, 72, 73, 37, 17, 52, 55, 40, 58, 24, 20, 85, 57, 45, 84, 96, 24, 
    75, 58, 98, 71, 36, 54, 34, 40, 53, 36, 41, 47, 67, 59, 80, 61, 33, 32, 68, 62, 49, 69, 45, 59, 103, 58, 60, 94, 86, 23, 
    90, 75, 95, 65, 36, 44, 36, 66, 63, 41, 37, 39, 45, 48, 54, 44, 54, 65, 58, 56, 54, 69, 53, 84, 84, 47, 53, 62, 63, 32, 
    93, 81, 75, 47, 33, 47, 47, 87, 64, 42, 36, 33, 30, 32, 33, 34, 48, 39, 0, 24, 41, 55, 36, 75, 62, 43, 47, 45, 63, 49, 
    87, 76, 69, 69, 67, 69, 45, 89, 63, 45, 43, 38, 30, 31, 33, 30, 35, 34, 27, 76, 92, 87, 62, 94, 63, 39, 41, 45, 77, 60, 
    80, 82, 91, 96, 87, 79, 46, 90, 65, 55, 50, 37, 25, 25, 28, 25, 28, 42, 57, 90, 92, 83, 63, 92, 52, 32, 37, 52, 86, 63, 
    89, 97, 100, 92, 79, 78, 61, 86, 64, 60, 51, 37, 27, 27, 32, 37, 46, 54, 61, 69, 69, 72, 60, 81, 45, 33, 38, 58, 84, 59, 
    106, 104, 100, 93, 79, 78, 77, 72, 59, 59, 52, 40, 35, 33, 35, 38, 44, 48, 54, 62, 67, 75, 63, 68, 48, 34, 38, 62, 70, 61, 
    108, 101, 99, 91, 83, 78, 84, 57, 55, 59, 50, 38, 39, 36, 38, 42, 45, 43, 47, 55, 59, 63, 59, 58, 52, 34, 40, 52, 51, 69, 
    
    -- channel=147
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=148
    128, 128, 118, 126, 124, 121, 114, 123, 122, 109, 107, 104, 116, 106, 97, 113, 124, 137, 148, 148, 140, 150, 152, 151, 126, 107, 116, 144, 126, 107, 
    132, 131, 128, 126, 136, 126, 102, 103, 111, 115, 106, 114, 129, 133, 146, 156, 155, 151, 151, 160, 161, 153, 146, 151, 142, 137, 135, 160, 136, 117, 
    142, 141, 140, 138, 145, 141, 117, 104, 100, 94, 97, 96, 94, 111, 128, 131, 149, 151, 154, 161, 161, 147, 137, 145, 153, 149, 146, 152, 150, 146, 
    144, 145, 144, 144, 146, 135, 83, 74, 72, 37, 52, 46, 30, 44, 40, 48, 82, 85, 112, 140, 141, 130, 136, 138, 145, 153, 149, 143, 162, 168, 
    144, 145, 144, 145, 154, 139, 55, 28, 28, 0, 5, 5, 0, 4, 0, 0, 9, 10, 23, 63, 109, 131, 147, 136, 133, 153, 146, 132, 148, 166, 
    145, 145, 141, 145, 149, 146, 77, 24, 23, 11, 18, 12, 9, 26, 26, 18, 11, 9, 12, 6, 58, 138, 169, 151, 146, 139, 127, 106, 116, 152, 
    143, 144, 145, 144, 124, 125, 96, 22, 34, 59, 90, 81, 57, 51, 43, 37, 34, 27, 36, 34, 39, 96, 144, 155, 147, 121, 120, 120, 124, 135, 
    145, 144, 149, 137, 112, 134, 98, 16, 38, 60, 72, 96, 76, 39, 33, 31, 40, 38, 33, 59, 45, 49, 109, 132, 121, 128, 128, 123, 103, 86, 
    147, 146, 146, 132, 126, 137, 72, 13, 44, 43, 30, 72, 65, 34, 33, 33, 40, 52, 39, 54, 60, 38, 91, 133, 140, 145, 140, 108, 83, 84, 
    152, 148, 146, 141, 100, 67, 32, 9, 65, 61, 33, 45, 42, 32, 29, 32, 41, 56, 42, 54, 71, 48, 81, 136, 149, 145, 147, 128, 123, 131, 
    148, 148, 152, 155, 91, 67, 26, 0, 41, 43, 30, 16, 9, 24, 31, 35, 40, 37, 23, 32, 64, 74, 76, 95, 116, 142, 145, 143, 144, 145, 
    140, 150, 157, 143, 113, 115, 61, 0, 0, 0, 15, 18, 0, 0, 10, 15, 9, 0, 0, 5, 30, 57, 60, 81, 134, 172, 169, 155, 145, 144, 
    122, 132, 144, 119, 104, 114, 68, 15, 0, 8, 14, 39, 38, 18, 15, 18, 21, 31, 57, 60, 46, 51, 58, 85, 122, 143, 158, 168, 154, 144, 
    113, 125, 132, 128, 103, 85, 34, 44, 35, 29, 39, 56, 70, 51, 34, 32, 38, 45, 65, 66, 52, 49, 53, 70, 94, 105, 104, 134, 152, 147, 
    140, 135, 99, 102, 93, 91, 85, 72, 31, 21, 10, 0, 0, 1, 3, 21, 43, 44, 48, 34, 17, 35, 48, 65, 72, 60, 42, 72, 129, 145, 
    124, 108, 58, 47, 64, 100, 146, 85, 29, 23, 19, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 21, 105, 146, 
    107, 112, 67, 54, 68, 100, 105, 64, 22, 22, 55, 84, 61, 41, 44, 3, 0, 0, 0, 11, 28, 0, 0, 0, 0, 12, 38, 59, 115, 150, 
    113, 114, 60, 63, 92, 108, 34, 23, 40, 47, 51, 73, 65, 93, 72, 30, 50, 83, 70, 93, 103, 75, 77, 73, 63, 64, 77, 86, 86, 130, 
    120, 109, 49, 46, 106, 108, 13, 5, 52, 57, 27, 18, 26, 48, 36, 89, 91, 54, 49, 68, 68, 64, 67, 55, 84, 85, 46, 38, 47, 114, 
    125, 118, 55, 15, 64, 76, 21, 12, 31, 45, 41, 25, 8, 0, 8, 84, 86, 51, 48, 62, 56, 55, 50, 30, 88, 87, 16, 0, 28, 109, 
    119, 121, 72, 33, 23, 40, 33, 15, 3, 22, 41, 33, 14, 0, 0, 37, 59, 26, 14, 21, 15, 15, 20, 0, 21, 57, 26, 13, 37, 108, 
    109, 115, 67, 67, 53, 35, 21, 2, 0, 14, 16, 39, 56, 75, 49, 22, 37, 46, 37, 25, 18, 12, 42, 53, 26, 35, 71, 86, 55, 97, 
    102, 109, 50, 40, 84, 55, 19, 12, 7, 13, 5, 29, 40, 97, 69, 6, 32, 111, 98, 64, 68, 40, 70, 138, 54, 17, 68, 68, 30, 86, 
    93, 103, 29, 0, 21, 38, 47, 51, 18, 7, 10, 14, 13, 41, 30, 6, 28, 81, 42, 12, 25, 17, 33, 59, 23, 24, 39, 21, 8, 82, 
    89, 97, 30, 0, 0, 32, 72, 57, 26, 5, 1, 13, 18, 18, 18, 18, 12, 24, 54, 72, 87, 79, 75, 40, 22, 33, 31, 13, 10, 75, 
    74, 80, 72, 48, 34, 39, 71, 49, 35, 21, 10, 10, 14, 12, 12, 16, 0, 0, 88, 136, 139, 108, 111, 63, 23, 20, 20, 21, 23, 70, 
    63, 78, 92, 79, 48, 32, 79, 54, 37, 38, 22, 8, 11, 10, 10, 20, 23, 29, 79, 94, 87, 82, 83, 40, 18, 12, 17, 32, 29, 65, 
    78, 82, 72, 63, 52, 31, 78, 49, 37, 40, 27, 13, 13, 16, 13, 19, 32, 37, 47, 50, 57, 77, 89, 27, 9, 15, 21, 35, 27, 59, 
    75, 68, 61, 55, 50, 29, 52, 40, 36, 35, 32, 21, 14, 15, 14, 14, 16, 20, 24, 30, 42, 58, 86, 30, 6, 13, 21, 27, 12, 54, 
    57, 50, 46, 46, 53, 33, 18, 30, 43, 40, 28, 21, 14, 10, 9, 12, 13, 13, 11, 13, 19, 26, 48, 32, 0, 0, 13, 8, 9, 64, 
    
    -- channel=149
    0, 0, 0, 0, 0, 0, 9, 13, 5, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 5, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 11, 0, 0, 14, 7, 0, 13, 0, 5, 8, 5, 3, 4, 0, 4, 3, 0, 0, 9, 6, 0, 
    0, 0, 0, 0, 0, 0, 25, 13, 0, 21, 0, 7, 14, 0, 22, 30, 14, 31, 17, 10, 12, 6, 0, 0, 0, 2, 3, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 27, 14, 10, 7, 0, 7, 0, 0, 1, 0, 1, 19, 24, 21, 10, 0, 0, 0, 2, 1, 12, 8, 0, 2, 
    0, 0, 0, 0, 10, 14, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 5, 0, 0, 0, 0, 3, 8, 6, 5, 6, 
    0, 0, 0, 0, 19, 25, 15, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 2, 0, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 17, 0, 23, 39, 0, 0, 5, 0, 0, 0, 5, 10, 0, 0, 11, 0, 0, 0, 4, 5, 19, 2, 0, 0, 0, 0, 
    0, 0, 0, 8, 6, 0, 38, 18, 0, 0, 23, 10, 17, 11, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 27, 46, 19, 0, 0, 0, 4, 27, 9, 1, 0, 1, 0, 3, 0, 0, 1, 0, 0, 0, 0, 0, 6, 0, 0, 
    6, 0, 0, 0, 24, 13, 23, 10, 2, 19, 0, 2, 17, 6, 3, 2, 0, 14, 12, 4, 11, 0, 0, 5, 11, 0, 14, 5, 0, 0, 
    6, 0, 1, 35, 29, 0, 3, 0, 8, 14, 2, 0, 0, 1, 5, 5, 8, 14, 0, 0, 17, 10, 6, 11, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 41, 28, 10, 23, 5, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 13, 16, 0, 0, 5, 12, 3, 0, 0, 
    0, 0, 21, 22, 14, 24, 50, 7, 0, 0, 0, 7, 9, 10, 7, 8, 5, 1, 0, 10, 8, 0, 0, 0, 0, 14, 29, 17, 2, 0, 
    0, 0, 39, 29, 15, 12, 0, 0, 6, 7, 14, 22, 35, 36, 19, 9, 4, 7, 24, 42, 29, 9, 5, 4, 11, 6, 19, 26, 5, 0, 
    0, 4, 31, 38, 30, 0, 0, 10, 6, 0, 4, 0, 0, 2, 0, 9, 17, 20, 22, 21, 16, 14, 16, 14, 18, 11, 0, 6, 0, 0, 
    5, 8, 20, 4, 0, 0, 30, 51, 17, 14, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 2, 31, 0, 0, 0, 66, 48, 5, 0, 12, 9, 21, 0, 8, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 32, 14, 0, 6, 48, 5, 0, 0, 0, 26, 36, 17, 57, 0, 0, 8, 0, 0, 34, 24, 4, 7, 0, 0, 7, 14, 19, 0, 
    8, 2, 18, 8, 1, 42, 27, 0, 0, 20, 10, 0, 0, 24, 23, 0, 1, 14, 3, 0, 14, 13, 8, 25, 0, 11, 32, 13, 0, 0, 
    11, 2, 16, 0, 4, 35, 12, 0, 11, 21, 17, 4, 0, 0, 0, 19, 45, 20, 2, 15, 22, 20, 14, 0, 12, 46, 17, 0, 0, 0, 
    4, 9, 41, 0, 0, 5, 5, 0, 0, 0, 20, 13, 0, 0, 0, 0, 14, 0, 0, 2, 0, 7, 0, 0, 12, 36, 1, 0, 0, 0, 
    0, 0, 46, 37, 0, 0, 0, 0, 0, 0, 11, 6, 25, 0, 8, 28, 13, 0, 0, 0, 0, 0, 0, 0, 9, 14, 0, 11, 23, 0, 
    1, 3, 29, 33, 19, 17, 0, 0, 2, 0, 0, 0, 4, 25, 59, 19, 0, 2, 36, 10, 0, 0, 0, 23, 55, 0, 0, 47, 20, 0, 
    5, 9, 30, 0, 0, 8, 0, 4, 14, 0, 0, 0, 0, 13, 32, 0, 0, 16, 9, 0, 0, 0, 0, 38, 45, 0, 6, 11, 0, 0, 
    10, 30, 21, 0, 0, 0, 0, 31, 15, 0, 0, 4, 4, 3, 1, 0, 12, 25, 0, 0, 0, 0, 0, 8, 16, 10, 13, 0, 0, 0, 
    5, 17, 12, 0, 0, 0, 0, 26, 15, 0, 0, 4, 2, 2, 1, 1, 0, 0, 0, 10, 31, 18, 14, 47, 25, 8, 3, 0, 0, 0, 
    0, 0, 7, 19, 11, 8, 0, 28, 6, 7, 15, 8, 0, 0, 0, 6, 0, 0, 0, 19, 27, 7, 11, 50, 24, 1, 0, 0, 0, 0, 
    0, 3, 12, 14, 0, 0, 9, 31, 2, 12, 17, 8, 0, 0, 0, 0, 0, 1, 5, 9, 3, 9, 13, 40, 14, 0, 0, 0, 0, 0, 
    6, 8, 5, 2, 0, 0, 18, 20, 1, 10, 16, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 30, 31, 9, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 18, 6, 5, 11, 12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 15, 4, 0, 0, 0, 0, 0, 
    
    -- channel=150
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 24, 30, 22, 17, 5, 16, 34, 30, 17, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 3, 0, 4, 0, 0, 5, 7, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 21, 12, 0, 8, 6, 5, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 4, 9, 11, 17, 10, 0, 0, 0, 0, 1, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 6, 19, 11, 4, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 17, 0, 0, 0, 0, 15, 15, 19, 11, 20, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 18, 10, 0, 0, 
    0, 0, 0, 0, 17, 0, 0, 0, 0, 7, 24, 30, 31, 35, 30, 18, 14, 27, 15, 0, 0, 0, 0, 6, 19, 19, 19, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 24, 30, 24, 20, 27, 27, 7, 0, 0, 0, 0, 0, 0, 0, 22, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 30, 28, 26, 25, 9, 0, 0, 0, 0, 0, 0, 0, 4, 24, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 24, 22, 17, 10, 0, 0, 0, 5, 0, 0, 0, 0, 15, 19, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 16, 17, 12, 8, 12, 16, 9, 0, 0, 0, 0, 0, 13, 20, 13, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 12, 16, 14, 14, 11, 10, 5, 0, 0, 0, 0, 0, 4, 22, 18, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 7, 5, 6, 5, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 16, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 9, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=151
    128, 128, 132, 128, 109, 87, 100, 99, 92, 91, 89, 98, 107, 119, 122, 130, 126, 125, 124, 124, 126, 127, 126, 122, 128, 131, 132, 120, 134, 131, 
    130, 130, 131, 129, 111, 81, 97, 93, 76, 86, 71, 73, 86, 85, 89, 106, 101, 118, 115, 121, 125, 130, 127, 122, 122, 119, 122, 129, 138, 126, 
    123, 124, 125, 124, 103, 56, 68, 63, 42, 60, 43, 43, 55, 47, 53, 69, 60, 83, 97, 109, 127, 135, 120, 120, 120, 114, 121, 140, 140, 125, 
    121, 120, 122, 117, 103, 51, 54, 52, 29, 44, 31, 35, 44, 38, 42, 48, 41, 53, 77, 106, 124, 137, 117, 116, 116, 110, 115, 138, 141, 134, 
    121, 120, 119, 107, 102, 61, 51, 65, 37, 47, 36, 39, 47, 39, 42, 42, 40, 48, 59, 94, 117, 122, 116, 113, 107, 106, 107, 129, 141, 142, 
    120, 122, 113, 96, 103, 60, 41, 73, 49, 57, 55, 45, 46, 36, 30, 33, 28, 35, 49, 65, 94, 109, 108, 103, 106, 112, 116, 122, 133, 140, 
    121, 122, 109, 96, 111, 51, 34, 66, 37, 40, 51, 30, 35, 35, 30, 37, 33, 31, 47, 44, 66, 103, 108, 105, 115, 117, 106, 104, 109, 129, 
    120, 120, 109, 94, 96, 37, 29, 62, 30, 39, 59, 34, 37, 37, 28, 35, 37, 32, 52, 40, 52, 96, 106, 118, 127, 122, 106, 114, 124, 136, 
    118, 120, 106, 71, 75, 25, 27, 47, 19, 23, 35, 18, 26, 26, 22, 26, 28, 25, 45, 40, 42, 75, 92, 106, 117, 117, 117, 129, 135, 133, 
    112, 117, 101, 69, 81, 31, 20, 18, 9, 14, 18, 12, 19, 16, 17, 14, 14, 14, 27, 27, 29, 43, 64, 93, 109, 114, 118, 122, 120, 118, 
    105, 105, 85, 70, 78, 20, 11, 9, 21, 24, 26, 19, 15, 8, 7, 4, 9, 21, 22, 18, 22, 28, 61, 98, 114, 114, 121, 120, 120, 120, 
    93, 82, 66, 61, 64, 12, 26, 30, 52, 35, 30, 23, 13, 12, 16, 21, 31, 44, 34, 25, 35, 42, 63, 82, 85, 94, 112, 115, 119, 120, 
    85, 65, 60, 53, 57, 31, 41, 33, 38, 11, 12, 4, 0, 0, 8, 13, 12, 11, 1, 5, 28, 42, 56, 67, 71, 75, 97, 107, 110, 120, 
    69, 38, 45, 45, 64, 61, 47, 26, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 21, 29, 34, 42, 46, 69, 101, 100, 116, 
    53, 21, 44, 56, 74, 55, 27, 21, 16, 0, 20, 22, 27, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 21, 26, 44, 89, 94, 111, 
    73, 35, 61, 70, 68, 21, 13, 28, 25, 20, 50, 36, 50, 31, 21, 37, 46, 45, 71, 62, 40, 53, 46, 57, 63, 46, 45, 75, 94, 103, 
    74, 26, 53, 67, 46, 0, 28, 42, 29, 14, 29, 15, 32, 14, 41, 64, 71, 70, 85, 69, 53, 76, 75, 85, 70, 39, 32, 46, 88, 95, 
    75, 25, 50, 63, 29, 2, 46, 40, 22, 5, 22, 18, 24, 13, 55, 44, 30, 32, 43, 29, 27, 39, 32, 57, 33, 9, 22, 36, 97, 95, 
    80, 26, 40, 49, 21, 10, 43, 23, 14, 7, 20, 24, 26, 22, 49, 23, 24, 42, 42, 32, 30, 35, 35, 51, 27, 10, 31, 44, 97, 91, 
    81, 29, 43, 44, 31, 22, 29, 10, 13, 7, 12, 19, 29, 20, 22, 11, 10, 8, 5, 2, 2, 17, 13, 12, 7, 17, 38, 41, 94, 90, 
    82, 25, 43, 44, 29, 32, 24, 13, 22, 15, 28, 32, 49, 15, 12, 31, 38, 27, 32, 38, 28, 57, 55, 13, 36, 46, 32, 26, 90, 91, 
    76, 16, 29, 44, 25, 39, 39, 19, 25, 23, 29, 21, 29, 0, 0, 41, 63, 33, 43, 55, 39, 68, 55, 0, 32, 37, 5, 3, 88, 91, 
    62, 5, 20, 38, 34, 54, 37, 19, 21, 22, 24, 15, 19, 0, 7, 34, 39, 20, 33, 48, 36, 52, 25, 0, 27, 28, 9, 26, 100, 86, 
    51, 18, 36, 61, 58, 66, 23, 15, 21, 22, 22, 21, 22, 14, 21, 20, 34, 66, 85, 96, 82, 85, 31, 20, 32, 20, 25, 43, 95, 77, 
    50, 43, 52, 59, 56, 58, 13, 27, 28, 21, 21, 21, 19, 20, 23, 18, 41, 87, 74, 70, 64, 65, 11, 10, 18, 22, 37, 45, 84, 70, 
    56, 49, 40, 32, 31, 56, 10, 36, 26, 15, 15, 24, 25, 27, 33, 36, 51, 73, 47, 46, 53, 55, 1, 11, 23, 32, 43, 39, 74, 66, 
    58, 48, 38, 32, 28, 49, 9, 34, 22, 12, 14, 27, 30, 30, 32, 31, 34, 40, 32, 44, 54, 51, 0, 16, 27, 34, 38, 34, 73, 64, 
    46, 44, 44, 40, 28, 31, 14, 33, 20, 15, 17, 26, 32, 30, 30, 29, 28, 28, 26, 29, 30, 26, 0, 8, 27, 33, 33, 39, 78, 62, 
    43, 41, 44, 45, 31, 19, 21, 31, 19, 17, 21, 27, 34, 34, 32, 30, 32, 30, 28, 28, 24, 22, 1, 7, 27, 34, 37, 59, 85, 62, 
    52, 50, 50, 46, 32, 9, 27, 25, 18, 23, 29, 34, 40, 37, 34, 35, 41, 42, 41, 42, 39, 37, 24, 23, 38, 46, 59, 78, 82, 57, 
    
    -- channel=152
    157, 158, 160, 161, 148, 133, 145, 162, 137, 112, 112, 119, 116, 116, 128, 139, 158, 169, 175, 182, 189, 196, 188, 169, 154, 169, 198, 194, 176, 172, 
    150, 151, 148, 149, 141, 108, 97, 121, 111, 90, 90, 99, 113, 129, 132, 144, 154, 164, 193, 210, 206, 201, 200, 186, 174, 184, 208, 214, 199, 182, 
    143, 145, 146, 148, 144, 96, 57, 59, 36, 23, 22, 18, 39, 64, 71, 94, 107, 124, 169, 205, 210, 198, 195, 189, 191, 203, 218, 242, 238, 201, 
    143, 144, 144, 144, 131, 79, 23, 2, 0, 0, 0, 0, 0, 0, 0, 0, 4, 35, 107, 159, 192, 198, 184, 180, 200, 212, 225, 253, 265, 228, 
    143, 143, 145, 141, 120, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 150, 186, 177, 166, 186, 200, 215, 242, 271, 255, 
    144, 144, 143, 131, 119, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 95, 167, 190, 169, 166, 185, 198, 217, 251, 259, 
    143, 145, 139, 116, 112, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 121, 193, 174, 163, 171, 179, 182, 208, 246, 
    145, 147, 136, 106, 95, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 140, 164, 158, 160, 159, 160, 171, 199, 
    147, 147, 137, 101, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 78, 137, 143, 148, 126, 120, 131, 144, 
    153, 150, 134, 73, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 107, 141, 146, 133, 123, 128, 135, 
    163, 154, 132, 72, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 100, 145, 149, 142, 143, 144, 144, 
    158, 153, 128, 101, 77, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 96, 147, 160, 152, 148, 145, 144, 
    143, 139, 115, 106, 102, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 71, 107, 131, 139, 145, 146, 143, 
    140, 124, 107, 99, 89, 73, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 41, 48, 72, 120, 142, 143, 
    137, 105, 90, 112, 117, 110, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 132, 144, 
    130, 83, 45, 90, 131, 136, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 108, 145, 
    105, 57, 20, 68, 117, 101, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 90, 146, 
    95, 53, 24, 78, 103, 46, 1, 12, 0, 0, 2, 20, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 85, 145, 
    94, 43, 8, 68, 93, 28, 0, 3, 0, 0, 0, 0, 0, 2, 9, 7, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 62, 134, 
    102, 41, 0, 30, 66, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 131, 
    99, 47, 0, 0, 30, 14, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 134, 
    69, 32, 0, 16, 18, 0, 0, 0, 0, 18, 27, 26, 5, 0, 0, 0, 38, 9, 0, 0, 0, 0, 8, 0, 0, 26, 11, 0, 31, 133, 
    29, 0, 0, 41, 49, 0, 0, 0, 0, 7, 21, 40, 57, 43, 0, 16, 76, 62, 19, 12, 0, 8, 55, 2, 0, 30, 38, 3, 46, 111, 
    0, 0, 0, 0, 44, 24, 0, 0, 0, 0, 12, 23, 34, 38, 18, 18, 43, 61, 46, 22, 11, 0, 18, 0, 0, 12, 9, 0, 36, 80, 
    0, 0, 0, 0, 0, 11, 1, 0, 0, 0, 0, 17, 26, 23, 21, 16, 19, 57, 64, 24, 7, 1, 0, 0, 0, 20, 8, 0, 8, 44, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 13, 30, 26, 21, 10, 14, 71, 105, 75, 51, 39, 7, 0, 0, 28, 18, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 27, 24, 24, 25, 18, 37, 61, 49, 35, 16, 0, 0, 5, 26, 19, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 24, 24, 21, 25, 26, 21, 13, 4, 4, 0, 0, 0, 5, 27, 21, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 13, 8, 5, 4, 2, 0, 0, 1, 4, 0, 0, 0, 25, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 0, 0, 
    
    -- channel=153
    1, 4, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 13, 17, 9, 4, 0, 0, 0, 0, 0, 0, 0, 7, 6, 0, 0, 2, 0, 6, 
    1, 4, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 6, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 19, 0, 0, 27, 18, 26, 25, 24, 33, 24, 12, 18, 7, 0, 4, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 0, 0, 35, 33, 34, 21, 11, 23, 29, 27, 27, 26, 25, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 15, 5, 17, 14, 0, 4, 14, 18, 21, 12, 26, 18, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 15, 0, 0, 13, 10, 19, 11, 0, 34, 12, 0, 8, 8, 1, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 15, 0, 0, 12, 3, 0, 10, 7, 7, 13, 0, 21, 25, 0, 10, 4, 0, 8, 18, 18, 15, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 1, 1, 0, 2, 0, 0, 3, 0, 2, 17, 0, 0, 0, 4, 3, 11, 5, 1, 0, 
    0, 0, 0, 3, 0, 4, 0, 0, 0, 5, 9, 10, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 3, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 17, 10, 10, 15, 21, 14, 3, 2, 11, 21, 23, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 15, 5, 12, 0, 5, 12, 7, 6, 7, 5, 0, 4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 27, 31, 28, 15, 16, 3, 0, 12, 11, 20, 31, 7, 0, 0, 2, 6, 13, 4, 0, 7, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 3, 6, 13, 34, 46, 40, 40, 28, 41, 48, 35, 44, 26, 10, 2, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 17, 0, 0, 0, 0, 12, 0, 5, 6, 0, 0, 0, 0, 0, 18, 
    0, 3, 0, 0, 0, 12, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 10, 0, 0, 0, 6, 0, 0, 0, 0, 0, 4, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 6, 0, 0, 16, 
    0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 19, 12, 0, 0, 5, 3, 0, 0, 0, 3, 20, 0, 0, 14, 15, 0, 0, 15, 
    0, 1, 0, 0, 3, 2, 12, 5, 0, 0, 0, 0, 0, 6, 0, 0, 15, 25, 6, 11, 18, 3, 27, 7, 0, 0, 0, 0, 0, 16, 
    0, 7, 0, 0, 11, 15, 18, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 6, 0, 0, 0, 0, 0, 15, 
    0, 29, 5, 0, 5, 5, 5, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 32, 16, 20, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 47, 39, 14, 0, 0, 7, 2, 8, 3, 0, 0, 0, 0, 0, 0, 0, 10, 34, 15, 10, 9, 11, 0, 0, 0, 3, 0, 0, 11, 
    0, 17, 18, 3, 0, 0, 11, 0, 8, 7, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 3, 0, 0, 8, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 1, 6, 0, 0, 1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 13, 
    0, 3, 5, 10, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 6, 0, 12, 
    7, 11, 10, 9, 13, 0, 0, 0, 0, 0, 2, 3, 2, 5, 3, 2, 4, 7, 3, 0, 0, 0, 11, 12, 0, 0, 10, 16, 0, 10, 
    
    -- channel=154
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=155
    394, 384, 393, 396, 386, 347, 313, 293, 287, 279, 283, 298, 297, 313, 345, 375, 409, 422, 418, 410, 412, 408, 406, 386, 364, 363, 373, 345, 322, 316, 
    425, 420, 417, 424, 404, 350, 302, 290, 299, 288, 304, 320, 329, 360, 379, 394, 413, 418, 422, 417, 399, 398, 414, 410, 402, 392, 388, 357, 353, 362, 
    444, 443, 443, 449, 428, 352, 272, 242, 244, 251, 255, 258, 274, 296, 307, 333, 347, 357, 363, 379, 376, 382, 409, 419, 414, 401, 380, 370, 380, 382, 
    456, 455, 455, 454, 425, 327, 239, 186, 168, 194, 195, 183, 196, 203, 212, 242, 250, 273, 294, 313, 349, 387, 404, 411, 409, 388, 360, 365, 382, 388, 
    455, 454, 457, 451, 405, 290, 198, 144, 131, 163, 173, 166, 168, 167, 166, 176, 176, 186, 229, 276, 326, 387, 402, 404, 399, 364, 333, 336, 363, 393, 
    454, 453, 456, 435, 395, 308, 198, 146, 159, 208, 223, 231, 229, 213, 198, 185, 180, 175, 181, 253, 328, 375, 394, 400, 374, 346, 318, 316, 341, 379, 
    453, 456, 447, 407, 384, 333, 208, 175, 219, 270, 275, 281, 267, 246, 241, 235, 228, 228, 221, 239, 289, 345, 387, 387, 365, 358, 335, 302, 299, 346, 
    453, 457, 438, 396, 379, 304, 186, 179, 235, 280, 305, 297, 257, 234, 229, 239, 242, 246, 261, 256, 254, 299, 353, 381, 398, 394, 364, 310, 286, 333, 
    449, 452, 438, 399, 344, 250, 163, 167, 191, 208, 242, 240, 219, 210, 210, 224, 238, 233, 248, 263, 253, 288, 341, 386, 414, 416, 374, 337, 333, 361, 
    435, 448, 434, 357, 287, 222, 148, 154, 159, 166, 187, 189, 186, 186, 193, 203, 213, 205, 223, 247, 245, 274, 326, 370, 415, 440, 420, 406, 409, 418, 
    418, 440, 417, 316, 260, 199, 126, 107, 114, 138, 152, 158, 167, 160, 159, 160, 159, 162, 188, 218, 222, 222, 260, 333, 414, 447, 455, 455, 455, 455, 
    392, 411, 373, 310, 275, 201, 101, 63, 103, 142, 155, 152, 151, 143, 130, 121, 128, 153, 176, 185, 184, 180, 221, 306, 385, 418, 431, 444, 454, 456, 
    364, 367, 310, 265, 250, 189, 127, 106, 124, 147, 167, 164, 138, 117, 110, 116, 137, 169, 167, 141, 138, 156, 207, 276, 334, 371, 392, 411, 443, 455, 
    341, 315, 247, 191, 191, 183, 199, 168, 147, 140, 132, 128, 104, 87, 90, 104, 122, 142, 132, 105, 99, 115, 150, 192, 227, 257, 310, 366, 422, 452, 
    310, 249, 189, 158, 193, 228, 214, 152, 118, 89, 77, 84, 78, 74, 73, 60, 43, 40, 28, 31, 50, 47, 57, 76, 108, 149, 214, 310, 395, 447, 
    294, 217, 143, 146, 224, 261, 172, 103, 87, 80, 77, 82, 83, 81, 54, 20, 15, 20, 25, 43, 54, 35, 28, 46, 92, 135, 175, 281, 371, 434, 
    300, 214, 137, 141, 215, 197, 106, 71, 94, 132, 150, 125, 123, 113, 56, 52, 80, 76, 113, 135, 95, 76, 68, 97, 156, 185, 194, 249, 332, 412, 
    324, 232, 158, 156, 186, 101, 47, 71, 101, 117, 141, 133, 150, 118, 117, 174, 193, 173, 204, 226, 196, 180, 166, 178, 215, 215, 186, 195, 296, 396, 
    324, 230, 148, 142, 138, 56, 28, 61, 71, 57, 63, 69, 89, 100, 166, 196, 196, 198, 213, 214, 203, 198, 192, 228, 225, 166, 128, 141, 256, 376, 
    330, 234, 127, 107, 99, 54, 32, 25, 31, 27, 20, 19, 36, 69, 133, 138, 122, 121, 128, 120, 112, 108, 117, 164, 142, 87, 87, 131, 244, 364, 
    339, 249, 127, 65, 77, 60, 29, 2, 6, 12, 17, 31, 59, 77, 83, 71, 82, 117, 116, 97, 94, 105, 123, 146, 112, 81, 116, 145, 228, 352, 
    339, 250, 145, 69, 62, 61, 47, 20, 0, 0, 18, 52, 92, 75, 23, 22, 75, 116, 109, 102, 102, 135, 168, 125, 77, 104, 132, 109, 196, 343, 
    326, 224, 117, 82, 62, 76, 97, 59, 8, 0, 0, 28, 86, 53, 0, 22, 113, 134, 135, 155, 149, 196, 236, 116, 51, 83, 90, 73, 185, 334, 
    301, 193, 85, 69, 95, 141, 147, 80, 22, 0, 0, 0, 0, 0, 0, 0, 56, 88, 156, 215, 217, 224, 213, 108, 31, 13, 12, 42, 184, 325, 
    276, 199, 126, 103, 127, 172, 163, 99, 39, 7, 0, 0, 0, 0, 0, 0, 0, 84, 189, 253, 252, 240, 169, 65, 0, 0, 0, 54, 185, 309, 
    274, 261, 217, 174, 150, 172, 155, 109, 62, 27, 0, 0, 0, 0, 0, 0, 13, 155, 255, 291, 281, 282, 188, 55, 0, 0, 20, 74, 183, 296, 
    288, 292, 261, 209, 166, 178, 140, 106, 81, 41, 0, 0, 0, 0, 0, 0, 33, 117, 175, 207, 227, 236, 155, 37, 0, 0, 32, 77, 178, 291, 
    279, 267, 244, 211, 168, 170, 117, 93, 77, 45, 1, 0, 0, 0, 0, 18, 40, 68, 90, 120, 160, 180, 101, 19, 0, 0, 29, 70, 177, 291, 
    259, 244, 229, 217, 181, 147, 88, 71, 64, 43, 8, 0, 0, 0, 1, 9, 21, 40, 62, 91, 122, 148, 83, 15, 0, 0, 21, 70, 200, 303, 
    246, 243, 241, 232, 190, 124, 73, 57, 47, 29, 18, 11, 10, 16, 21, 21, 29, 45, 64, 81, 98, 117, 87, 24, 0, 5, 31, 112, 243, 309, 
    
    -- channel=156
    74, 72, 75, 77, 78, 69, 54, 46, 47, 46, 49, 51, 44, 48, 56, 59, 71, 74, 71, 71, 71, 69, 72, 70, 66, 61, 57, 52, 50, 48, 
    86, 85, 82, 84, 82, 79, 61, 55, 62, 53, 65, 65, 59, 67, 68, 70, 81, 74, 73, 67, 65, 67, 74, 74, 72, 64, 59, 52, 55, 61, 
    91, 91, 91, 92, 89, 81, 59, 55, 63, 61, 67, 68, 68, 72, 69, 69, 71, 60, 55, 58, 58, 63, 74, 76, 74, 67, 56, 49, 52, 62, 
    97, 96, 96, 97, 93, 87, 70, 58, 64, 76, 75, 74, 80, 79, 80, 81, 76, 72, 54, 46, 57, 66, 75, 79, 73, 61, 52, 43, 46, 59, 
    96, 96, 97, 97, 85, 74, 72, 55, 62, 74, 80, 77, 78, 78, 79, 83, 80, 79, 75, 55, 48, 64, 74, 78, 73, 58, 50, 43, 43, 57, 
    96, 96, 99, 95, 81, 80, 70, 49, 58, 73, 79, 91, 89, 80, 78, 73, 76, 74, 70, 77, 62, 54, 66, 75, 67, 62, 52, 47, 44, 50, 
    96, 96, 97, 92, 84, 96, 71, 56, 64, 67, 60, 83, 92, 91, 94, 87, 85, 88, 76, 76, 72, 67, 68, 70, 67, 64, 53, 38, 37, 45, 
    95, 96, 94, 89, 82, 86, 66, 61, 85, 98, 92, 99, 96, 91, 91, 89, 87, 94, 90, 88, 75, 63, 68, 77, 80, 75, 70, 55, 51, 58, 
    94, 96, 96, 96, 79, 82, 64, 58, 71, 81, 83, 87, 86, 84, 84, 84, 85, 87, 86, 91, 83, 70, 67, 71, 80, 85, 77, 70, 65, 68, 
    91, 94, 95, 94, 85, 90, 61, 53, 53, 64, 72, 75, 77, 78, 78, 79, 78, 79, 80, 84, 82, 77, 74, 72, 84, 92, 85, 79, 78, 83, 
    87, 92, 90, 70, 62, 76, 54, 44, 45, 56, 67, 75, 72, 67, 66, 66, 66, 69, 75, 77, 70, 64, 67, 75, 89, 95, 96, 96, 96, 97, 
    79, 86, 79, 64, 56, 64, 40, 48, 55, 60, 67, 72, 76, 69, 60, 59, 63, 68, 69, 63, 53, 42, 42, 49, 65, 76, 82, 92, 96, 96, 
    79, 81, 65, 57, 54, 53, 45, 54, 54, 63, 70, 69, 62, 59, 54, 51, 53, 57, 50, 41, 38, 34, 42, 52, 67, 75, 70, 76, 92, 96, 
    72, 69, 44, 26, 35, 45, 63, 65, 58, 57, 47, 47, 38, 39, 40, 42, 49, 56, 50, 41, 36, 38, 45, 51, 59, 68, 74, 70, 87, 96, 
    55, 57, 39, 21, 26, 41, 57, 63, 45, 49, 46, 50, 42, 36, 29, 16, 10, 10, 10, 16, 18, 8, 9, 16, 38, 56, 67, 69, 84, 96, 
    65, 60, 35, 23, 36, 52, 40, 43, 32, 32, 26, 38, 36, 38, 27, 18, 17, 22, 20, 28, 35, 22, 19, 28, 42, 52, 63, 67, 75, 93, 
    63, 54, 24, 12, 38, 47, 30, 24, 26, 33, 26, 23, 29, 33, 17, 21, 25, 20, 27, 27, 23, 22, 18, 29, 47, 53, 49, 50, 59, 85, 
    72, 65, 35, 15, 31, 27, 16, 19, 19, 34, 40, 33, 32, 25, 24, 40, 38, 29, 39, 48, 41, 32, 27, 28, 49, 57, 46, 48, 57, 83, 
    72, 66, 37, 15, 17, 16, 8, 15, 15, 23, 29, 26, 31, 33, 34, 48, 68, 71, 73, 70, 68, 67, 65, 68, 64, 57, 46, 41, 47, 78, 
    71, 66, 38, 24, 16, 14, 7, 4, 4, 2, 6, 12, 21, 27, 37, 35, 34, 38, 39, 37, 36, 33, 38, 46, 39, 34, 40, 44, 42, 71, 
    76, 68, 29, 10, 21, 13, 7, 1, 0, 0, 0, 9, 22, 33, 29, 15, 24, 48, 48, 41, 42, 38, 44, 62, 35, 22, 41, 43, 38, 68, 
    80, 70, 34, 0, 9, 20, 18, 9, 0, 0, 0, 0, 5, 9, 4, 0, 1, 22, 26, 25, 29, 26, 28, 31, 15, 14, 21, 21, 32, 70, 
    85, 69, 33, 7, 0, 19, 34, 18, 1, 0, 0, 0, 11, 5, 0, 0, 6, 11, 23, 31, 34, 44, 49, 23, 12, 17, 21, 22, 33, 72, 
    87, 67, 41, 24, 24, 31, 40, 24, 8, 0, 0, 0, 0, 0, 0, 0, 5, 19, 53, 72, 69, 68, 76, 40, 5, 0, 0, 13, 36, 76, 
    82, 67, 52, 39, 33, 38, 49, 33, 14, 3, 0, 0, 0, 0, 0, 0, 0, 0, 24, 43, 46, 49, 42, 15, 0, 0, 0, 15, 41, 79, 
    76, 73, 61, 52, 44, 39, 49, 33, 19, 6, 0, 0, 0, 0, 0, 0, 0, 23, 43, 57, 62, 67, 51, 12, 0, 0, 0, 20, 44, 78, 
    81, 80, 74, 66, 54, 42, 38, 29, 23, 10, 0, 0, 0, 0, 0, 0, 0, 19, 43, 57, 64, 67, 52, 11, 0, 0, 3, 19, 45, 80, 
    81, 82, 74, 64, 50, 44, 32, 26, 22, 10, 0, 0, 0, 0, 0, 0, 5, 14, 22, 31, 41, 47, 31, 12, 0, 0, 3, 16, 46, 81, 
    81, 79, 73, 70, 61, 44, 23, 18, 17, 8, 0, 0, 0, 0, 0, 0, 1, 8, 16, 23, 32, 39, 23, 7, 0, 0, 0, 19, 58, 88, 
    81, 82, 80, 76, 64, 48, 23, 9, 7, 2, 1, 0, 0, 3, 4, 4, 6, 13, 21, 26, 30, 34, 27, 9, 0, 0, 4, 33, 69, 89, 
    
    -- channel=157
    468, 462, 465, 469, 461, 408, 342, 305, 320, 345, 350, 360, 382, 410, 436, 465, 473, 477, 470, 459, 446, 439, 449, 454, 450, 424, 400, 371, 364, 360, 
    511, 507, 508, 513, 498, 426, 350, 294, 284, 313, 312, 318, 327, 341, 375, 404, 417, 439, 422, 412, 406, 417, 438, 459, 465, 440, 402, 377, 388, 406, 
    532, 530, 530, 529, 495, 395, 298, 227, 217, 238, 234, 238, 230, 224, 238, 259, 281, 312, 323, 336, 358, 400, 433, 457, 453, 422, 381, 359, 380, 420, 
    537, 534, 537, 530, 501, 384, 259, 178, 174, 218, 218, 228, 231, 217, 211, 205, 202, 204, 210, 261, 327, 405, 447, 460, 434, 395, 343, 318, 340, 401, 
    536, 535, 533, 516, 490, 401, 293, 224, 215, 294, 305, 312, 323, 318, 318, 297, 268, 261, 232, 243, 313, 405, 464, 472, 430, 376, 312, 281, 293, 367, 
    535, 535, 525, 493, 465, 389, 314, 278, 289, 392, 433, 421, 394, 371, 364, 363, 348, 340, 340, 314, 307, 354, 417, 452, 435, 388, 342, 300, 280, 330, 
    535, 535, 521, 486, 460, 385, 311, 272, 275, 362, 414, 416, 401, 358, 342, 354, 361, 359, 367, 364, 340, 327, 358, 422, 436, 424, 380, 322, 277, 292, 
    533, 533, 518, 476, 434, 359, 278, 263, 263, 310, 327, 337, 352, 333, 329, 343, 355, 356, 373, 368, 360, 366, 378, 438, 477, 477, 431, 371, 336, 353, 
    526, 531, 512, 436, 373, 276, 230, 237, 248, 293, 294, 284, 296, 299, 307, 318, 326, 328, 346, 362, 369, 376, 387, 439, 498, 509, 501, 478, 467, 477, 
    502, 523, 507, 441, 368, 268, 211, 171, 171, 219, 246, 245, 249, 258, 266, 268, 266, 264, 277, 307, 327, 336, 343, 384, 460, 513, 529, 530, 533, 533, 
    467, 494, 470, 418, 381, 312, 224, 134, 109, 161, 232, 245, 239, 221, 209, 206, 207, 224, 237, 246, 247, 255, 297, 354, 447, 515, 538, 536, 537, 537, 
    431, 436, 407, 348, 318, 273, 236, 179, 180, 206, 255, 280, 274, 240, 204, 207, 232, 276, 289, 267, 222, 200, 245, 312, 383, 438, 485, 514, 533, 536, 
    412, 390, 352, 290, 266, 235, 229, 224, 249, 245, 250, 245, 242, 222, 187, 184, 203, 230, 228, 203, 166, 147, 179, 225, 274, 309, 368, 442, 506, 537, 
    404, 338, 260, 217, 254, 279, 273, 254, 212, 179, 145, 113, 106, 115, 112, 114, 117, 119, 98, 79, 76, 77, 100, 121, 161, 198, 254, 351, 454, 528, 
    369, 277, 191, 149, 224, 287, 284, 227, 173, 166, 148, 121, 109, 97, 66, 30, 0, 0, 1, 4, 1, 0, 0, 15, 76, 146, 225, 313, 416, 511, 
    373, 280, 217, 170, 219, 214, 183, 145, 147, 181, 212, 216, 226, 176, 130, 82, 56, 61, 109, 136, 135, 93, 42, 71, 137, 219, 287, 335, 415, 489, 
    401, 295, 228, 194, 213, 149, 82, 63, 134, 171, 170, 182, 224, 209, 221, 215, 237, 255, 280, 295, 304, 276, 235, 266, 285, 290, 289, 290, 367, 447, 
    417, 297, 206, 161, 166, 112, 51, 25, 91, 119, 93, 64, 93, 126, 205, 245, 277, 247, 255, 260, 257, 251, 235, 285, 292, 264, 206, 184, 295, 412, 
    424, 309, 193, 103, 86, 70, 46, 16, 36, 58, 63, 46, 49, 52, 132, 196, 230, 211, 200, 202, 198, 189, 185, 210, 218, 195, 145, 141, 271, 401, 
    421, 327, 221, 95, 51, 45, 39, 2, 0, 0, 33, 54, 81, 77, 84, 81, 120, 146, 141, 127, 117, 135, 139, 149, 138, 138, 167, 181, 281, 390, 
    420, 320, 229, 130, 78, 67, 41, 5, 0, 0, 0, 55, 154, 140, 97, 52, 93, 155, 168, 147, 133, 179, 217, 181, 136, 123, 186, 216, 279, 366, 
    421, 307, 185, 97, 90, 119, 97, 55, 4, 0, 0, 0, 79, 90, 62, 20, 87, 182, 231, 214, 202, 249, 264, 217, 142, 61, 99, 139, 228, 347, 
    408, 286, 153, 30, 43, 150, 174, 132, 41, 0, 0, 0, 0, 0, 0, 0, 14, 85, 153, 190, 208, 235, 195, 126, 62, 10, 9, 44, 183, 340, 
    393, 313, 205, 109, 85, 172, 203, 168, 68, 0, 0, 0, 0, 0, 0, 0, 0, 72, 204, 319, 331, 341, 239, 109, 7, 0, 0, 43, 190, 340, 
    378, 359, 323, 256, 204, 216, 192, 173, 96, 30, 0, 0, 0, 0, 0, 0, 0, 87, 244, 379, 393, 375, 269, 135, 0, 0, 0, 67, 216, 346, 
    377, 378, 365, 319, 247, 234, 183, 177, 108, 62, 0, 0, 0, 0, 0, 0, 16, 98, 173, 254, 285, 300, 208, 91, 0, 0, 0, 79, 224, 344, 
    377, 374, 346, 306, 246, 218, 160, 152, 102, 67, 7, 0, 0, 0, 0, 0, 17, 73, 106, 154, 207, 254, 175, 66, 0, 0, 0, 76, 220, 339, 
    367, 348, 325, 299, 251, 196, 123, 104, 83, 58, 13, 0, 0, 0, 0, 0, 0, 26, 61, 106, 155, 199, 150, 60, 0, 0, 0, 70, 218, 343, 
    344, 333, 327, 314, 264, 185, 101, 62, 63, 44, 13, 0, 0, 0, 0, 0, 9, 28, 53, 81, 110, 138, 107, 51, 0, 0, 0, 99, 247, 371, 
    355, 359, 360, 345, 304, 197, 103, 29, 29, 29, 20, 17, 24, 29, 35, 40, 55, 79, 103, 120, 130, 141, 117, 78, 29, 7, 61, 174, 314, 408, 
    
    -- channel=158
    44, 32, 47, 64, 48, 17, 40, 65, 55, 48, 46, 43, 26, 19, 27, 40, 61, 65, 59, 48, 60, 74, 71, 35, 6, 13, 36, 16, 5, 20, 
    55, 50, 50, 62, 43, 2, 29, 86, 96, 98, 109, 107, 125, 135, 122, 124, 113, 91, 82, 71, 69, 81, 88, 68, 48, 31, 38, 34, 37, 44, 
    73, 71, 72, 78, 57, 8, 45, 118, 114, 136, 142, 121, 161, 179, 168, 189, 165, 140, 116, 85, 80, 92, 89, 80, 76, 47, 29, 52, 69, 54, 
    88, 87, 87, 86, 60, 0, 35, 135, 123, 132, 134, 103, 125, 130, 133, 175, 172, 170, 158, 111, 90, 100, 83, 69, 74, 47, 26, 65, 95, 73, 
    88, 89, 91, 87, 57, 0, 0, 78, 101, 84, 78, 62, 70, 58, 49, 76, 91, 101, 124, 130, 117, 109, 78, 57, 59, 44, 28, 60, 104, 103, 
    88, 89, 90, 80, 79, 11, 0, 49, 102, 67, 42, 40, 70, 78, 62, 54, 57, 62, 65, 101, 135, 143, 107, 67, 41, 29, 6, 22, 85, 126, 
    86, 90, 80, 57, 81, 52, 0, 94, 162, 133, 104, 73, 83, 120, 125, 111, 97, 96, 96, 80, 96, 146, 143, 87, 46, 25, 0, 0, 55, 126, 
    88, 92, 71, 46, 84, 57, 8, 121, 181, 166, 188, 140, 92, 121, 131, 131, 121, 108, 137, 114, 62, 103, 129, 83, 60, 38, 5, 0, 22, 82, 
    93, 91, 71, 55, 97, 79, 40, 129, 145, 111, 162, 150, 112, 125, 132, 134, 136, 116, 137, 142, 85, 101, 128, 103, 83, 57, 0, 0, 0, 29, 
    107, 94, 69, 23, 53, 68, 48, 140, 167, 128, 136, 138, 131, 134, 138, 141, 146, 139, 156, 169, 132, 128, 165, 165, 131, 89, 43, 32, 43, 54, 
    126, 108, 72, 7, 26, 25, 12, 99, 161, 146, 119, 105, 108, 121, 133, 135, 133, 134, 140, 153, 155, 138, 151, 172, 153, 106, 87, 89, 89, 88, 
    134, 121, 81, 60, 87, 38, 0, 32, 89, 109, 106, 95, 74, 83, 105, 106, 98, 99, 80, 71, 107, 116, 125, 162, 165, 133, 113, 101, 90, 88, 
    118, 103, 69, 69, 100, 57, 18, 38, 70, 91, 116, 129, 89, 70, 88, 102, 112, 129, 105, 61, 76, 108, 144, 181, 187, 173, 170, 147, 105, 88, 
    87, 64, 70, 74, 74, 36, 29, 76, 116, 113, 127, 163, 146, 113, 111, 131, 152, 170, 158, 118, 108, 120, 143, 168, 179, 176, 202, 207, 144, 92, 
    81, 31, 56, 101, 102, 62, 23, 56, 110, 91, 71, 87, 97, 89, 79, 100, 118, 117, 116, 102, 97, 112, 132, 155, 176, 153, 166, 220, 181, 106, 
    61, 0, 0, 83, 136, 107, 50, 68, 81, 44, 14, 0, 0, 13, 0, 15, 35, 22, 29, 16, 0, 11, 42, 69, 109, 100, 100, 175, 186, 123, 
    37, 0, 0, 75, 112, 53, 55, 116, 95, 73, 97, 70, 52, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 61, 84, 153, 197, 151, 
    50, 0, 7, 111, 96, 0, 16, 132, 125, 88, 121, 139, 149, 103, 71, 65, 42, 51, 105, 109, 51, 43, 45, 64, 77, 67, 110, 165, 221, 181, 
    46, 0, 0, 120, 108, 0, 0, 103, 128, 81, 59, 84, 126, 123, 171, 162, 100, 116, 152, 145, 128, 135, 133, 163, 135, 56, 77, 137, 215, 193, 
    63, 0, 0, 67, 95, 22, 13, 52, 92, 92, 61, 45, 54, 71, 146, 165, 106, 87, 109, 112, 102, 104, 98, 129, 130, 62, 45, 91, 194, 201, 
    80, 0, 0, 8, 43, 35, 23, 9, 46, 82, 88, 70, 50, 14, 34, 120, 130, 78, 63, 78, 72, 83, 71, 34, 73, 104, 65, 56, 177, 213, 
    85, 0, 0, 45, 35, 20, 16, 0, 0, 34, 84, 113, 121, 41, 0, 66, 119, 39, 0, 20, 12, 46, 57, 0, 0, 140, 128, 77, 188, 225, 
    95, 0, 0, 91, 89, 42, 15, 0, 0, 9, 60, 110, 168, 108, 17, 75, 177, 129, 62, 78, 55, 92, 134, 4, 5, 129, 132, 102, 209, 232, 
    104, 0, 0, 25, 94, 100, 48, 0, 0, 0, 17, 42, 80, 71, 42, 67, 144, 150, 88, 54, 30, 46, 48, 0, 24, 66, 63, 82, 205, 231, 
    108, 10, 0, 0, 35, 111, 68, 0, 0, 0, 0, 14, 26, 32, 39, 34, 65, 134, 101, 31, 13, 18, 0, 0, 14, 56, 62, 83, 187, 219, 
    106, 73, 13, 0, 29, 95, 54, 17, 24, 0, 0, 3, 23, 27, 33, 17, 45, 174, 209, 161, 127, 114, 1, 0, 4, 54, 86, 101, 178, 210, 
    106, 107, 85, 53, 38, 92, 55, 33, 57, 10, 0, 0, 11, 18, 32, 41, 59, 135, 174, 165, 154, 127, 0, 0, 1, 50, 96, 109, 180, 205, 
    109, 101, 85, 62, 33, 73, 61, 56, 65, 26, 0, 0, 14, 23, 38, 63, 82, 100, 110, 123, 141, 129, 0, 0, 3, 57, 92, 109, 184, 195, 
    108, 99, 86, 74, 34, 27, 48, 71, 59, 33, 13, 7, 17, 27, 29, 36, 52, 68, 82, 104, 126, 134, 33, 0, 0, 55, 79, 104, 180, 175, 
    98, 90, 80, 73, 34, 0, 19, 72, 61, 37, 24, 15, 17, 24, 22, 24, 34, 40, 44, 57, 71, 83, 40, 0, 0, 30, 58, 100, 159, 144, 
    
    -- channel=159
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end gold_package;
