library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -5828, 151, 1948, 1856, 25, -2849, 4756, 864, -3720, -2174,

    -- weights
    -- filter=0 channel=0
    2, 0, -13, 1, 1, -3, -9, -1, -8, 4, -4, 0, -10, -8, -5, -6, -16, -19, -19, -14, 0, -6, -6, -6, -5, -10, 6, -6, -6, 4, -9, -15, -16, -1, -11, -14, -6, -14, -2, -8, 5, 7, -6, -9, -7, -15, -11, -7, -8, -8, -3, 1, -13, -7, -3, -8, -9, 3, -6, 4, -17, -9, 0, -14, -2, -13, -16, -13, -20, -11, -8, 5, 5, 4, -3, -14, -10, -10, -4, -6, -3, -12, -14, -5, -19, -11, -5, 4, -1, -4, -11, -5, -8, -7, -10, -19, -9, -14, -28, -15, -21, -10, 1, -4, 0, -1, -22, -2, -14, -14, -16, -17, -20, -33, -17, -20, -2, -3, 1, 5, -17, -5, -16, 0, -12, -14, -7, -11, -16, -25, -14, 0, -3, -2, -7, -3, -10, -16, -4, -16, -5, -15, -11, -21, -12, -19, -9, -8, 4, -9, -5, -18, -17, -14, -15, -6, -10, -19, -22, -22, -5, -8, -2, -7, 7, -10, -12, -21, -11, -7, -13, 0, -12, -8, -9, -10, 5, 10, 4, 1, -3, -19, -18, -2, -1, -16, -11, 0, -9, 3, -10, 9, 9, 1, -3, -12, -21, -10, -14, -17, -16, 2, 1, -6, -7, -1, 8, -7, 1, -2, 1, -15, -17, -13, -11, -5, -11, -4, -4, 3, 2, -5, -8, 1, 2, 11, 10, 8, 3, 1, 9, 16, 16, 12, 9, 11, 3, 7, 10, 11, 2, 14, 15, 14, 8, 5, 12, 24, 11, 14, 21, 19, 17, 10, 1, 14, 19, 16, 11, 19, 20, 16, 9, 6, 19, 17, 14, 20, 12, 12, 2, 10, 25, 24, 9, 5, 13, 6, 3, 18, 25, 26, 16, 12, 19, 5, 18, 15, 17, 23, 18, 3, 3, 8, 11, 20, 28, 24, 19, 10, 9, 5, 21, 16, 18, 6, 6, -3, 5, 2, 14, 22, 27, 12, 22, 7, 13, 21, 17, 28, 14, -1, -1, -13, -3, 9, 17, 21, 17, 21, 10, 9, 20, 23, 24, 16, 6, -7, -20, -11, 1, 19, 21, 30, 23, 3, 22, 16, 17, 28, 11, 10, -16, -14, -4, 8, 18, 28, 16, 7, 18, 6, 12, 13, 29, 22, 1, -3, 0, -7, 13, 18, 27, 17, 6, 19, 11, 13, 21, 9, 17, 8, -1, 10, 0, 9, 15, 30, 15, 12, 12, 19, 28, 27, 14, 15, 6, -1, 5, 19, 28, 14, 20, 17, 13, 9, 6, 18, 23, 20, 4, 13, 16, 4, 10, 23, 34, 20, 11, 11, 9, 16, 13, 18, 21, 19, 6, 18, 10, 28, 22, 30, 16, 2, 5, 9, 16, 21, 3, 12, 5, 4, 6, 3, 13, 10, 5, 1, 2, 4, -1, 2, 7, 1, -6, -9, 1, -8, 0, 8, 4, 5, -4, -3, 4, 6, -5, -2, 8, 3, 6, 2, 0, 10, 3, 10, -8, 7, 8, -5, 6, 0, 4, -7, -4, -6, -5, -1, -1, 5, 3, -3, -1, 6, -2, -7, -10, 1, 8, 0, 5, 4, 0, 4, -3, 1, -5, -6, 0, -1, 0, -3, -5, -7, 0, -9, 4, 0, 4, -4, 2, 5, -3, -9, -7, -8, 3, 7, -2, 0, 3, -11, -5, 1, -7, -6, -3, -1, 0, 1, 4, -7, 1, -5, -6, 0, 4, -12, 0, -14, -3, 7, 3, 9, 2, -7, -6, 0, 2, 1, 0, -8, 1, -10, -13, -1, 4, 2, -2, 5, -5, 4, 0, -9, 7, 4, -3, -6, -13, -10, -10, -7, -8, 3, 1, -1, 3, -10, 2, 4, 6, -7, -8, 3, -10, -5, -8, 9, 6, -4, -7, -1, -1, 7, 6, 3, -6, 3, -7, -9, 5, -9, 9, 3, -5, 8, -7, -6, 7, 7, 8, -8, 0, -9, 3, -4, 0, 6, -2, -8, -9, 1, 6, -6, -8, -1, 2, -5, -6, -4, 5, 7, -5, -6, 3, 9, -8, 5, 4, -1, -6, 3, 2, -3, -7, -6, 3, -8, -8, 2, -5, 7, 0, -3, -8, 7, -8, 1, -4, 0, 6, -2, 3, -8, 6,
    -- filter=0 channel=1
    13, 1, 13, 0, 0, 14, 12, 3, 8, -4, 5, 5, -1, 15, 13, 5, 12, 5, 8, 6, 12, 14, 13, 1, 3, -5, 3, 9, 12, 5, 0, 9, 10, 10, 0, -4, 6, 1, 1, -4, -8, -5, -8, -2, 10, 2, 12, 6, 4, -9, -6, 14, 2, 3, -9, -17, -20, -11, -5, 0, 8, 14, 3, -6, -8, -11, 10, 3, 7, -3, -11, -20, -7, -5, -6, 11, 0, 8, -9, -17, -4, 8, 9, -6, -5, -9, -14, -12, -19, -8, 15, 0, 9, -10, -7, -6, 0, 9, 5, -15, -8, -13, -27, -14, -7, 8, 10, -2, -7, -26, -9, -5, 3, 2, -10, -20, -21, -24, -6, -4, 2, 3, 3, 0, -19, -9, -6, 5, 0, -9, -21, -14, -23, -9, -11, 10, 9, -3, -6, -20, -18, -6, 16, 4, -11, -20, -25, -10, -16, 3, 12, 2, -5, -10, -17, 0, -7, 13, -4, -1, -6, -9, -18, -10, -5, 18, 1, 0, -6, -7, -1, 5, 12, 5, -17, -9, -18, -12, -13, 7, 11, 17, 16, 0, 0, -5, 11, 6, 0, -13, -12, -15, -6, -1, 13, 6, 14, 17, 14, 3, 4, 1, 2, 3, -7, -12, -13, -5, 1, 17, 6, 0, 3, 8, 8, 1, 8, 11, 4, -6, -8, 3, -4, 10, 12, -16, -5, -6, -15, 0, 2, -6, -5, -6, 5, 0, 6, -4, -1, 14, 0, -18, -9, -16, -3, -4, 0, 14, 15, 8, -4, -5, 1, -1, 14, -7, -9, -8, -4, -11, 10, 21, 14, 8, 10, 2, 0, -4, 4, 15, -8, -15, -21, -16, -5, 2, 29, 27, 26, 7, 0, -5, -3, -8, 0, -6, -11, -15, -18, 1, 19, 23, 27, 28, 3, 10, 0, -1, 1, 4, -7, -5, -9, -1, -5, 12, 34, 30, 23, 25, 0, -1, -17, -6, 5, -7, -3, -9, -5, 2, 22, 44, 43, 43, 14, 5, -8, -15, -3, -2, -4, -21, -9, 5, 10, 26, 38, 51, 41, 26, 15, -1, -9, -16, -9, -1, -9, -7, 4, 4, 28, 39, 42, 33, 22, -4, -4, -9, -5, -3, -3, -5, -9, -5, 0, 29, 47, 39, 39, 21, 9, -9, -14, -14, -11, -1, -17, -13, -5, 0, 11, 36, 36, 33, 7, 9, -10, -8, -15, 0, -9, -4, -3, -19, 3, 1, 19, 36, 17, 13, 4, 0, -3, 0, 7, -7, -15, -5, -13, -8, 1, 27, 24, 11, 7, -4, -2, -8, -5, 6, -4, -12, -20, -5, -8, -7, 15, 22, 19, 10, -5, 6, 4, 6, 7, -7, 0, -19, -11, -9, -1, 3, 4, 10, 1, 8, 5, 9, 2, 13, 2, -4, 2, -1, 2, 1, 7, -2, 8, 2, 5, 0, 1, 6, 11, 9, 10, 5, 6, 5, -2, -1, 7, -2, 7, -2, 2, 7, -4, 11, 0, -5, 5, 0, 3, 6, 4, 6, -2, -8, -12, 0, -9, 5, 0, -6, 4, 6, -3, -12, 4, 6, 0, -3, -7, -5, -9, -1, -10, -5, 9, 10, 3, -6, 2, -5, 0, 7, -9, -3, 4, 0, -2, 1, -1, 7, -6, -5, -1, 0, 0, -2, -6, 4, -10, 2, 2, 0, -4, -10, -6, -5, 2, 0, -14, -15, 5, -2, -1, -10, 5, 3, -1, -6, 0, 9, 8, -1, -5, -18, -7, 4, 2, -2, -6, -8, -7, -11, -6, -11, 2, 10, 4, -5, -9, -8, -1, 2, -8, 0, 3, -15, -11, -12, -11, 9, 0, -6, -5, -4, -14, -4, 0, 8, 3, -12, -5, -8, 0, -2, -7, -4, -4, 4, 1, -3, -5, -7, 2, -9, 0, -10, -8, -13, 2, 6, -6, 2, -3, 1, -4, 4, 1, 3, 5, -6, -3, -11, -6, -5, 0, 8, -3, -3, -11, -6, 9, -4, 5, 4, -13, -15, -13, 3, 8, -5, 5, 8, 0, 1, 0, 3, 6, -3, -1, -9, -11, -4, -9, -5, -5, -3, -1, -6, 3, 2, 4, -3, 5, 4, -10, 7, -6, 0, -1,
    -- filter=0 channel=2
    -8, 9, 3, 0, 5, 1, -3, 6, -8, 4, -7, 9, 7, 0, 0, 7, -5, -6, 1, -4, -5, -7, 3, 0, 4, -7, 0, 9, -4, 6, -1, 3, 5, -8, 3, -6, -6, 0, 5, -5, 0, 7, -4, -5, -6, -5, -1, -4, -7, -2, 5, 0, 5, 7, 8, -2, 4, 0, -6, -7, 5, 8, 3, -2, 2, 5, -4, -7, 1, -3, -5, 7, -1, -8, -8, -8, -5, 0, -4, 4, 7, -3, -6, -10, -8, -10, -1, 0, 9, -9, 7, -1, 8, 2, -4, -5, -3, 0, 0, 0, -1, -6, 5, -8, 1, -6, -4, 7, 0, 0, 7, 0, 7, 2, -1, 4, -2, -9, -4, -6, -5, -2, 2, -4, -9, 2, -10, 2, 0, -5, -7, 5, 5, 5, -4, 0, -1, 0, -3, 2, 6, 3, -10, -3, 7, 0, -6, 0, 3, -4, 5, 4, 8, 0, -8, 5, 5, -2, -3, -9, -5, 2, 1, -3, 0, 8, 5, -2, -8, -4, -2, -6, -5, -5, 5, -3, -3, 9, 7, 0, 9, 0, -2, -7, 0, -3, -5, -1, -8, -1, -8, 1, 0, -8, -2, 9, 2, -4, 9, 8, 0, 4, -3, 6, 8, 0, -5, 3, -6, 1, -1, -3, 2, -8, -6, 3, -7, 9, 3, 2, -8, 6, -3, 1, 0, -2, -4, 2, 2, -8, -12, 1, -11, -6, -6, -6, 2, -9, 1, -2, -3, 5, 5, 0, -1, -12, -6, -5, -3, -6, -13, -10, 3, -4, 2, -11, 2, 0, 5, -1, -10, -5, 5, 6, 4, 0, -12, 1, -7, -9, -10, -8, -2, -4, -10, 2, -4, 5, 1, -4, 5, -8, 1, 0, -11, 2, -3, -4, -10, -12, 2, 0, 1, -11, -3, -1, 2, -10, -3, -11, 2, -5, 1, 0, -3, -3, 4, -3, 1, 2, -9, 2, -8, -8, 6, 4, 1, -13, 6, 4, -4, -7, 6, -8, -10, -2, 5, -7, -4, -6, -9, -6, -2, 2, 7, 6, 5, -9, -7, 5, -6, 0, -1, -7, -10, 4, -10, -5, -8, 4, -11, -5, 0, 4, 0, 3, -6, 2, 4, -4, -6, -13, -8, -1, -2, -4, 3, 7, -11, -1, 6, 1, 4, 0, -2, 6, -9, 0, 2, -11, -5, -11, 5, 2, -10, 1, 0, -11, -10, -4, 2, -11, -13, -4, -6, -9, -9, 3, 4, -5, 2, 5, -9, -3, -2, -9, -10, -9, -5, -4, -1, 2, -5, 4, -4, 2, 0, -3, -9, -11, -6, -5, -13, -6, 2, 3, -12, 0, 3, 1, 1, -6, -4, -6, 5, 1, -6, -10, 4, -6, 0, -5, 3, -10, -3, -5, 4, -10, -6, -8, 8, -1, 0, 2, 1, -3, -9, -2, -5, 4, -6, -1, -8, -2, -6, -4, 0, 4, -7, -1, -2, 0, 6, -3, 7, 5, -3, -5, 8, 6, 0, 7, -1, -3, 3, -6, 6, 3, 3, 2, 1, -8, -5, -6, 2, -8, -7, 7, 5, 6, 5, 0, 7, 1, 7, -9, 6, 0, 6, -2, -8, 7, -6, 0, -7, -2, 1, -8, -1, 0, -9, 1, -1, -2, 0, -5, 1, 4, 0, -5, -5, 3, -9, 1, -4, 1, -4, 1, -3, 0, -5, -3, 9, -1, -3, -1, 3, -10, 2, 7, -8, -2, -4, 1, 7, 5, -6, -6, 4, 0, -6, -10, -7, -2, -3, 1, 4, -6, -5, -3, 3, 7, 3, -3, 2, -8, -5, -4, -9, 4, -6, -9, -7, 9, 0, 1, 4, -8, 5, -5, 0, 8, 3, -2, 7, 1, 7, 0, -2, 6, -6, -2, -6, -6, 2, 6, 3, 5, -1, -9, -7, 5, 5, -4, -2, -5, 8, 0, -9, 2, -9, -8, 0, 3, -3, -10, 5, 7, -4, 0, -2, -4, 0, -2, -4, 8, 2, -7, 4, 1, 3, 6, 1, 6, 4, 5, 2, -9, -7, 5, 1, -5, -1, 2, 5, -1, -1, -1, 6, -8, -3, -7, 0, 0, 9, 7, -1, 8, 0, -6, 6, 6, 3, -4, -7,
    -- filter=0 channel=3
    11, 9, 8, 2, 14, 10, 7, 5, -2, 0, -1, -9, -7, -6, -8, 2, -1, 5, -1, 17, 11, 9, -4, 9, -3, -6, 9, -2, 0, -4, -6, 0, 1, 3, 1, 9, 11, 8, 3, 9, -3, 2, 0, 7, -6, 8, 9, 2, 2, 13, 12, -5, -6, 5, 9, -3, -6, 1, 5, -1, -1, 5, -1, 8, 2, 0, -6, -5, -1, 1, 8, 2, -3, 12, 0, -5, 0, -6, -2, 0, -7, -4, -11, 6, 5, 10, -2, 8, 4, 8, 6, 4, -9, -8, -2, -3, -1, 3, 6, 8, 6, 6, 8, 6, 6, -9, -4, 2, -13, -15, -7, -8, 5, 0, 9, 9, 12, -2, 3, 2, -8, -10, -13, -15, -15, 1, -7, -11, 6, -5, 10, 11, -2, 8, 5, 7, -5, -2, 3, -1, -8, 1, 4, 5, 0, -3, 7, 0, -3, 12, 9, 1, -2, 4, -8, 4, 0, -8, 5, -5, -1, 7, -3, 0, -4, 0, 4, 5, -5, -4, 9, -5, 2, -6, 9, 0, 6, -3, 8, -4, 4, -3, 11, 14, 9, -1, -6, -9, -7, -7, -5, 10, -4, 8, 5, -2, 1, 6, 16, 7, 5, -3, -6, 5, -2, -1, 0, -3, -4, -4, -3, 13, 12, 4, 15, 0, 6, 0, 0, -4, 1, 5, 3, -11, -1, 1, -4, -5, 3, -5, 0, 5, 9, -7, -3, -4, 1, 9, 6, 0, -4, 1, 8, -1, 7, 12, -6, 0, 12, -5, 9, 7, 17, 7, 3, 1, -14, 6, 8, 3, 7, -2, 7, -7, 1, 8, 0, 0, 13, 1, -10, -8, -5, 2, 0, -5, 6, 0, -6, -1, 7, 0, 3, 11, 10, 0, -6, -15, -5, -12, 0, 2, -7, -6, 4, -2, 11, 0, 19, 17, -17, -5, -12, -12, -6, -2, -16, -11, 2, -2, 0, 5, 3, 18, 5, -11, -8, -14, -13, -12, -4, -14, 0, -10, 4, -2, -1, 15, 13, 22, -18, -6, -12, -25, -15, -17, -12, 3, -6, 7, 2, -3, 16, 16, 10, -12, -5, -22, -19, -16, -3, 0, 0, 7, 9, -1, 3, 13, 8, 12, -1, -9, -14, -11, -9, -14, -6, -6, -2, -2, 3, 5, 7, 8, 17, -14, -15, -10, -14, -14, -9, -3, -8, -9, 2, 1, 10, 12, 2, 13, -2, -14, 0, 1, -2, -4, 2, -8, -6, 2, 11, 10, 3, 7, 6, -8, -10, -4, -5, 8, 1, -11, 0, -3, -3, 11, -1, 15, 6, 10, -7, -5, 7, 0, 4, 5, 10, 5, -1, 10, 9, -3, 10, 6, 7, -3, -5, 6, 7, 0, 2, 5, -5, 9, 9, 1, -5, 4, 5, 1, 9, 3, 6, 8, 1, -2, -5, 3, 0, 3, 0, 0, 3, -1, -3, 6, 7, 12, -4, -5, -4, -5, -6, 6, 6, -3, -9, 0, -3, -4, -7, -5, 2, 7, -4, 6, -1, 9, -7, 0, 8, -7, 3, 0, 9, -6, -5, 8, -3, -6, 3, 1, 8, -4, 6, 1, 1, -4, 1, 8, 7, -6, -8, 1, 4, -8, -6, 4, -1, 0, 5, 2, 0, 9, 5, -3, -7, -5, 3, -8, 5, -5, 8, 2, -2, 4, 7, 1, -7, 9, 6, 2, 2, 5, 6, -9, -8, 0, 2, -8, 0, -8, 7, -1, 9, -3, 0, -7, -10, 4, 5, 7, -4, -1, -2, 7, 1, 8, -1, 2, -7, 3, 2, -4, -11, 5, -7, -3, -6, -9, -2, 6, 3, -5, -3, 7, -3, -2, 6, -5, 0, 2, -8, 7, 4, 5, -1, 9, 0, 9, -2, 10, 0, 6, 2, -4, -10, 0, 0, -11, 1, -3, -2, 0, 6, 2, -4, 11, 10, 10, 3, 0, -5, -3, 8, 1, -3, -4, 9, 1, 3, -1, 6, 7, 11, 2, 4, 0, -2, -9, -6, 6, -2, -7, -7, -6, 12, 3, -3, 3, 10, 0, -4, 0, 2, 1, -6, -5, 0, -5, -2, -4, 4, 4, 5, 9, -4, 0, 7, 3, 6, -4, 6, 4, 2,
    -- filter=0 channel=4
    2, -3, -14, 0, 1, 3, 12, 14, 8, 2, 5, 9, 12, 16, 19, -7, -14, 1, -2, -2, 0, -6, 14, 4, 8, 5, 7, 6, 20, 21, 3, -1, -11, -1, 0, -2, 3, 1, 11, 8, 6, 20, 3, 6, 9, 6, 2, -7, 1, 6, 9, 12, 9, 12, 14, 13, 12, 17, 20, 6, -5, -6, 2, 9, -4, 3, 12, 13, 17, 11, 14, 2, 7, 5, 17, 2, -3, -11, -2, 3, -4, 2, 4, 6, 1, -3, 14, 20, 21, 11, 0, -1, -7, 5, 6, 1, 1, -7, 5, 6, 7, 6, 14, 8, 20, 1, -13, -2, 2, 4, 0, 1, -7, -9, -6, -13, 9, 9, 15, 9, 1, 6, -4, -9, -6, 2, 0, -5, -11, 3, -9, -7, 11, 5, 15, -8, -6, -8, 5, 0, -2, 8, -2, 2, 1, 0, 2, 18, 23, 8, 6, -8, 6, -5, 7, 8, 13, -1, -2, 10, -1, 10, 11, 18, 8, -8, -11, -8, -4, -2, 7, 5, 14, 4, 9, 15, 14, 14, 8, 19, -5, -2, 0, -4, 2, -6, 8, 7, 18, 7, 7, 18, 25, 13, 18, -5, -12, -2, -7, 5, 3, 6, 5, 17, 8, 7, 21, 8, 9, 4, -11, 5, -7, -2, -3, 8, 12, 6, 10, 16, 10, 15, 20, 13, 16, -8, -8, -13, -4, -11, -13, -2, 0, 2, 0, -10, -10, 0, -4, 4, -14, -9, -19, -6, -6, -13, -8, -9, -6, -11, 1, 1, -13, -12, -2, -9, -14, -17, -3, -7, 0, -7, -14, 0, -4, -2, 0, -18, -3, 0, -17, -3, -3, 0, -12, 2, -12, -12, -1, -13, -5, -7, -16, -15, -10, -14, -14, -14, -12, 2, -1, -11, -12, -17, -7, -15, 0, 1, -6, -9, -14, -9, -12, 2, -7, -9, 0, -8, -12, 0, -18, -5, -4, -14, 0, -4, -3, -15, 0, -13, -12, -10, -14, -18, -20, -21, -10, -1, -8, 0, -11, -14, -5, 0, -10, 0, -6, -9, -3, -9, -19, -9, -15, -11, -6, -5, -6, -10, -11, 2, 3, -17, -17, -9, -20, -22, -13, 0, -13, -4, -7, -10, 0, -8, -8, -14, -14, -7, -3, -2, -3, -12, -5, -13, -9, -16, -8, -13, 0, 0, -1, -7, -13, -14, -8, -4, -7, -12, -12, -5, -4, -9, -17, -7, 4, 4, 1, -8, -14, 4, -14, -13, -7, -6, -4, -4, -13, -1, -11, -3, -15, 0, -8, -4, 0, -7, -1, -13, -14, -3, -2, -17, -6, 0, -12, -17, -4, -8, 0, -7, -12, -8, -7, -17, -16, -11, -6, -8, -9, -14, -6, 1, -8, -6, 0, -8, -1, -4, -2, -10, 4, 1, 0, 1, 2, 0, 7, -8, -8, -5, 8, -4, -5, 8, -3, 5, -8, 2, -11, -9, -11, 3, 8, 3, 5, -3, 0, -5, 4, 8, -10, -1, 3, -6, -1, -10, -2, -1, 7, 0, 0, 1, -2, 10, 12, 7, -4, 0, -9, 1, -8, 7, 10, -6, 11, 0, 7, 2, 8, -4, -2, -8, 6, -1, 4, 6, 6, -8, -7, -6, 9, -5, 12, 8, 7, 7, -6, -3, -3, 0, -7, 0, -2, -6, -1, 8, -1, 0, -3, -5, -7, -11, 0, -10, 5, -3, -10, 6, -10, 0, 6, -6, 7, 12, 12, -4, -5, -8, -2, -11, -8, 1, 6, -2, -13, -3, -3, 3, 5, 0, 0, 2, 4, 4, 3, -3, 7, -5, -2, 4, 0, -9, 2, 1, 7, 4, -8, 0, 6, -9, -8, -3, -8, -9, 3, 6, -3, 6, 1, 0, -8, -7, -3, 1, -10, -8, 3, -9, -6, -6, 0, -5, 4, 8, 8, 4, -3, 1, 5, -6, -9, -9, 9, -6, 8, 4, 10, 11, 6, 1, -7, 3, -5, 0, -2, 0, -6, -8, 0, 4, 4, -4, -1, 8, 7, -6, -11, 2, 2, -2, 7, 1, 2, -4, 4, 7, 11, 6, -2, 12, 2, -2, -2, -6, 7, 8, 6, -8, -6, -5, -2, 11, -3, -7, -2,
    -- filter=0 channel=5
    7, -6, -1, 0, 7, 8, 4, 2, 8, 8, -4, -9, -1, -1, 4, -4, -6, -1, -15, -10, -2, -4, -13, -16, -9, -8, -14, -5, -10, -7, -6, -12, -14, -16, -9, 1, -16, 0, 0, -1, -11, -14, -17, -6, -4, 2, -2, -16, -9, -7, -5, 2, -5, 0, -7, -2, -1, 4, -12, 7, 11, 0, 9, 8, 4, 5, -2, 5, 4, -3, 12, 0, 11, -10, 2, 13, -4, 12, 14, 14, 11, -2, 1, 4, 11, 18, 9, 4, 3, 6, 1, 17, 6, 16, 11, -4, 3, -3, 13, 8, 21, 21, 3, 0, 3, 4, 8, 11, 25, 8, 5, 3, -9, 6, 5, 2, 5, 3, 9, 0, 14, 10, 20, 24, 9, 7, 5, 3, -3, 4, 0, 19, 14, 3, -1, 11, 11, 5, 7, 13, 7, 1, -9, -5, 11, 7, 4, 5, -2, 7, 16, 0, 8, 1, 6, 10, -2, 0, 10, 3, 19, 15, 14, -2, 16, 13, -9, -8, 7, 0, 2, -6, -1, 5, -1, 12, 0, 0, -3, 9, 0, -2, -14, -8, -5, -9, -7, 1, -2, 8, -7, 1, -13, -5, -8, 1, -4, -15, 0, -3, -9, -6, -1, -14, -7, -14, -11, -4, -2, -5, 2, -7, -15, -11, -4, -5, -2, -4, -16, -4, -8, -7, -1, -15, -4, -8, -12, -1, -2, 4, 0, -8, -7, 0, -4, 7, -5, 6, 0, 7, 1, -14, -20, -15, -14, -9, -9, -16, -7, -10, 0, -2, -10, -11, 2, -14, -6, -28, -15, -9, -8, -9, -2, 1, 2, -11, 2, -5, -6, 8, -1, -10, -12, -6, -2, -2, 3, -6, 1, 9, 0, -1, 9, 7, 9, 0, -2, -10, 5, -5, -1, -1, -4, -6, 11, 11, 18, 6, 4, 1, -3, -16, -3, 5, 1, 4, 3, 1, 1, 6, 13, 8, 14, 9, 5, 1, -2, 4, 15, -3, 2, 0, 4, 6, 7, 11, 19, 5, 14, 3, 3, -1, -2, 5, 0, -2, 7, -1, 6, 12, 24, 14, 5, 10, 7, -8, -5, -6, 1, 1, 1, -3, 5, 2, 13, 7, 8, 16, 4, 17, -4, -11, 6, 9, 10, 0, 4, 6, 10, 8, 8, 24, 2, 10, 15, -9, -9, -6, -2, -1, 6, 2, -4, 10, 9, 21, 6, 1, -2, 5, 2, -9, -21, 2, -5, 0, -11, -6, 0, 7, 6, 17, 14, 11, 3, -11, -19, -23, -16, -10, 1, -5, -11, -4, 2, 0, -2, 0, -2, -4, -11, -18, -22, -23, -18, -21, -18, -10, -3, -12, -5, -1, -6, -9, 7, 2, -16, -6, -5, 0, -3, -8, -14, 0, -7, 0, 4, -5, 7, 0, 9, -3, 2, -1, -3, -5, 0, -6, 3, 8, -4, -2, 2, 0, 5, -3, 3, -2, 1, -7, 0, 5, 5, -6, 7, 1, 4, -9, -5, 5, -6, -9, -5, 10, 7, 8, -2, -1, -8, -8, -6, -8, -6, 2, 9, 7, 0, -3, 6, -2, 1, 5, 2, -6, -2, 13, -1, -1, 6, 3, 11, 4, 10, 0, -3, 4, 8, -1, 5, 7, 1, -2, -5, -2, 6, 10, -3, 4, 8, 15, 6, 9, 1, -5, 7, 12, -1, 8, -1, 12, 10, 2, 0, 18, 2, 5, -5, 6, -2, 12, 0, 0, 14, 8, -3, -3, 2, 13, 16, 6, 7, 1, -4, 0, 3, 12, 0, -3, 5, 5, -2, 14, 2, 18, 2, 7, -4, 2, -6, 6, -4, 12, 7, 0, 0, 0, 12, 8, 14, 6, 13, 9, -9, 3, 0, 1, 6, 9, 5, -1, 9, 3, 6, 9, 0, -1, -5, 3, -4, 14, 0, 0, 7, 8, 6, 8, -3, 6, -4, 3, 1, 3, 4, 4, 2, 8, -3, -3, -8, 5, 0, 7, 9, 1, -7, 6, -5, 9, -2, 0, 11, 1, 6, 3, 10, 0, 5, 0, 1, 0, -7, -8, -3, 5, 4, 6, -9, -9, 4, 3, 0, -3, -2, 7, 9, 1, -6, -1, -2, 4, -3, 10, -7, 7, 1,
    -- filter=0 channel=6
    6, 0, 15, 12, 2, 4, -6, 9, -4, 4, -3, 7, -2, 11, 9, 3, 6, 10, 0, 3, 6, -6, 2, -6, 1, -2, -4, 11, 11, 9, 10, 3, 9, 16, -1, -3, -9, -3, -1, -11, 0, 4, 6, -7, 9, -3, -1, 9, 2, 9, 8, -6, -6, 0, -13, -9, 3, -5, -7, -1, 12, 0, 0, 16, 15, 18, 12, 0, -1, 7, 2, 0, 7, -6, -2, -3, 11, 10, 13, 8, 19, 8, 20, 2, 10, 8, 3, -5, -2, 0, 5, 10, 9, 16, 16, 13, 26, 34, 26, 23, 8, -3, 3, 1, 2, 8, 9, 1, 0, 10, 28, 33, 34, 38, 18, 20, 2, -10, 6, 4, -1, 1, -5, 6, 16, 30, 32, 36, 34, 16, 19, -4, -11, -7, 0, -4, -4, 0, -1, 6, 14, 22, 21, 23, 14, 11, -7, -4, -4, -10, 8, 13, 0, 1, 14, 23, 9, 6, 4, -1, 5, 0, 4, -8, -6, 0, 2, 3, 2, 5, 7, 3, 9, 3, -8, -7, -2, -8, 7, 3, 14, 0, 0, 15, 11, 7, 7, -14, -9, 1, -5, 6, 3, -3, 5, -1, 7, 5, 12, 1, 1, 1, -2, -15, -4, 6, 10, 12, -4, 4, 2, 3, 16, -2, 3, 9, -5, 0, -8, -5, 10, 11, 14, 10, 5, -16, -5, -9, -7, 0, 9, 6, -5, 8, -8, -2, 0, 1, 10, 4, -11, 0, -4, 0, -11, 2, -15, -6, 1, -2, 1, 1, 3, 2, 11, -3, -17, -20, -3, -16, -1, -10, -20, -8, 0, 2, 0, 6, 6, 3, -7, -24, -17, -18, -11, -9, -16, -27, -13, -19, -11, 0, 6, 5, 3, -16, -20, -26, -21, -27, -13, -15, -21, -16, -18, -5, -9, -1, 0, -5, -19, -13, -29, -19, -27, -21, -19, -11, -17, -9, -6, -22, -18, -14, -4, -9, -14, -25, -23, -32, -22, -10, -15, -11, -4, -10, -13, -15, -2, 1, -10, -19, -30, -26, -24, -23, -21, -15, -13, -9, -11, -14, -9, -1, -14, -18, -11, -18, -23, -36, -19, -24, -11, 0, -13, -8, -25, -6, -13, -2, -15, -15, -29, -17, -26, -25, -12, -7, -2, -5, -12, -10, -20, -6, -3, -3, -19, -10, -14, -24, -14, -24, -10, -8, -23, -21, -6, 1, 1, 2, -14, -20, -14, -21, -12, -8, -12, -12, -19, -9, -17, -5, -4, -10, 0, -10, -15, -8, -16, -19, -20, -7, -11, -15, -11, 0, 4, 6, 4, 1, -6, -7, -14, -13, -13, -8, -12, -5, 0, 2, -10, -3, -3, 0, 15, -11, -9, -16, -4, 0, 0, 4, 3, 5, 6, 4, 1, 13, 0, 4, 2, -1, -1, -6, -3, 10, 3, -8, 0, -9, 7, 4, 8, 6, 0, -6, 1, 0, -2, 10, -6, 3, -4, -6, 6, 3, 1, 1, -4, -6, 2, 3, -3, 4, 4, -4, 6, -12, -8, -9, -6, -6, 5, -7, 0, 10, 11, -7, 0, -4, -1, -7, 2, -12, -3, -9, -1, -4, 6, 6, 3, -4, 5, 3, 2, -6, 0, 0, -6, -2, 8, 0, -7, 4, -10, 0, 3, 2, 4, 7, 0, 6, -2, -1, -2, -9, -10, 1, 7, -4, -4, 6, -7, 2, 14, -1, 2, 15, 16, 13, 10, -4, -5, -2, -8, 0, -1, 8, 12, 2, 15, 15, 9, 4, 3, -4, 3, -2, 0, -7, 9, 9, 6, 6, -1, 15, 6, 11, 0, 9, -5, -6, -6, 7, -3, 3, -4, 3, 0, 0, 1, 16, 10, 6, 11, 2, -8, -1, 6, -2, 8, -5, -3, -5, -2, 4, 1, -2, -4, 0, -6, 8, 5, -3, -6, 0, -5, 1, 7, 4, 3, 7, -10, 5, -10, 1, 3, 2, 2, -9, -4, 3, -6, 1, 6, 0, 3, -1, -9, -5, -4, 8, -7, 1, 0, 10, 10, -4, 9, -1, -5, 7, 0, -5, 0, -8, -6, 9, 9, 5, 6, 6, -1, 1, -5, 5, -5, -9, -4, -7, -7, -2, -3, -7, 0,
    -- filter=0 channel=7
    0, 4, -12, 4, 3, 2, 0, 9, 8, 10, 7, 11, 11, 5, 6, -2, -6, -8, 2, 7, 3, 13, 18, 9, 20, 15, 23, 16, 11, 5, -11, 3, -7, -5, -2, -6, 5, 9, 14, 20, 16, 10, 23, 9, 2, -8, -5, 0, -6, -2, 5, 5, -5, 1, 4, 18, 12, 19, 12, 10, -6, -8, 1, -12, -5, -11, -11, -4, -8, -6, 10, 20, 18, 26, 10, -1, -9, 4, 4, 2, -3, -6, -22, -26, 0, 19, 28, 11, 8, 10, -7, -7, -3, -5, 8, 0, -7, -27, -37, -6, 9, 26, 19, 23, 18, -11, -8, -1, -6, -4, 6, 0, -30, -33, -15, 22, 21, 31, 7, 15, 3, 2, 9, -3, 1, -8, -9, -23, -39, -4, 19, 21, 28, 18, 5, -14, -1, 4, -4, 2, -10, -17, -18, -27, -8, 9, 20, 12, 8, 0, 0, -10, -11, -3, -7, -1, -11, -18, -15, -6, 17, 27, 20, 23, 8, -9, -10, -7, 0, -2, -4, -4, -10, -12, -1, 13, 17, 14, 15, 1, -11, -7, 1, -12, 0, -5, -2, -3, -2, 15, 7, 27, 25, 13, 4, -13, -8, 3, -12, 3, 3, 7, 8, 8, 10, 19, 16, 12, 17, 18, 4, -2, 2, -7, -8, 6, 15, 8, 16, 10, 12, 7, 10, 9, 1, 9, 15, 9, -7, -8, 0, -5, -2, 3, -2, -4, -23, -17, -10, -23, 1, 2, 8, -3, -3, -5, 0, 0, 2, 1, -4, -19, -26, -17, -19, 6, 17, 5, -7, -6, 0, -5, -10, 3, -14, -16, -13, -18, -27, -31, 16, 11, 15, -6, -13, -1, -12, -6, -1, 0, -11, -11, -6, -17, -14, 14, 15, 0, 6, -12, -14, -5, -12, -11, -2, -13, -4, -1, -22, -31, 10, 24, 14, -5, 0, -11, -14, -17, -28, -14, 3, 1, -5, -15, -29, 14, 11, 19, 0, 10, 5, -14, -26, -25, -14, -14, 5, -15, -5, -29, 18, 25, 15, 15, 10, 5, -15, -13, -26, -24, -10, 5, 1, -21, -15, 15, 26, 8, 2, 4, -4, -15, -17, -25, -16, 2, -4, -3, -14, -15, 14, 24, 11, 8, -4, -13, -12, -18, -20, -21, 4, 5, -7, -11, -31, 9, 27, 12, -1, -12, -5, -18, -13, -20, -7, 7, -9, -10, -5, -22, 19, 5, 6, 3, -8, -7, -17, -6, -7, -9, 0, -7, -13, -24, -24, 17, 4, 14, 0, -10, 1, -10, 2, 0, -1, 0, -2, -14, -15, -21, 4, 3, 11, -1, -8, 2, 6, 0, -5, -14, -13, -6, -8, -17, -17, 11, 11, 5, -2, -13, -7, -1, -6, 0, -11, 0, -17, -10, -25, -26, 2, -10, -7, -9, 1, 3, 0, 0, 4, 1, 1, 6, -5, -2, 8, -10, 2, -10, -4, 8, -3, 0, 4, 9, -2, 8, 2, 10, -2, 10, -11, -1, 5, -4, 2, 6, 0, 7, -3, 3, -4, 1, 4, -3, 7, -1, 3, -11, 0, -9, -10, 4, -1, -8, -1, -5, 12, -2, -2, -3, -9, -4, -2, 7, -10, 4, -3, 5, -3, -8, -4, 10, 6, -3, 11, 5, 0, 0, -6, 8, -5, -1, -6, -5, -8, 3, 14, 7, 7, -3, -11, 5, -2, 7, 0, 5, -2, -2, -5, -10, 13, 3, 16, 7, 5, -11, 6, 1, 5, 4, -7, -3, -15, -5, -10, 7, 2, 14, 12, -2, 1, -3, 0, 10, -2, 10, 5, -14, -9, -11, 0, 2, 3, 11, -4, -3, 1, -5, -5, 3, 9, -7, -8, 0, -6, -1, 10, 6, -3, 10, -2, -9, -8, 6, -4, 0, 4, -11, -1, 1, 5, -1, 4, 6, 4, 3, -1, 4, -2, 5, 6, -9, -3, -3, 8, 10, 10, 8, 15, -5, 5, 4, 5, -11, -9, 0, 0, -3, 1, -4, 3, -2, 3, -2, -5, 3, -5, -6, -9, 1, 6, -2, 2, 13, 9, 13, 0, 15, 8, 2, -1, -1, 2, -4, 4, -5, -1, 10, -3, 3, 8, 2, 5, 7, 6,
    -- filter=0 channel=8
    -6, 4, 2, 5, 4, 0, 1, -15, -13, -7, 3, -16, -22, -30, -36, -9, -11, 0, -14, -2, -5, -2, -14, -16, -7, 0, -7, -26, -26, -28, -6, -14, 0, -16, -9, -5, -11, 0, 3, -1, 5, -16, -10, -21, -31, -7, 0, -7, -13, -13, 4, -11, -5, -3, 3, -2, -14, -7, -27, -28, -12, -4, 1, -13, -4, 0, 9, 2, 9, 15, -1, 2, -18, -33, -38, -5, -8, -9, -6, 2, 6, 15, 2, 1, 15, 0, 1, 0, -13, -37, 0, -5, -3, 2, 11, 10, 7, -6, 5, 7, 4, -5, -13, -27, -28, -8, 0, -3, 4, 13, 20, 0, -4, 12, 14, 8, -7, -2, -23, -22, -1, 0, -3, 5, 4, 2, 2, 7, -1, 15, 3, 0, -7, -19, -20, -2, -13, 0, -5, 14, 16, 13, 2, -1, 0, 7, 0, -14, -15, -28, -7, -8, 0, -1, 2, -2, -3, -2, 11, 9, 7, -1, -15, -16, -38, -2, 0, -4, -3, 4, 3, 7, -6, -2, 6, -7, 5, -6, -23, -24, 3, -3, -6, 1, -13, -8, 0, 0, -9, 3, -2, -13, -16, -28, -38, 0, -12, -12, -9, -5, -16, -7, -3, -7, -5, -7, -7, -18, -18, -25, -3, 4, 2, -7, 3, -7, -10, -3, -3, -13, -10, -11, -19, -34, -33, 8, 10, 9, 5, 17, 13, 19, 9, 18, 23, 11, 12, 19, 14, 3, 12, 15, 14, 28, 20, 10, 14, 18, 10, 17, 20, 19, 19, 15, 8, 3, 23, 17, 13, 8, 16, 17, 3, 1, -1, 8, 10, 18, 7, 12, 15, 15, 20, 18, 12, 13, 19, 18, 8, -7, -1, 4, 7, 12, -5, 21, 20, 9, 22, 27, 13, 16, 0, -2, -3, 1, -1, 0, 0, 4, 21, 18, 14, 9, 27, 23, 2, 1, -4, -4, -4, -2, 12, 6, 7, 20, 13, 20, 14, 11, 6, 11, 2, 7, 5, 6, 6, 11, 3, 5, 7, 11, 10, 16, 13, 10, 6, 2, -2, 11, 1, 1, 7, -3, 1, 13, 24, 9, 16, 23, 16, -7, 1, -2, -1, -5, 1, -3, -7, -4, 11, 24, 19, 8, 15, 21, 2, 7, 10, 10, -6, -1, 5, 11, -3, 5, 9, 15, 11, 23, 16, 9, -7, 0, 6, -1, -5, 8, 6, 3, 5, 20, 11, 7, 15, 14, 18, 9, 10, 8, 8, -3, 10, 11, -3, 19, 25, 12, 24, 19, 7, 13, 7, -4, -6, 5, 16, 3, 2, 13, 16, 12, 22, 17, 8, 12, 23, 5, 6, 13, 12, 5, 12, 7, 1, 14, 18, 25, 22, 16, 15, 14, 21, 15, 16, 16, 26, 19, 19, 5, 1, -2, 8, -5, -7, -10, 0, 0, 0, -4, -3, -1, -3, 0, 0, -9, -1, 1, -2, -3, 3, -4, -10, -4, 0, -9, 0, -2, -13, -4, 6, -6, 0, 3, 1, 2, 2, 0, 3, -9, -5, 6, 3, -17, -9, 6, -1, -5, 7, 8, -2, -5, 1, 8, 9, 6, 2, 0, -12, -15, 6, 1, -2, 5, 5, 9, 9, 7, -3, -2, 6, 2, -9, -16, -10, -2, 0, -6, 8, -7, -4, 4, -6, 6, 5, 6, 7, -8, -9, 0, -7, 1, -10, 1, 8, -3, 0, -6, -5, 5, 7, 1, -4, -6, -18, 3, 0, 2, 0, -4, 8, -3, 8, -3, 6, -1, -1, 6, -4, -14, 3, 6, -8, 4, 2, 6, -5, 2, 0, 10, 12, -6, 0, -11, -2, -7, 1, -3, -8, 4, 3, 2, -8, 6, 4, 6, 6, -2, -8, -11, 8, 5, 1, -1, 4, 5, -6, -3, -4, 11, 9, 0, -3, 0, -15, -5, -7, -6, -4, 2, 0, 5, 7, 9, 2, 3, -3, -6, -11, -12, -10, -10, -2, 3, -8, 0, 4, -6, 1, 7, 8, 0, -1, -9, -2, -8, 5, 0, 0, 4, 0, -5, 0, -13, 1, 1, -2, -12, -3, -17, -2, -3, -3, -12, -9, -11, 3, 3, -11, -6, 2, 1, -10, -1, -19,
    -- filter=0 channel=9
    2, 7, -2, 4, -5, -5, -4, -19, -16, -17, -13, -12, -8, 6, 8, 7, 14, 2, 3, 3, 4, -5, 1, 3, 0, -8, -6, 0, -1, 0, 3, 16, 9, 17, 4, -4, 4, 3, 5, -11, -9, -7, -4, 11, 7, 3, 12, 4, 9, 5, -1, 5, -6, 0, -2, -12, -25, -16, -4, 6, -3, 2, 14, 7, -4, -8, -8, 7, 12, -7, -7, -12, -6, -7, -7, 4, 5, 1, -9, -2, 0, -1, 6, 0, 0, -18, -11, -11, -17, -8, 6, -3, 0, -4, -10, -8, -7, 3, 10, 11, -4, -16, -16, -1, 4, 5, 5, 4, -10, -5, -10, -3, 8, 18, 19, -16, -25, -8, 0, -4, 0, 6, 5, -6, -8, 3, -4, 4, 25, 17, -8, -10, -23, 0, -8, 0, 4, 10, 0, -1, -5, -1, 2, 22, 16, -1, -23, -12, -5, -1, -4, 6, -2, 10, -9, -5, -8, 5, 10, 10, -7, -12, -11, -14, -2, 7, -1, 14, 13, -5, 2, -2, 3, 7, 0, -18, -12, -10, -11, 6, 4, 17, 5, 3, 12, -2, -2, 6, 7, -5, -10, -16, -4, 2, -4, -3, 4, 15, 8, 6, 8, -4, 8, -7, -2, -4, -13, -2, 6, 3, 0, -2, 4, 11, 0, -3, 1, -3, -14, -2, -18, -2, -2, 7, 0, 4, 0, 4, 8, -1, -18, -21, -11, -18, -9, -12, -4, -16, -13, -6, 9, 7, 22, 11, 5, 11, 5, -8, 0, -20, -17, -22, -11, 0, 6, 13, 20, 35, 15, 20, 10, 2, -4, -12, -1, -16, -14, -14, -7, -8, 11, 31, 25, 25, 14, 2, -1, -1, 3, -10, -1, -2, -18, -3, -1, 16, 18, 17, 7, 3, 2, -8, -3, 4, -2, -13, -15, -5, 1, 3, 13, 24, 12, 1, -6, 6, 2, 0, 1, -2, -10, -16, -8, -1, -9, 6, 22, 11, 9, -1, -7, -3, -3, 5, -2, 3, -13, -4, -1, 3, 9, 14, 11, -6, 2, 5, -2, -3, 9, 6, 3, -7, -8, 3, -6, 3, 18, 11, 2, -2, 2, 8, 5, 16, 1, 3, -9, -7, -12, 3, -4, 8, 6, 4, -5, -7, -12, 6, 5, 8, -2, -3, -5, -15, 4, -2, 13, 18, 7, -2, 3, -7, 0, -3, 0, -6, -12, -3, -5, -2, 15, 17, 26, 17, 7, 7, -2, -7, -4, -14, -7, -17, -2, -11, 0, 11, 17, 29, 10, 10, -3, -5, -8, 6, -11, -23, -18, -6, 2, -2, 6, 15, 28, 10, 7, -2, -4, -3, -2, -7, -23, -6, -5, -7, 0, 9, 18, 9, 16, 8, 0, -8, -9, -12, -28, -21, -23, -13, -3, 5, -10, 0, 5, 3, -11, 4, 4, -4, -12, -10, -13, 5, -10, 7, 1, -2, 8, 11, 4, -8, 5, -4, 0, -1, -6, -1, -7, 4, 0, 5, -8, -5, -5, -6, 0, 0, 6, -2, 9, -2, 0, -4, 0, 0, -4, -6, 7, -7, 3, -4, 6, 4, -7, -1, -6, -5, 3, -10, -3, -6, 5, -3, 5, -3, 0, -1, -7, -6, 6, -3, -12, -5, -15, -5, -8, 3, 9, 7, 4, -2, 4, -9, -2, -3, -2, -2, -5, 0, -8, 5, 4, 3, -10, 2, -6, -5, -4, -2, 0, 10, 1, -14, -5, 0, 6, -11, 6, -7, -4, -6, -4, 10, 3, 6, 5, -5, -12, -15, 4, 4, 1, 5, 4, -7, -8, 1, -5, -2, 13, 10, -7, 2, -10, -9, -4, 0, 9, 8, -3, 1, -11, -7, 1, 14, 8, 5, -5, 2, -12, 1, -3, 4, 7, 3, -1, -2, -4, 4, 7, -5, -7, -5, -1, 0, 8, -3, -1, -5, 0, 8, 4, -2, -5, 11, -1, -9, -15, -10, -6, 5, 6, 10, 11, 10, -5, -2, 2, -2, -3, -6, -9, 0, -1, -5, 5, 3, 8, 0, 4, 8, 4, 0, 0, 0, 7, 0, -10, 0, 10, 4, -3, -10, 4, -5, 0, -11, 1, -10, -10, -8, -7, 1, 3, -5, 0,

    others => 0);
end iwght_package;
