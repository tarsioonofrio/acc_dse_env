LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE inmem_package is
		type padroes is array(0 to 4000000) of integer;

		constant input_mem: padroes := ( 
					-- bias

					-- weights

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 221, 0, 
			0, 0, 0, 
			

			399, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 123, 
			0, 0, 0, 
			

			0, 133, 249, 
			0, 0, 252, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 506, 383, 
			

			4, 0, 0, 
			0, 0, 134, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 39, 
			0, 0, 0, 
			

			0, 0, 0, 
			273, 0, 0, 
			0, 0, 0, 
			

			0, 372, 0, 
			129, 766, 0, 
			0, 0, 0, 
			

			251, 0, 0, 
			0, 0, 861, 
			0, 0, 0, 
			

			698, 518, 294, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 498, 0, 
			0, 0, 0, 
			0, 823, 157, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 25, 0, 
			

			0, 0, 501, 
			0, 0, 162, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			468, 0, 0, 
			0, 121, 0, 
			781, 0, 123, 
			

			0, 0, 0, 
			0, 0, 264, 
			0, 270, 983, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 54, 0, 
			0, 0, 0, 
			

			267, 0, 207, 
			193, 0, 701, 
			193, 0, 0, 
			

			0, 0, 0, 
			0, 571, 368, 
			453, 0, 504, 
			

			0, 142, 0, 
			0, 0, 9, 
			0, 0, 0, 
			

			184, 141, 346, 
			575, 898, 1005, 
			867, 765, 0, 
			

			0, 449, 0, 
			318, 657, 694, 
			0, 0, 0, 
			

			517, 1139, 0, 
			0, 0, 751, 
			793, 0, 97, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 193, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			235, 968, 489, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			153, 0, 0, 
			206, 757, 547, 
			0, 0, 0, 
			

			0, 652, 0, 
			0, 0, 0, 
			0, 821, 1487, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			490, 531, 827, 
			0, 0, 0, 
			0, 0, 0, 
			

			235, 0, 415, 
			144, 459, 0, 
			0, 0, 0, 
			

			0, 767, 0, 
			103, 147, 0, 
			0, 0, 414, 
			

			512, 0, 350, 
			0, 0, 0, 
			0, 0, 209, 
			

			0, 0, 0, 
			0, 505, 0, 
			0, 0, 0, 
			

			300, 732, 0, 
			0, 0, 8, 
			0, 0, 437, 
			

			286, 0, 0, 
			839, 376, 540, 
			0, 0, 0, 
			

			171, 68, 987, 
			0, 0, 0, 
			0, 0, 187, 
			

			0, 0, 49, 
			0, 0, 0, 
			0, 0, 0, 
			

			382, 0, 219, 
			0, 154, 0, 
			847, 0, 0, 
			

			0, 0, 0, 
			0, 38, 655, 
			325, 65, 362, 
			

			179, 0, 0, 
			0, 435, 873, 
			622, 0, 0, 
			

			169, 0, 0, 
			0, 141, 0, 
			0, 372, 0, 
			

			635, 0, 0, 
			0, 39, 505, 
			0, 0, 0, 
			

			0, 0, 0, 
			829, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 270, 
			

			0, 30, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 1073, 
			343, 0, 0, 
			644, 216, 996, 
			

			0, 0, 0, 
			0, 0, 0, 
			899, 1369, 1442, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 341, 285, 
			

			0, 0, 359, 
			0, 121, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			879, 0, 427, 
			196, 407, 462, 
			507, 0, 0, 
			

			460, 651, 837, 
			250, 782, 1087, 
			0, 1738, 755, 
			
