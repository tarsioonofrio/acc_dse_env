library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -- layer=3
    -3470, -5491, -1783, 4491, 6233, -3455, 7750, -6763, 2614, -1997,

    -- weights
    -- layer=3 filter=0 channel=0
    4, 9, 24, 29, 1, -3, 17, -12, -2, 23, 1, -8, -6, -39, 19, 4, -45, -4, -6, 12, -4, -6, -6, -2, 40, 17, -6, 2, 30, -37, -22, -1, 2, 22, 1, 4, 8, -6, -2, -117, -3, 6, 0, -3, 4, -13, -9, 15, 13, 1, 0, 9, -3, 8, -8, -8, -13, 11, 0, 19, -17, -1, -4, 2, -16, -9, -49, -27, 2, 2, 6, -10, -7, -5, -2, -1, 3, 10, -25, -6, 23, -5, -2, -6, -3, 0, 2, -1, 0, -13, -6, -64, 23, -14, -10, -7, 1, -8, -21, 27, 12, -5, -43, 18, 0, -4, -41, 4, 21, -12, 2, -6, 0, -12, -4, 2, 3, -35, -9, 7, 3, 3, 54, -16, -32, 4, 8, 11, 1, -6, -11, 25, 0, -103, 8, -4, -8, -5, -74, 0, 0, 10, -7, -9, -19, -23, -54, -16, 0, 1, -8, -12, 6, 21, 25, 5, 1, -24, 55, -8, 19, 5, -32, -22, -9, 3, 24, 7, 30, 18, 16, -9, -3, -4, 6, 0, -63, 29, -11, -36, 1, 13, 33, -1, -13, -3, -5, -52, 7, -3, 7, -29, -17, 25, -13, -7, 2, -18, -30, 24, 6, -15, 4, 7, 12, 37, 11, 3, -4, -36, -2, -4, 58, 0, -13, 2, 4, 15, -7, -41, -5, -19, -1, 1, 5, 18, -23, -1, 17, 4, 19, -47, 7, 1, -5, 1, -1, 1, 10, 5, -12, -4, -8, -10, 6, 8, 11, -14, 61, 31, 61, -33, -36, 66, -3, -30, -63, -3, 6, -5, 24, -59, 14, -6, -34, 13, -2, -15, 8, -2, 4, -4, -32, -27, -7, 31, 14, -8, 4, 5, -3, 7, 5, 7, -41, 29, 8, -57, 0, -14, 1, -49, 3, 38, -23, 6, 19, 9, 2, -15, 0, -8, 36, -36, 2, 6, -2, -4, 3, 12, 14, 17, -20, 17, -15, 8, 23, -13, -29, -3, -33, 19, -7, 7, 1, -21, -6, -15, 2, -33, -8, 25, 22, -8, -6, -5, 3, 17, 13, 30, 31, 4, 7, -2, -16, -1, -5, 1, -1, 5, 7, 24, 10, 0, 5, 9, 2, -5, 4, -4, -5, -6, 13, -3, 8, -6, 10, 1, 4, -13, -7, 0, -5, 23, 1, -40, -33, -25, -12, -18, 20, 5, 2, -56, 2, 0, 15, -7, -1, 8, -27, -6, -16, 8, -15, -12, 3, 12, 32, 4, -10, 3, -17, 2, 34, -10, 6, -37, -13, 27, -7, -6, -22, 2, 22, -7, 29, -60, -30, -7, -46, -10, -19, 9, -8, -5, -7, -7, -34, 6, -27, 3, 34, -14, 2, 7, 41, 33, -6, 0, -11, -25, -54, -10, -8, -8, 0, -9, 16, -7, 9, 5, -11, -2, 4, 2, -8, -7, -6, -15, -6, -7, 0, -6, -4, 5, -18, -4, -7, 47, -9, -3, -15, 16, -6, 1, 5, -8, 9, -5, -13, 0, -2, -44, -6, 10, -4, -17, -3, -14, 7, 48, -3, 9, 20, -14, 0, 4, 3, -6, 5, 9, -15, -4, 6, 2, 2, -51, 23, -1, 5, 31, 1, -2, 4, -19, -2, -7, 9, -19, 12, 22, 8, 0, -14, 8, 18, 9, 29, 11, 19, 14, -7, 1, 16, 0, 11, 0, -11, 8, -4, -15, 27, 28, -4, 14, 34, -25, -1, -6, 7, 5, -6, 8, -21, 1, 7, -1, -28, -2, 33, -1, -5, 11, -7, 8, 23, 19, 15, 0, 0, 16, -15, -19, 22, 5, -21, 9, -36, -16, -6, 26, 5, -6, -5, 3, 9, -6, -9, -27, -1, -3, 6, -2, 2, -2, 7, 1, 5, -7, -5, -2, -13, 10, 23, -24, -4, 0, 0, 1, 9, 1, -15, 6, 31, 10, 30, -16, -38, -19, 25, -13, -23, -3, 6, 6, 5, 0, -7, -1, 0, -17, -5, 5, 2, 17, -27, -4, 18, -2, 0, -10, 5, 17, -1, -27, -4, 3, 0, -4, -16, 8, -1, -3, 0, -8, 15, 2, 19, 28, -1, -16, 6, -2, -6, 17, 3, 5, 2, 14, -6, 1, 27, 4, -38, 16, -2, 4, -5, -9, -21, 1, 18, -9, 3, -5, 2, -8, 2, -25, -12, 2, 5, 5, -26, -8, -6, -6, -4, -34, 8, 0, 0, -44, -22, 0, -6, 1, -7, 9, 4, -10, -9, 1, -5, -2, -3, 20, 9, 2, -13, -40, -75, -27, 13, 9, 4, 2, -5, 19, 7, 0, 0, 0, 25, 26, -1, 19, 18, -17, -27, -50, 10, -78, 10, 0, -5, -2, 5, -1, -19, 4, -1, 9, -2, -19, 5, 3, 15, 2, 31, -19, 8, -17, -9, 0, 0, 0, -47, 9, 16, 29, 0, -16, -16, -5, -2, -21, 8, -6, -2, -16, -1, 7, -28, -38, 27, 11, -12, -13, -16, 0, 3, -10, -2, -41, -17, -8, 2, -60, -7, -7, 4, -42, -3, -27, -22, -7, 26, 5, -9, -22, 1, 3, 5, -19, 1, 2, -9, 25, 42, 22, -3, -25, -16, 8, -8, -7, -12, 26, -7, -5, -13, -34, -11, -7, -5, 35, 9, 13, -2, 12, 9, 2, 23, 0, 20, -2, -4, -4, 19, 26, 13, 5, -1, -6, -7, 7, -5, -11, -3, 5, -31, -43, -2, -4, 0, 0, 0, 3, -3, 7, -1, 0, -2, 1, 0, 7, -16, -3, 1, 0, 0, 0, -3, -1, -3, -7, -7, -1, 3, -13, -8, -6, -1, 10, -4, 20, 14, 0, -6, 30, 22, 4, 11, 0, 1, -15, 11, 6, -20, -2, 32, 2, 36, -2, 20, 0, -8, -7, -27, 11, -2, -27, -10, 6, 7, 4, 22, 3, -1, -14, 15, -8, 14, 16, 21, -5, -3, -8, -16, -6, -32, 2, -7, 0, -7, 12, -34, 43, 5, 0, -3, -2, -28, -8, 0, 1, -2, -29, -13, 3, 15, 18, 25, 4, 16, 4, 0, -5, -3, 1, -1, 3, 3, 2, 1, 1, 4, -6, -20, 27, -6, 7, -2, -1, 0, 8, 25, -15, -7, -3, 34, -14, -20, -18, -7, 3, -6, 10, -7, -41, 14, 40, 15, 1, 2, 13, 9, -11, 1, 8, 3, 3, 31, -1, -3, 2, 3, 14, 20, 11, 3, 1, -26, -2, -11, -14, -6, 4, 0, 21, -3, 28, 2, 5, -9, -19, -21, 3, -22, 20, 23, -15, -7, 3, 14, -3, 36, 8, 0, 0, 23, -60, -8, 1, -2, -9, 45, -30, -6, -5, 0, -20, -1, 1, -11, -7, 10, -14, 23, 30, 6, -16, -2, 0, 4, 3, -16, -10, 16, 0, 1, -6, -36, -22, -15, 0, 5, -8, 46, 44, -5, -68, 0, 1, -4, -7, -3, 0, -4, -28, -41, 0, -3, -8, -20, -6, 1, 20, -3, -10, 1, -8, 15, 5, 17, -24, 13, 0, 0, -4, -29, 8, 18, -1, -51, -31, 5, 0, 22, -4, 49, -14, 5, 0, -5, 7, -7, -8, -1, -28, -3, -16, -9, -4, -22, -34, -4, 2, 6, 17, -23, 25, 8, 73, 2, -25, -2, 4, 0, 8, 16, -1, -5, -4, -12, 3, 14, 5, -26, 14, 8, -8, 5, -5, 2, -1, 14, 3, 1, 14, 16, -2, -8, 5, -61, -18, 0, 1, 8, 5, -4, 9, 1, 12, -25, -6, -8, -6, -20, -7, -56, 24, -1, 0, 20, 2, -14, 6, 0, -4, 18, 0, -6, -70, -15, 8, 12, -8, 5, -4, -30, 0, 12, -8, 5, 7, 1, 32, 11, 1, 3, -22, 0, 14, -1, 13, -11, -36, 6, 5, 6, -4, 10, -8, 18, 23, -9, 3, -17, 7, -18, 9, 10, -22, 9, -3, 10, -6, 2, 11, -52, 1, 2, 9, -6, -2, 3, 6, -6, 0, 7, -36, -53, -18, -3, 3, 9, 3, -41, 5, -11, -1, 19, -68, -6, -3, -24, -11, 4, -10, 8, -13, 7, 0, -19, 6, 0, 26, -16, 36, -8, 0, -6, -36, -14, -12, -2, 0, -5, -28, 40, -14, -1, 4, 4, -50, -46, -6, -4, 4, 5, 14, -9, 1, -34, 22, -9, -13, 2, 26, 8, 18, -25, -7, -15, 14, -1, -1, 6, -21, -26, -6, 26, 6, -29, 25, -13, -36, -5, 52, -5, 35, -11, -14, -29, -1, -12, -7, -5, 10, 0, 40, 17, 4, -12, 5, -18, 6, 0, -2, 1, 1, -20, -1, 7, 5, 0, 0, 25, -5, -4, 1, -1, 7, -22, -3, 0, 10, -21, 0, 6, 6, -1, 3, 5, -6, -6, -27, 15, -15, 4, 9, 14, 3, 25, 40, -2, 21, 0, 2, -2, -15, 5, 3, 0, 7, 10, -5, -10, -12, -54, -2, 20, 4, -19, 7, -8, 11, 25, -5, -23, -9, 8, -2, -62, -6, -2, -1, 6, -13, -13, -28, -2, 0, 17, 1, -6, -3, 0, -6, 18, 1, -18, 5, 8, 1, -3, 6, 17, -63, -7, 1, 1, 5, -20, -3, -5, -2, 3, -43, -39, -6, 8, -12, -6, 8, 28, 3, -4, -6, -6, -16, 6, 3, 4, 2, -7, -5, -4, 6, -21, 7, 4, -5, 13, 18, 6, 3, -18, -23, 10, 3, -27, -17, 0, -5, 4, -25, -4, 2, 2, -8, -10, 12, 12, 0, 14, -11, 9, -8, -1, 9, 4, 5, 7, -7, 9, 6, 5, 22, 1, -1, 3, 21, 48, 4, 7, 6, -3, 6, 22, 12, 14, -38, -4, -1, -7, 16, -12, 6, 0, 39, -5, 40, 6, 8, -28, 29, -22, 15, -10, 0, -33, -47, 36, 7, 0, -53, 4, 11, 3, 7, -1, -43, -4, -14, -4, 0, -8, -8, -13, 8, 29, -2, 3, 17, -8, 8, 0, -29, -38, -2, -10, -15, -61, 1, 35, 5, -7, 1, 9, -31, 2, 9, 2, 0, 0, -1, 0, 9, 4, 1, -16, 0, -28, 0, -3, -5, 0, 16, 1, -5, 4, -3, -20, -34, -3, 0, -13, -3, 3, 3, 21, 27, 16, -8, -13, -5, 15, -22, -32, -4, 17, -24, -3, -2, 1, 20, -5, -6, 2, 1, 8, 42, -2, -6, -21, -11, -26, -6, -12, -18, 2, 16, -37, 19, -11, -47, 0, 1, -1, 0, -18, -1, -3, 5, 7, -5, -23, -4, -41, -36, -1, 33, 4, -8, 1, -6, 15, -9, 4, -48, 7, 2, 21, -1, -63, -2, 0, 0, 4, -2, -6, 33, 0, -28, 0, -6, -3, -9, -39, -45, 16, -20, 3, -2, 2, 6, -2, -2, 4, -19, 14, 7, 3, -24, -2, 19, -15, -4, -9, -7, -6, 22, -25, -22, 9, 0, 20, 41, 10, -6, -10, -22, 13, -12, -5, 3, 5, -12, 8, 11, -4, -21, -5, -4, -25, 7, -3, 4, 0, -6, 42, 9, 46, -22, -3, 10, -1, -1, 7, -44, 10, -6, -11, 0, 0, 26, -6, 29, -35, -2, 27, 10, -35, 1, -8, -17, 9, -3, 35, -3, 12, 16, 24, -17, -18, -8, -22, -23, -7, -6, 6, 4, 6, 10, 26, -11, -33, -21, -10, -13, 3, -2, -3, 1, 24, 17, 19, -10, -2, -36, -39, -9, 2, -43, -2, 30, 9, -2, 7, 6, 5, -34, -47, -2, -2, 22, 5, -11, 5, -41, -44, 22, -19, -43, -26, -4, -2, 4, -12, 36, 5, -4, -3, -16, -43, 13, -17, 10, 3, -11, 8, -39, -12, -3, 4, -12, 3, 7, 10, 4, -3, -11, 26, 4, -2, 12, 16, -8, 0, -13, -12, 3, -7, 63, 0, 0, 0, -7, -29, -9, 4, 1, 7, 6, -2, 9, -11, -21, -6, -6, -6, 27, 3, 6, 8, 0, -6, 15, 18, -52, 4, 0, -24, -2, 25, 32, -7, 0, -22, -3, 8, 0, -44, 3, 50, 19, 8, -9, 52, 21, 40, -16, -12, -1, -14, 2, -29, -11, -17, -66, 21, -6, 1, -37, -9, -5, -4, -9, -1, 14, -11, 17, -26, 3, 8, 7, -11, -16, 2, 7, 1, 0, 16, -7, 49, -8, -7, -42, 5, 29, -2, -6, -13, 7, 16, 0, 0, -13, -1, 15, 1, -1, -8, 9, -27, -25, -4, -7, 2, -10, -6, 4, 1, -8, -10, -4, -10, -9, 8, -7, 18, -6, -8, 6, -27, -63, 4, 2, 7, 24, 6, -4, 0, 20, -22, -16, 9, 24, -7, -12, -7, -9, 4, 58, 2, 1, -18, 6, -19, -7, -8, 1, -2, 3, -6, -6, -5, 9, 3, -98, -14, -3, -5, 34, -14, -8, -40, -8, 6, -4, 12, -17, -31, -8, 1, -2, -12, 33, 24, -1, 61, -4, -38, -22, -8, -4, -26, 10, -22, -11, 3, 3, 11, -14, 8, -30, 8, -18, 10, 3, -1, -3, 8, 37, 4, -9, -27, 3, -16, -1, 28, 10, -56, 12, 0, 8, 2, 3, 4, -31, 10, -5, 1, -10, -16, -26, -16, 2, -10, 28, 0, 4, 3, -24, 4, 7, -5, -4, -5, -2, 9, 14, 16, 2, -13, 4, 3, 7, 0, 13, 0, -3, 4, -1, 14, -24, -43, 1, -12, 2, 2, 7, 7, -28, 25, 5, 24, 23, -4, 3, 8, -4, -13, 3, 1, 2, 6, 1, 2, -4, 1, -21, 5, 0, 0, -6, 4, -21, 20, 1, -25, -24, 2, 20, -15, -11, 1, -3, 20, 6, -9, -8, 18, -18, -6, -11, -13, -2, 3, -2, 0, -2, 3, -6, 13, 1, -1, -3, 6, 0, 7, -6, -31, -9, 9, -3, -17, 13, -2, -2, -3, -3, -18, -21, -37, -36, -11, 4, -6, -4, 27, -4, 33, 7, 4, -7, -7, 6, -6, 5, -7, -3, 16, 0, -12, -14, 17, 10, 20, 4, 0, -22, -6, 7, -15, -3, 1, 0, 13, -44, 11, -3, -9, -10, 45, 22, -28, 6, -18, 39, -7, -17, -6, 1, 4, -4, 13, 45, 7, 6, -3, -17, 14, 2, 3, -32, -6, 5, -1, 4, -3, -13, 31, -2, -10, 9, 0, 10, 1, 5, 9, -13, 21, -51, -7, 22, -40, 35, 2, -34, -23, 16, 29, 13, -19, -41, -11, 0, 25, 34, -1, -3, -4, -17, -3, 1, 42, -6, -14, 66, -5, -5, -2, -1, 5, 12, 24, -38, 24, 13, -7, 15, -45, -14, 1, 5, 1, 23, 35, 4, 25, 8, 0, 34, 8, 8, -31, 38, 6, 19, -3, -46, -7, 5, -14, 11, 21, -5, 1, -4, 30, -27, -21, -1, -26, 0, 8, -1, -10, 4, 0, -26, -1, -26, 27, 3, 16, -12, -6, 6, 8, -26, 20, 41, -44, 6, 1, 6, -29, 0, 6, -11, -6, -6, -45, -9, 4, -5, 7, -6, 6, 2, 0, 9, -7, 0, -12, -6, -1, 19, 1, 0, 3, 22, 0, 0, 6, -4, -4, -29, -30, -22, 4, 10, 2, 0, -24, 32, 3, 0, -37, 1, 4, -17, -9, 0, -2, 3, 0, -11, 13, 0, 5, 1, 2, -9, 27, -3, 22, 1, 13, -18, 38, -23, 8, 26, -39, -5, 2, -8, 3, -7, -27, 42, 12, -8, -9, -15, -8, -6, 4, 6, -7, 3, -21, -8, -2, -19, -1, 17, -10, -17, -1, 6, 9, -13, -9, -1, 0, 8, -2, 4, -8, 7, -6, 10, -32, -9, -2, 5, -4, -5, 0, -18, 3, 5, 7, 8, 2, -2, 2, 5, 0, 17, -3, 4, 4, -44, -6, 7, -1, 9, 7, 3, 48, -35, -18, 50, 7, 28, -4, 16, -10, 0, -5, 15, 11, 4, -15, 24, 5, 6, 4, 1, 6, 2, -30, 6, -5, 7, 1, 2, -19, -7, 0, -39, -53, 0, -15, -23, 1, -3, -15, 31, -14, -18, -1, 1, -4, 11, 17, -6, -42, 2, 21, -3, -4, -6, -25, -12, 3, 46, 0, -9, -4, -21, -2, 16, -5, 2, 19, -20, 0, 2, 7, -71, -6, -3, -10, 0, 15, 5, 30, 17, 8, 0, 0, -31, 0, 0, -2, -5, 8, -3, -5, -7, -26, 5, -7, 6, -3, -12, 2, 12, -13, -58, -6, -6, -8, 4, -1, 1, 0, -53, -19, -6, 10, 1, -42, -4, -1, -39, -12, -4, -2, -6, 7, -84, -30, -60, 20, 4, 2, -3, -23, -19, -3, 0, -61, 18, 14, -16, 38, 3, 22, 17, -26, -1, 1, 0, 0, 0, -2, -50, -2, -2, -10, -9, -1, -16, 25, 5, 2, -1, 32, -7, -2, 7, 0, -15, -11, 2, -1, -1, -33, 4, 0, 3, 0, -2, 15, -14, -18, 4, 8, 11, 13, -4, 4, -15, -9, -3, -6, 6, -8, 6, -17, -5, -30, -73, 0, 4, 5, -1, 28, 11, 12, 28, 20, 0, -4, 7, -87, 28, -16, 23, 2, -10, -10, 5, -2, 4, 18, 43, 25, 1, 3, -20, -19, 25, 25, -1, -3, 10, 42, 1, 7, -25, -3, 0, 14, -22, 2, 2, -19, 0, -9, 12, -12, 6, -15, 4, 2, -26, -6, -30, 11, -10, 11, 9, 3, 18, 10, -39, -7, 20, 24, 7, -2, -6, 2, -7, -3, -4, -90, -6, 10, -7, 2, -13, 0, 23, -14, -29, -16, -55, -82, 9, 14, 0, 3, -9, -8, -3, -47, 25, -36, -31, 0, 16, 2, 0, 2, -10, 7, -33, 0, -7, 14, 10, -31, 15, -10, 38, -19, -8, 2, -4, 36, -20, 6, -8, 5, 8, -14, -8, -3, 10, -7, 16, -15, 3, 3, 0, 10, 49, -27, -2, -4, 9, 30, 30, 7, -12, -27, -5, -32, -7, -5, -63, 9, 9, -18, 5, 13, -7, 30, 27, 2, -1, -12, -9, -6, -49, 2, 33, -28, 0, -4, 9, -31, 6, -6, 13, 35, 9, -68, 3, -6, -4, 35, -6, -3, 0, 10, 2, -49, 6, -11, 5, -5, 5, 30, 3, -5, 0, 6, -7, -28, 9, 4, -5, -12, -4, 2, 0, 3, 11, -2, -15, -7, 16, 9, -47, 1, -6, 2, -3, -6, 15, -3, -30, -87, -6, -7, -11, 14, 0, 12, -5, -46, -52, 3, 9, 13, -5, -45, -7, 3, 2, -17, 16, 12, 24, -30, 10, 6, -31, 4, -2, -21, 5, -12, 36, -59, 11, 25, -7, 7, -13, -32, -5, -8, 8, 9, -4, -4, 6, 15, 32, -2, 37, -23, -79, -1, 11, -4, 8, 35, 4, -1, -6, 0, 19, -45, -4, 10, -3, -11, -11, 0, -9, -8, 4, -14, -41, 3, -10, 0, 2, -10, -6, -33, -2, 23, 12, -8, 9, 13, -30, -9, 0, -32, 24, 9, 8, -14, -74, -12, -21, 9, 18, 10, 20, -4, 11, -25, 1, 5, 8, 4, -9, 42, -1, -5, 5, -7, -1, 33, 9, 4, -7, 0, -70, 28, -4, 9, -10, 48, 9, 0, -47, 5, 6, 0, 7, 28, 6, -5, -6, -8, 33, 1, 2, -20, 37, 6, 36, 3, 7, 17, 13, 13, 8, 3, 0, -41, -43, 25, -21, -3, -14, 0, 22, -1, 6, -7, -33, 6, -24, 36, 0, -2, -3, 19, -2, 2, 27, -4, -16, -7, 4, -20, 1, -37, 5, 3, -16, -24, -13, -20, 7, 6, 32, 77, 31, -4, -1, 3, 1, 7, -5, 7, -5, -7, 34, 18, -7, 22, -6, 0, -4, -9, -2, -18, -1, 0, -3, -21, -3, -22, -19, 20, 2, -2, -4, -14, -53, -12, 0, 41, 39, 7, 10, -26, -2, 12, 0, -4, 7, -5, 35, 1, 3, -5, 1, 5, 18, 5, 1, 42, 11, 24, -7, 34, 0, 18, 14, 20, 60, 3, -17, -21, 2, 7, 1, 27, -3, 0, 15, -5, -7, 7, 51, -29, 3, 6, -33, 12, 3, -2, -8, -32, -1, 11, 26, -49, 2, 23, -8, -69, -49, 3, 8, 15, -7, 23, 11, -21, 15, 16, 4, -8, -4, 21, 5, 32, -2, -41, 0, -14, 1, -13, 5, 1, -16, 3, -4, 6, -14, 31, 7, 7, 6, 17, 9, -5, 11, -6, 12, 5, -7, 17, -22, 3, -2, -1, -27, 28, -8, -35, 2, -17, 3, -2, -19, 10, 9, -7, -12, 17, 15, 1, 4, 35, -4, 31, 10, -3, -40, 1, 5, 0, -3, 7, -8, 8, -1, 2, 8, -2, -8, -4, -12, -26, -34, -17, 21, -31, 4, 2, 18, 7, 15, 9, -2, -12, -27, 78, 15, 0, 5, -10, 25, 7, -9, -2, 14, 6, -7, 10, 19, 20, 10, -5, 20, 20, 6, 0, -5, -13, 18, 1, -17, 5, -15, 23, -20, -5, -43, -7, -8, 29, 2, -14, 2, -4, 19, -3, -3, 12, -20, 25, -1, 5, -11, 2, 20, 28, 14, 18, -8, -3, -7, 10, -14, -39, -2, 25, 8, -30, -5, 10, -21, 0, -13, -6, -31, 17, -16, -1, 1, 30, -1, 11, -29, -32, 2, 40, -7, -6, 2, -7, 2, -4, -2, 11, -5, 13, -1, -16, -6, -4, -10, -27, -2, -8, 5, 0, -8, -17, 0, -7, -1, 13, 8, -11, -18, 4, -14, -6, -33, -5, 0, 24, 2, -1, -8, -23, -2, 39, -29, 0, -23, -62, 2, 10, 28, 19, -9, 25, -17, -17, 0, 0, -3, 17, -10, 44, 3, -17, 1, -15, 0, 4, -28, 7, 19, -8, 0, 0, -8, 28, 4, -3, 2, 2, -4, -60, 4, -24, -3, 1, -16, 4, -3, -34, -8, 5, -5, 31, -19, 0, -15, -27, 23, 5, -2, 40, -5, -22, 6, -2, 7, 7, -10, 9, 1, -1, 0, -3, -22, 16, -2, -5, 0, 3, -14, -3, -9, 1, -7, -5, 2, 50, 1, -21, -22, -5, -6, 12, -5, -2, -6, -41, -34, -1, 0, 39, -76, 5, 36, 0, 4, 6, -11, 6, -10, 20, 25, 14, -6, -29, -6, 21, -1, 1, -7, 3, -5, -2, -6, 5, -1, -1, -61, -24, 6, 9, -45, -13, -6, -20, -22, 5, -1, -30, -3, 14, 3, 2, -5, -3, 10, -19, 4, 8, -7, 16, -17, -6, 7, 22, -4, -20, 0, 4, 2, 60, -19, 6, -6, -4, 0, 14, -18, 3, 9, 4, 24, 2, -24, 34, -5, 6, 4, -16, -9, 33, 18, -1, 35, -13, -6, -7, 23, 20, 11, 1, 37, -15, -44, -6, -7, -16, 25, 25, 7, -10, 34, -5, 0, 5, -3, -7, 9, 6, 41, -7, 0, -10, 4, 7, -3, 3, -17, -1, -2, 4, -8, 9, -6, -33, -2, 2, 2, 3, 7, 1, -38, -4, 8, 9, 31, -18, 4, 3, -18, 13, 13, 6, 9, -6, -32, 9, -10, -1, -20, 3, -13, 4, -7, -13, 13, -35, 5, 17, -15, 9, -18, 12, 0, 4, -4, -38, 3, -9, -4, 0, 8, 0, 6, 2, -2, -18, 29, 22, 30, -1, -32, -22, 0, -4, -18, -1, -2, 11, 16, -9, 7, 32, -1, -49, -7, -1, -6, -18, -1, -94, 56, -21, 5, 23, 3, 0, 0, 26, 2, 25, 14, -6, -8, 8, 2, -11, 2, 6, -14, 17, -5, 9, 4, -23, -49, -31, -3, 14, 17, 11, -13, -7, -63, -8, -4, 3, -55, 6, -5, 0, 10, -24, -29, 21, -18, -16, 3, 0, 8, 1, 14, -9, -13, -7, 16, 3, -5, 18, 46, 16, 63, 5, -7, -7, 0, -2, -3, 8, -7, -1, -9, 0, 5, -3, -13, -8, -20, -39, 43, -8, 39, 11, -5, 24, 3, 1, 32, -6, -6, 19, 15, 14, -25, -18, 29, 13, 0, -5, -7, -2, 65, 4, -3, -7, -5, 40, 1, 2, -20, 42, 1, 8, 0, -15, 12, 28, -16, 0, -23, 21, 3, 1, 14, 0, -32, 38, -11, 9, -3, 0, -7, 34, -5, 4, -31, -5, 8, -4, -24, -31, 12, -1, -3, 45, -26, -6, -14, -25, -28, -15, 5, -11, -34, 6, -14, 18, -22, 0, -29, 8, 9, 5, 5, 4, 8, -10, 10, 0, 5, 5, -3, 7, -7, 7, -2, -33, 0, 4, -14, 3, -2, -8, -31, 4, 0, -4, -9, 20, 0, -6, 0, -7, 0, 20, 2, -3, 3, 42, 9, -12, -6, 5, -1, 6, -39, -6, -24, -17, 0, -12, 22, 29, 6, -18, 17, -2, 11, -26, 3, 8, 1, 8, -2, 15, 4, -3, -30, 2, 4, 18, -12, 12, 4, -13, -4, 12, 0, 37, -2, 19, 13, 3, -3, -11, -6, -13, 6, 22, 32, -23, 18, -20, 1, 10, -15, -25, 12, 1, -2, 3, 3, -6, 0, -15, -10, 4, 3, -7, 33, 5, 1, 20, 14, -47, 7, 7, -6, 1, 52, -19, 3, -8, 3, 2, 9, -31, -7, -1, 6, -9, 1, 0, -4, 0, -6, 5, -7, 52, 1, -5, -9, -11, -4, -6, -17, -9, -6, -14, 5, -6, -2, 44, -17, -1, 31, -5, 12, 3, -4, 5, -11, 13, 43, 0, 5, -16, 19, 33, -4, -1, 0, 6, -4, -15, 9, 6, 0, 7, -3, -20, 4, -7, -28, -10, 0, -5, -28, 5, -1, -1, 21, 17, -27, 1, 1, -13, -3, 11, -6, -36, -24, -24, -25, 5, 0, -58, 20, -11, 1, -2, -10, 22, -55, 2, -17, 4, -13, -47, -57, -7, -3, 0, -3, -4, -15, 21, -5, 0, -20, 27, -14, 18, 8, 0, 12, -6, 3, 36, -10, 50, 4, 5, -12, 34, 39, -26, -1, -13, 30, 20, -16, -20, -26, -8, -6, -1, -2, -1, 3, -8, -7, 11, -9, 11, 4, 10, -9, 0, -21, 1, -6, 4, 1, -62, -37, -1, -34, -2, 3, 6, -11, -11, -37, -12, -6, 1, -23, 0, 33, 0, 1, 4, 1, -32, 4, -8, 3, -1, -1, 0, -20, 0, -15, -5, -6, 27, -26, 26, -6, 0, 14, -4, -56, 21, 13, -4, -5, -2, -17, 0, 0, 0, -23, -6, 0, 4, 3, -23, -28, 42, -18, -5, 28, 9, -7, 4, 14, -21, -3, 5, -19, -52, -5, -22, -9, 3, -14, -1, 4, 15, -2, -13, 46, -18, -28, -8, -5, -5, -5, -4, -29, 25, 9, -19, 17, -8, -1, -15, -4, -3, -42, -16, 5, -6, 4, -30, 45, 0, -4, 7, 21, -49, 26, 3, -11, 0, -5, 17, 17, 5, 0, -3, -37, 40, 2, -29, 13, 1, 19, -5, 20, 2, -24, 2, -8, -7, -13, 4, 16, -24, 2, -6, -15, -1, 29, -7, 6, 7, -4, 0, 7, -10, 7, 15, -4, -9, -32, 1, 27, 41, -12, 16, 14, -17, 17, -44, 7, 2, 1, -33, 9, 19, 5, 3, -50, -9, 15, -18, 2, 0, -7, -3, 15, 5, 1, -32, -9, 20, 11, -5, -36, -22, 6, -2, 22, 8, 5, 29, 15, -3, 7, -47, -5, -6, 40, -5, 19, -30, 4, -10, 0, 4, -12, 29, 7, 28, -44, -30, 25, -5, 6, 26, 32, 24, 0, -2, -24, -2, -3, 40, 9, 0, 6, -1, 47, -20, -36, 5, 16, -5, 6, 0, -31, -12, -13, 24, -6, -5, 6, 4, 36, -6, -6, -20, 7, -19, 3, 2, -8, 0, -14, 0, 6, -21, 34, -10, -9, 4, 4, 20, -5, -3, 6, -15, 1, -1, 1, 0, 7, 21, 0, 6, 27, 7, 3, -5, -2, 6, -14, -4, 20, -3, 1, 30, -10, -45, -33, -3, 24, -102, -5, -4, 27, 43, -7, 15, 6, -17, -36, 0, -2, -75, -5, 0, 3, -62, -11, 46, 10, 5, 2, -40, 26, 2, 0, -5, 4, 54, -11, -28, 6, -6, 9, 17, 1, -4, -8, -10, -1, -2, 5, -32, -1, -40, 4, 0, 19, 5, -21, -38, -8, 0, -5, 19, -8, -40, -6, -3, 0, 2, 30, -5, -8, 6, 4, -7, 21, -9, 5, -5, -9, -15, -10, 6, -7, -3, 3, 3, 4, -7, 3, 9, -28, 0, 8, -8, 29, -5, -5, 65, 33, -4, 5, 1, -8, 9, -17, 7, 41, -3, -4, -8, 50, 4, 18, -2, -6, 24, -1, 6, -3, -9, -7, -1, 8, -43, 0, 6, 5, 9, -27, 25, -1, -3, -2,
    -- layer=3 filter=0 channel=1
    -1, -5, 6, -7, 5, 8, 6, 30, -7, 16, 0, 10, -2, 29, 0, 2, 39, -20, -11, 14, -5, -5, 20, -26, 65, -16, -8, 1, -3, 2, 27, -10, -4, -4, -28, -4, 9, -8, 5, 10, -4, -8, 4, -1, -12, -12, -27, -19, -1, 8, -4, -2, -1, 8, 16, -44, 3, 0, -3, 9, 33, 6, 63, 8, -4, 6, 27, -4, 3, -21, -4, -5, 2, 6, -1, 13, -3, -28, 9, -4, 6, -2, 11, -7, 4, 16, 13, -6, 9, 6, 8, 8, -32, -13, -25, -4, 0, 3, 6, 22, 13, 7, 15, 11, 23, -39, 51, 0, -21, -8, 10, -11, -9, 5, -5, 0, -5, -12, 4, -3, -4, -6, 19, 15, -1, 3, 15, -16, 14, 22, -13, 6, -9, 1, -1, -1, 1, 6, 49, -7, 1, -3, 2, 7, -12, -6, 16, 17, -9, -33, -16, -8, -11, 24, -29, -4, -10, 1, 0, -2, -20, 0, -16, 0, -8, 2, -22, -2, 0, 1, 48, 17, 13, -6, 0, 4, -2, 67, -9, 30, -26, -13, -13, -7, -8, 3, -13, -5, -16, -2, -4, 27, 6, -18, -23, -4, 2, -18, 4, -35, 24, 40, -2, 0, 19, 12, -26, 3, -6, 8, 4, -23, -8, -11, -11, -4, 3, -1, 2, 16, -8, -12, 19, -20, -1, -8, -4, 18, 15, -3, 12, 12, -3, -1, -8, -9, 6, 15, -7, -5, -24, -4, -3, 15, 4, -18, -24, 8, -43, 60, 7, 9, 11, -23, -6, -5, -35, -3, 1, -2, 8, 69, -15, 0, 8, 0, -6, 6, -2, -11, -6, 3, -18, -41, 5, -14, -12, -2, -2, 8, 3, 6, -24, 1, 0, 9, -2, -8, -27, 0, -2, 11, -2, 1, 8, -4, -23, -1, 4, 22, -16, 3, 13, 2, -39, -4, -2, -1, -4, 0, -42, 48, 0, 12, 2, 5, -43, -40, -1, -2, 6, 11, -39, -14, -25, -12, -4, -26, -7, -24, 13, -28, 0, 1, -16, 1, 8, -35, -7, -22, 19, 8, -14, -1, -54, 1, -4, 8, -17, 7, 35, -15, 2, -2, -7, -2, -22, -3, -3, -3, -3, -2, -34, -10, 4, -15, 9, -8, -15, 13, -7, -13, 5, -17, -7, -9, 10, -19, 4, -1, 3, -5, 15, -8, -2, -6, 38, 9, 4, 9, -40, 9, 4, 2, -24, -1, -7, -13, 35, 2, 12, 6, -36, 0, 22, 0, 16, 45, -41, -14, 3, -16, 17, -1, -7, -7, -17, 26, -32, 23, -8, -4, 17, 8, 20, -8, -5, -6, -1, 2, 15, -4, -31, -12, 7, -22, -17, 12, 5, 4, -10, -1, 57, -5, 5, 5, -4, -84, 22, 2, -18, 11, -51, 22, -10, 4, 0, 1, -2, -19, -3, -7, -5, 1, -6, 5, 7, 0, 13, -10, 1, -6, -28, 6, 9, 4, 5, -8, 7, 7, 2, 15, 2, -11, -6, -4, 3, 2, -5, 27, 8, 6, -2, -1, 19, 2, 14, 4, 3, 0, -6, 1, 18, -4, 1, -8, -6, -14, -14, -2, 2, -30, -24, -5, 2, -8, 7, 8, -3, -16, -15, -2, -4, 4, -6, -13, 2, 0, 13, -48, -2, -37, 4, -8, 17, 10, 2, -32, -6, 4, 19, 3, 15, 1, 7, -43, 2, -40, -5, -1, 3, 6, 6, 4, 11, 6, -11, -16, 6, -5, -17, 18, -6, -2, 0, 8, -5, -37, -1, 9, 7, 18, -30, 0, 13, -4, -5, 18, 18, -44, 1, 18, 5, -4, -5, 2, 0, 3, 0, 5, -8, -9, 1, 3, 15, 0, 6, 28, -12, -2, -1, -9, 25, -1, -30, -22, 4, 3, 8, 5, -22, -27, 21, 6, -22, -3, -7, -7, -10, 9, 1, -22, 6, -10, -1, 0, 4, 4, 1, 23, -5, -2, -1, 5, -4, 9, -59, 0, 0, -8, -5, 8, 5, 29, -6, -2, -17, -16, -4, 1, 33, -8, 3, 7, 0, -1, 20, -9, 26, -28, -3, 24, -4, -2, -14, 18, -5, -3, -7, -9, -3, 4, -19, 0, 15, -20, 1, 4, -59, 0, -25, -27, 10, -47, 9, -3, -2, -2, 12, -36, -41, -27, -3, 4, 3, -1, 3, -5, -19, 10, 19, 6, 6, 38, 10, -36, -10, -9, 3, -20, 4, 0, 7, 10, 0, 1, 36, -8, -16, 3, -8, -17, 0, -6, 12, 8, 5, -23, 4, -22, 4, 20, -6, -15, -26, -4, 8, -7, -22, -42, 23, -11, -2, -27, -9, -1, 2, 0, -10, -21, -19, -1, 13, 2, 6, 0, 4, 17, 13, -6, -42, 31, 8, -55, -29, -28, -5, 30, 20, -15, -36, -21, -28, 5, -12, 2, 3, 23, 7, -7, 6, 14, 1, 0, -19, -7, -19, 17, -1, 1, -9, -5, -3, 33, 27, -12, -19, 0, -5, 3, -10, -1, -3, -2, -6, 36, -3, -8, -17, -6, -5, 38, 25, -6, -49, -38, 3, 29, -2, -48, -27, -24, -3, 34, 5, -23, 1, 1, -3, 24, 14, 2, 3, 11, -12, 28, -15, -14, -4, 0, -7, -4, 9, 3, -15, -4, -11, 13, 4, -9, -3, 5, -23, -1, 6, 3, 21, 3, 0, 0, 4, 0, -18, -48, -10, 8, -11, -5, 16, 4, 9, 3, -6, -6, 21, -4, 5, 21, -24, -4, 7, 35, -8, -1, 8, -20, 7, -56, 13, 23, 3, 4, -31, -1, 24, 21, 6, -16, -16, 0, 0, -47, -15, 2, -16, 14, -18, 0, 13, -13, -1, 15, -5, -6, 16, 2, -12, 6, -37, -7, -37, 32, -2, -25, 26, -5, -27, 2, -13, -8, -5, 42, -10, -5, 6, 11, -18, -5, 3, -5, -11, -7, 1, 10, -5, -19, -1, 3, 6, 0, 0, -2, 7, 8, 3, 10, -3, -5, -4, 5, 21, -6, -6, 13, -29, 29, -20, -7, -5, -6, -8, -4, 5, 5, 0, 4, 3, 3, -40, 2, 38, 4, -2, 2, -33, -21, -5, 0, -5, 14, -7, 5, -2, -28, 17, -52, -8, 16, -7, 3, -3, 12, 5, 0, -6, -3, -22, 19, -23, -1, 2, 7, 5, 0, -13, -8, 2, -5, 0, -10, -24, -13, 0, -33, -29, -2, 23, 15, -1, 5, 1, -23, 11, 33, 2, -6, -5, 11, -8, 0, 13, -24, -11, 43, 0, -4, 6, -8, 2, 3, -6, 7, -31, -4, -8, -21, 3, -34, 15, -1, 6, -3, -1, 26, 1, -12, -1, -6, 3, -1, -17, -27, 6, 7, -4, 31, -3, -2, 2, -9, 9, -1, -9, -4, 16, 3, 7, 4, -4, 10, -27, -20, -10, -36, 0, 0, 0, 6, 2, -6, 10, -25, 15, -6, -12, -5, 1, 3, -3, 23, -4, -5, -1, -2, 44, -20, -26, 19, -20, -2, 4, 6, 20, 11, 6, -4, 25, -20, 7, 9, 1, 7, 1, -59, -4, -5, -4, 17, -2, -8, 5, -12, 3, -12, 0, -7, 50, 23, -21, -3, 31, -14, -13, -12, 14, 10, -13, -2, -12, -8, -6, 5, -41, -24, -5, -6, -2, -6, 10, 17, 23, 0, 1, -9, -3, -7, -13, -28, -20, -5, -8, 2, 12, 4, -30, -1, 3, -8, 2, 0, -4, 2, -16, 3, 27, 0, 7, 6, 2, 0, 0, 12, 1, -14, -6, -17, -7, -4, -13, -1, -16, 9, 13, -6, -7, 2, -13, 14, -43, 3, 1, -3, -61, -9, -16, 46, -3, 5, -13, -34, -7, 9, 0, -23, -17, 12, -6, -8, -25, 11, 0, 3, 0, 6, -6, 4, 12, 19, -7, 0, 43, 32, 9, -11, 23, -8, 5, 5, -7, -1, 4, -11, 17, -7, -39, 1, 5, 12, -1, 9, 1, 20, 18, -13, -43, -41, 9, 53, -3, 11, 4, 0, 10, 19, -14, -20, -30, 1, 11, 43, -5, 0, 4, -20, -1, 1, 12, 27, -42, 25, 4, -38, -17, -4, 8, 0, 22, 56, -6, -2, 0, 25, 8, 2, 3, -18, -4, 9, 16, -6, -31, -1, -8, 20, -13, 6, 5, 4, -3, 0, -4, -32, 42, -33, -16, 43, -13, 12, 6, 5, 19, -27, -27, 4, 30, -12, -25, 5, -12, 14, -4, -35, 9, -24, 27, -2, 7, 0, 16, 2, 8, 17, 7, -14, 31, 7, -3, -1, 39, -4, -3, 1, 9, 3, -3, 9, 8, 9, 4, 5, -8, 1, 10, -2, 8, -5, 6, -1, 4, -14, -15, 5, 4, 4, 0, 0, 3, -8, -8, -17, 2, -8, 4, -3, -13, -1, -14, -2, -4, 58, 34, 0, -7, 30, 7, -1, -7, 9, -8, 0, -19, -4, -67, 7, -11, 6, -33, -9, -6, -13, -1, 35, -13, -23, -8, 24, 0, 4, 0, 2, -8, -5, 7, 24, -17, -5, -23, -18, -18, -2, 5, -8, -31, 0, 5, 6, -13, -2, -1, 2, 16, -4, -3, 3, -3, 2, -22, 2, -3, 14, -6, -11, 37, 10, -11, 0, -14, 38, -20, -6, 0, -1, -21, -10, -10, -6, 5, 10, -4, 4, 12, -6, -2, 20, 0, -6, -31, -14, -3, -6, 11, -13, 0, -1, 12, 14, 35, -46, 9, -9, -1, -37, 2, 34, 18, -11, -1, 7, 29, 6, -22, 0, -5, -6, -2, 0, -9, -9, -9, 5, 5, -18, 19, -3, 1, -35, -36, -8, -64, 18, 4, -1, 16, 6, -39, -37, 5, -3, -3, 32, 0, 3, -18, 32, -15, 3, -4, 0, -7, -29, 11, 0, 5, 3, 24, 42, 9, 17, 0, -2, 15, 32, 2, -2, 4, 14, 5, -24, 2, -2, 0, -18, 47, -12, -30, 35, 7, 28, 0, 0, -18, 25, -27, -4, -5, 13, -3, -25, 27, -6, 0, 1, 40, -40, 1, 40, 1, 0, 5, -6, 1, 5, 0, 4, 28, -12, -11, -1, 4, -8, -5, -2, 3, 8, 7, 5, 6, -7, 19, -25, -5, 0, -2, 6, 5, -11, 2, 0, -26, -6, 13, 8, 14, 9, -13, -4, -49, 14, -10, -6, 2, -3, 7, 45, -4, 28, 0, -2, -4, -8, -32, 3, -36, 13, 9, 9, 13, 29, 0, -10, -30, -4, 1, 3, -57, -10, 9, 8, 0, 0, -24, -24, -4, -28, 7, -24, -38, 4, 0, 37, -26, 4, -5, 26, 22, -6, 9, 4, 14, 17, -10, -5, -14, -1, 0, 22, -43, -6, -54, 2, 1, 4, 22, -12, 20, 38, -16, -17, 5, -5, 1, -2, -2, -67, 11, -9, 17, -11, -15, -60, 0, -1, -5, 13, 1, -12, 12, -20, 6, 6, 3, -39, -6, -8, 2, 3, 24, 6, -31, 29, -31, 6, 3, -3, 8, 3, -9, -5, 0, 26, -3, -6, -35, -15, 3, 10, 5, 0, -4, -6, 0, -7, -6, 0, -9, 3, 14, 0, 4, 7, 3, 25, 14, 8, -28, -13, 36, 46, -20, 17, -2, -18, -17, -7, -24, 28, -9, -11, -33, -2, 32, 21, 1, -8, 0, 28, 8, 7, 7, -48, 14, 7, -11, 16, -35, -4, 14, -1, -16, -46, 0, 2, -8, 24, -3, 7, 10, 12, -4, 15, 26, 5, 31, -6, -5, -7, -5, -1, 12, -13, -31, -13, -1, -20, 39, -4, 19, 49, -4, -27, -5, -9, 10, 27, 0, -6, -21, 2, -19, 14, -1, -10, -6, 24, 4, 34, 17, 16, -9, 5, 22, 5, -6, 7, 3, 4, 1, 6, 0, 0, -74, -4, -4, 17, 20, 2, 30, -54, 16, 0, -9, 1, -2, 6, 3, -3, -10, 7, -25, 7, 4, 18, -1, -1, 19, -35, 0, -4, -1, 16, 5, 11, -17, -23, 2, -10, -31, 7, 0, -32, -6, -23, 47, 6, -1, -21, -22, 0, 29, 18, 5, 33, -33, -10, -71, 2, -2, 3, -28, -1, -44, -4, -29, 51, -15, 0, -2, 10, 24, 2, 22, 7, -2, -5, -33, 27, 3, -10, -22, 10, 1, -9, 0, 0, 26, 3, 7, -5, -8, 21, -7, -4, -53, -8, -2, 3, -5, 30, -11, 1, 0, -3, 6, 13, 4, -8, -3, 11, 0, 17, 4, -3, -3, 0, 5, -18, 0, 5, 6, -6, -9, -5, 17, 7, -11, 12, -5, -4, 21, -29, -3, -8, 33, -2, -7, 0, -29, -9, -37, 33, -4, 10, 8, -13, 2, 45, 1, -16, 6, -9, -26, -12, -32, -9, 10, 2, 7, -1, 5, -2, 2, 5, -2, -11, 46, -8, 1, -3, -15, -5, -73, 23, -5, -6, -5, 13, -12, -2, -2, -1, -2, -36, 30, -4, 31, -7, 11, 12, -4, -3, -64, 25, 24, -7, 4, 1, -31, 8, -37, 37, 6, -6, -22, -30, -3, 1, -4, 39, -7, -11, -34, -6, -7, -2, 22, -5, 18, 0, 7, -5, -5, -6, -21, 4, -7, -5, 5, 9, -46, 39, -49, 5, -17, -14, -7, 5, -6, -23, 4, -1, 2, 0, -4, -1, 7, 37, -58, 2, 13, -2, -20, -4, 9, -24, 3, -2, 0, -5, 8, -35, 21, -93, 4, -6, 4, 2, -4, -37, 17, 4, -2, 2, 17, 34, -41, 6, 5, 3, -87, -4, 2, -31, 6, 5, 0, -1, 4, 13, -6, 1, 0, 20, -28, 6, -12, 0, 8, 36, -11, 55, 8, 0, -18, -17, 0, 3, -43, -11, 11, -5, -1, -4, 0, -24, -5, 6, 1, -11, -9, -2, -2, 18, -5, 7, 1, 35, 18, -9, 14, 6, -30, 9, -1, -6, 20, 0, -14, 10, -53, -2, 10, 3, -2, -7, -9, -22, 25, 10, -2, -11, 16, -2, -4, 5, 10, -24, 28, 6, -3, -13, 15, 8, -6, 9, 8, 9, 60, 22, 2, -41, 1, -4, 22, -29, -16, 1, 5, -27, 28, 6, 8, 33, -6, -43, -5, -18, 9, 17, 3, 6, -22, 2, 1, 10, 6, 24, 3, -2, -9, -13, -4, -3, 3, -3, 2, -44, 1, -7, 31, 0, 8, 1, -9, -32, 43, -29, 6, -42, 32, -18, 0, -6, 6, 4, -16, 4, -29, -51, 10, -38, -20, -6, 23, -3, 17, -9, -1, 5, 0, -5, -46, -15, -41, -2, -11, 2, -66, 0, 1, -1, 24, 6, 14, 25, 3, 55, 24, 3, 0, 0, 2, 1, -24, 0, 20, 2, -1, 0, -24, -6, 14, -16, -15, 15, -4, -27, -5, -7, -2, 33, -13, -55, 1, 3, 1, 7, -25, 3, 6, 10, 6, -1, -11, -33, 0, -25, 2, 21, -4, 23, -38, -12, 12, -7, 1, -5, 8, -3, 2, 0, 5, 1, -41, 7, 10, 3, 11, 5, -45, 57, 11, -4, 2, -12, 0, -1, 5, 3, -12, 6, -40, 3, 4, 23, 13, 4, -8, 15, 1, -7, 2, 4, 1, 12, -56, 14, 8, -8, 41, 5, -8, -17, -3, -38, 9, 10, -10, 10, 0, -4, 12, 36, -16, 15, -45, -4, -33, -1, 19, -11, 3, -9, -5, -12, 20, -45, -5, -9, 1, 9, 8, -4, -16, -3, -9, 3, -8, 7, -37, -1, -58, 31, -96, -15, -5, -5, -15, 5, -14, 7, 14, -5, -2, 35, -15, 8, 0, 3, -7, -12, -18, -8, 3, -12, 1, 32, -65, 0, -8, -1, 4, -19, 28, -3, -3, 6, -1, -21, -7, 5, 0, -9, -8, 6, 0, 2, 17, 22, -3, -2, 0, -32, -6, -8, -15, 8, -6, -2, -45, 12, -43, -9, -8, 28, 0, -7, -6, -2, 7, 23, -8, -1, -40, 35, -27, 4, -7, 4, 2, -1, 3, 10, 8, 8, 0, -5, 36, -6, -6, -15, 21, 9, -58, 27, -7, -7, -14, -9, -3, -14, 8, 0, -2, -11, 14, -5, 18, 0, -27, 19, -2, -5, -42, -5, 9, -34, 8, 4, -33, 47, -11, 8, 0, 2, -18, 26, 1, 11, 4, 26, -1, -27, -46, 0, 7, -17, -65, 48, -18, -63, 5, 24, -1, 0, -16, 14, -28, -11, -7, 28, 19, -12, -26, 2, 6, 41, 17, -9, 0, -37, 5, 1, -4, -4, 0, 0, -2, 41, -9, 0, -32, 6, 15, 4, -7, -57, -6, 2, 10, -9, 54, -59, -28, -41, 1, -3, -8, -7, -11, 6, -10, -3, -57, -17, 8, 17, 1, -1, 26, -8, -39, 7, -2, 7, -1, -3, 7, -8, 5, 0, 6, 4, -4, -1, 5, -4, -50, -1, -23, 24, -28, 10, -19, 4, -34, -14, -8, 2, -28, 7, 4, 11, -7, 3, 11, -8, 33, -8, 10, 3, -14, -6, -11, 52, -28, 8, -1, 0, 8, -7, 0, -4, -58, 12, 5, -1, -11, 4, -20, -3, -4, 31, -8, -5, 1, -5, 18, 12, -5, -39, 12, -19, -1, 9, -9, 2, -7, 34, 0, 0, -9, 7, 2, -42, 0, -4, 1, 12, 3, 28, -28, 11, 6, -6, 8, -81, -14, 9, -8, -2, -3, -23, -52, 4, -28, 35, 5, -6, 2, -21, 0, 0, -1, 39, 3, 10, -26, 23, 24, 21, 4, 11, -3, -5, 5, -6, 0, -12, 5, -5, -36, 9, 3, 14, -1, -40, 13, -30, -34, -6, -51, -7, -18, 43, -8, -19, -25, -1, -3, -62, 44, -20, -6, 2, -18, -3, 0, -5, -7, 11, 0, 4, -46, 13, -15, -14, -1, 16, 25, 5, -4, 40, 1, 6, 28, 27, 4, 37, 3, -1, -3, -37, 2, 7, 54, 8, -68, -1, -5, 2, 19, -7, -46, -35, -13, 3, -7, -4, -2, -8, -15, -29, 11, -70, -12, 1, 4, -41, -44, -6, 14, 9, -33, -10, -18, -60, -2, -3, -1, 2, 4, 43, -60, 3, -12, 7, 1, -46, 8, 26, -16, 1, 4, -4, 10, -5, -3, -23, 1, 0, -29, -58, 17, -2, -15, 7, -12, -6, -1, 2, 1, 8, -40, 8, 4, 18, -28, -4, 4, -21, -4, -10, -3, 25, -8, -2, -2, -24, -3, -27, -13, -4, -28, -48, 0, 24, 23, 3, -4, 24, 0, -7, 35, -16, -27, -2, -12, -3, -9, -2, 20, 6, 24, -9, 52, -8, 25, -56, 12, 1, 4, 25, 1, -7, -28, 7, -24, 8, -59, -14, -11, -6, -32, -7, -66, 4, 0, -3, 11, 8, -25, -7, 18, 16, -5, 29, -21, 20, -4, -4, 3, 5, -16, 5, -4, -18, -3, -15, -15, 8, -5, -7, -42, -9, -22, 2, -9, -4, -8, -12, 9, 0, 2, -2, -12, 6, -15, -7, -22, 12, 2, -2, 4, -24, 7, 7, -33, -4, 0, -3, 7, -25, -10, -40, -5, 41, 4, 17, -8, -8, -1, -24, 0, 1, 17, -1, -39, 0, -6, -2, -4, -7, -21, 0, -4, -6, -7, -10, -25, -3, -4, -57, -34, 6, 3, 11, -1, -5, 14, 16, -9, -6, 3, 3, -8, -7, -29, -6, 53, -27, -24, -29, 1, 8, -13, 0, -58, 9, 4, 0, 32, -23, 0, 47, -2, -50, 17, -5, -4, -5, 3, -73, 8, -6, -24, -4, 8, 0, 13, -10, 0, 2, 5, -10, 0, -3, 11, -25, -2, 0, -9, -27, -3, -37, 9, -2, -21, 22, -24, -31, 0, 21, 0, -1, -3, 9, 7, 2, -3, -15, -25, 6, -10, 5, 7, 9, -1, -1, 4, -6, 8, 0, 0, -21, 9, -8, 13, 2, 3, -3, -17, -27, 15, 4, 1, 16, 18, -19, -17, 4, 15, 3, -36, 0, 0, -53, 3, -5, 6, 8, 10, -9, -6, -7, -45, -5, 12, 5, -20, -3, -39, -23, -60, -13, -7, 29, -21, -12, -5, -12, -51, 8, 2, -8, -7, 5, -30, -77, -19, 1, 1, 23, -4, 0, -4, -17, -20, 0, -4, -30, 35, 3, -17, -1, 17, -36, 8, 5, -14, 6, 0, 19, -16, -56, -12, 7, 1, 9, 35, 16, 18, 30, 37, -14, 1, 5, -13, -2, 2, -42, 4, 1, -5, 10, -60, 56, 32, 8, -1, -10, 24, 2, 1, -38, 0, 6, -24, -30, -9, 6, -1, 15, -18, -13, -22, 34, -22, 9, -7, 19, -1, -32, -6, -1, 11, 35, -2, -4, -57, 13, -28, -19, 23, 41, 4, -5, -4, -6, 0, -54, 22, -3, -40, -4, -6, 21, 4, 29, 0, -43, -11, -17, 44, 23, -4, -11, 4, -43, -70, -13, -39, 20, 9, -48, -14, 6, 17, -26, 0, -6, -1, 14, 0, 4, 20, -13, 56, 20, -10, -76, 10, 3, 2, -38, -7, -10, 5, -25, 6, 59, -37, 0, -7, 38, -11, 8, -65, -8, -44, -11, 1, 0, -48, -5, -35, 35, -28, 11, -1, -29, 13, -29, -21, 36, -15, -15, 1, -3, -57, 3, -34, 7, -25, 9, 2, 6, 8, 26, -3, -5, 5, -17, -13, 0, 26, -4, 3, -5, -8, -50, 1, -3, -3, 0, 16, -9, -66, -6, -3, 16, -40, -7, 11, -9, 14, 8, -4, 0, 16, -7, -2, -2, 3, -5, -29, 4, 4, 14, -17, -8, 9, 6, 0, 12, 1, 40, -3, -33, 11, -15, -4, 5, 17, -5, -50, -85, -6, -30, -22, 6, 4, -22, -8, -4, 27, -15, -40, 6, 17, -3, -41, 10, 0, -4, -37, -4, -29, -5, 15, 5, -13, -32, -2, -3, 4, 0, 21, 4, -17, 0, -51, 47, -1, 5, 13, 0, -37, -18, -7, -6, 21, -8, 19, 6, 8, -27, 0, 20, -6, -26, 2, -13, -29, -6, -16, -7, -4, -15, 5, -11, -42, 6, -9, -4, -69, 19, -20, 1, -2, -2, 1, 0, 1, -9, -6, 0, 0, -12, -15, 4, 17, 24, -5, 5, -43, 5, 1, 0, 27, -2, 3, -5, 33, -18, 23, 0, 3, 29, 1, -39, -8, 74, -3, 3, 0, 9, 6, -55, -23, -3, -2, -5, 4, 0, -22, -9, 2, -1, 3, 20, 34, 4, 1, 35, 37, -5, -21, 37, 3, -4, -48, 14, -21, -27, 7, 0, 2, -28, 23, 7, 36, 29, -25, -10, 6, 7, 6, -2, -73, 42, 4, -6, -30, 46, 6, 24, 1, -8, 29, -18, -2, 3, -6, 26, 4, 43, -33, 2, -2, 4, -35, 14, -15, -18, -4, 0, -8, -1, 29, -38, 9, -16, -5, -7, -16, -84, -15, -2, -16, 9, -18, -19, 0, -1, -7, 5, 19, 8, -6, -6, -3, 67, -5, -5, -1, 8, -1, -4, 0, -35, 0, 4, 1, 7, 29, 0, 9, 21, 21, -3, -3, 3, 0, -38, 25, -1, -29, -23, 20, -22, 14, 17, 11, 31, 10, -8, -6, 26, 4, -6, -4, -7, -3, -61, -10, 3, 33, 22, 32, -9, -16, 10, 24, -25, -53, -14, 3, 6, 4, 4, 4, 1, 6, -25, -6, 3, -8, -8, 22, -30, -13, -47, 6, -17, -31, -7, 2, 5, 5, 7, -4, 9, 33, 7, -8, 0, -3, -29, -1, 9, 23, 0, -7, -8, 6, -23, -25, 5, 2, -2, -14, 17, 23, 3, 44, 0, 39, 4, -13, -7, 4, 18, -14, -1, 1, -33, 26, 3, 15, 0, -7, 34, 0, 9, 4, -5, -1, -3, -25, -47, -13, 3, 15, 12, 11, 8, -27, 2, -5, 5, 0, -2, 5, -12, -2, -4, -50, 20, 6, -15, -19, -14, -25, 38, -11, 12, 0, -8, 4, -3, 3, 27, -19, -5, 10, 6, -3, 7, -2, 16, 23, 3, 29, 4, -6, -31, 4, 34, 6, -35, 16, 2, -25, -49, -16, -30, -13, -5, -24, -11, 3, -4, 1, 48, 3, -9, 43, 38, -9, -2, -5, 43, -22, 0, -6, -2, -9, -32, 11, 30, 0, 20, -73, -8, 0, -21, -1, 43, -19, 5, 16, 0, -4, 9, -24, -8, 15, 34, 20, 22, 7, 28, -12, -13, -31, -25, -15, 12, 2, 1, -9, -24, -34, 1, 7, -20, -17, -21, 11, 13, 8, -10, 0, 1, -29, 21, 31, 4, 20, 1, 7, -29, 3, 40, 23, -4, 14, 4, -15, 3, -9, 6, -8, -7, -36, 31, -9, 1, 9, -11, 2, 0, -8, -4, 0, 3, -44, -8, -3, 10, -14, -6, -15, 20, -3, 3, -11, 45, 3, 27, 11, -33, 0, -21, -31, 2, 17, 12, -4, -5, 16, -1, 1, -49, -23, -2, 11, 20, 19, 25, -3, -1, -9, 9, 9, 4, 29, 6, -30, 5, 21, -5, -43, 15, 1, 13, -6, -2, 5, -7, -50, -30, -47, -7, 18, -6, 23, 33, -17, -13, -6, -4, -19, -1, -23, 3, -16, 11, 0, 18, 20, -30, 3, 2, -31, -3, -11, -7, 9, -13, 1, 0, -14, 2, 0, 21, 29, 4, -33, 0, -2, -9, -3, -14, -5, 5, 0, 1, -1, -9, -36, 4, 3, 16, -10, -1, -9, -67, 4, 3, 10, -7, 1, 1, -9, -10, -16, -7, -6, 45, -1, 7, -1, -4, 0, -24, -7, -3, -39, 6, -23, 0, 5, 5, 3, 3, 2, -3, -2, 6, 7, -37, 9, 8, 6, 62, 17, 0, 9, 39, -6, 0, -10, -6, -48, -53, -6, -4, 1, -11, -17, -6, -8, 32, 5, 3, 7, 5, 2, -6, -29, 41, -8, 4, 27, 15, 15, 49, 7, -19, 23, 22, -5, 13, 5, 4, 10, -4, -20, -5, 3, -15, 8, 32, -9, -51, 4, -15, -4, 1, -33, 10, -15, -4, -8, 48, -20, 35, -28, 7, 22, -82, -14, 60, 0, -5, -4, 0, 2, 0, 7, 3, -9, 23, 4, 6, -22, 6, -4, -7, -6, -34, 0, 13, 7, -2, 41, -24, -36, 6, 27, 9, -7, 0, 2, -11, 2, -7, -34, -48, -37, -48, 35, 14, 25, -1, -20, 0, -9, -43, 0, 3, 0, -55, 1, -1, 5, 2, 14, 11, 17, -5, -31, -12, -30, -32, -3, 7, 1, 23, -29, 6, 6, -5, -16, -16, -3, 8, 0, -2, -5, 0, -8, 12, -9, -39, 8, -10, 2, -23, 9, 0, 1, -30, 30, -2, -42, 0, 4, -4, 2, -2, 19, -5, -5, -11, 18, -10, 8, 4, 3, 1, 5, -16, -10, 5, 50, -15, -1, 1, -6, 6, -7, 22, 23, -1, 5, -32, 5, -18, 17, 5, -7, -26, 22, -16, 7, -29, 7, 0, -19, -44, -2, -4, 8, 56, 28, 27, 24, 16, -4, 11, -2, 16, 8, 13, 1, -8, -48, -1, 2, -9, 8, 0, 41, 35, 16, -5, -14, -3, -1, 4, 3, 29, 1, -5, -18, 5, 1, 14, 5, -48, -13, 41, -20, 22, 57, -19, 7, 3, 2, -56, -6, 1, -42, 8, 11, 8, -20, -12, -5, -6, -18, 0, -9, 24, -1, 0, -30, -13, -21, -47, -5, 21, 5, 3, -3, -42, 10, -32, 17, 30, 4, -2, 2, 12, 2, -16, 2, 7, -11, -1, 13, 0, 0, -54, -25, 8, -39, 17, 25, -2, 7, 31, -40, -33, -67, 8, -14, 36, -1, 4, -33, -10, -21, 2, 5, -4, -14, -13, -12, -43, -1, -28, -5, -29, -15, 26, -56, 5, -18, -6, -7, -75, -44, 10, -17, -5, 17, -6, 17, 8, -3, 0, -36, 4, -54, -44, 4, -2, 1, -9, 23, 7, 1, 1, -1, -2, -14, -4, -9, 18, -43, -7, 9, -37, -8, 2, 3, 5, 6, 27, -16, -40, 6, -18, -48, -1, 30, 6, 5, 8, -4, 5, 0, 2, -40, -7, 8, 11, -5, 3, 5, 2, 6, 8, -12, 3, 53, -4, -36, 23, 17, 16, -64, -40, -2, 53, -20, -6, 5, -5, -35, 4, -15, -11, -31, -3, 16, 0, -7, -11, -3, 0, 26, 8, -10, 5, 35, -29, -2, 0, 1, -11, -5, -3, -19, -24, 3, 0, 0, -5, 3, -13, 9, 0, -3, 0, 10, 4, -16, -9, 0, -8, 5, -49, 9, -6, 2, 4, -3, 1, 4, -9, -61, 13, 2, -8, -60, 12, -4, -8, -20, -31, -5, -3, -30, -51, 7, 0, -9, -19, -3, 38, 7, 11, 1, -23, 9, -4, -60, -27, 27, 1, -3, -2, -6, 4, 32, 5, 9, -1, -1, 2, -17, -1, -6, 8,
    -- layer=3 filter=0 channel=2
    -4, -3, 14, -34, -1, -4, 12, 13, 1, -5, -10, 4, 3, 4, -26, 8, -64, -1, -14, 13, 9, 0, 12, -3, -8, 9, -8, -5, -50, -55, 10, 10, -6, -15, -25, -8, -9, -9, -7, 15, -1, -18, 10, 3, -2, -4, 41, 3, 17, 3, -4, 1, 10, 4, -12, -13, -30, -5, 8, -20, -9, 24, 18, 2, -17, -33, -4, 14, -16, 22, -5, -13, -3, -5, -2, -6, 1, 6, 10, 1, 1, 8, 18, -10, 4, 13, 14, 2, -3, -4, -3, -4, -17, -36, 10, -2, 0, 5, -31, -22, 22, 2, -4, -2, 14, 30, -22, 2, -4, -13, -32, -4, -7, -6, 3, -4, 4, 11, -4, 0, 3, -1, -40, -25, 5, 6, -6, -14, -15, -49, -9, -5, -12, 21, -34, 5, -1, 12, 11, 0, -10, -6, 0, 5, 10, 19, 6, 20, 6, 37, 1, -9, -8, -31, -12, -2, -5, -2, -51, 3, -6, 0, 11, 22, -2, -9, -9, 8, -31, -1, 9, -3, -18, 0, -9, 2, 3, -7, 18, -38, -13, -3, -26, -5, -12, -1, -24, -9, -1, -5, -2, -10, 31, -55, -6, 0, -10, 0, -9, -20, -13, 14, 0, -5, 15, 19, -1, -1, -8, -1, -17, -25, -19, 15, 21, -39, 0, 9, 0, 50, 6, -8, 20, -46, -10, -3, 21, -29, 11, -14, 30, 7, 14, -6, 3, 5, 2, -17, -50, 1, 7, 0, 0, -23, -6, 35, -14, -23, -2, 17, 17, -12, -9, -9, 9, -6, 9, -5, -34, -9, 5, 20, 1, -17, -3, -5, -4, 0, -3, -4, -2, 2, 35, 8, 16, 0, -2, -6, 9, -2, -3, 4, 9, 6, -7, -7, -1, -31, -1, 9, 2, -17, 9, 21, -19, -3, 8, -11, -6, 33, 18, -3, -11, -25, 12, -11, -3, 9, 34, 20, 24, 5, 5, -32, -12, 4, -4, -9, 0, 7, -43, -4, 1, -19, -2, -7, 0, 11, 0, 33, -2, -20, 26, 4, 10, -5, -3, -9, -7, -46, 21, 6, 0, 1, 16, -5, 3, -7, -8, 1, -3, 23, -15, 0, 1, 0, 37, -3, 9, 7, 6, 3, 14, 8, 0, 8, -14, 0, -7, 14, 11, -2, -4, -9, 3, 11, 3, 13, -5, 4, -32, 0, -2, 53, 6, -36, 0, -5, 2, -2, 7, 10, 24, -13, -6, -33, -24, 10, -50, 5, 19, 7, 25, -1, -46, 0, 19, 1, -31, -21, -10, -17, 36, 2, -25, 12, -23, -11, 15, -18, -2, 4, 17, 0, 7, -10, 1, -5, -20, 5, 22, -4, -32, -17, -9, 2, 14, -47, -2, -3, 10, -26, -4, -5, 2, -8, 1, 33, -17, -6, -17, -9, -7, -41, 8, -4, -3, 5, 0, -15, 7, -3, -7, -6, -9, 3, -19, 1, 20, -41, -3, 4, -2, 4, 2, 1, 0, 4, -8, -3, 21, 5, 49, -9, -18, -20, 4, -29, 0, -13, -6, -21, 16, -9, -33, 17, -7, -1, 5, -7, -6, 4, -13, 6, 8, 2, -5, 10, -23, 2, -5, -5, -3, -3, 28, -54, -5, -8, -18, -21, 1, 0, -8, 6, 10, 2, -26, -7, -65, -28, 14, -23, 6, 4, 17, 0, -3, -1, -3, 1, -25, -14, -8, -59, -2, 21, -10, 18, -1, 1, -6, -9, 3, 33, 9, 3, -4, 11, 8, -6, 9, -27, 1, -34, -5, -3, -2, -7, 7, 0, -2, 4, -40, 0, 20, -1, -9, 14, 56, -26, -4, 14, -10, 6, -6, -6, 7, -2, -5, -10, -21, 4, 15, 4, 14, 5, -8, -11, 6, 2, 7, -15, 17, 33, -4, -14, -15, 7, -3, 1, 5, 34, 16, 4, -6, -32, -3, 1, 11, 2, 10, 5, 0, -6, -1, -22, 6, 1, -1, 28, 1, 50, 9, 1, 62, 14, -10, -2, 2, -7, 7, 3, 14, 23, -15, -1, -17, 7, 3, 10, -1, -16, -6, 6, 0, -4, 0, 0, -22, 34, -1, 45, 6, 4, -8, -9, -16, 0, 3, -16, -27, 6, 9, 0, -7, -15, -8, -7, -20, -1, 7, -11, -4, 15, -12, 5, -10, 1, 17, -55, 0, -46, -7, -8, -3, 6, -3, -4, 17, 26, -13, -1, -11, 5, -16, -27, -16, 2, -9, -3, -43, 0, 8, -17, 3, 1, -14, -15, -17, 1, 4, 6, 13, 10, 2, -14, -6, -16, -3, 13, -8, -21, -8, -14, -4, 7, 6, -2, 8, 35, 23, -41, -11, 5, -11, 4, 2, -7, -2, 21, -25, -9, -30, -2, -2, -29, 3, -7, -23, -17, 7, 26, -16, -18, 23, 27, 1, -68, 20, -11, 19, -22, -19, -44, -25, -1, 14, 3, 7, -8, 6, -8, -1, 5, 51, 5, -29, 23, 0, 10, 17, -1, -4, 25, 31, 8, -15, 25, -10, -14, -40, 17, -1, 31, 5, -8, 17, 9, 11, -3, -5, -4, 3, -2, -27, 14, 4, -9, 1, -14, -42, 0, -14, -27, -10, 14, -8, 4, 21, 0, 9, 10, 1, 2, 45, 5, -9, -24, 8, -25, -4, -16, -24, -22, -10, 8, -15, -1, -4, 9, 0, -8, 6, 1, 1, 2, -5, -6, -6, 12, 12, -1, 0, 1, -12, 6, 10, 6, 2, -6, -8, -7, 4, 9, 41, -9, 3, 10, 25, 8, -23, -9, -6, 4, 2, 8, -6, -19, 25, 15, -9, 0, 10, 5, 11, -33, -5, 14, -17, 7, 0, 2, -32, 1, 34, 14, 4, 18, 37, 0, -23, 6, -6, 6, -14, -1, -12, -17, 6, -1, 32, -23, -2, -7, -20, -7, -16, 2, -13, 11, 2, -12, 17, -3, -21, -7, -33, -14, -7, 4, 9, 4, 27, 0, 14, 11, -4, 0, 0, 12, 1, 10, 14, -11, -47, -1, 4, -22, 2, 6, -36, -2, -5, -12, 11, -1, -3, 4, -2, -7, 2, -30, 1, -6, -3, -3, 20, 3, -13, 9, 0, -29, 7, -4, -6, 15, -11, -8, -25, -3, -6, -10, -1, -22, 18, -18, 10, -19, 2, -23, 4, -4, -14, -23, 7, -7, 24, -15, -4, 1, -1, -1, 0, -1, 6, -3, 0, 1, -7, 1, 27, 9, -6, -8, 5, -7, 3, 0, -1, 0, -14, -11, 3, -3, 4, -7, -13, -34, -10, 6, 0, -8, 12, -23, -3, 2, -13, -33, -67, -1, -2, -5, -19, -36, 25, -49, -2, -22, -8, 25, -9, 6, -3, 31, -5, -15, 10, -8, 7, 0, 10, -34, 12, 1, 7, -5, 4, 9, 10, -18, -14, -7, -3, -16, -5, 12, -8, -3, 1, -5, 34, 36, -7, 27, -6, -5, -3, -1, 5, 4, 4, 14, -2, 4, 0, 5, -39, -5, 9, 33, 8, -5, 4, -11, -12, -14, -35, -19, 11, 3, 9, 0, 27, -30, 21, -1, 17, 11, -27, -4, -15, 6, -10, 26, 16, -1, -5, -23, 7, 0, 5, -10, -8, 4, 4, 4, -36, 9, 20, 6, 19, -10, 9, 29, 12, -18, 8, 4, -19, -1, 0, 8, -7, -3, 0, -1, -4, -6, 8, 3, 4, -19, 2, 31, -8, -13, 1, 20, -17, 2, -8, 18, 49, -5, 10, -3, 41, -15, 3, -2, 29, -9, 21, 6, -17, -33, -15, 2, 1, 1, 13, 4, 10, -54, -14, 1, 30, -2, -10, -6, -30, -19, -11, -6, -2, 1, -31, 22, -13, -2, -2, -16, 8, 23, -3, -14, -7, -7, 2, 9, -15, 7, 7, 46, -2, -3, -1, 13, 7, -3, 7, -7, 7, -39, -6, 0, 5, -16, 2, -2, -2, -45, 16, -8, -36, 15, 0, -1, 2, 1, 4, 18, 4, 2, 33, 5, -6, -10, -3, 6, -16, 7, 2, 18, 18, 37, 19, -37, 2, -21, -11, 2, -9, -21, 23, 12, -16, 5, -18, -22, -3, -10, 6, -8, 3, -1, 36, -27, 18, -14, 0, -9, -30, 3, 0, -15, -8, -4, -22, -1, 4, -53, -1, 8, 5, -11, 2, 15, 22, 0, 2, -7, -7, 9, -26, -5, 3, -44, -12, 31, -4, 21, -2, -21, 63, 27, 12, 4, 0, 1, 2, 10, 34, -5, -18, 1, 0, -27, 1, 1, 2, 0, -11, -4, 5, -5, -4, 3, 14, -9, -4, -25, -15, -6, -5, 5, 11, -4, 10, 10, 5, -1, -34, -1, 19, 4, -2, 1, 4, 0, 11, 4, -2, 7, 4, -4, 11, -10, 2, -23, 18, 2, 5, 0, 3, 3, 6, -21, -5, -24, 22, -4, 1, -20, 13, -4, 26, -46, 2, -75, 9, 6, -4, 13, 0, 5, -24, -11, -23, 25, 14, -5, -32, 9, 9, 7, 16, 4, -34, 1, -28, 6, 7, -9, 6, -45, 37, -1, -14, 7, -10, -31, -2, 0, 50, -8, -4, 7, -18, -5, 3, -1, 10, 5, 17, 2, -41, 22, -9, -6, -5, 16, -2, -6, 12, -6, -2, -3, -5, -12, 6, 19, -5, -5, -6, -24, 4, -20, -14, -7, 8, 0, 12, -20, 7, 6, -6, 0, 0, -6, -7, 1, -5, -14, 0, 5, -6, 14, 6, -7, 8, 1, 0, -9, 16, 23, 36, 13, -9, 10, -5, 33, 4, 22, 4, -9, 9, 0, 44, -6, 4, 6, -4, -2, -9, 0, -45, -6, 7, 5, -7, 0, -3, -8, 6, -18, 11, 8, 30, -40, 4, -3, 47, -38, 30, 30, -4, -3, -7, -2, -9, -3, 19, 3, -13, -20, -3, 6, -6, 19, 6, 7, 0, 7, -1, -4, 29, -8, 5, -28, 18, -17, -2, 4, 4, 0, 3, 21, 31, -9, -11, -23, 26, -4, 1, 28, 6, -19, -9, 9, -2, -18, 25, -4, -4, -6, -1, -17, -2, 0, -3, 32, -59, 9, -12, 16, -12, -6, -6, -6, 10, -1, 8, -2, 21, -1, 6, 3, -8, -8, 4, 2, 1, 1, 1, -11, -10, 40, 0, -19, -21, 5, 8, 14, -13, 11, -2, -1, -6, 36, 18, 12, 0, -15, -16, -12, 2, -4, -7, 55, 2, -1, -9, -1, -9, 0, -7, -9, 1, -18, -6, -8, 47, 0, -2, 11, -7, 17, 7, 17, -20, -10, 2, 7, 9, -9, 1, -11, -6, 7, 6, -19, -43, 8, -5, -32, -2, 7, -2, -23, 22, -10, -7, -7, 3, -8, -6, -13, 4, -11, -2, -2, 7, 0, -10, 15, -14, 23, 43, -6, 0, -1, -1, -23, 3, -65, 17, -2, 0, 4, 0, 6, 9, 58, -11, -1, -7, 2, 12, 13, 10, -4, 1, -1, -12, 2, 1, 15, 4, -4, -19, 8, 5, -9, -4, -53, -10, -66, 31, -27, -25, -6, 9, 29, 3, -14, -7, -19, 31, 18, -3, 5, 33, 32, -7, 0, 6, 13, 0, 5, -8, -2, 1, 11, 36, 1, 8, 6, -1, -14, -6, -7, -24, 4, 12, -33, 35, -40, 48, -10, -6, -12, 13, 12, 28, 14, 7, -34, 7, 10, -53, 30, -12, -10, -7, 3, -6, 0, -18, 25, 26, -8, 0, 22, 28, -4, -3, -29, -3, 1, 17, -68, -9, 12, 1, -6, 2, -42, 6, 28, 19, -7, -24, -9, 0, 27, 15, -1, 23, 0, -12, -5, -4, 2, 26, 17, -9, 32, 17, 7, -6, 9, 7, -14, -7, 6, 11, 10, -21, -25, -16, -3, 1, 1, 5, -13, 0, -18, 16, -4, -6, 1, 2, -4, 43, 24, 5, -4, 4, -2, -3, 4, 6, 2, 31, 2, 13, -29, -12, -4, 1, 1, 7, 1, 4, -7, 6, 7, 2, 10, -5, 5, -34, -1, -18, -11, -13, -1, -6, 13, 6, 13, 29, 53, 1, 22, -7, 0, -10, 14, 0, 5, -46, 4, -1, 12, -27, 3, 5, -3, -41, -15, 7, -1, 40, 0, 52, -3, 8, 3, 5, -25, -21, -7, 15, 10, -6, -32, 6, 4, 21, 7, 2, -24, -34, 2, 11, -8, 22, -2, 24, -12, -5, 0, -28, 0, 50, -5, -3, -10, 6, -40, 5, 22, -5, -2, -18, -2, 23, -5, 3, 1, 5, 2, -31, 4, -9, -3, -30, 0, 18, 5, -4, 1, 7, 0, -5, -1, -4, -1, -19, -4, 5, -7, 28, -14, 4, -8, 1, -4, 8, 4, 20, -7, 7, -1, 28, -21, -19, 13, -9, -55, 4, 6, -3, 5, 0, -17, 7, 3, 10, -12, 24, 0, 2, -2, -5, -1, -23, -10, 1, 2, 7, -11, -5, 7, 7, -7, 17, 9, -32, -29, 5, 2, -77, -39, -41, -2, -6, -6, 2, 9, -23, 1, 1, 13, 4, 36, 1, -4, 20, 8, 42, 19, -4, -4, 28, -24, -15, -56, -5, -17, 7, 35, 2, 1, 3, -1, -2, -22, -64, -10, 2, -4, -15, 24, -44, -56, -6, -12, -4, 7, 2, -34, -21, -2, 7, 28, -7, 24, 41, -12, -20, 59, 17, 23, 0, 59, -3, -8, -4, 4, -7, -4, 0, 0, -23, 10, -12, -4, -8, 3, 0, 0, 12, -6, -2, -4, -2, 18, -20, 7, -6, 6, 5, -4, 33, -10, -3, 3, -22, -27, 14, 8, 5, -12, 16, -28, -14, -1, -8, -41, -2, -6, 4, 14, -8, 4, 9, -1, 10, -29, 39, -5, -42, 15, -57, -73, -7, 55, 7, -22, -16, -1, -7, -3, 3, -21, 8, 8, -2, -2, 39, 20, -30, -17, 6, 0, -1, 0, 2, -30, -1, -7, 1, 10, -25, 1, -1, -3, 4, 15, -9, -2, -11, 3, 27, -19, -16, 0, 5, 1, 6, -4, -7, 28, -31, -3, -8, -1, -4, -2, -5, -7, -11, 50, -3, -2, 7, 0, -46, -24, -50, -3, -6, -54, -43, -20, -5, -12, 8, -4, -18, 15, -7, 5, 0, 18, 0, -24, 19, -15, 1, -22, -7, -24, 7, -28, 7, -12, -20, 5, 0, -11, -4, -17, -6, -51, -42, 15, 1, 0, -4, -4, 1, -13, -1, -2, -28, 0, 6, -13, 1, -1, -21, 3, 10, -11, 48, -43, 33, 3, -11, -17, 8, 0, 14, 21, 32, -43, -3, -8, -51, -7, -7, -6, 0, 20, 5, 6, -30, 17, -27, -47, 7, 0, -12, 7, 0, -19, 15, 0, -41, -1, -7, -13, 9, 0, 9, -8, -6, -13, -12, 3, 10, -8, -6, -42, -37, -7, -39, -3, 19, 2, -12, 8, -68, 6, -13, 13, -36, 6, -7, 0, -13, 31, 71, 7, -23, -8, -61, -21, -4, -9, -5, 14, 3, -18, -57, 11, -28, -5, 19, -11, -1, -4, 12, -48, -5, -7, 15, -1, 20, -9, -3, 16, -15, -5, 54, -2, -24, 7, 7, 7, 25, 7, 4, -3, 6, 0, -2, 6, 0, -35, 38, 0, 12, -52, 0, 6, 8, -5, 1, 37, 35, -69, -9, -31, 17, 5, -33, 2, -5, 55, -25, 2, 9, -9, 44, -4, 41, 37, -17, -35, 38, -3, -3, -4, -20, 1, -2, -8, -23, -12, -18, -26, 10, -4, -8, -33, -12, 0, -21, -5, -43, 2, -30, 26, -48, 2, 1, 2, 25, -1, 1, 5, -1, -5, 24, 8, 18, 43, 4, 7, -16, 3, -10, -1, -40, 22, -28, 4, 7, -22, -3, -32, 17, 4, -17, -22, 12, -5, 19, 8, 1, 1, 1, -9, -9, 6, 1, 2, 0, -3, -12, 3, -1, -51, -2, 3, -39, 15, 6, 7, 30, -7, -1, -2, -20, -31, -22, -43, -5, -15, 6, 5, 3, 16, -10, -7, 6, 9, 55, -39, 10, 5, 0, -2, 1, 0, 13, -3, -7, 7, -9, -53, -11, -8, 0, 23, 18, -6, -13, 11, -10, 1, -21, -22, 6, -22, -4, -7, -6, -48, 7, -2, -27, 17, 2, 23, -5, -6, 27, -3, 0, -49, 2, -2, 29, -40, 14, -17, -1, -25, -5, -30, -1, -3, -2, -8, 1, 10, 0, 5, -12, -5, 30, 35, 13, 7, -1, -1, 0, 1, -10, 17, 18, -8, 2, 22, -54, 5, 21, -11, 0, -21, 9, -20, -10, 2, 2, 2, -11, 0, -3, -10, 0, 28, -35, 0, 28, -4, -36, -4, -6, 14, 2, -7, -6, -7, -32, -16, 7, 14, -11, -9, 0, -4, 37, -15, 24, -5, -6, 7, -5, 18, 18, 0, -22, 19, -5, -10, -7, 9, 0, -3, -7, 39, 7, 0, 1, -7, -2, -27, -1, 0, 24, 15, -30, -3, 33, 29, -3, -8, -4, -1, -9, -4, 1, -16, -4, 0, -4, -4, 7, -13, 19, -28, 4, 13, -30, -2, -5, 15, -8, 2, -9, -9, -1, 2, -12, -5, 9, 3, 5, -7, -5, 1, -38, -12, 4, -31, 21, 0, -1, -2, -38, -23, -7, -66, 22, 2, -3, -7, -3, 2, 3, -10, 0, 1, -16, 9, 27, 11, 11, 5, -11, 0, 12, -11, -4, -53, 0, -3, -4, 13, -10, 7, -11, -25, -29, 44, -13, 8, -5, -19, 3, -6, 7, 7, -3, -4, -6, 28, -1, -2, 13, 2, -34, 0, -22, 54, 4, 9, -4, -1, 4, 25, 9, 7, 5, -5, -1, -18, -7, -6, -32, 61, 48, -23, -4, 1, 25, 23, 0, 3, 18, 0, 14, 22, -45, -39, 1, -1, -26, -15, -3, -10, -4, -6, -2, -1, 23, -36, 8, -37, 13, -42, -9, 0, -5, 23, 7, 2, -7, -63, -1, -46, 6, 2, -7, -3, 0, -2, -41, 4, 5, -5, -8, -15, -15, -2, -3, -37, 22, 38, 6, 34, 26, 29, 2, -16, 13, 6, 0, -5, -15, 1, 39, 3, -11, -36, -31, -4, 1, 17, 0, 44, -4, -14, 0, 22, 11, -5, 49, 3, 3, -25, 24, 16, 16, 10, -2, -6, 5, -3, -3, 0, 4, -5, -23, 34, -12, -4, 6, 6, 31, -6, 9, 0, -2, -2, -47, -8, -1, -1, 21, -2, 1, 40, -6, -2, 4, -18, 2, -56, -5, 28, 4, -22, 17, -6, 6, 20, 3, 56, 7, 8, 0, -22, 16, 9, 12, 19, 1, -25, 24, -3, -73, 1, -20, 8, 3, 0, -13, 8, 2, -44, -29, 28, -9, -21, -10, -4, 4, 6, -1, 28, 48, 2, -33, 3, -20, 29, 39, -14, 5, 3, 45, 11, 11, 3, 18, 22, 6, 0, -4, -41, 7, -1, 33, 20, -12, 7, 3, 5, 7, 13, 26, -6, -12, 0, 27, 0, 23, 5, -1, -6, -1, -4, 1, 5, 5, -10, -1, 0, -20, 6, -46, -37, -6, -2, 15, 1, -1, 4, -18, -3, 3, -6, -1, 12, -12, 32, -16, -96, 5, -12, 0, -18, 9, 4, 9, -8, 36, 31, 9, 4, -1, 0, -5, 5, -13, -2, 1, 8, -1, -24, 47, -6, -3, 4, 25, 0, -24, 8, 6, -3, 31, -50, 35, 20, 5, -6, 2, 21, 36, -6, -18, 6, 36, -42, 3, 5, -21, -11, 28, -3, -1, -5, -18, -4, 0, -11, 3, 21, 12, -7, -10, 2, 5, -45, -7, -2, 2, 5, 1, -3, 63, -44, 16, 40, 6, 18, 0, 2, 6, 24, -9, 1, -1, 35, -18, 12, -7, -2, 0, -11, 17, -18, -19, -15, -9, -4, 4, -6, -10, 8, 10, -5, -17, 0, -52, -4, -70, -6, 0, 4, -4, -9, 0, -8, -18, -16, 50, -25, 11, 7, 3, 6, -6, 8, -7, -4, -7, -2, 27, 4, -51, 4, 5, 27, 5, 0, 7, 19, 0, -8, -1, 36, 4, 6, 1, 0, -20, -27, 24, 7, 1, -2, 27, -2, -2, 32, 6, 16, -12, 2, 1, 6, 31, -39, 5, -13, -3, 3, -11, 17, 5, 15, -1, 17, -15, -7, -7, 2, 15, 2, -8, -6, -61, 2, 24, 0, 15, 12, 8, -11, -1, 4, 25, -3, 11, 26, 14, -3, 6, 2, -6, -27, -29, -51, -43, -4, 22, -5, -2, 2, 9, 3, 51, 0, 4, -19, -58, -40, 0, 1, 0, 10, -4, 7, -6, 12, -1, -2, 7, 2, 0, 5, -14, 5, -8, 38, 26, -26, -17, 23, -3, -41, -8, 28, 0, -18, 31, -44, 0, -7, 8, 6, 18, 25, -43, -23, 0, -3, 5, -6, 5, -17, 16, 3, 1, -8, -3, 19, 10, 35, 55, -28, 32, -2, -5, -11, -62, -61, -4, -25, 53, 1, 1, -15, 0, 31, 0, 7, -13, 11, -11, -3, 3, 19, 10, 3, 23, 19, 0, 7, -14, 22, -8, -4, 0, 22, 4, -17, 29, -19, -9, -37, 27, 6, 6, 16, 9, -7, 18, 4, -7, -2, -3, 3, -8, -1, 3, 0, -5, 2, -2, -30, 6, 40, 4, -5, -7, 5, -2, 9, 1, 4, -20, -2, -2, 20, -8, 6, -11, 12, 5, -15, -5, 28, 12, -20, -45, 5, -3, -16, -3, 26, -13, -6, 18, 0, 18, -7, 29, 0, 0, 20, -21, 1, -24, -4, -10, -2, -7, 0, 9, 0, -3, -4, -13, 0, 27, 6, -7, -17, -39, -5, 10, 11, -10, -2, 0, -43, -2, -40, 13, -10, -6, -16, 39, -3, 6, 33, 3, 0, 48, -4, -5, 4, 28, -5, 3, -10, -5, -47, -13, -20, 40, 3, 35, -7, 38, -4, -3, -5, -21, -71, 5, 13, 0, -12, 1, 6, 12, 0, 40, -45, -2, -49, -18, 2, -19, 19, 9, -6, 2, -4, -16, -3, 9, -3, 4, -28, 1, -7, 3, -12, -9, 8, 15, 11, 2, -3, 2, -16, -8, -34, -42, -4, -8, -3, -5, 8, 22, 0, -5, -13, 13, -4, 5, -7, -9, 0, 10, 7, -2, 10, -20, -27, -2, 10, 27, 1, -5, -4, -26, 0, 6, 0, 10, 15, -1, 24, 1, -33, 7, 9, 0, 7, -13, -13, 10, -4, -21, 24, -13, -1, 2, -3, 7, 8, 12, 0, 8, 7, 3, -33, -9, -4, 0, -45, -2, -6, -15, -27, 5, 5, -17, 7, -26, -10, 2, 4, -8, -8, 8, -1, -17, -12, 30, 25, 2, 5, -12, 9, 19, 20, -3, -5, 59, 7, -18, -34, 3, 59, -15, 44, 3, 0, -3, -56, -10, -39, -19, -4, -2, -8, -73, 8, 29, -5, -3, -5, 0, 6, -1, 47, -32, 5, -1, -25, -4, 6, 19, -1, 2, -18, 7, 5, -5, -31, 7, -5, 3, -9, -2, 0, -5, -8, -105, -6, -51, -4, -8, 5, -5, -26, 4, -1, 7, -1, -18, 29, -2, -45, 0, -8, -4, 8, -13, 16, -78, 2, 24, 28, -24, 10, -29, 6, -6, 15, -22, 7, -4, 23, -4, -10, -9, 31, -1, -27, 6, 0, -16, -58, 63, -7, 4, 15, 41, 5, -25, 37, -16, -16, 12, 0, 2, -6, -11, -18, 3, -3, 1, 0, -15, -8, 2, -13, -4, -17, -29, -9, -7, 3, -10, -4, -5, 29, 13, 3, 21, 0, 22, -33, -1, 0, 36, -9, 23, 11, -25, 30, 48, -5, -2, -10, 16, 33, -41, -20, 5, 9, -53, -4, -15, 3, 10, 11, 20, -3, -16, -32, 0, 29, 0, -2, -2, -31, -4, 10, -30, 10, 7, 10, 7, 3, 0, -11, -12, 22, -13, 5, 21, -42, 3, -9, -6, 6, 1, 12, 6, -5, 12, -38, -8, 5, 36, -46, 17, 2, 22, -21, -1, 0, 6, -2, 5, -21, 19, 6, 11, -4, -11, 7, 0, 7, -24, -34, -10, 15, -16, -9, -47, -38, -3, -17, -1, 2, 32, 33, -7, 9, -26, 6, -12, 58, -7, -14, 5, -4, 6, -4, -3, -11, 9, -59, 0, -17, 25, -3, -7, -34, -19, 7, -44, -22, 2, -25, 23, -2, 6, 7, -3, -53, 19, -4, 10, -5, -5, 2, -27, 9, 10, -51, 11, 3, 8, -45, -38, 15, 7, -2, 0, 13, 6, 7, 22, -2, 24, -6, -9, 12, 31, 35, -7, 5, -6, -5, -3, 27, 29, -33, -15, 7, -5, -9, -8, -32, 24, -61, -24, -3, 7, -3, 31, 4, -4, 10, -1, -8, -18, -66, -10, 5, 5, -1, 13, -8, -3, -3, -9, -1, 9, -3, -2, -19, -8, 7, 14, -25, -6, -4, 2, 21, 1, -11, -19, -57, 2, 8, 55, 3, -54, -34, 0, 5, -38, 0, 0, 34, -18, 6, 19, -7, -19, 11, 10, -2, 16, 20, -40, -4, 35, -11, 3, 6, -34, -43, -23, -18, -8, 19, 0, 3, 29, 7, 14, -6, 21, -21, -21, 3, 9, -39, 25, -8, 1, 0, -30, 8, 39, 8, 8, 10, 1, 9, 11, 18, -1, -1, 9, -17, 40, -7, 0, 4, -7, -36, 22, -7, -6, -11, -11, -5, 9, 7, -11, -3, 7, -11, -4, -3, 2, 0, -9, -3, 18, -3, -41, 13, -3, 3, 28, 0, 1, -1, -41, 33, 0, 8, -29, -4, 0, 10, 11, -58, -1, -1, 2, -12, -5, -25, 1, 2, 37, -60, 21, 0, 0, 4, -9, -3, -46, -7, 2, -3, 0, 14, -16, -4, 3, 12, 0, -6, 16, 28, -3, 0, 17, -5, 12, 27, -11, 7, -8, 0, 45, -6, -56, 4, -53, -49, 4, 6, 9, -12, 28, -18, -10, 3, -26, 12, -39, -35, -7, 3, -58, -48, 0, -1, 8, -42, 2, 7, -14, -2, 5, -3, -45, -11, 3, -5, 0, 22, 4, 0, -24, 21, -22, 7, -1, -13, -14, 38, -9, 4, -1, -5, 8, 37, 6, 8, -4, -7, -9, 8, 6, -5, -2, 4, -41, -8, 65, -5, -45, -2, -3, 3, 8, 2, 0, -5, 36, -24, 7, -42, 5, 1, -3, 0, 0, 10, 6, -5, -10, 10, -12, -10, -30, 5, -15, 18, -15, -5, -4, 23, 0, 0, -3, 44, 4, 29, -7, -5, -33, -54, -17, -9, 37, -1, 11, 14, 4, 5, 0, -39, -37, 12, 7, -6, -28, -21, -4, 6, -2, 0, -39, 6, 15, 39, 4, -9, -3, -7, -1, 22, -15, 0, -6, 17, -22, 7, 3, 6, 3, 10, -7, 8, 11, -10, 19, -7, -3, 27, 24, 3, -4, -14, -65, 44, -64, -33, -48, 8, 7, -8, 3, -2, 0, 5, -8, -4, -10, -15, -5, 4, 10, -3, -9, 13, 15, 25, -9, -37, 4, -1, -21, -9, 2, 0, 3, 42, -14, -37, 12, -11, -13, 19, -1, 32, 2, 1, 0, -2, -9, -29, 10, -14, -2, -36, 0, 19, -13, 18, 9, -7, -1, 2, 5, 0, 25, 5, 11, -2, 0, 0, -5, 4, 25, -1, 17, -2, -9, 19, 14, -54, -3, 3, 6, 2, 33, 28, 48, 32, -26, -13, -6, 31, -11, 2, -1, -13, 4, -9, 40, 0, 15, -8, 14, -3, 44, -5, -13, 36, 7, -39, 8, -46, 6, 11, -14, -6, 2, -1, -6, -3, 2, -6, 11, -13, -1, 15, 1, 5, 56, 60, -19, -7, 6, 19, -8, 5, 14, -35, 8, -16, 0, 5, -3, 11, 22, -7, 0, -8, -17, -49, 4, -10, 6, -6, 3, 0, 25, -8, 11, -9, 46, -4, 0, -30, 41, 30, -32, 5, 6, 7, -15, 0, -7, 3, -17, 5, -30, -11, -7, 1, 5, 2, 10, 4, 0, -5, 0, 9, -11, 2, -4, -19, 2, -6, 0, 33, -10, -8, -8, -4, 7, -43, -4, 1, -10, 7, 19, 0, -22, 17, -3, -38, -5, 3, -7, -3, -5, -6, -19, -16, 5, 23, 14, 7, 20, 11, 26, 3, -31, 17, 65, -5, -46, -13, -7, -24, -9, -51, -37, 0, 2, -7, 5, 42, 3, -19, -23, -6, -2, 31, -31, -12, -4, -2, 16, -5, 31, 6, -33, 15, 1, 17, -41, 9, -7, -4, 1, -25, 10, 10, -8, -8, -3, -51, 34, 3, -9, 4, 11, -24, -4, 0, -2, 12, 9, -15, 6, 0, 4, -2, 12, 0, 5, -10, 4, -35, -10, 5, -17, 15, -5, -1, 11, 9, 5, 4, -14, 11, -13, 24, -7, -13, 0, 16, 5, -49, -16, 47, 1, 10, 27, 46, 43, 3, 10, -3, -3, 1, -50, -6, 3, 9, -5, -10, 35, 3, -1, 13,
    -- layer=3 filter=0 channel=3
    19, -8, -22, 1, -3, -5, -38, 13, 12, 29, 7, 8, -8, 3, -12, -6, -2, 29, -2, 0, -5, -8, 24, -9, -18, -32, 3, -3, 50, -10, 8, -24, 2, -6, 34, 21, -6, -13, 6, -29, 7, 27, -39, 7, 0, 1, -10, 15, -11, -11, 0, 1, -3, 5, 34, 7, -8, 5, 3, -30, 6, 12, -19, 0, 4, 15, 12, -40, 8, 18, 2, 3, 0, -2, 3, 7, 4, -21, -41, -2, 17, -4, -11, 0, 6, -8, 19, -3, 11, 0, -15, -9, -11, 32, -8, 3, -4, -2, 14, -20, 24, -3, -4, -25, -7, -40, 12, -9, 26, -17, 8, 0, 1, -7, -4, -7, -2, 13, -17, 12, 0, 1, 32, -17, 12, 9, 0, 17, -12, -11, 5, 0, 4, -24, 2, -4, 5, 2, -12, -3, 5, 3, 2, -2, 29, -7, -55, -14, -5, -31, 4, 10, -4, -5, -16, 4, -3, -9, -15, -8, 16, -7, 10, 5, -2, 0, 37, -4, -14, -9, 3, 15, 18, -3, -4, -8, -18, -2, -23, -32, 3, 9, 37, 7, -8, 5, -6, 25, -8, -4, -4, -2, 4, 10, -10, 6, 14, 29, 0, -5, -21, 8, -4, 4, -18, 14, -20, -5, 13, -9, -5, 3, -28, -19, 5, -6, -2, 42, -3, 8, -5, 8, -4, 23, -16, 1, 2, 17, -37, -30, -23, -23, -7, -5, -5, 0, 5, 27, 58, 10, 0, -6, 4, 10, 6, -11, -41, 0, -6, -24, 11, -2, 1, 12, 3, 3, -42, -6, 5, 22, -15, -24, -6, 12, 12, 13, -4, -4, 9, -46, -10, 8, 1, -42, 0, -32, -3, 2, 38, -7, -8, -15, 14, 18, -27, -38, 5, 0, 5, -11, -3, -28, 0, -5, -6, -2, -7, 2, -7, -11, 9, -2, -11, 21, 28, -3, -6, 25, 36, -10, -40, 19, -27, 5, -1, 0, -9, -1, 13, -5, 11, -9, 23, 6, -8, -30, 6, 25, -3, 12, -16, 18, 8, 4, -41, -2, -4, -14, -26, 0, -4, 10, -7, -9, 29, 6, -3, 3, -18, 5, 9, 14, 5, 2, -3, 4, 5, 7, -4, 4, 2, 5, 1, -1, -7, -36, -45, -3, -3, 22, 10, 4, 4, -43, 2, 18, 16, 9, -5, 2, -19, -4, -13, -9, -6, -16, -6, -5, 4, 0, 37, -8, -4, 16, 1, 24, -17, 3, 18, -3, -3, -2, -29, -3, -31, 5, -2, 25, 39, -20, 6, 24, -20, 0, -2, 9, -14, 23, 17, -33, -20, -2, 2, 41, 12, 2, 9, -9, 0, -4, 15, 5, -13, 17, 5, 4, 14, 24, -6, 0, -7, 12, -1, -1, 0, -17, -4, 2, 8, -9, 5, -21, 2, 5, 2, 5, -2, 8, -5, -1, 10, 5, -3, -1, -4, -2, 18, -1, -35, 11, -3, -6, -45, 17, -7, 2, 10, 21, -10, 0, 3, 3, 21, 7, -11, -29, 8, -8, 1, -11, -15, -29, -6, -5, 39, -8, -24, -9, 3, -2, -1, -1, 10, 6, -9, 4, -1, 11, -27, -3, 1, 26, 14, -6, -11, 29, -1, 2, 21, -3, -23, 0, 7, -7, -3, 2, 9, -6, 2, 23, 11, 0, 7, -4, -6, 26, -59, 1, -7, 3, 33, 17, 18, -26, 5, 18, -3, 18, 9, -3, 6, 12, -1, -9, 37, -3, 10, -3, -8, 24, -15, 17, -10, -17, 2, 7, -56, -15, -17, 2, -2, -24, -19, 3, 10, -3, -4, -3, 2, 12, -6, 5, -4, 9, 6, -4, 0, 0, -3, -33, 49, 4, -3, -3, 16, -5, 7, 14, -7, 1, -11, -5, -24, 22, 11, 28, -18, 4, 4, -11, -9, -25, 9, 2, 19, -57, -55, 46, 15, -2, -40, -13, 26, 12, 7, -45, 3, -10, -5, 2, 0, -4, -2, 5, 32, -12, 58, -5, -41, 2, 11, -22, 3, -48, 12, 0, 0, 9, 6, 0, -14, 41, -6, 0, -8, -5, 11, 12, -30, -9, -9, -46, 7, -5, 3, 9, 17, -1, 0, 15, 11, 3, 12, 0, 16, -20, 2, 6, -7, 9, -30, -23, 0, -39, 19, 0, -9, 8, -8, 11, -10, 1, 7, 5, 22, -1, -1, 5, -13, 1, 16, 1, 12, 22, 31, -26, 0, -3, -1, -30, 47, 1, -22, 26, 3, -7, -43, -5, 3, -4, 1, -20, -3, 15, -24, -57, 20, 24, 1, 29, 5, 26, -1, 3, 3, -29, 6, -12, 0, 39, -37, -3, -5, 6, -3, -11, 0, -1, -1, 0, -2, -8, 0, 1, -7, -11, -4, -6, -11, 17, -34, -19, -16, -4, 7, -17, 1, 31, 11, -1, 0, 23, 23, 13, -16, 10, -22, 12, -7, -4, 2, -11, -4, 9, 16, -5, 15, -13, -6, -32, -19, -3, 4, 12, -48, 35, 21, -7, -4, 32, 42, 7, -6, -1, 2, -15, 21, -7, 40, -17, 3, 0, -5, 4, 9, -52, 17, -22, 6, -1, -28, -17, 0, 19, 23, 3, 3, 6, -28, 33, 14, 8, 10, 14, -40, 17, 3, 16, 7, -9, -5, -19, -14, -20, 16, 3, -23, -5, 0, 12, -19, -18, 9, -2, 8, 1, 1, -5, 8, -7, -16, 3, 36, 10, 1, -9, 3, 1, 10, -3, 5, 5, 0, -1, -3, 5, 7, -20, 34, -2, 0, -2, -8, 12, 4, 13, -4, 10, -12, 2, 2, 28, -1, -4, -13, 0, 0, -9, 13, 6, 3, 12, 3, 3, 13, -12, -14, -42, -40, 1, -16, 10, -94, 6, 3, 11, -6, 4, -9, -8, 35, -3, 3, 35, -16, -3, 13, -11, -33, 25, 13, -12, 9, 1, 36, -28, 25, -12, 1, -5, -17, -6, 29, 6, 7, 19, 3, -4, 18, 10, 0, -1, -16, 22, 13, -5, 9, -6, -7, -62, 19, -14, -4, -10, 4, 1, -32, 9, 0, 3, 4, -28, 4, -6, -5, 2, -5, 0, 19, 5, -30, -1, 8, -2, 12, -13, 0, 5, 24, -1, 1, -6, -31, 11, 34, 32, -9, 0, 5, 0, 5, 6, -42, -20, 9, 1, -17, 10, -22, 2, 0, -7, -5, -9, -18, -6, -8, -6, 1, 22, -4, -5, 8, -21, -33, -5, -4, 58, 7, 2, 14, -1, -7, -25, -7, 4, 4, 12, -20, 4, -5, -33, -9, -38, -7, 3, -20, -39, 47, -4, 6, 8, 45, -14, 26, 7, 1, -3, -23, 16, -1, -12, 6, -28, -6, -1, -31, 7, -6, 8, -56, -5, -1, 14, 3, -8, -4, -4, -13, 12, -17, 0, -5, -47, 30, -21, 26, 0, 7, 65, 1, -8, -10, 4, 8, -6, -1, 5, 5, -3, -3, 0, -32, -4, -18, 6, 13, 0, 0, -26, -10, -2, 2, -4, 4, 23, -26, -39, -42, 0, -7, 6, -59, -11, 1, 5, 11, -9, 1, 14, 13, -7, -12, -6, 5, 9, 7, 7, 7, -8, 6, -14, 1, 25, 0, 1, 19, -18, 10, 8, -19, 7, 23, 17, 21, -58, -13, 31, 1, -1, -1, 0, 7, 0, 0, 4, -15, -4, 26, -24, -24, 26, 0, -14, 13, 6, 2, -24, 11, -8, -3, 10, 2, -5, 1, 3, 6, -26, -5, -6, 8, -3, -46, -48, 13, -8, -10, -3, -2, 8, -43, 18, 17, 7, -40, 5, 46, 4, -12, -7, 22, -17, -26, -8, -20, 13, 31, 37, -11, -4, 2, -34, 8, -10, 2, 3, -4, 1, -12, 0, -4, 7, 0, -6, 13, 3, 27, -59, 10, 1, 9, 0, -4, 7, 4, 2, 19, -18, -9, -12, -4, 43, 10, -6, -28, 27, -9, -6, 9, 3, 5, 13, -29, -2, -26, 1, 1, -38, 8, -5, 8, 24, -25, -38, -40, -2, 37, -17, -3, -17, 28, -8, 24, 0, 4, 1, -12, 20, 2, -11, 9, 0, -5, -36, -8, -1, 3, 21, -7, -4, -2, -8, 2, -3, 8, -3, -31, 39, 4, -28, -5, -14, -23, -13, -3, 44, -4, -21, -20, 3, -29, 0, 2, 9, 9, 1, 8, 15, 18, -1, 10, 22, -18, 1, -38, -26, 3, 4, -12, 11, -21, 33, 12, 1, 2, 32, -11, 15, -12, 8, -5, 12, 0, 2, 15, 14, 7, -2, -33, -3, -1, -29, -3, -17, -20, 9, 0, -3, 3, 0, 9, -11, -7, -5, -15, -23, 5, -6, 5, -2, -48, -6, 3, 2, 6, 2, -2, 8, 3, 14, 9, 3, -6, -45, -11, 2, -2, 2, -5, 14, 34, 36, -8, 32, -21, -8, 8, 16, 0, -24, -18, -5, 5, -19, 14, -10, -20, -20, -3, 16, 8, 9, 42, 0, -29, 0, -23, -2, 28, 12, 13, 9, 31, -37, -1, -22, -20, -6, -4, 0, -14, 0, 23, -5, -5, -4, 8, -29, 16, -3, 6, -9, 0, -5, 13, 4, 0, 29, 5, 40, 21, -35, 5, 4, -53, -27, 16, 1, 0, -2, -10, 4, 45, 7, 3, 9, 13, 39, 19, -1, -6, -4, -2, 29, 0, 0, 2, -1, -3, 2, -26, 0, -8, 30, 5, 7, -25, 0, -7, -9, -13, -1, -1, -3, 20, -6, 50, -18, -16, -39, 2, 19, 2, -1, 7, -10, 15, -9, -6, 8, 12, 4, -9, 5, 5, 0, -11, 6, -2, -5, -2, -9, 4, 0, -3, 1, 24, -6, 32, -21, -2, 6, 19, -5, -14, -65, -1, -2, 7, -27, -21, 5, 0, -6, 12, 34, 6, -8, 35, -13, -14, -8, -5, -2, 9, -17, -1, 57, -5, 30, -32, -11, 1, -4, 1, 11, 7, -4, -64, 0, -9, 6, -15, 13, 19, -51, -4, 14, -1, -1, -21, -9, -6, -4, 8, -18, -28, 32, 35, 9, 14, -13, 8, 1, -13, 6, -10, -1, -6, 0, -2, -2, 1, 17, -9, 6, -28, -4, 26, 1, -6, 13, 6, -4, -13, -6, 21, 23, 2, -5, 8, 5, -1, -1, -13, -18, -5, 8, 1, 8, -6, 56, 0, 4, 24, 20, 3, 0, 7, -17, -7, 5, 9, -16, 8, -42, -5, -9, 6, -12, -10, -6, -18, 11, 22, -14, 43, -16, -5, -4, -3, 0, -5, -7, -6, 7, 0, -4, 3, -4, 8, 36, -12, 18, -6, 14, 0, 8, -8, -32, -6, -9, -8, -13, -35, 4, 4, 0, 5, -11, 6, 5, -9, 4, -4, -5, 6, -15, 9, -6, 5, -3, 22, 18, -14, 21, 3, -9, -17, 7, -16, 2, -7, -21, -38, -4, 4, 4, 24, 45, 11, -6, 8, -25, -40, -38, -1, -26, 1, 0, -7, -12, 7, -5, 14, -10, -27, 13, 4, -17, 2, 18, -1, 14, -4, -3, 6, 5, -1, -44, 2, 2, -34, -38, 3, -27, -12, -10, -13, -8, 4, 3, 0, -5, 7, -6, 22, -3, 0, 20, 4, -10, 24, 28, -11, 31, 3, 10, -17, -4, 4, -10, -24, -20, 6, -7, -7, 6, -35, 14, -12, 15, -3, 0, 4, -38, -6, 4, -2, -21, -23, 24, -7, -7, -21, -5, -8, -3, 8, 0, -18, -30, 7, -12, -4, 14, 2, 1, 10, -35, 8, 6, -4, -4, -5, 17, 3, 0, 17, -33, -9, -60, 0, -2, 15, 1, 52, -4, 8, -2, -18, 0, 15, -1, 22, 2, -27, 5, -19, -29, -17, -18, -3, -50, 6, 2, -40, -24, -3, 7, 12, 5, 0, 37, -48, -55, 11, -3, 0, -1, -1, -3, 2, 3, -14, 8, 7, 2, 0, -2, -6, 4, 0, 0, -9, 5, 0, -5, -44, -5, 4, 35, 22, 9, 1, -58, -2, -5, 1, -15, 2, -17, 1, 21, -2, -14, 13, -5, 2, 1, -10, 37, 1, 2, -1, 2, 18, -2, -27, -15, -55, -3, 17, 0, -1, -3, -5, -3, 13, -3, 36, 4, 9, 3, -32, -5, 0, 2, -6, -2, -1, 1, 0, 11, 48, -42, 14, -2, 18, -7, 30, -22, 9, 0, 22, 6, -24, -2, -27, -2, 0, -1, -2, 1, 8, 6, 63, 5, 2, 1, 3, -14, 0, -13, -8, 10, -2, -4, 7, 28, -14, 4, 4, 0, 0, -29, 2, -7, -2, 0, 11, 11, 19, 8, -28, 15, -3, 0, 22, 4, -13, 3, -21, 13, -2, 0, 23, 7, 3, 15, 1, -26, 0, 11, 10, -4, 9, 9, 11, -1, 7, 10, 25, -6, 2, -3, 2, 5, 14, 7, -3, 0, 7, -24, -16, 5, 3, -42, -15, -2, 11, -16, 0, 7, -4, 23, 65, 43, 9, 1, 4, 17, -7, 3, -9, -33, -7, 17, 5, -4, 6, -26, 23, -13, 3, -1, 0, 17, -11, -53, -5, 8, -26, 0, 4, 8, 0, 31, 4, -10, 10, -5, -2, -12, -37, -42, 15, 3, -5, 13, -4, -2, 4, -6, -23, -9, -7, 27, 30, 38, -16, 6, 2, -23, -15, 27, 3, -10, -2, 4, 0, 3, 0, 11, -9, -1, 54, 3, 43, -7, 1, 0, -1, -24, -18, -9, 2, 0, -60, 14, 11, -9, 31, 4, 4, 0, -18, -18, -6, -6, -23, 2, 34, -14, -17, 0, 26, 10, 15, 4, -9, 8, 0, -1, -5, 43, -1, -23, -1, 3, 21, 5, 27, -6, -17, 11, -25, 20, 4, -42, -11, 22, 14, -17, -1, 0, 8, -17, 7, 9, 5, 0, -48, 54, 32, 21, 1, -4, -16, 2, -5, -60, 9, -5, 13, -14, -21, 7, -30, -4, 10, 29, 0, 6, -18, 1, -14, -3, 24, -15, -3, 7, -2, -4, 13, 17, 21, -11, -33, -5, -46, -1, -18, -9, 16, 1, -33, -9, -2, -11, -8, 30, -24, -10, -2, 0, -102, 5, -8, 26, 5, 1, -76, 14, -6, 9, 3, 30, -28, -18, -2, -37, 8, 20, 0, -26, 2, 28, 0, 2, 29, -81, 0, -4, -47, 8, -35, 30, 20, 11, -11, 3, 9, 5, 6, 26, 33, 5, -1, 0, -1, 10, 1, 45, -32, -7, -29, -24, 23, 16, -28, 3, 0, -20, 37, -15, -21, -18, -5, 13, -1, 11, -5, 12, 3, -2, 7, -49, 7, 6, 51, -13, -34, -1, 1, -27, 15, -3, -1, -61, -26, -8, 23, 0, 3, 17, 35, 3, 0, -42, -7, -31, 9, 4, -21, -3, -3, 3, 48, 0, 18, 19, 1, 3, -4, -6, 17, 4, 5, 12, -3, -7, -4, 4, -21, -7, 17, 8, 2, -15, 43, 38, -17, 12, 8, 7, -4, 18, 8, 13, -4, -2, -20, 2, 6, 43, -39, -19, 2, 0, -10, -5, 3, -9, -4, 3, 11, -10, -14, 8, -8, 6, 3, 5, 20, -1, 2, 4, -3, 2, 10, 6, -2, 7, 32, -1, 0, -14, 6, -5, 0, 10, 7, -17, -12, 7, 10, 11, -8, 6, 6, 31, 1, -13, -6, -2, -3, 6, -32, 3, -9, -37, 3, -3, -14, -10, 38, 10, -4, 0, 23, -9, 19, -2, 34, 15, -19, 61, -4, 0, 5, 4, 28, -6, -2, -17, 20, -15, -16, 7, -3, -3, 39, -1, -1, -2, 7, 1, 5, 9, -39, -87, -1, -31, 0, 10, 1, -3, 12, -8, 10, 2, -7, -7, 5, 3, 38, -1, -11, 0, 0, -12, 8, 1, 6, -4, -2, 31, 3, 9, -2, 7, 4, 5, 11, -4, -12, -27, -4, 9, 12, -11, 4, 2, -10, 1, 7, 0, -20, 35, -16, 11, -15, -40, -1, -3, 5, -46, -9, 30, 0, 2, -2, 4, 1, -4, 0, -5, -2, 0, -6, 0, -5, 8, -5, 40, -15, -6, -8, 6, 22, -7, 3, -10, 0, -4, 15, -13, -20, 13, 8, -2, -2, 40, -25, 6, 15, 28, 0, -24, -1, 5, -4, -19, -8, 36, 0, 8, 7, -18, -18, 12, 9, -9, -16, 12, -4, 7, 8, 0, 3, -21, -3, 2, -17, 0, 43, -30, 5, -35, 4, -11, -7, -2, 20, 0, -1, -4, -3, 9, 4, 24, 1, -4, 12, 10, -42, 35, -5, 12, -5, 3, -11, 0, -8, 4, -4, 44, 39, 0, -3, -5, -1, 3, 7, 30, -6, 11, 5, 3, 8, 34, -21, 13, 2, -4, 2, -4, -13, 30, -46, 13, -21, 8, -10, 21, -19, -10, -4, -25, 0, 7, -3, 9, -4, -3, 1, 5, -1, 20, 4, -9, -10, 2, 19, 4, -3, -14, 0, -11, 7, -11, 4, 7, -9, -6, -7, -3, 13, 24, -5, -4, -4, 0, -4, 8, 3, -3, 5, -3, 14, -2, 0, -44, 10, 3, 8, -18, -10, 0, -8, -10, -11, 5, 0, 3, -13, 7, 5, -12, 2, -39, -10, 7, 5, 0, 10, 2, 18, -15, 14, 3, 23, 0, -2, 8, 3, -30, 10, -3, 8, 23, 6, 25, -34, -4, 6, -7, -79, 28, -9, 1, 0, -8, 12, -15, -12, 0, 8, 30, 25, 7, 32, -31, -8, 25, -5, 12, -1, -13, 18, -8, 6, -31, 3, -19, -4, -17, 19, -26, 0, -8, -2, -6, 7, 1, -4, 20, 14, 9, -89, -2, 6, -47, -5, 20, 29, -38, -2, 9, 17, 24, -13, -26, 6, 0, 0, -14, 17, 19, -11, 11, -30, -5, 42, 20, -8, -4, 6, 2, -9, 3, 28, 42, 27, -5, -1, -60, 13, -9, -4, -16, -1, 0, -9, -7, 9, 7, -24, -21, 0, 10, -8, -15, 23, 2, 5, 0, 3, -8, 25, 4, 1, 20, 4, -21, 0, -3, -2, -25, -30, -2, 5, 14, 15, 5, -12, 11, 0, 4, -14, 9, 2, 39, -19, 32, 0, 18, 1, 8, 8, -40, -16, -2, -7, -2, -6, -12, -34, -59, 6, -7, -11, -6, 5, 6, -3, 1, 5, 11, 24, -15, 7, 7, 0, -9, 15, -2, 8, -1, -2, -5, 25, 0, -4, -50, -18, 5, 1, -14, 3, 3, -6, -14, -6, 23, 13, 25, 6, 5, 26, -8, 10, -2, 4, -8, -15, 2, 9, -3, 7, 6, -9, -6, -5, -3, 19, 12, 17, 10, -3, 1, -25, 8, -9, -16, -8, 5, 18, 23, 6, -31, -19, -2, -2, -6, 3, -16, 29, -2, -18, 7, -7, -15, -16, 3, 2, -7, 10, 3, -11, -4, -41, 3, -7, 11, 5, 8, 2, 5, -2, 15, -17, -3, 6, 12, -4, 10, 25, 7, -3, -1, 23, 0, 4, -1, -9, -6, 7, -18, 4, 3, -2, 7, 6, -7, 2, -6, 24, -23, -2, 2, 4, -11, 0, 5, 20, 27, 3, 6, -8, 26, -32, -3, 27, -43, -8, -27, 0, -14, 4, 1, 13, 7, 18, -6, -10, -3, -6, 5, -6, -2, 17, 7, 7, -4, 5, 21, -14, 8, 9, 16, 0, 5, 11, 8, -8, -3, -22, -11, -14, -13, -7, -7, -8, 13, 22, -1, -3, 5, 0, -17, -4, 0, 12, -1, -30, -8, 6, -6, -22, 9, 7, -16, -9, 13, -11, 15, -5, 3, -6, -2, 3, 27, -10, 6, -6, -10, -27, 58, -7, -8, 6, 46, 1, 5, 14, 43, 37, -8, -8, -30, -19, -33, 0, 7, 7, 15, -40, -20, -9, 20, 0, 0, 7, 5, 0, -4, -6, -11, -15, -2, -22, -2, 36, -3, -5, -11, -5, 5, 14, -1, 9, -17, -9, 43, 46, -7, 7, 4, 19, 31, 31, 9, -19, 0, 25, 26, 4, -7, -1, 23, 8, 1, -8, 6, -1, -2, 0, -44, -11, 4, 0, 4, -37, -26, -7, 4, -10, -4, -11, 22, 12, -7, 0, -17, 6, -4, -1, 3, 3, 20, 0, 6, 2, 1, -9, 0, -1, 15, -4, 25, 8, 12, 2, 9, -14, -3, -12, 12, -14, 7, 31, -3, 36, 38, 5, -8, 16, 6, 47, -28, 12, -16, -36, 0, 8, 7, 6, 27, -36, -26, -1, -12, 0, -5, 0, -2, -8, 32, -18, -5, -7, -26, -8, -7, -1, 3, 4, 15, -27, -4, -9, -6, -1, 5, -2, -10, 1, -5, 5, -7, -25, -6, -28, 13, 17, 2, -7, 8, -3, 11, 3, 0, -15, -2, -4, 2, 14, 14, 22, -18, -12, 33, 0, -3, 2, -5, 0, 13, 5, 10, -14, -5, 6, -28, 3, 0, 4, 18, 12, 3, 25, -29, 0, -17, -10, 26, -6, -12, 14, 28, -32, 25, -40, 0, -17, -2, 1, 4, -1, -8, -2, 1, 17, -36, -25, -15, 7, 26, 0, -7, -3, -48, -2, 9, -12, 8, 2, -25, -12, 8, 10, -11, -9, 2, 2, 0, -4, -11, -5, -41, -32, 9, -16, -28, -2, 11, 5, 8, -10, 27, -6, -13, -11, 2, 2, -8, 50, 11, 24, 3, 4, -11, -21, 12, -9, -18, 6, 7, -11, 33, 33, 24, -5, 0, -73, 4, 2, -44, 27, 23, -11, 4, -32, -8, 25, 8, -3, 0, 34, 0, -13, -9, 8, -2, -4, -6, -13, 6, -1, -10, 0, -7, 19, -3, -9, 41, 12, -1, 12, -1, -1, 5, -3, 35, 2, -21, -10, -21, 7, -5, -6, -10, 5, 9, 0, 2, 0, 2, 1, 7, -30, 0, -22, -4, 21, 12, 17, 9, 10, 0, -68, 0, 7, 6, -38, -23, -36, -21, -18, -13, 0, 33, 1, 1, 28, -2, 10, 9, -20, -2, -5, -3, -26, -26, -35, 16, -2, 0, -8, 3, -2, 3, 32, -19, 4, -11, 15, -10, 9, 6, -16, -5, -16, 8, -2, -9, -6, -5, 2, 4, -3, -30, 0, -3, -22, 1, -11, 2, -11, -33, 0, -9, 5, -1, -13, 2, 0, -8, 23, 2, 2, 9, 30, -19, -4, -7, -24, 1, -4, -9, -15, 28, -42, -24, 2, -36, -6, 30, 3, -21, 6, 0, -10, 0, 42, 11, 0, 4, 8, 2, 9, -6, -10, -8, -5, 1, -3, -6, -36, 4, -4, 9, -15, 3, 1, -16, 1, 3, 0, -7, 0, -3, -4, -1, -11, -4, 1, 5, 34, 3, 25, 27, 2, 3, 4, 5, -26, -43, -5, -3, -34, -2, -44, -32, 0, -27, 2, -8, 7, -5, 0, 41, -2, -19, -1, -1, -10, -4, -9, -11, 32, 0, 6, 54, 3, -4, 18, 13, 19, -9, 0, -17, 7, -11, -14, -2, 0, 14, 22, 13, -11, -36, -2, -1, 3, 2, 8, 8, -8, -27, 45, 5, 40, -2, -3, 1, 3, 20, -5, 7, -1, -12, -53, 15, -19, 5, 26, -5, -2, 2, -21, 14, 21, -3, 24, -23, 9, -19, 5, -9, 15, 2, 7, 1, 2, 24, -3, 0, 3, 2, 0, 5, 6, -9, 10, 9, -19, 5, -4, 12, -49, 13, 27, -20, -5, -1, -4, 3, -4, -3, -29, -10, -6, -10, 1, -6, 9, 33, 22, 0, 4, -4, -17, -3, 0, -11, 23, -1, 7, -20, 0, -7, 22, 6, 16, 14, 3, 6, -23, -4, -65, -12, 9, -24, 3, 6, 2, 5, -18, -18, -6, 9, -35, -15, -1, 1, -10, -4, -5, 14, 0, 3, 5, 14, 11, 60, 14, -2, -11, -7, -6, -4, 13, -2, -4, 9, -3, -9, 2, 3, -5, -29, 15, -41, -8, 36, -7, 8, -4, -21, 3, -59, -17, -4, 14, -17, 0, -10, -15, 35, 29, -27, -5, -15, 1, 0, 3, 5, 10, 14, 8, -6, 5, 2, -7, 10, 3, 5, -5, 29, 19, -24, -5, -1, -28, -32, 6, -14, 20, -3, -11, -13, -8, 38, -19, -18, -84, -29, 3, -5, 5, -18, 0, 3, 23, 11, -25, 30, -16, -9, 0, 3, -2, 40, -29, 4, 18, -25, -4, -36, -14, -2, -2, 13, -4, -3, 4, -1, -1, -2, 8, 3, 26, 8, -34, 18, -11, 46, 8, 29, 1, 17, -18, -9, -20, -3, -6, 6, -27, -32, -1, 2, 5, -9, -31, 33, -26, -25, 0, -20, 5, 0, 15, -18, 0, 3, -44, -5, 6, -5, 3, 0, 13, -5, 0, -11, -43, 6, -3, 9, 12, -1, 0, 13, -4, 5, 4, 7, -30, 6, 5, -5, -9, 3, -14, 6, -9, -14, 11, 2, -11, 32, -9, 10, 1, -13, 7, -14, 7, -64, 11, 30, -16, 0, 0, 8, -11, -49, 28, 0, 5, 0, 2, -7, 5, 22, -14, 19, -22, -13, 6, 7, 6, -2, -18, -3, 10, -14, 7, 21, 6, 1, -1, -4, -4, -5, 25, -2, -10, -9, 21, 11, -34, -6, -37, -36, 0, -1, 1, -1, 9, 0, 17, -4, 7, -2, -4, -11, -10, -3, 0, -4, 1, 0, -26, 10, 5, -21, 7, -19, -34, 4, 15, 3, -11, -15, 17, 0, 2, -4, 3, -8, -7, -2, -1, 0, 3, 7, -7, 2, 3, -48, -2, -1, -25, 7, 3, -6, -20, -2, 7, 1, -4, 3, -63, -27, -4, -34, 1, -8, -8, 11, 0, 29, 1, 7, 7, 33, 23, 0, 0, 6, 0, 5, 2, -6, -4, 1, -8, 3, -13, 5, 0, -8, -12, 8, 6, -29, 0, 0, 20, 8, 22, -35, 4, 4, -3, 11, 12, 8, 19, 17, 43, 4, 0, -8, 8, -41, 3, -12, -7, -7, -60, -7, -28, -8, -3, 3, 12, 22, 9, -2, 0, 1, 6, -21, -3, -3, -16, -7, 46, -30, 8, -6, 3, 2, -6, 8, -2, -25, 33, -1, -7, -33, -30, -9, 38, 2, 5, -12, -7, -51, 4, -5, -4, -2, 3, -3, 8, -4, -5, 35, 33, -11, 7, 2, 14, 0, 0, -3, 7, 0, 0, -1, -23, -13, 5, 0, -17, -5, 1, -4, 8, -3, -36, 5, 21, 25, 32, 3, -5, -12, -45, -1, -4, 9, 4, 5, 9, 5, 0, 10, 1, 42, -5, 0, 7, 2, -14, -4, 14, -4, 7, 15, 0, -34, -2, -6, 15, -10, -3, -11, 27, 0, 2, 0, 4, 5, -10, 28, -14, -14, 8, 40, 17, 5, 1, -23, 6, 8, -1, 12, -25, 0, -4, 10, 6, -18, -4, 10, -32, -4, -45, 0, 16, 33, 12, -4, -2, 0, 30, 1, 13, -7, -20, -9, -18, 7, 1, 7, 3, 13, 6, 3, 2, -13, 23, -14, 8, -1, -11, 10, -8, -10, 4, -19, 0, -4, 33, -22, 14, -12, -6, -40, 8, -30, 44, 13, -3, -21, -2, -18, -1, -28, 1, 0, 12, 12, 10, -1, -43, 59, -29, -13, -30, -53, 2, -10, -6, -7, 6, -19, -5, 8, 7, 3, 0, -13, 5, 7, -12, -20, -27, 21, -24, 22, -36, 13, 3, 7, -2, -21, 0, -11, -52, -34, -18, 0, 33, -3, -10, -1, -4, 25, 7, -7, -35, 3, -17, 17, 1, 8, -18, 2, -13, -23, 17, -5, -10, -5, 3, -62, 0, 12, 1, -17, -9, -14, 0, 0, 35, -16, -4, -1, 9, 4, 3, -9, 6, -9, -7, 16, -9, 17, -8, -13, 2, 22, -9, -4, 3, -22, 17, 7, 1, -21, -12, 41, 1, 21, -6, 24, 0, 0, -20, 4, -8, 1, 4, 2, 0, 29, -29, -27, 32, 4, 1, 0, -9, 6, -3, 3, 24, -9, 10, 1, 7, 2, -2, 1, -19, 1, 8, 12, -8, 0, 20, 0, 5, -17, 4, -6, -3, 0, 4, -5, 0, -19, 9, -54, -19, -1, -1, 6, 7, -7, -6, 5, -7, 27, -5, 0, -1, -14, 4, -6, 17, 19, -8, 22, 9, -4, -6, 7, 50, -1, 40, 0, -13, -15, 17, 13, 7, 16, 2, 24, 2, 7, -3, 5, 12, 4, 2, -12, -13, 4, -5, 29, 6, 2, -5, 5, -11, -3, 12, 5, -10, 24, -5, -61, -35, 2, -4, 0, 29, -23, -18, 0, 2, 3, 1, 20, -59, 2, 15, 2, 2, -61, 29, 2, 0, -7, 0, -20, 8, -8, -1, 6, -3, 2, -30, -4, 4, -9, 0, -3, 24, -10, 15, 6, 4, -31, 7, 7, 10, -11, 9, -48, -4, -27, 6, -16, -1, -10, 3, -46, -6, -3, -12, -13, 24, -4, 1, 0, -1, 0, 4, 8, 9, -3, -8, -22, -4, 5, 0, 23,
    -- layer=3 filter=0 channel=4
    32, -2, -35, -7, -8, 4, -34, -38, -7, -15, -8, 7, 10, -29, 13, -7, 38, -31, -35, 27, 6, -2, 26, 17, -26, 4, 4, -3, -29, 41, -30, -21, 8, 10, 0, -19, 6, -10, -6, 41, -6, -39, -12, 3, -4, -22, 19, -21, -26, -1, 1, 15, 6, -10, -17, -9, -22, -1, -4, -23, 6, 25, -31, -7, -6, 9, -46, 1, 2, 0, -4, -8, 0, 4, 6, -3, 3, 0, -2, -1, -2, 1, -34, -11, 6, -11, -6, 0, -11, -6, 12, 38, 15, -7, -9, 6, -9, 0, 47, 26, 0, 0, 32, -7, -6, -33, -11, -8, -18, -12, 32, 3, -7, 4, 3, -5, -4, -7, -5, -5, -8, -2, 35, -7, -3, 2, 0, -21, -20, -52, 5, -16, -4, -1, -22, 13, -7, 1, -46, -26, -2, -3, 0, -10, -29, 13, -18, 20, -9, -19, -19, 4, -2, 28, 0, -10, 1, 29, 10, -2, 4, -3, -39, 18, 0, 5, -25, 2, -49, -3, -12, 0, -10, -3, -5, -2, -19, -13, 15, -11, -19, -11, 12, 2, 1, -10, 16, -63, -12, -3, 3, 19, -13, 26, 7, -10, -9, -3, -20, -13, -24, 18, -7, 2, -3, -12, 2, 6, 3, 5, -10, -14, 16, 9, -19, -8, -6, -2, 6, 5, -7, 4, -34, -29, -5, 12, -20, -31, 17, 2, -18, 32, 3, -3, -3, -7, 0, 24, 32, 3, -3, 6, -4, -26, -3, -2, 0, -18, 0, 22, 27, -6, 3, -36, 3, -10, 42, 13, 13, -4, 13, -5, -5, 2, 5, 8, 0, -9, 4, 13, -6, -8, 29, 32, 11, -20, 0, -31, -2, 3, -4, 26, 12, 8, 29, 5, 4, -24, 20, 6, 2, -22, 4, 4, 12, -1, 7, -7, 3, -21, -16, -5, 9, -8, -42, 11, 6, -39, -15, -21, -1, 41, 1, -7, -9, 10, -9, -16, -18, -10, -11, -3, 15, -24, -2, 29, -4, 7, -6, 2, -12, 0, 14, 0, 12, 0, -5, 4, -11, 24, 6, -5, -3, -4, -24, -1, 0, -10, 22, -1, -2, -29, 11, 6, 0, -3, 2, 0, -8, -9, -9, -1, -4, 6, 1, -13, 30, -8, -5, 17, -2, 0, 0, -13, 2, -18, -25, 12, -6, 5, 8, 6, -37, -4, 7, 19, -24, -5, 4, -18, -33, -6, 18, 14, -34, 31, 30, -1, -19, 6, -7, 0, -27, 2, -12, -19, -20, 20, -1, 36, -3, 62, -6, -8, 1, -8, -6, -2, -6, 11, -1, 4, 1, 7, -10, -2, 5, 4, 1, -8, -57, -1, 30, 18, 2, -63, 18, 10, -8, 3, 1, -11, 0, -7, -5, 13, 4, 22, 31, -6, -3, 15, 8, -24, 23, -1, 1, -5, 0, -31, -4, -1, -7, 8, -6, 0, 20, 4, -11, 3, -3, 0, 17, -12, 6, 5, -29, -9, -5, 9, -16, 35, -60, -6, 0, -18, -8, -9, 6, -38, 16, 3, 10, 1, -5, -18, 7, -10, 2, -4, -1, -10, 5, -2, -7, -8, -9, -3, -3, -3, -3, -1, 27, -1, 6, 22, 0, -6, -3, -25, 0, 2, 7, 4, 10, -4, -28, 2, -38, 14, -28, 46, 1, -9, -20, -6, -20, 4, -7, -1, -3, 21, 13, 35, 1, -5, 16, -24, 2, 0, -6, -4, -9, -18, -4, -5, -7, -8, 19, -34, -20, 17, 3, -18, 8, 2, -17, 0, -1, 0, 2, -11, 41, 13, -23, 4, 1, 5, -41, 32, -6, -15, -5, -5, -3, -6, -2, 0, 3, 29, 28, 1, 12, 6, -35, -8, -2, 8, 12, 2, -10, 7, -15, 0, 29, 0, 36, 7, -4, -9, 32, -4, 15, 8, 2, 36, 16, 1, -20, -16, -30, 34, 27, 0, 6, -28, -2, 0, -4, 13, -6, -18, 5, 5, 32, 20, -9, 0, 6, -23, -9, -2, -27, 35, 0, 12, -34, -10, -1, 9, -19, -36, 3, 9, 2, -4, -7, 4, -60, 0, 3, -44, -5, -2, -6, 21, -24, -2, -2, -21, 5, 2, -12, 2, 29, 1, 6, 2, -3, 3, 25, -7, 7, 6, -3, 3, 3, 0, -26, 6, -13, -12, -14, 4, 2, 0, 0, -3, 11, -36, -46, 6, -8, -2, -14, 43, 77, -9, 2, 11, 37, 6, -8, 4, 8, -4, 33, 4, 5, -4, 1, 22, -18, -4, 32, 15, -14, 16, 4, -20, -3, 32, 13, 0, -24, -10, 0, 10, 1, -54, -3, 30, -16, 41, 0, 4, -6, 6, 0, 9, 14, 9, -12, -2, 2, -6, -12, -7, -4, -29, -40, 43, 45, 38, 49, -27, -8, -21, 50, 5, -17, -3, 30, 18, -7, -9, 6, -44, -3, 1, 7, 11, -4, 0, -25, 28, 30, -18, -11, -34, 33, 0, -7, -3, 19, -30, -6, 0, -4, -13, -17, 0, -8, 6, 4, 16, 1, -7, 27, -4, -4, -7, -3, 6, 9, -33, -26, -6, 7, -5, 26, -11, 38, 50, 39, 25, 0, -3, -2, -39, -33, 7, 4, -19, 17, 9, 4, -14, 8, 31, -3, 2, 13, -5, 13, -2, 1, 0, -11, -5, -23, -21, 9, -5, 0, 3, -10, 2, -6, -3, 18, 13, -20, 9, 4, 0, 0, 6, -15, 8, 6, 5, -7, 2, 2, 7, 4, 0, -40, 0, -5, -12, 6, 7, 2, -19, 2, 12, 6, 15, -2, 0, -2, 3, -15, 41, 3, -36, 24, 0, 3, -51, -23, 4, -20, -20, -14, -1, 0, -11, 8, 5, 0, 5, -32, -8, 44, -4, 23, -22, -8, 12, -3, -8, 13, -9, 0, 2, 2, -23, 27, -43, -5, -1, -6, 15, 43, -5, -5, -6, -2, 3, -42, 1, -44, -2, 3, 43, 13, -75, -4, -6, -3, -6, 28, -6, 3, 14, 2, -1, -19, -9, 0, -4, 14, -50, 16, -1, -9, -5, 12, 3, 2, 1, 2, 0, -4, 2, -38, -4, -4, 39, 4, -9, 0, -18, 0, 5, -18, -36, -2, -3, -46, 36, -5, 6, 3, 12, 7, -1, 0, -30, -2, 32, -3, -7, 16, 3, 31, 9, 7, 6, 5, 5, 13, 0, 3, 4, 1, -12, -52, -10, -4, 32, 18, 5, -5, -14, -9, -2, 9, -60, 0, 3, -9, 1, -9, -12, -26, -8, -26, -11, -20, -7, -3, 5, 0, 7, 10, 26, -7, 7, 4, 49, 24, -4, 0, 19, 37, -31, -2, -5, -9, 32, -2, -13, 10, -7, -14, 16, 44, -13, -12, -18, -7, -67, 0, -8, -29, 4, -18, -6, 3, 3, -28, -7, -18, -6, 3, -11, -27, 42, 6, -32, 1, 8, 8, -4, -4, 4, 7, 37, -6, 5, 14, 0, -17, -10, -3, -21, -3, 8, 3, 1, -42, 17, 42, 9, 35, -8, -1, -1, 28, 15, -37, -6, 7, 21, 3, 11, 16, -12, -23, 11, -8, -2, -3, -26, 1, 2, -4, -48, 8, -14, 0, 4, 10, 0, -31, 7, -17, -24, -1, -19, -40, 58, 3, 42, 9, 2, 0, 13, 32, -5, 0, 9, 0, 0, -22, 6, -28, -2, 8, -71, -26, 7, -5, -28, 33, -2, 1, -22, 13, 2, -10, -3, 22, 32, -7, -6, -37, -2, 30, -3, -32, 22, 51, -1, -4, -1, 3, 26, -27, -1, -3, -7, -5, -3, -5, -3, 10, -15, 21, 1, -17, -2, -19, -53, 11, 6, 4, 8, 0, 4, -22, -21, 9, 15, 40, -4, 8, 7, 6, 2, -27, -46, 11, 29, -11, 12, 0, -10, 4, -7, -10, 2, 17, 6, -9, 17, -10, -51, 26, 1, -5, -3, -10, -3, 4, 6, 8, -13, -5, -2, 22, 5, 4, -21, -10, 2, 7, -35, -57, 5, 3, 5, 4, 43, -4, 21, 30, 8, -9, 7, -80, 22, 17, 0, -56, -15, -4, -12, -6, -2, -5, 4, 29, 33, -21, -30, -11, 12, -23, 6, 0, -4, 0, 1, 0, 32, -4, 10, 8, 0, 0, -18, -4, -26, -9, -8, 11, -14, -7, 37, -14, -3, 8, -10, -18, -9, 10, -61, 13, -22, 29, -5, 1, -10, -7, -5, 3, 23, -36, 2, 34, -3, 16, -7, -11, -30, 0, -3, 8, 13, -28, 15, -10, -7, -25, -4, 2, 1, -2, 6, 0, 0, 6, 1, 19, -4, 0, 4, 26, 3, -31, -17, 4, 4, -20, -5, 34, 7, 4, -5, -7, 0, -3, -7, -2, -28, -46, 6, 2, 10, -3, 0, 9, -21, 0, -11, -19, 12, 5, -7, 43, 0, 23, 0, 0, -42, -14, 0, 9, -9, 24, -9, 5, -12, -2, -20, 6, 9, 4, 0, -18, 0, 19, 5, 40, -15, 49, -27, -45, 6, -11, -14, 16, 4, -8, -4, -9, -16, 21, -38, -6, 5, -40, 34, -6, 2, -5, 5, -26, -7, -24, 5, 19, -52, -1, 0, -21, 3, -3, -2, 12, -21, -11, -5, -10, 9, -10, -33, -26, -5, -5, 4, 0, -44, 13, 5, 7, -7, -2, -5, 1, 0, 3, -7, -6, 1, -25, -8, 35, 7, 3, 1, 16, 10, -12, -3, -57, -11, -4, -1, -40, -15, -3, 38, 6, -11, -2, 27, 8, -42, 1, 20, 3, 1, -42, -27, 38, -1, -9, -5, -8, -2, 20, -9, 7, -5, 4, 26, 1, 1, -5, 24, -10, -3, -7, 49, 1, -5, -27, -32, 32, 30, -9, -3, 7, -22, -8, -7, 21, -1, 0, -14, 6, -7, 2, -9, -5, -9, -1, -8, -12, 5, -9, -56, -3, -6, -17, 35, -7, -4, -10, -5, -6, 5, 8, -5, 0, 1, -43, -37, -15, 9, -5, -27, -5, -7, 15, 0, 39, 3, 3, 22, 7, 7, -14, 1, -26, -15, 0, -15, 0, -20, -2, 2, 11, -11, 0, -5, 0, 4, -33, -3, 50, -6, 7, -6, -5, -14, 19, -9, -9, 4, 0, -37, -8, 14, 9, -6, 5, -1, -33, 2, 8, -15, -1, -6, 20, -31, -12, 10, -22, 6, -5, 6, -4, 15, 0, -8, -2, -1, 1, -15, 4, 1, 23, 19, -15, 3, -3, 2, 8, -12, -18, -46, -7, 6, 13, 9, -8, -5, -15, 4, 3, -14, -6, 6, 6, -18, 11, 3, 0, 49, -10, -12, 3, 25, -28, 4, -13, 25, -41, -10, 18, 3, 15, 29, -2, 6, 18, -6, 15, -6, 1, -6, -11, -1, 1, -9, -10, 9, -4, -4, -21, -7, 0, 4, -14, 5, 7, 15, 19, 5, -1, -8, 17, -48, -23, -4, 2, 35, -3, 65, -13, 6, -6, 2, -18, -13, -4, -5, 5, 5, 27, -51, 12, -29, 12, -9, 4, 3, 6, 9, -6, 2, 6, 11, -10, 3, 25, 19, 7, 11, -50, -29, -9, 5, 9, -4, 7, -16, -21, 0, 0, -3, -4, -34, 5, 27, -21, -60, 20, 30, -7, -20, 0, -69, -1, -37, 6, 3, -5, -18, 30, -10, 12, 4, 13, -2, -1, 5, -7, -2, -4, 5, -5, 29, 29, -30, -14, 7, -32, 4, -12, 55, 10, 37, 7, 4, -8, -67, 1, -8, -6, -6, -3, -21, -16, -4, 0, -5, -4, -1, 13, 0, -18, -13, 27, -3, -5, -35, 32, -31, 9, -7, -7, -17, 3, 3, 21, -20, -88, -5, -17, 12, -13, -2, 2, 12, -6, 19, 6, 6, -23, 23, 26, -8, -7, -3, -2, -9, -14, -17, -9, 4, -6, 0, 19, -1, -2, -12, 14, -5, 10, -78, -2, -1, -12, -2, -1, -6, -2, -5, -4, 1, 28, 5, -6, -48, 18, 4, -9, -1, 6, 11, 3, 17, -2, 8, -2, 13, 3, -14, -25, 4, -61, 19, -4, -7, 7, 2, 1, 34, 15, -4, 8, -15, -38, -18, 36, -6, -27, -14, -50, 3, 20, -3, -2, -20, 5, -11, 34, 9, 3, -49, -3, -10, -5, -12, 15, 11, 27, 24, 26, -6, -12, 4, -20, -15, 3, -7, -13, 1, -67, -5, 23, 17, 4, 34, 34, 1, -8, 1, 58, -9, -4, 4, -5, -3, 0, -23, 8, 4, -7, -16, -6, 21, -29, 6, -2, 6, 13, 9, -6, -1, -10, 3, -3, 9, -17, -6, -30, -29, -2, 0, -36, -21, 7, -8, 20, 8, -2, -8, 20, -7, 2, -24, 4, 75, -6, -6, -8, -38, -15, 3, 5, -8, -6, 25, -19, 5, -9, -2, 0, -4, -7, 0, 0, -10, -1, 1, -23, -1, 2, 18, 4, -5, -24, -21, -6, 0, 62, 12, -4, -18, -10, 2, 5, -6, -41, 0, -44, 12, -24, -38, 6, 6, 8, 19, 18, 26, -5, -5, -23, -48, -2, 25, -1, 15, -38, -19, 2, 2, -2, -27, -6, 26, 19, -2, -16, -1, -52, -38, -12, -39, 0, -45, -5, 4, -17, 32, 11, -6, -3, 27, 7, -9, 27, 3, 5, -64, 7, 7, 0, -24, 7, -1, -5, 0, 4, 1, 0, -22, -15, 6, 4, -3, 38, 0, -2, -4, -2, 5, 3, -5, -22, -7, -1, -32, 15, 6, 6, -2, -4, 8, -4, -4, -21, -36, -32, 2, -5, -20, -31, -6, 1, -4, -1, -16, -3, -1, 4, -36, 2, 6, -4, -6, 13, 11, -19, -1, 1, -9, 43, -28, -17, -62, -3, 21, -42, -17, -1, 10, 37, 10, 7, -6, -6, 2, 1, -18, -76, 1, 3, 25, -11, -1, -5, -37, -3, -6, 0, -10, 11, -8, -11, 7, 3, -17, 1, 2, 21, 6, -35, -39, -14, 23, 19, -5, 5, 8, -41, 13, -24, 23, 51, -17, 14, 7, -10, -6, 16, 5, -38, 2, -5, 31, -45, 35, -16, 4, 2, -21, 1, -40, -15, 6, -3, 0, -10, 23, 0, -9, 10, -12, 39, 40, -34, -34, -12, -4, 4, 32, -3, -32, 0, 3, -49, -12, -1, -10, 10, -9, -8, -3, -25, -86, 0, 6, -4, 1, -3, -25, -44, -3, -77, 8, -8, -17, 4, -49, 2, -19, -21, 9, -35, -33, 16, -44, -6, -28, -6, 0, 0, 2, 21, 22, 11, 7, -8, -37, -2, -2, -3, 30, 5, -1, -27, -28, -12, -38, -16, 25, -25, 7, 0, -92, -23, 4, -49, 35, -4, -8, 26, -14, -1, 28, -7, -47, -25, -9, 0, -22, -1, -27, -26, 0, 10, -26, 5, -9, -3, -3, 21, 1, -3, -21, -5, 12, 9, -2, 41, -1, -29, -3, -15, 3, -6, -12, 12, 4, -2, -23, 1, 37, -67, -43, 5, -3, -29, -1, 5, -7, -8, -37, -26, 5, 2, -5, 36, 2, 0, 2, -3, -3, 6, -13, 22, 8, 5, 2, -17, 9, 0, -9, 4, 4, 28, -3, -1, 9, 19, 0, -4, -68, 2, -9, 6, -28, -2, -22, -33, 45, 5, -24, -20, 1, 8, -25, -6, -12, 44, -10, 0, 21, 25, -7, 8, -3, -12, -34, -29, 1, 26, -11, -13, -7, 14, 11, 5, 11, -28, 1, -23, -6, 2, -37, -21, 1, -18, -3, 34, -4, -7, -28, 28, -8, 4, -18, -49, 0, 4, 2, 18, -1, -25, 8, 36, 43, 8, -15, 0, -28, 0, 0, -1, -23, 14, 0, 8, -1, -2, -57, 6, 3, 1, -18, -33, 33, -7, -1, -9, -1, 0, -6, 3, -2, 0, -10, 1, -5, 39, 4, -52, 8, -3, 2, -19, 23, -6, 2, 89, -20, -5, 5, -48, 3, -16, -1, 22, 37, 0, 21, 3, -8, -6, -28, -10, -10, -10, -45, -62, -1, 2, -8, -3, -9, 7, 4, 1, 5, -7, -30, -4, 6, -4, -6, -13, -9, 5, -16, -3, 3, 22, -5, 0, -4, 4, 0, -1, -10, 34, -1, -21, 28, 14, -41, -9, -6, 6, 14, -15, 0, -7, -11, 1, 0, 12, 21, 2, 18, -20, 8, 1, -1, 2, 15, 6, 7, -26, -3, -4, -2, -9, -26, -21, 26, -3, -15, -5, -9, -13, -18, -29, -4, -10, 16, 1, 3, -7, 3, -19, -45, 20, 0, -12, -25, -6, 8, -1, -5, -9, 2, 5, -20, -33, -8, 7, -10, 5, -6, -7, -12, -4, -5, 4, 5, -19, -7, 2, 48, 51, -1, -5, -4, -27, -12, 69, -13, 24, 2, -29, 42, -7, -16, -6, -10, -6, 0, 0, -33, 1, 5, 10, 6, 2, 2, -5, 1, 7, -22, -27, -4, -59, -3, -5, -10, 22, 19, -6, 6, -35, 4, -4, 4, 0, -41, -9, -2, 6, 0, -55, -7, -16, 10, 5, -28, -7, 2, -5, -22, 12, 6, 0, 6, -12, 4, 15, 2, -11, -15, -8, -9, 23, 4, -2, 22, -11, 81, 5, -4, -2, -7, 5, -7, 0, -4, 1, -18, 10, 6, -2, -2, 10, 6, 0, -2, 0, -37, -14, -66, 8, -8, 7, -27, 21, -26, -14, 24, 6, 5, -19, 17, 6, -12, -2, 37, 8, -4, 9, 26, 5, -30, -2, -14, -3, 14, 2, 6, 41, 7, -1, 11, 21, 1, -33, 1, -37, -72, -1, -19, 0, -7, -5, -18, 5, -4, 44, -7, 4, 10, -6, -19, 1, 18, -27, -31, 8, -9, -32, -3, -7, 12, -14, 4, 16, 1, -38, 4, -2, -9, 2, -26, -4, -2, -4, 48, 0, 1, -36, -41, 2, -2, -3, 12, -8, 2, -7, -19, -23, -24, 20, 22, -7, -22, 15, 11, -4, 18, -4, -34, -9, 4, 15, -11, 1, 24, -2, 6, 24, -2, -23, 19, 0, 16, -5, 21, 27, 32, -1, 14, -3, 8, 15, 3, -19, 5, -11, -13, 25, 7, -6, -7, 3, -11, 5, -14, 14, -12, 15, -2, -14, 9, -10, -14, -4, 7, 2, 6, -28, -9, -24, -3, 5, -19, -9, -5, 27, 45, 16, -6, 8, 2, -24, 0, 2, -14, -6, -6, 15, 2, -1, 39, 20, -4, -11, 29, -8, 8, 3, 15, 3, 7, -6, -8, -1, 19, 24, 6, 12, 3, 0, -26, 2, 0, 4, -5, 15, 0, 4, 9, -22, 25, -18, 0, -13, 0, 56, -2, 0, -2, 0, -7, -7, 28, -39, -53, -6, 0, 4, 7, -4, 0, -14, 24, 20, -15, 28, -2, -15, -7, 8, 13, -7, 5, -21, -6, -22, -3, -23, 28, 2, -20, -12, 19, -6, 7, 44, 2, 0, 3, -6, -15, -7, -22, 36, 6, -3, 2, -4, -15, -1, 3, -3, -6, -13, -16, -7, 10, -1, 5, 11, 3, 3, -6, 16, 6, 6, -8, 22, 8, -7, 3, 45, -18, 0, -5, 30, 1, 6, 9, -15, 52, -5, -20, -4, 27, 13, -22, 4, -8, 1, 24, -19, -8, 5, -6, 3, 7, 0, -4, -7, -8, -5, 9, -8, 1, -4, -7, -25, -3, 19, 0, 5, 0, 1, 17, -31, 19, -6, -5, -1, 11, 26, 0, -16, 6, 34, -19, 0, 0, 0, 13, 17, 22, 0, 6, -22, 23, 9, -7, -7, -5, -55, -17, -1, -10, 5, 36, -7, 6, -5, -9, -9, -8, -41, -6, -8, 24, -6, -3, 9, -3, 25, 49, 20, -4, 7, 39, 20, 45, 18, 3, -7, 2, 18, 40, -5, -33, -6, -8, -10, -3, -6, -5, -7, -5, -4, -5, -37, -2, -34, 1, -7, 8, 6, -9, 0, 9, 31, 18, -51, 1, 33, -7, 2, -6, -10, 32, -84, -2, 0, -52, -5, -3, 16, -4, -29, -6, -6, 5, 3, 12, 10, -6, 0, 11, -2, 25, -6, -7, -14, -31, -36, -3, -25, 6, 1, 24, 4, -58, -1, 2, 11, 6, 7, -1, 5, 1, 0, 4, -3, -1, 5, -4, 9, 21, -9, 28, -7, -8, 3, -8, 12, 3, -1, -54, -39, 8, -35, 6, 0, 30, 8, -5, 13, -1, -61, -5, 27, -24, 0, 4, -8, -4, -25, 16, 22, -5, 3, 8, 3, -9, -5, -6, 7, 21, 34, -3, -9, 0, 38, -14, 12, 1, -7, 6, -22, 12, -5, 23, 6, 7, 35, 11, -1, 1, -3, -3, 11, -46, 19, 3, 6, 22, -1, -10, 5, 38, 1, -2, 21, -9, -2, 2, 2, -25, 4, 0, 14, -44, 11, -15, -4, -6, -2, 34, -6, -8, -17, -4, 2, -28, 3, -26, 30, 9, -4, 0, -12, 32, -47, 13, -3, 20, 8, -1, 23, -1, -71, 7, -10, -9, -16, -35, 2, -7, -5, 6, -10, -2, 15, 37, 8, -11, -8, 30, -5, 5, 7, 57, -3, -21, -4, 46, -3, -31, 5, -26, -7, 9, -6, -14, -20, -1, -5, 19, -3, -7, 64, -7, 8, -31, 14, 13, -6, 5, -19, 3, -12, -14, 17, -1, -14, 6, -23, -23, -43, 6, -16, 10, -25, -22, -2, -24, -3, 13, 2, 0, 10, 14, -15, -5, -17, 5, -9, 18, 13, 4, 0, 3, -7, 7, -13, 2, 10, -14, -10, 3, 23, 22, -1, 5, -3, 6, -43, -7, 4, -6, -3, -7, 14, 5, -3, 3, 59, 0, -11, -3, 0, 13, -2, 26, 3, 32, -23, -13, 5, 19, -20, 5, 17, -10, 2, -8, 37, 6, 0, 42, 0, -2, -27, 22, -6, -15, -2, -7, -15, -6, -4, 9, -23, 3, 24, 17, 23, 39, 24, -12, 0, -28, -25, -9, -16, -3, -14, 4, 9, -20, 22, -5, 0, -27, -2, -7, -7, -7, 29, -8, -21, 5, -52, 20, -6, -2, -17, 9, -4, 0, 0, 6, -7, 1, 3, 8, 4, 11, 0, 0, 3, 6, 35, 11, 2, -6, 2, -12, -3, 10, -2, 3, 7, -7, 1, -1, 1, 7, -24, -29, -7, 5, -27, 21, -9, -4, -49, 7, 9, -7, 19, -10, 23, 23, 8, 18, 6, 16, 3, -12, 25, -65, 3, 4, -67, 28, 10, 3, 0, -6, 1, -4, -6, 0, -4, 6, 2, 33, 3, 15, 0, -18, -31, 7, 10, -67, 5, 3, 39, -16, 4, 30, -1, -1, 4, 14, -24, 2, -19, -27, 0, -40, 2, -10, -19, -8, -15, 11, 1, -8, 18, -12, 11, 4, -1, 23, -18, 8, 2, -5, -11, 32, -3, 4, 7, -1, 0, -12, -18, -30, -3, -19, 2, -46, 7, 5, -34, -25, -28, 2, 4, 2, 2, -4, 29, -7, -28, 45, -7, 5, -1, 13, -2, -1, -12, 0, -5, 4, 4, 8, 11, -1, -55, -3, -11, 6, -1, 20, 11, -4, -7, -8, 7, -12, -23, 13, -32, 6, -3, 6, 27, 37, -75, 0, -8, -23, -3, -40, 3, -13, -46, -9, 0, 6, -2, 9, 0, 2, -1, -5, -4, -15, -6, -4, -3, -18, 20, -3, -16, -19, -34, 34, -33, -53, -10, -1, -27, -7, -4, 0, 0, -29, 4, -1, 4, 1, 2, 53, 32, 28, 1, 41, 12, -6, 1, -47, 24, 0, 2, -48, -17, 1, -23, -3, 3, -12, 0, 7, 46, -5, 23, 5, 29, -45, -17, -3, -6, 6, -47, -12, -9, -63, -38, -9, 0, 0, -11, 3, 2, 30, -16, 6, -20, -8, -53, -4, -41, -6, 5, -6, 27, -34, -3, 12, 4, 13, -22, 7, -14, -5, -3, -50, -2, 34, -1, -12, -5, 28, -1, 28, -4, 41, 0, 5, 32, -3, -3, -2, -12, -9, 24, -21, -29, -51, -8, 2, -1, -1, 4, 9, -6, -10, -15, 5, -2, -10, 3, -7, 54, 23, 36, -7, 0, -17, -23, -40, -3, 25, -11, -3, 23, 28, 4, -9, -15, -24, -16, -28, 1, 0, -1, -6, 2, -6, 5, -9, -22, -13, -1, -36, 22, -7, 1, -13, -38, 46, -55, 12, -4, 44, -17, 0, 6, -9, 5, 6, 8, 1, 26, 18, -3, -1, -12, 0, 23, -52, 18, -21, -5, 25, -1, -4, -17, 35, -12, 2, -2, 2, -4, 2, 4, 0, 7, 18, -15, -9, 15, 2, -4, 1, -2, 31, -32, 25, -14, -6, -34, 0, -10, 17, 1, -31, 6, 0, -1, -3, 46, -9, 7, -21, 0, 2, 15, 21, 9, -7, -6, -3, -13, 1, 6, 13, -5, 5, 19, -1, -8, -24, 34, 4, -12, -8, -10, -11, 11, 2, 0, 13, 15, 83, -7, -21, -32, -3, 13, 4, 6, 3, 5, 0, -4, -26, 29, 4, 4, -35, 5, -39, -49, -14, -14, -12, 0, 1, -15, -8, -30, -16, -31, 8, 16, 13, -4, -131, -24, 2, -3, 3, 0, -5, 2, 25, 17, 7, 64, 0, -1, 2, -8, -1, 28, -2, -7, 2, -50, 1, 0, 12, -2, 6, 0, -4, 28, 17, 1, 0, 0, -5, 3, 52, 26, 0, -4, 15, 39, -18, 8, 0, 1, -1, 5, -3, 0, 0, 0, -2, 4, 2, 35, 7, -21, -24, 0, 0, 0, 31, -14, 5, -24, -14, 8, 7, 23, -18, 45, -21, -2, 13, 3, 29, 10, 46, 0, -17, 10, -5, -21, -47, -35, -5, 4, -9, 2, -7, -27, 8, 6, 7, -6, 7, -52, -6, 0, -45, 17, 3, 21, 8, 5, -10, -2, 11, 3, 4, 0, -9, -7, -21, 26, -6, -5, 8, -19, 1, 0, -7, -12, 5, 0, -13, -6, -7, -3, 48, 17, 0, 0, 32, -43, -5, -3, -1, -4, 34, 2, 19, -1, 2, -2, 18, -47, -10, 0, 18, 8, 23, 2, 7, -6, 24, -25, -1, 10, -16, 13, -10, 18, -8, -16, 5, 11, 7, -8, 37, 0, 0, 5, 4, 5, -8, -3, 0, -15, -6, -9, 9, 8, -2, -3, 0, 7, -7, 3, 11, -22, 36, 17, 39, 14, 4, 6, -3, -47, 39, -19, 4, -16, 34, -15, 7, -47, -11, -44, 20, -5, -12, 7, 25, 0, -6, 2, 23, 2, -29, 9, 0, -83, 27, -32, -4, 8, -20, 10, 5, -17, -23, -5, -1, -45, -11, -2, -3, 2, 0, -4, 1, -6, 5, 25, 24, -3, -9, -8, -4, -12, -13, 9, -51, 5, 0, 6, 22, -36, 7, 26, -9, -4, -5, -8, 3, 43, 3, 2, 26, 16, 10, -15, -4, -9, -8, 22, -2, 12, -11, -40, -24, 0, -6, -1, -6, 22, 21, -27, 8, 2, 25, 7, -49, 16, 3, 0, -4, 10, -15, -29, -4, 10, 5, -9, 12, -2, -6, 2, 4, 15, 21, -10, -14, 4, 28, -4, 13, -3, 26, -14, 2, -4, 0, -10, -4, 5, -49, -12, -3, -8, -42, -2, -2, 4, 1, -4, 23, 20, 2, 28, 5, 2, -1, 0, 24, -23, -26, -16, -13, -8, 48, -4, -18, 0, 1, -33, -1, -12, 21, 4, -12, -1, 4, 49, 0, -3, 4, 4, -9, 2, -3, 11, -6, 4, 12, -4, -25, 2, 7, 0, -29, -7, -5, -3, 38, -7, 19, -6, -26, -3, -12, -6, -2, 13, -1, -2, -1, 1, 0, 22, 7, 13, -32, -11, 29, 6, 26, -15, -1, -14, 26, -19, -6, -11, 5, 22, 6, -34, 4, -9, -51, 18, 25, -3, 29, -2, -10, -1, 51, 33, 19, -27, 7, -17, 1, -6, -5, 36, -27, 2, -6, 7, 0, 13, -7, -3, -15, -41, 3, 41, -5, 25, -3, 1, 8, -56, 0, -5, -10, -6, -4, -13, 0, -8, 27, 23, 7, -1, -2, 0, 3, -4, 28, -1, 50, 29, -10, -4, -19, -5, -6, -12, -27, -8, 13, 11, 5, 0, 13, -16, 2, 0, 2, -36, -34, -30, 23, 14, 10, -8, 9, -24, 0, 0, -9, 9, -47, 14, -45, -2, -35, -13, 7, -7, 0, -1, -16, 26, 24, 36, -2, 7, -42, -4, -11, -5, 3, 4, 6, 1, 2, -51, 20, 9, -4, 9, -17, -3, 7, 15, -3, -23, -3, 0, -9, -4, 0, 18, -5, 8, -13, 11, -1, 25, 0, 6, -8, 10, -36, -3, 7, -8, 0, 3, 9, 51, -6, -7, -51, -2, 4, -20, -17, -5, -2, -3, -19, -1, 0, 44, -13, 18, 28, -12, -3, 0, -13, 11, 19, 17, 8, 1, 6, 25, -38, -8, -7, -6, 0, 6, 0, -63, 4, 0, -4, 1, 10, -15, -6, -8, -24,
    -- layer=3 filter=0 channel=5
    3, -3, -12, -41, 5, -1, -1, 10, -11, -18, -8, 0, 0, -28, 2, -8, 62, -13, 27, 12, 0, -5, -46, -29, -12, 12, 5, 3, -36, 18, -10, 32, 3, 26, 7, 32, -8, 1, -4, 22, 6, -24, 15, -2, 7, 8, -1, 37, -25, -15, 0, -25, 7, 4, -6, 2, -28, 0, 2, -15, 12, -41, 18, -8, 15, -2, -5, 3, -2, 20, 0, -8, -8, 3, -7, -7, 0, 2, -6, 7, -15, 8, 25, 0, -8, -12, -2, -7, 1, 5, 3, 26, -18, -23, 15, 2, -1, -5, -17, 14, -48, 4, -3, 0, -82, 27, 18, -9, -31, 3, -25, -6, -2, -22, -1, 2, -10, -14, 0, 6, 1, 3, -16, -9, 13, -2, -14, -18, -10, -3, 31, 13, 8, 21, 7, -2, -2, -3, 21, -7, -6, 1, -9, 6, 12, -17, 7, -6, -4, 30, 18, 0, 8, 8, 6, -2, -3, 20, 46, -2, -16, 7, 35, -13, -3, 3, 14, -2, -28, -50, -29, -1, 11, -9, -7, 3, 27, 9, 20, 6, -16, 2, 5, -2, 0, 0, 12, 14, 32, 5, -5, 6, -26, -18, -20, 9, 3, -41, 27, 14, 4, 12, -1, -5, -21, -13, -12, -9, -3, -18, -7, -10, 11, 31, -16, 67, -8, 6, 1, -39, -3, 1, 1, 15, 13, -5, -23, 50, -24, 29, -30, 45, 6, 8, 4, -5, 7, -7, -4, 3, 29, -9, 5, 5, 0, -22, -6, 49, -51, -15, -60, 17, 31, 17, -5, 9, 39, 8, -38, 5, -11, 29, -24, 4, -55, -14, -7, 8, 1, -26, 4, -8, 4, 9, -43, -16, 0, 31, 11, -4, -5, 9, -39, 31, 16, -13, -4, 73, -5, 26, 0, 13, 2, -35, 42, -3, 34, -7, 3, 30, -39, -1, -5, 0, 4, 3, 8, 33, -79, -49, 15, -18, -13, -29, -3, 0, 24, 10, 36, -3, 14, 21, -9, 0, -15, 28, 0, -5, -6, 18, 8, 3, -11, 0, 2, 3, 0, -9, -21, -1, 12, 2, -6, 0, 38, 6, -3, 1, 14, -4, -38, 16, 2, -7, 9, -5, -6, 6, -4, -1, -10, 5, -73, -3, 1, 9, 23, 0, 5, -8, 1, 7, 8, -2, 3, 40, 5, 27, -4, -10, -28, 5, 0, -16, -4, 18, -50, -6, -2, -12, 24, -5, -22, -40, -15, -41, -4, -11, -44, -5, -69, 5, 29, 2, 13, -14, -9, -15, 18, 31, -1, -25, -22, -4, -11, -4, 5, 42, -22, 24, 79, -5, 15, -58, 20, -4, 0, 0, -7, 0, 27, 4, -20, 28, -2, 8, 10, 6, -7, 8, -18, 8, -2, 6, 6, 2, -10, -2, -19, -4, 0, -11, 10, 17, -11, 7, -8, 5, 0, 7, -5, 7, 5, -8, 0, 0, 1, 0, 31, -5, -5, -3, -40, -25, -3, -4, 18, -17, 0, -7, 1, -37, -3, -4, -3, 52, 7, 4, -10, -46, -2, -34, -9, -10, -19, 20, -15, -11, -5, 4, -1, 2, 8, 6, 0, 7, 5, -17, -38, -12, 5, 13, 14, 7, -18, -15, 2, -5, -57, 50, 33, 6, 3, -3, 3, 1, -13, -2, 23, 30, 2, -32, 1, 6, 21, -10, 21, -27, 0, -8, -25, -1, -24, -4, -3, -8, 5, 3, 5, 8, -5, -21, -4, 0, -21, 7, -12, 20, -17, -35, 16, -6, -2, -8, 6, -2, -1, 27, 6, 3, -4, -16, 3, -8, -5, -15, -1, -14, -16, 9, -8, 12, 11, 6, 4, 0, -8, -13, 3, 55, -63, -3, 9, 0, 4, -7, -3, -20, 6, 2, 3, 7, 44, -14, 15, 48, 10, -9, 0, 2, 24, -8, -25, 3, -15, 2, -1, 46, 50, -2, -12, -36, -11, -3, -2, 5, -8, -10, 2, 17, -4, 0, -1, -9, -26, 26, 25, 6, -16, 5, 16, 37, 15, -31, -8, -21, -3, 0, 8, 10, 2, 2, 7, 2, -4, -7, -8, -32, 18, -51, 0, 40, -4, 0, 3, -45, 2, -7, -7, 18, 21, -7, -4, 0, 20, -5, 0, 1, 28, 2, 22, -1, -18, 45, -45, 9, 1, 0, 14, 42, 54, 3, 22, 2, -3, 1, -1, 2, -14, 21, 9, 1, 3, -28, 11, 4, -21, -3, -2, -12, 8, 10, 7, -5, -2, -8, -14, 5, -19, 3, -2, 16, 29, -20, -8, -5, -9, 13, 6, -20, 9, -33, 4, 0, 4, 5, -3, 2, -7, 15, -8, -5, -43, -9, 1, -1, 1, -8, -1, 4, 6, 0, 63, 4, 5, 20, -9, 15, -8, 4, 2, -19, -29, 12, -27, -18, 4, 6, -39, 11, 1, -60, -13, 2, -13, 0, 7, -5, 8, 2, -6, 15, 5, -3, -12, 9, 17, -26, -19, -4, -27, 0, 7, -10, -28, 18, 19, 1, -1, -7, 13, -11, 5, 23, 6, 12, -18, -1, -56, 7, -7, 6, -13, 0, 55, 44, -4, -9, 4, -6, 7, -5, 20, -35, -19, -9, -16, 7, 25, 23, 51, 0, 18, 21, -27, -41, 1, 43, 1, 28, -1, 16, 22, 11, 14, 0, 17, -4, -1, 0, 4, -9, 6, 2, -16, 0, 35, 6, 1, 13, 48, 1, 8, 14, -1, 2, 1, 0, 26, 7, 0, -7, 3, -5, -5, 2, 3, -39, -17, -3, -19, 9, 0, -13, -2, -6, -2, 29, -13, 11, -7, -39, -13, -5, 11, -32, 3, 8, -6, 4, 8, 6, 15, -7, -25, 17, -23, -8, -25, 3, 3, -15, 40, -2, 49, 4, -16, -9, -17, 26, 36, 16, 4, -75, -30, 1, -36, 5, 0, 0, -68, 56, 51, -8, -28, 27, -34, -1, -12, -6, 41, 4, 23, 6, -17, 1, 6, -13, -3, -26, 8, -4, 33, -1, 17, -2, -6, 1, -5, 10, 18, -7, -6, -1, -19, 7, 39, 0, 4, 2, -2, 8, -6, 3, 4, 6, -13, 8, 41, 1, -42, -7, -6, 5, -11, 3, 8, 4, 1, 26, 0, 9, 22, -17, -4, 17, 2, 13, 1, 52, 6, 31, -8, -28, -18, 0, -4, -6, 4, -10, 1, 10, -6, 2, -13, 1, 3, -9, -1, -12, -25, 0, -1, 10, 23, -4, -34, 8, 1, 9, -18, 5, 10, 4, 6, -1, -9, 59, 29, 1, 26, 16, 4, 38, 6, -8, 0, -8, -31, -5, -7, -6, -1, -5, -17, 0, 4, 5, -7, -11, -3, 7, -10, -10, -2, 13, 3, -5, -10, -10, 2, 3, -8, 3, -9, -10, -4, -4, -13, -4, 11, 4, -7, -8, -25, 8, -16, -9, 7, -23, -5, -2, -8, 21, -6, 6, 2, -6, 2, 5, -5, -9, -5, 0, -29, 10, -18, 9, -5, -8, 11, -8, -2, 1, -8, 11, 12, -7, 15, -4, -9, 3, 49, 6, 29, -8, -7, -18, -45, 19, 33, -1, 11, -5, -5, 5, 0, -17, 0, -3, 6, 19, 2, 0, 8, 8, 30, -13, 16, -4, 4, 3, -55, -38, 9, -33, -7, -44, 3, -8, 2, -8, 20, -16, 6, -1, 1, -2, -49, -17, 18, 1, 7, 37, 0, -5, -2, 24, 26, -3, -4, -35, -21, 3, 4, 3, 1, 25, -3, -10, 4, 3, 17, 31, 22, 1, -17, -7, 6, 2, 31, -31, 19, 8, -15, 9, -23, 1, 1, -1, -7, 1, -19, -7, 11, -19, -41, -35, -56, -6, -9, 19, 66, -20, 7, 16, 7, -3, -52, 1, -20, 1, 0, -30, 35, 19, -17, -51, 8, -1, 1, -16, -4, 34, 3, -4, 22, 25, 2, -4, 7, 33, -42, 3, 16, 0, -5, 3, -1, -12, 4, -16, 28, 0, 6, 5, 5, 11, -3, -19, 19, 8, -20, 2, 52, -1, -53, 29, 1, -29, -31, 16, 8, 18, -15, -42, -2, -24, -3, -25, -9, 2, -7, 5, 1, 1, -44, -32, 31, -31, 0, -12, 18, -7, 5, -2, -16, -29, 25, 0, 9, 48, 24, -11, -5, 22, -4, 15, -47, -2, -4, 0, -5, -39, -22, 4, 43, -66, 50, -35, 8, 16, -53, 3, -30, 0, 1, -15, 5, -7, 15, -18, -4, -1, 14, 2, 16, -11, 8, 8, -8, 13, -15, -3, -1, -10, 21, 0, 17, -1, -8, 26, -43, -17, -1, -2, 0, 8, 17, 0, 5, 3, 44, -9, 41, -10, 1, 0, 12, -6, 25, 4, -3, -12, -1, 2, -11, -2, -1, -35, -11, 1, 1, 1, 1, 2, -4, 3, 0, 14, -24, 42, 5, -17, 17, 7, -6, 11, 0, 8, 38, 4, 0, 24, 8, -3, 17, 12, -52, -15, 6, -5, -10, -6, -30, 0, 17, -2, -37, -2, -56, -15, 7, 44, -3, 7, -6, 3, 12, 3, 14, 0, -34, 21, 4, -6, -18, -14, 13, -5, 6, -4, 15, 1, 17, -4, -12, 3, 2, -49, -24, 31, 1, 0, -32, 3, -1, 5, 2, -7, 0, 29, -35, 6, -5, -5, 42, -15, 9, -1, 3, -3, 0, -46, -4, -4, 7, 3, 9, -2, -21, -3, 30, 12, -5, 7, 22, 13, 7, -4, -1, 5, 4, 5, -16, 21, -31, -32, 0, 20, -4, 22, -1, 24, -36, 2, 0, 0, 7, -8, -26, -2, 3, -4, -6, 0, -40, 6, 4, -3, 3, 4, 4, 0, -2, -32, -44, 6, 16, -28, 5, 8, 13, 18, -22, 15, 0, -6, -8, 7, -14, 2, -4, 0, -6, -17, 4, 7, -15, 20, 0, -15, -8, -6, -27, 7, 20, -14, -2, -10, 6, 18, 9, -2, 0, -7, 2, -24, 40, -11, -12, 15, 1, -13, 32, 9, -4, 32, -7, 6, 24, 14, -8, 7, -7, 7, 28, -51, -21, 0, -1, -23, -39, -18, -2, -2, 1, -1, 2, 6, -7, -4, -6, 15, -4, 4, -9, -13, -27, -7, 5, 0, -13, -6, 2, -8, 27, 12, -9, 6, -1, -2, -2, 4, -1, -10, 9, -2, -15, 30, -14, -19, 25, -10, -64, -25, -2, 2, -3, -28, -6, -7, 7, -25, 0, -13, -2, 0, 9, -12, 0, -5, 14, -3, -23, 15, 17, -18, -4, 6, -10, -9, -7, -4, 5, -36, -4, 0, 5, -7, 5, 1, -21, 4, 10, -57, 8, -5, 3, 50, -15, -2, 2, -4, 12, 0, -12, 0, 29, -8, 0, 0, -7, 2, -17, 29, 10, 0, -35, -2, 8, 3, -9, 37, 7, -8, -16, 3, 0, 5, 16, -1, -15, 12, -23, -11, 0, 18, -25, -11, -3, 6, 6, -9, 15, 14, -12, 23, -9, 5, 25, -21, -15, 5, -9, 14, -1, -11, -11, 19, -9, -2, 9, 19, 3, -12, -1, -6, 3, 0, 0, 0, -15, -21, -81, 26, -45, 44, -9, 2, -1, -2, -4, 20, -11, 3, -18, 5, 0, -68, 7, 20, -15, 0, -9, -33, -15, -19, 22, 16, 2, 39, 25, 3, -21, 7, -12, -3, -22, -12, -42, 3, -8, 3, 10, 6, 2, 3, 21, -8, -7, -37, -2, 22, -9, 6, -4, -9, -32, 4, 15, 35, 6, 9, 26, 0, 0, 8, 7, -53, -13, 7, 8, -5, 4, 0, -3, 6, 3, 6, 18, -26, -6, 14, 12, -37, -58, 6, 12, 11, -13, -5, -34, -2, 26, -3, 4, -6, 15, -21, 16, 7, -3, -14, 2, 26, 43, 3, 7, 11, 12, 4, -8, -17, 16, -6, 5, 7, 3, 11, 7, -1, -1, -8, 3, -5, -25, 4, 6, -6, 16, 0, -12, -3, 7, -8, -1, 5, -15, 1, -8, -12, 8, 10, 3, 41, 10, -14, 7, -11, 6, -19, 12, -41, -5, -8, 24, -3, 20, -33, -10, -75, -8, 1, -7, -12, -12, 5, -15, -14, 48, 3, -33, -9, 22, 0, -24, -11, -27, 6, 1, -5, 35, -29, -28, 2, 5, 12, -7, -8, 9, -1, -23, -25, -10, 3, -7, 5, 7, -32, 10, -7, 0, -3, -47, -5, 50, 3, -40, -32, -4, 39, 1, 14, -4, 0, -13, -6, -19, 5, -3, 11, -7, -46, 15, 0, 16, -4, 29, -5, -7, -2, 3, 0, 3, 0, 6, 1, 8, -11, 3, 10, 17, -10, -46, 35, 2, -5, -23, 27, -7, 4, -30, -25, -1, -5, -46, 16, 1, 15, 1, -22, 8, -12, -5, -10, -13, 27, -7, -1, 12, -4, 10, -9, 7, 4, -6, 0, 2, -4, 2, -6, -6, 4, -90, 6, 4, -7, 0, -10, 10, -36, -5, 1, -12, -27, -12, -17, -7, 6, 3, -16, -36, 2, 12, -49, -7, 19, -4, -1, 19, -21, -23, -26, -5, 3, 14, 36, -5, 3, -1, 1, 12, 14, -1, 4, 6, 0, 2, -41, -12, -15, 8, 9, 23, -56, -27, 0, -6, 21, 0, -8, -44, -9, 7, -4, -3, -34, -5, -28, 7, 0, -3, -60, -25, 13, -11, -19, 4, -3, -6, 1, 0, 2, -1, -36, -30, -6, -22, -6, 4, 0, -5, -25, 8, 0, -9, -2, 14, 11, -41, -29, -3, 7, -6, 8, 4, -30, -27, 0, 36, 10, -15, 0, 28, 1, -50, -5, 22, 5, -3, 9, -1, -9, -3, 18, 2, -23, 4, 0, 12, 8, 24, 1, 10, 15, 22, 4, -19, -78, 4, 25, -20, 2, 9, -4, 9, 5, 3, 1, 3, -4, -8, -27, -10, -2, -4, -6, 13, 2, 7, -23, 19, 0, 8, -22, -29, -3, -22, 5, 26, -12, 0, -1, -9, 6, 31, -43, 5, -4, 0, -3, -9, 1, -3, -9, 33, -27, 28, -6, 3, 2, 0, 4, -12, -6, 18, 8, -2, 24, 34, -25, 5, 2, -8, 32, -19, -55, 0, 3, -9, -2, -22, -27, -8, 1, -1, 5, -5, -12, -37, -4, 10, -12, 2, -7, 2, 11, 5, -3, 0, 46, -2, -1, 39, -15, -24, -34, -4, 6, 5, 4, 6, 5, 5, -19, -20, -10, 5, 10, -5, -2, -6, -3, -45, 29, 3, 29, -62, -18, 9, -26, 9, -29, 2, 1, -18, -14, -12, -10, 0, -2, 28, -6, -2, 12, 7, -27, -4, 0, 6, -29, 13, 45, -6, -27, 0, -9, -5, 26, 24, 4, 3, 19, 9, -18, -37, 8, -5, 35, -10, -36, -33, -7, -20, 9, -9, 4, 5, -3, 22, -31, 7, -46, 3, -1, 6, -12, -46, 4, -71, -5, -2, -11, 5, -15, 1, 3, 7, 20, -15, 9, 8, 3, 7, 0, -7, 9, 0, -64, 20, -7, 7, 4, 0, -29, 14, -35, 23, 0, -2, -2, 23, -9, -6, -15, 16, -8, -4, -18, 21, -1, 15, -9, -7, -10, 1, -11, -5, 1, 7, 2, 3, 2, -2, 3, -14, -25, -8, -6, -5, 21, 9, -27, 12, 12, 8, -5, 7, -6, 10, 3, -2, 13, 9, -5, 1, -48, -6, 1, -10, -22, 25, -3, -6, 3, -108, -6, -11, -2, 16, -5, -5, -2, 44, 14, -2, -29, -2, 26, 57, -7, 11, 2, -24, 8, -1, 34, -9, 1, 12, -3, -9, 1, 4, 7, -27, 6, 18, -8, -67, -5, 1, -24, 25, -1, 7, 0, 8, 6, 40, 3, 7, 4, -2, -17, 4, 6, -1, 8, -29, 7, -11, 6, 4, -5, 0, -30, -4, 7, 5, 6, -5, -5, 2, -9, -46, 17, 2, -2, 26, -4, -1, -5, -28, 13, 3, -7, 19, 39, 23, 0, 0, -36, 8, -1, -6, -11, -9, 4, 4, -2, 10, -5, 4, -5, -9, -3, -6, 2, 8, 7, 2, 3, -5, -2, -11, -6, 4, 0, -8, -7, 5, 0, -7, -4, -8, -27, 3, 7, 5, 3, 0, 7, -9, -9, 28, -2, -20, 14, -9, 4, 29, -57, 22, -45, -7, 2, -6, 19, -9, -31, 2, -19, -34, 20, 2, 9, -7, 10, -3, -3, -2, -5, -2, -3, -8, -39, 24, 6, 4, 40, -5, -2, -14, -3, 13, 10, -5, -37, -8, 22, 16, 7, -9, 24, 22, -19, -2, 6, 1, -7, 0, -5, 8, 6, -1, 22, -30, -8, 17, 2, 38, 4, 4, -16, 9, 8, -12, 5, -34, -15, 27, -21, 0, 7, 7, 0, -39, 6, -18, -2, 32, -1, 10, -46, 22, -3, -32, 24, 15, 0, 0, 1, -4, -1, -8, 12, -1, -32, 4, -8, -19, 1, 45, 0, 3, 8, -18, 31, -30, -47, -7, 15, 13, -18, 5, 2, 16, -9, -2, 4, 6, 2, 20, 11, -11, 6, -9, 28, -19, -14, 0, -28, 34, 0, -4, 0, -12, 0, 30, 0, 3, -12, 8, -3, 7, 0, 28, -45, -4, -30, -8, 3, -6, -6, 2, 7, 13, 45, -44, 4, 15, 6, 14, -4, -17, -8, -23, 3, -8, 2, -46, 5, 3, 7, 0, -6, 29, 11, -14, 2, -1, -7, 0, 7, -19, 5, -3, -4, -10, -3, 1, -53, -2, -33, -4, 7, -3, -19, 3, 6, 30, -41, 0, 10, -3, 26, -27, -50, -29, -70, -4, -6, -1, -6, -1, -15, 11, -4, 13, -7, -2, -9, -7, -3, 2, 18, -32, 16, 6, 10, -50, -1, -10, 0, 7, 0, 14, 22, 5, 20, 10, -2, 3, -2, 7, 3, -3, 1, -11, 7, 21, 6, 25, 33, 0, -12, 16, -7, 6, -37, -50, -8, 32, 13, 4, -6, 12, 0, -1, -18, -7, -3, -42, 6, 30, 10, -4, -4, -2, 1, 13, -46, 9, -57, -4, -23, -1, 14, -1, 0, -26, 35, -1, 7, -33, 9, 2, 6, 0, -12, -5, -17, 1, 18, 0, 1, 5, -37, 8, -5, 47, -2, -13, 8, -5, 12, -20, -32, -6, -3, 8, 14, 13, 0, 7, -3, -7, -9, 25, -33, -1, -4, 19, -2, -2, 4, -1, -2, 4, 6, 44, 1, -2, 6, 20, -3, -3, -5, 7, -3, 0, 21, -4, 37, -22, 14, 9, 2, -42, -1, -27, 25, -4, 10, 17, 0, -5, -29, 13, 4, -15, -4, -32, -8, -76, -3, -10, -4, -3, -1, -18, 8, -21, 10, -17, 1, 43, 15, 3, 56, -19, 4, 35, -2, -8, 14, -28, 1, -8, 2, 16, -34, 2, -8, -8, 1, -9, 6, 9, 6, -18, -6, 3, -30, 21, -8, 8, 0, -32, -40, 6, 0, -4, -6, 0, -25, -34, 3, -2, 16, 0, 1, -2, -7, 9, 3, -9, 19, 8, 1, -3, 5, 2, -5, -3, -2, -18, 41, -9, 2, 3, 37, 5, -7, -15, -9, 4, 4, 17, 13, 22, -2, -11, 0, 2, 39, -4, 31, -25, -21, -16, -2, 3, 5, -1, -8, 0, 7, -9, 6, 5, -5, -1, 6, -5, 22, -1, -3, 5, 6, -48, 0, 1, -18, 0, 0, 20, -23, -13, -23, 1, -5, -4, -28, -23, 0, -10, 0, 17, -6, -9, -3, -6, 0, -5, 7, 1, 4, -45, -15, -10, -12, -5, 29, -30, 1, -6, 4, -3, 19, 7, -7, 0, -13, 4, 2, -9, -4, 27, -49, -2, 23, 3, -3, -15, -22, 31, 5, 0, 19, -3, -17, 23, -6, -12, 4, 24, -3, -9, -1, -8, -3, 0, 1, 0, 4, 2, 14, -23, -2, 24, 0, -15, -9, 0, 24, 4, 6, 6, 4, -57, -7, 0, 4, -17, 2, -4, 9, 30, 9, 24, 6, -5, 35, -26, -19, 0, -2, -1, -43, -24, -3, 1, -2, 5, 7, 3, -19, -5, -41, -5, 0, 26, 17, -11, 5, -2, -6, -24, 24, 8, 6, 8, -16, -1, -6, 0, -6, 1, -4, 6, 0, -5, 0, 30, 21, 26, -12, 10, 35, -2, -15, 4, 18, -1, -8, 6, 5, 0, -6, 11, -7, -16, -26, 4, -7, -6, 1, 14, -2, 19, -1, 6, 8, 0, -5, -2, -29, -21, 21, 11, -13, -27, -6, 0, 0, 7, -12, -60, 2, 2, 21, -6, -8, 17, -4, 1, 0, 38, -27, 9, 7, 2, -7, 7, 13, -15, 3, -2, -14, -39, 13, 32, 25, -3, 1, -2, 16, -6, -42, 0, -13, -7, -9, 3, 4, 21, 16, -17, 20, -20, 0, -2, -14, -1, 4, 2, 33, -20, -6, 10, 9, 3, -36, -5, -2, 4, 17, 23, -11, -9, 20, 13, 27, 1, 18, 10, 6, -1, -14, -21, -45, -18, 12, 19, 25, -4, -8, -4, 18, -6, 1, 7, 16, 16, -18, -19, 19, -24, -4, 2, 5, -11, 0, -50, -19, 8, 23, -10, 5, 9, -15, -3, -46, 16, 7, 0, 16, 6, 29, 29, -9, 18, 1, 16, -20, 1, 32, 7, -35, -6, 0, 4, 15, 8, 4, 0, 17, 36, -4, -3, 5, 33, 31, -9, -42, 1, -3, 6, -25, -10, 10, -20, -4, 7, 1, 6, -3, -9, -8, 15, 4, -5, 14, 16, 4, 0, 12, -5, -6, 0, 0, 11, -5, 10, -3, -39, -5, -7, 0, -7, 0, 0, -4, -2, 11, -39, 9, -2, 30, -2, -4, 0, -19, 8, -35, -1, 6, 3, 14, 17, -2, -11, 14, -1, 21, -35, -6, 0, -22, -6, 0, -31, -9, 2, -9, -21, -4, -31, -2, -36, 2, 18, 17, 6, 9, 7, 18, 3, -7, -10, -15, -7, -8, -16, 0, 14, 36, 20, -26, 52, 9, 36, 2, 33, 9, -2, 0, -5, -9, 0, -7, -26, 2, 7, -1, 27, 18, 5, -4, 12, -12, -40, 4, -5, 17, -4, -4, -26, 7, 4, -3, 20, -1, 5, -8, 6, -4, 0, 2, 9, -4, -3, 4, 1, -4, 0, -7, 1, 23, -2, 8, 12, -11, -4, -10, -2, 2, 0, -2, -17, -4, 4, -15, -8, 9, -4, -5, 4, -38, -26, -1, -3, -1, 37, 0, 29, -9, -8, -4, 5, 7, 23, 10, 0, 4, -3, -1, 12, 7, -2, -15, -15, 1, 32, -39, 2, -2, -16, -9, -5, 1, -2, 3, -5, 31, 32, -6, 24, -8, 15, -13, 6, -9, 23, -52, 27, -24, 5, 0, -44, 18, -3, -7, 6, -19, -32, 4, 0, 8, -7, 0, 4, 37, -42, -3, 0, -2, 32, 0, -1, 12, -3, -7, 5, 6, 30, 8, 19, 4, -6, 3, -35, 28, -46, 6, -12, 9, 2, 3, -7, -43, -2, -6, 3, -1, -3, 11, 2, -67, 28, -9, 21, 7, -12, -1, 4, 0, -6, -6, -4, -1, 69, 2, 19, -12, 2, -2, -2, 3, 5, -4, 12, 1, -12, -6, -8, 34, -24, -13, -16, -26, 21, -5, 8, -4, 0, 0, 5, 5, -11, 0, 1, -4, 5, 20, -32, 3, 9, -5, 1, -29, -45, -59, -3, 25, 3, -23, -4, 0, -27, -12, -4, -6, -12, 7, 7, -30, -38, 6, -6, -14, 6, 3, 4, 37, -19, -5, 5, 30, -8, 0, 4, -4, -24, 7, -4, 2, -30, 7, 69, -52, 23, 35, -14, -1, -7, 6, 22, -46, 0, 8, 20, -18, -15, 5, -2, 3, -15, -17, -22, 6, -4, 8, -10, -59, 7, -1, 10, 0, -35, -42, -8, -15, 5, -12, -31, 24, -6, 0, 4, 13, 4, -13, -17, 12, 11, -11, 1, -7, 6, -12, -3, -7, -34, 39, 0, 10, -49, -35, 4, -88, -25, -11, -3, -9, -4, 8, 1, -13, 6, 0, -3, -2, -2, -46, 4, 6, 17, -6, -22, -31, 12, -49, 9, 6, 0, 21, -11, 9, -27, -12, -15, -9, 5, 20, 51, 17, 6, -7, 7, -16, 4, 5, -28, 0, -32, 53, 2, -30, -7, 2, 7, -47, 15, 14, -22, 12, 3, 9, 8, 3, -10, -15, -4, -33, -16, 6, -6, 5, 0, 0, 41, 1, 1, 10, -9, -88, 9, 0, 3, 11, 10, -2, -1, 3, -3, 9, 0, 19, 7, 6, -1, 15, 6, -33, 23, -5, 0, 24, 4, -29, 21, -41, -31, -7, 28, 0, 4, -20, 0, -10, -24, -5, -17, 12, -31, 1, -1, -5, 23, -2, 13, -8, 6, -10, 6, 2, -39, 4, 6, -11, 2, 8, -5, -2, 6, 22, -49, -7, -3, -34, -1, -8, -2, 10, 2, -8, 2, -44, 0, -12, 25, 0, 18, -17, 6, 36, 0, -1, 0, 17, 24, 5, -11, 29, 8, -22, -7, 1, -56, 7, -9, -4, -8, -10, 10, 3, 19, 18, -12, -36, -3, -3, 5, 7, -24, 6, 41, -24, 20, 13, -15, 2, -7, -5, -4, -11, -5, -3, -6, -2, 0, -3, -36, 5, 0, -44, 21, 18, -7, 0, -33, 0, -36, 5, -5, 16, 0, 15, -8, -11, 5, -22, -26, 26, 7, -7, -3, -1, -17, 8, 2, -8, 3, 0, -2, -1, -17, 0, 4, 18, -7, 6, -11, -4, 14, 6, -12, -16, 1, 7, 6, 17, 4, -22, -3, 19, 0, -9, 6, -73, -1, -8, -9, 4, 0, 17, -12, -7, 0, 4, 0, 0, 28, -7, 0, 5, -2, 21, -11, -2, -6, 4, 28, 8, 9, 12, 4, 2, 22, -49, -3, 2, -1, -8, -7, 35, 3, -7, -5, -19, 24, 21, 4, -2, 25, -10, 5, 1, -7, 8, -48, -34, -11, -24, 3, 15, -24, 7, -5, 2, -7, 16, -4, 23, -21, 7, -11, -8, -12, 7, -6, 15, -7, -15, 1, 1, 3, 36, 9, 0, 2, 19, -23, 18, 4, -1, -36, 26, 9, 5, -5, -11, -5, 4, -9, 6, 9, 4, 0, -17, -39, 3, -34, -5, -12, -9, 3, 16, 13, -6, 2, 2, -54, -11, 6, -4, -18, 1, -4, 0, -30, -2, 14, -5, 2, -39, -43, -5, -16, 0, -9, -21, 45, -3, -5, -23, 1, 1, 9, 3, -1, 15, 7, 4, 14, 35, 18, 0, -25, 23, -30, 23, -12, 3, 12, -7, 8, -1, -1, -2, -1, 0, -10, -10, 3, -7, -10, 8, -8, 27, -5, -5, -8, 1, 5, 19, -5, 4, 9, -1, -18, -8, 25, -2, -17, 26, 7, 7, -3, -3, 33, -1, 14, -9, -39, -5, -1, -9, -12, -26, 13, 28, -2, 9, -26, -3, -14, 3, -23, 10, -32, 0, 4, -11, -11, -1, -17, -4, 7, 11, -31, 9, -13, 28, -4, -11, -19, -21, -19, -13, 4, 8, -99, 20, -36, 21, -1, 0, -9, 10, 7, -9, 0, 0, 6, -28, -7, 6, 14, 14, -61, -57, 0, 0, -2, -7, 2, 6, 4, 28, 23, 0, -18, 10, 1, -16, 6, -10, 2, -10, 15, 27, 31, -57, -20, 27, -1, 0, -12, 4, 24, -8, -4, -20, -21, -1, -51, 5, -5, -5, 5, 5, 0, 8, -26, -5, 4, -13, -1, -10, -3, -1, 0, 5, -18, 32, -41, 3, 6, -15, 1, -6, 7, -26, 0, -6, -64, -3, 7, 2, 1, 21, -14, 2, -24, 8, 12, -38, -7, -18, 19, -20, -22, -3, 25, 6, 9, -7, 26, -3, 35, 4, -1, 3, -34, -5, 1, -11, -3, 21, 1, 7, -21, -13, 5, -1, 1, 7, 3, -28, 33, 23, -16, -5, -12, 12, -17, 6, -5, -3, 28, -6, 20, -2, 2, -5, 1, 0, -54, -5, -4, -4, 3, 6, 20, -1, -4, -23, 1, -4, 12, -45, -4, -17, 4, 2, -5, -34, 32, 12, -10, 7, -24, -6, -10, -12, -9, -19, 6, -4, 2, 17, 11, 3, -59, 6, 8, -36, -15, -4, -19, -7, -4, -1, -24, -7, -31, 3, -11, 9, -7, -13, -6, 9, 54, -7, -4, 3, 0, -20, -12, -8, -2, -2, 0, -51, 24, 2, -11, -8, 28, -2, -26, 7, 0, 7, -7, 19, 8, 17, -5, 0, -8, 23, -11, 2, 7, 6, -1, -46, 7, -3, -13, -11, -45, 18, 0, 6, -5, 7, -6, 12, 0, -9, -5, -2, -10, -2, -19, -4, 27, -1, -4, 1, 27, -2, -2, -5, -5, 34, 2, 0, -10, -1, -5, -20, 7, -1, 8, -12, -7, -22, -14, 0, 3, -3, -7, -10, -54, -8, 2, 9, 1, 0, 20, -2, -8, 6, 1, 36, 24, -9, 4, 13,
    -- layer=3 filter=0 channel=6
    -4, -3, -2, 7, 0, -4, -1, 30, 16, 7, 3, -6, 0, 23, 22, 1, -51, 25, 8, -29, -5, -6, -3, -43, -9, -43, 6, 7, -14, -24, 25, -31, 4, 13, -7, -2, -2, 3, 1, -23, 5, -34, 13, 9, -17, 0, -24, 20, -21, -60, 0, -7, -7, -8, -59, -11, -1, 0, 3, -23, 9, -3, 0, 3, -29, -20, 11, 47, -18, -13, 5, -3, -2, -3, 5, 6, 1, -4, 0, 7, -16, -8, 29, -1, -3, 11, -14, 1, 2, -3, -7, 3, 11, -4, -44, 6, 0, 0, -2, 5, -23, -1, -21, -11, -27, 11, 4, 8, -5, 18, -4, 1, -5, -27, 2, -3, 6, -12, 4, -4, 1, 0, 16, 13, 1, 7, -59, -8, -26, 30, 7, 18, -14, 24, -8, 28, -5, -6, 19, -19, 7, 6, -2, -10, -8, 32, 12, 17, 0, 13, 1, -6, -7, -39, -12, -9, -3, 16, -10, -5, -25, -5, -4, -20, 6, -2, -30, -3, 38, -5, -12, 56, 18, 4, 0, 5, -28, 0, -7, 40, -41, -5, -1, -5, -7, 5, -1, 28, -23, 6, -1, 9, 9, -28, 18, 8, 15, 24, 30, -14, 5, 4, 6, 5, -57, -19, 0, 10, -8, 35, 20, 48, 14, -29, 0, 36, -7, -29, -13, -23, 8, 0, -8, 15, 9, 2, 15, 3, -36, 16, 9, 18, 0, -6, -1, 1, 7, -9, -28, 0, -26, 5, 7, 14, 0, -2, -59, -28, -61, -28, -3, 21, 16, -2, 1, 15, 30, -1, 14, 22, -7, 19, -12, -1, 3, -28, 3, 12, 3, 24, 2, 6, 0, -6, -7, 16, -6, 23, -14, -10, 3, -63, -5, -28, 26, -21, -1, -34, -11, -15, 0, 31, -9, 26, 0, 7, -12, 17, 0, -16, 0, 9, -2, 4, -8, -33, 1, 0, -29, -8, -17, -19, 6, 30, -11, -3, -27, 29, -3, 0, 7, 26, -8, 11, 4, -16, 7, 18, -2, -38, -33, -26, 6, -9, -1, -1, -9, 12, 3, 18, -16, -4, -2, 2, -15, 0, -3, -17, -21, -11, -2, -12, -8, -8, -6, -4, -64, 7, 0, 0, 5, 4, 27, 6, 3, 0, -30, 7, 0, -18, 6, -1, 0, 0, 3, -19, 12, -12, 0, -2, 20, -8, 39, 31, 0, -23, 1, -4, -6, -10, -9, 10, -21, -46, -20, 8, -2, -6, -23, 0, 37, 6, 15, -13, 5, -10, 22, -6, -32, -56, 6, -10, 26, -2, -10, 0, -14, 1, 18, -26, -14, 4, -18, -57, -5, -9, -3, -7, 62, -1, 19, -3, 24, 7, 5, 27, -41, -20, 1, -7, 8, -16, 12, 8, -7, 3, 0, -30, -9, 1, 0, 11, 13, 27, 13, -6, 0, -9, -7, -1, 4, 1, 6, -8, 4, 0, -52, -7, -30, 8, 5, -6, 48, 13, -3, -6, 29, -11, 4, 5, -7, 5, 51, 33, 3, 0, 2, 23, -6, 23, 18, -8, -2, 1, -22, -40, -10, -10, 4, 1, -10, 0, -4, 0, -7, -1, -2, -6, 30, 4, 2, -34, -1, 2, -10, -36, -7, 5, 23, -10, -61, 5, -3, 2, -6, -16, 49, 2, -11, 2, 8, -1, 0, -2, 0, -26, 48, -11, -2, 2, 7, -9, 26, -22, -1, 6, -17, -13, -1, 3, 4, 17, 2, -49, -7, 0, -6, 12, 10, 24, -25, -15, -10, -45, -7, 5, 46, 0, -28, -9, 2, 16, 36, 29, -2, 1, -12, 0, -4, 10, -10, -1, -6, 3, 5, -5, 2, 0, 2, 4, -24, -3, -15, 3, 12, -4, 4, -19, -3, -3, 0, 0, -16, 0, -1, -39, -70, 4, 0, -2, 11, 2, -42, 9, 12, 51, 12, 2, -24, 8, -19, -2, -29, 7, 3, 6, -2, -3, -9, -11, 5, 4, 7, -9, -62, -39, -44, 4, 2, -15, 20, -19, -34, 21, 5, 39, -8, 12, -5, 6, -29, -32, -8, -3, -7, 5, 18, 7, 14, -7, -9, -20, 0, -6, -8, 8, 3, -6, 1, -41, -7, 2, 0, -3, 12, 32, 4, 3, 0, -6, 11, 35, -11, -10, 10, 4, 1, 7, -14, 16, 18, 25, -5, -3, 31, 5, -12, 7, -19, 36, -4, -5, 1, 21, -1, 25, -19, 6, 10, 0, -13, 45, 1, -12, -3, -1, -24, -2, 11, -3, -16, 63, 6, -13, 11, -21, -8, 5, -5, -27, -4, 2, -6, -18, 13, 16, -5, 9, 13, 0, -37, 12, 0, -34, -13, 4, -2, -4, 6, -22, 30, 1, 23, -10, 8, 13, 4, -55, 29, -10, 23, -31, 15, -1, -51, 53, 5, -2, 0, -9, -12, 20, -13, 16, 0, -8, -4, -37, -2, 1, 0, 23, 3, 7, -7, -16, 1, 0, 0, 23, 0, 6, -10, 15, -1, -12, 25, -22, 6, -19, -17, -27, 3, -41, 0, -5, -1, 0, -47, 0, 4, 4, 51, -5, -4, -46, -37, -33, 2, 11, 30, -59, 0, 15, -18, -36, -6, 5, -37, -49, -41, -8, -40, -44, 3, 15, 3, -31, -1, 12, -1, -4, 5, -10, -63, 1, -25, -9, -7, -46, 21, 11, -7, 0, -5, 2, 8, 8, 7, -3, -46, -13, 20, -1, -18, -7, 1, -1, -12, 1, 6, -3, 1, 5, -16, 0, -2, -14, 28, -1, -12, 22, 0, -6, 5, 3, -5, -23, -18, -57, -3, 0, -39, 0, -33, -14, 5, -46, 4, 5, 0, 2, -6, -1, 2, -25, 15, -34, -36, -7, 15, -6, -19, -1, -45, -3, 6, -11, -10, 2, -24, -55, -7, 43, -18, 0, 4, -5, 8, -37, 37, -31, -36, 0, -29, 7, -37, 1, 5, -4, -29, 6, -21, 6, -23, 5, -10, -43, -87, 16, 6, -10, 40, -12, -31, 8, 0, -13, 2, -10, 36, -3, 14, -5, 24, 27, -9, 6, -4, 10, -4, -16, -6, -7, -9, -6, 11, 11, 24, 5, -11, 12, -2, -8, 13, -14, -1, 9, 12, -7, -7, -10, 13, -12, -9, -11, 4, 8, -6, -43, 1, 0, 32, 24, -15, 4, 5, 8, -42, -5, -7, 1, -4, -5, -14, 3, 0, -7, 3, -9, 2, 0, 7, -39, 2, -6, 8, -15, 6, -6, 4, -11, -37, 0, 6, 9, 16, -55, 28, 4, 13, 13, 17, -1, 0, 0, 36, -44, 1, -86, 7, 9, -13, -9, -26, -27, 4, -25, -39, -23, -6, 3, 0, -18, 3, -41, 16, 11, 5, -7, -75, 20, 2, 14, -11, -5, -8, -1, -3, 19, -34, 0, 7, 37, 30, 38, 17, -7, -16, 23, 4, -12, -6, 8, -9, -6, 0, 0, -4, -10, 7, -6, 8, -1, -16, 6, 39, -1, -2, 0, -11, 10, 8, 3, -10, -1, -2, 25, 14, 0, -11, -11, 9, 9, 0, 6, 19, -6, -32, -20, -29, 5, -10, 2, -3, -5, 0, -42, 6, 1, 1, 34, 3, 43, 0, -1, -12, -39, -8, 4, 1, -16, 7, -7, -12, 19, -10, 14, -13, 6, 0, 8, -22, -12, -1, -7, -10, -10, -51, 3, 5, 12, 7, -29, -4, -11, 0, -23, -20, -6, -2, -24, -30, 4, 6, 2, 1, 18, -3, -5, -31, -10, -7, -7, -5, 0, 1, 3, 5, 0, 8, 22, -16, -10, 13, -9, -14, -5, -5, 5, -15, -1, 20, 5, -7, 30, 32, -18, 17, -4, 17, -14, -32, -11, -4, 23, 6, -2, -20, -12, 15, -7, -9, -18, 8, 21, 25, 7, 1, 16, -3, 5, -10, 29, 3, -6, -77, -7, -2, 8, -14, -25, 7, -3, -22, 11, 5, 0, 3, 5, 5, 7, 41, -4, -8, 3, -10, -7, 13, -10, -12, -8, 13, 22, 33, 21, 21, -35, -7, -14, 20, -3, 48, 12, 41, 15, -4, -20, 22, -35, 0, 10, 2, 14, 4, -6, 19, 10, 6, 0, 0, -55, 9, 7, -5, 36, 10, 0, -53, -9, 4, 23, -18, -12, 3, -37, -1, -12, 37, -4, -38, 8, 2, -5, 4, -2, 3, 3, -53, 22, 5, -24, 11, 43, -50, -26, 16, 12, -3, 3, -1, -53, -38, -2, -38, -14, 25, -6, -1, 24, 3, 10, -8, -45, -14, -18, 27, -8, 16, 6, -2, -28, 5, -22, 37, 9, 16, 0, -50, 1, -4, -7, -17, -11, 22, 38, -7, 0, -15, -3, -61, 3, 0, -7, 1, 4, 38, 0, 1, 18, 32, 3, 3, 9, -8, -2, -4, -7, 3, -38, -29, -16, 6, 5, -49, 0, -8, -4, -4, 76, -1, 5, 3, -29, -9, -3, 22, -23, 4, -40, -14, 3, -31, 8, -1, 6, -18, 0, -22, -2, -7, 25, 18, 7, 3, 24, 18, -7, -33, -8, 22, 41, 22, -18, -30, -1, -7, 12, -7, -10, 1, 1, -14, -6, 34, -5, 1, -17, 3, 11, 0, 38, 0, -5, 8, 24, 28, -1, 0, -11, -9, 11, 12, 7, 5, 5, -6, 14, -10, 5, 1, -1, -11, -6, 5, 4, -8, 2, 5, -1, 30, -5, -26, -21, -9, 0, 21, 1, -13, -9, 36, 24, 6, 3, -10, 16, -45, 1, 12, 25, 6, -38, -7, 12, 2, -16, -16, 3, 1, -16, -23, -5, 1, 1, -1, 7, 33, -8, -9, 6, 6, -7, -13, 5, 6, -79, 4, 6, -6, 1, -1, 0, -40, 16, 8, 16, 2, 3, 6, 19, 3, -5, -34, -39, -3, -45, 7, 1, 19, -25, 0, -8, -5, 0, -35, -32, -12, -61, -9, 18, -3, 12, -5, 0, -2, 8, 6, -12, -14, 0, 5, 5, -50, 39, -7, 8, -6, -45, 8, 2, -13, 12, -10, 0, 5, -46, 2, 6, -17, 4, -15, 9, 31, 24, -21, 3, -9, 4, -8, -7, -5, -10, -7, -22, 9, 0, 22, 0, 6, -2, 3, 15, -1, -7, -1, -6, 13, 12, -26, 16, -62, 1, -1, -2, 11, 11, -8, -8, 1, 8, -88, -48, -25, 1, -3, 18, -2, -1, 5, -17, 0, 1, -6, -2, -5, 5, 1, -5, -16, 22, 8, -10, -10, -8, -80, 0, 0, -6, 0, -22, -17, 8, 5, -2, 5, 14, -1, -1, 1, -1, -21, 41, -15, 0, 5, -9, -1, 3, -13, -52, 2, 2, 1, 23, 0, 3, -11, 1, -3, 5, 0, 3, -35, -8, -24, -32, -28, 5, 24, 6, -8, -6, -40, -14, -28, 4, -36, 18, -16, 0, 0, -8, -2, 10, -45, -1, -1, -5, -16, -19, 27, 0, 4, 24, -35, -28, -2, -28, -4, 0, 40, 6, -2, -6, -5, 40, -21, 22, 3, 52, -7, 24, -7, -17, 2, 24, -21, -6, 25, -23, 0, -7, -6, 49, 37, -35, -14, -71, 3, 5, -5, 6, -8, 5, 26, -7, 14, -1, -4, 32, -4, -26, -1, -53, -38, 2, 9, 7, -14, 24, 0, -2, 6, 7, 0, -17, 47, 32, -5, -21, 22, -20, 5, 5, -7, -32, 6, -6, -5, -14, -10, -35, -8, -4, 47, -4, 3, 22, -14, -10, -58, -2, 2, 12, 42, -16, 4, 37, 8, -29, -24, 0, -24, 16, 7, -47, -8, -5, 18, -37, -4, -29, 5, 8, -37, 31, 3, -24, -8, 38, -3, 4, -14, 9, 22, 0, -11, 8, 22, 0, 20, 0, 0, 12, -3, 6, 5, -9, 11, 0, -14, 1, -4, -46, -4, 0, -18, 4, 0, -6, 26, 4, -2, 7, -20, 0, -3, 23, -5, -5, -1, -5, -30, 2, -5, 6, 4, -3, 12, 1, 0, -47, 21, 4, 2, 0, -10, -2, -4, -2, 4, -27, -4, -50, -6, -15, 18, -2, 7, 19, 3, -25, -14, -1, 4, -77, 2, -4, -39, -26, -6, -64, -22, -7, -88, -4, -3, -6, 28, 9, -7, 2, -16, 38, -18, 60, 0, 27, -17, -2, 18, 6, -1, -3, 0, -23, -11, 4, 2, -45, -15, -6, -6, 6, 14, -4, 4, -7, 7, -26, -3, -34, 0, -12, -5, 0, 2, -9, 10, 0, -8, 11, 6, -1, 19, -4, 4, -5, 25, -66, 8, 0, -9, -6, -4, 9, -7, 0, 4, -2, 13, 0, -32, -7, 27, 1, -5, 0, 54, -3, -10, -5, -6, 10, -7, 7, -11, 0, 33, -19, 5, -1, 0, 8, 0, -21, -3, -12, 0, 5, 67, 2, -30, 0, -3, -4, 1, 1, -46, 4, 0, 5, 2, 0, 29, -12, -6, 9, 42, 6, 34, 37, 0, 2, -24, -6, -14, 11, 4, -5, -3, 11, -14, -9, -15, 35, -11, 0, 2, 7, -2, -56, 4, -19, 5, -5, 23, -57, -26, -37, -9, 4, 9, 10, 0, 5, -4, 3, -5, -17, 53, -5, 5, -5, 20, -8, 76, 51, 5, -32, 4, -2, 12, 0, 39, 4, 0, -13, 36, 22, 13, -9, -24, 15, 19, -28, -16, 39, -6, 6, 8, -2, -10, -4, -4, 54, -9, 1, -1, 0, -35, -9, -4, 28, 6, -4, 6, 10, 40, -10, 5, 18, -37, 6, 0, -13, -53, 7, 30, -3, 34, 7, -2, -30, 6, -1, -12, 51, -19, 0, -9, -5, 7, 8, -9, 39, 3, 31, 4, 0, -20, -38, -33, -9, 36, -1, -12, -11, 33, 46, -13, 37, -32, 11, -3, 0, -19, 1, -2, -6, 2, 2, -1, 27, 38, -25, 5, -38, 2, 1, -6, 41, -66, -4, 10, -29, 18, -3, 63, 5, 31, 13, -2, 3, -16, 1, -25, 47, 13, 19, 32, 0, 4, -2, 5, 15, -4, -40, -16, -2, 28, -6, -5, -5, -15, 14, -75, 0, -3, -3, 31, 5, -4, -7, 14, -75, 62, -20, 5, -46, -3, 9, -18, 15, -5, -13, 0, -26, -20, -14, 55, 9, -6, 18, -10, 2, 0, 6, -9, -10, 67, -11, 3, -5, 50, 16, -37, 40, -32, 37, -3, 4, -7, -8, -8, -10, -1, 8, 0, -4, 5, 5, 6, 36, 12, 47, 52, 44, 29, 38, 15, -16, -3, 30, 25, 13, 21, 7, -31, 47, -16, -15, -18, -4, 0, -7, 7, 49, -5, 7, 25, 17, 27, -19, 1, 15, 3, -10, 3, 19, 5, -16, 30, -82, -4, 0, 9, -13, 3, -5, -6, 17, 18, -4, -47, 14, -10, 36, -8, -4, 10, -20, -39, -35, -6, 15, 35, -99, 27, 3, 66, -5, -5, 5, 45, 23, -52, -1, -15, -39, -12, -12, 2, -18, -4, 29, 6, -17, 15, 15, -5, 3, -38, -1, 7, -41, -1, -32, 22, -5, 21, -5, 9, -6, -6, 12, -25, -4, 20, 16, -7, -10, 0, -5, 1, -2, -5, -3, -2, 0, -5, -9, -10, -18, -6, -4, 0, 16, -5, 11, 6, -31, 3, -20, 5, 24, -5, -2, 14, -5, -32, -18, -10, 13, -55, -7, -6, 40, 22, 4, -11, -79, -73, 19, -19, -13, -37, 5, -2, -5, 19, -2, 45, -15, -31, -24, 1, -11, 5, 10, 0, -2, -33, 5, -33, -1, 7, -6, 10, 4, -50, -66, -27, -13, 5, 8, -5, -8, 18, -6, -14, 18, 5, -48, -33, 39, -5, -9, -30, -38, -18, 1, 7, 0, 0, 36, -1, 0, -10, 9, 70, -14, 4, 7, 2, 5, 8, -6, 2, 7, -1, 3, -3, -3, 30, -4, 24, 31, -9, 2, -11, -11, -1, 5, -25, -13, 5, 3, 3, 17, 33, 19, -7, -17, -9, -49, -3, 2, 9, -17, -8, 7, 27, 13, -70, 5, -6, 0, -2, -3, -12, 6, -1, 5, -2, 63, -36, -9, -1, -64, 11, 4, 22, 13, -8, 2, 13, 19, 20, 24, 7, -2, -14, 8, -30, -3, -13, -37, -1, 4, -4, 4, -6, -26, 3, 27, -7, 0, -45, -47, -22, -57, -7, 12, 15, -4, 1, -10, 4, -6, -3, -49, 3, 0, 5, -10, -42, -26, 0, 32, -11, 10, -2, 1, -30, -15, 1, 8, -6, 3, 44, 5, 11, 4, -5, -19, -4, 9, -15, 30, -5, -8, 0, -3, 0, -8, -4, 14, -4, -1, -27, 7, -31, -6, -7, -16, -3, -2, -3, 5, 16, 21, -23, -14, -36, -7, -7, -1, 19, 30, 13, -9, 31, 25, -25, 13, -15, -5, 7, -13, 13, 0, 3, -22, 4, 2, -1, 35, 9, 29, -1, -3, 19, 3, 0, -9, 0, -6, -32, -25, 15, 22, -5, -1, -18, -2, -9, -2, 12, -11, 1, -8, 4, 3, 4, 25, 21, 11, 3, -56, -6, 1, 7, -16, -1, -7, -4, -4, 2, -2, -11, 1, 22, 12, 6, 5, -57, -9, -27, 10, 0, -3, -1, -8, -8, -4, 3, -10, 0, 5, -18, 14, -27, 2, 7, 0, -13, 12, -15, 6, -1, -34, -17, -21, -24, -7, 7, -3, 10, -38, -2, 30, -4, -11, -80, 10, 4, 1, -5, -23, -47, 4, 4, 21, 10, -1, -3, -16, -9, -10, 0, -10, -17, -32, -6, 4, 7, -25, -51, 28, 47, 7, -9, 5, 2, 2, 7, -7, 0, -4, 1, 3, -14, 12, -4, -21, -2, 21, 15, 14, 35, -38, -56, 10, 4, -1, 35, -3, -34, 22, -17, 11, -15, -16, -36, -48, 3, 5, 0, -27, 5, 4, -24, 9, 12, -9, -8, -6, -23, -8, 3, -22, 8, -1, -66, -26, 0, 1, 25, -9, -2, -27, -6, -7, 50, -9, -24, 18, -4, 26, -16, 3, 16, 43, -35, -9, -1, 20, 24, -13, -30, 51, -11, -15, -1, -13, 39, 3, 27, -3, 15, 41, -28, -4, -5, -8, -4, -22, 5, -10, -10, 10, 13, -6, 35, 7, 4, -120, -63, -74, -23, -5, -11, -10, 20, -4, 6, 4, 8, 0, 13, 23, 2, 0, 1, 3, -16, 7, 2, 2, 2, 1, 11, 0, 4, 25, -15, -7, -1, -37, -1, -3, 9, -44, 2, -34, 1, -12, 7, 2, 58, 4, 15, -21, 2, 22, 8, -10, -3, 47, -1, -5, -8, -84, -15, 26, 9, -9, -46, 3, -5, 0, 14, -6, 23, -24, -45, 56, -4, -34, -3, 32, 40, -6, 9, -6, 27, 4, 16, -2, -19, -1, 22, -12, 21, -9, 3, 2, -21, 3, 34, 6, -32, -17, -5, -13, -14, -27, -7, 5, 33, -4, 23, -7, 9, -15, 6, -16, -36, -4, 6, -5, -20, -22, -16, -6, -2, 0, -3, 11, -7, 9, 0, -2, -6, 4, 54, 2, -8, -14, 0, 2, -5, -29, -8, 0, -33, -5, -5, 6, -37, 0, 5, -11, 13, -58, 1, 26, -8, -45, -20, 9, -13, -7, -24, -35, -32, -7, -8, -7, -3, 7, 17, 5, -13, -3, -7, 29, -17, 4, -3, -23, -5, 2, 15, 29, 1, -8, 12, -7, 35, -9, -6, 0, 9, -28, -37, -6, 18, -18, -1, -18, -4, -10, -1, 21, 35, -5, -2, -7, -27, 15, -14, -22, 4, -21, 30, 24, 0, -8, -8, -8, 4, 6, -2, -3, 5, -26, 22, 4, 4, -9, -6, -68, -4, -4, 54, -26, 4, 6, -2, -36, 11, 38, -13, -5, -27, -26, -37, 21, 6, -12, 0, -10, 5, -7, 0, -7, 6, 5, 7, 0, 4, -4, 1, -10, 2, -9, 0, -6, 2, 4, -19, 33, -18, -29, 25, -5, -5, -5, 3, -17, -16, 0, -6, 37, -26, 5, -34, 1, -66, 1, 23, 0, -3, -6, -3, -5, -1, -3, -3, -38, 0, 0, -12, -12, 21, 6, 31, 10, -44, 11, 17, -4, -6, -19, -20, 8, 5, 0, -21, 17, 1, -7, 0, -4, -23, -20, -17, -4, 1, -54, -8, -4, -9, 20, 2, 7, -2, -9, 9, -2, 19, 0, 9, -36, 7, 1, -27, 0, -9, -27, 0, -14, -23, -6, 2, -11, -3, 4, -6, -1, -15, 2, 0, 6, -8, -4, -4, -28, -2, 8, 11, -11, -2, 0, 43, -1, 2, 35, 19, 39, 9, 24, 3, -8, 0, -17, 9, -5, -12, -32, 14, 18, -3, 47, -11, -20, -5, 11, -1, -16, 10, -8, -7, -12, 4, 11, -1, 12, -25, -7, -39, -12, -10, 1, 6, 1, -4, -2, -13, -5, 22, 0, -1, 31, 5, 10, -35, 6, 24, 23, 10, -6, -35, -8, 0, -10, 26, 5, 10, 4, 1, 18, -38, -19, -60, -16, -1, -4, 5, -13, 2, -5, -10, 13, -2, 27, 4, -40, -2, -4, 6, 15, 8, 32, 3, 1, -5, 8, 2, 0, 6, -35, -4, 9, 14, 5, 27, 2, -9, -14, -13, 5, 17, 29, -5, 22, 1, -15, 5, -1, 30, 26, 5, -4, -5, 2, -23, -13, 4, -7, -19, -17, 18, -7, 19, 43, -9, -36, -5, -4, -13, -3, 15, -13, 23, -7, 0, -44, 8, -17, -2, 8, 6, 5, 1, -6, 3, 2, 32, 3, 31, -23, -11, -3, -3, 7, -29, 2, -8, 3, -3, 7, -21, -10, 1, 2, -75, 4, 15, -26, 0, -17, -3, 0, -1, -9, 18, 16, -1, 13, -39, 0, -29, -6, 0, -15, -49, 2, 0, 2, -11, -4, -35, -13, -14, -49, 15, 2, -20, -9, 47, 0, -9, -3, 1, 5, -40, 12, 3, 4, -2, 0, 23, 0, 30, 6, -21, -33, 40, -20, -21, -2, 10, -30, 0, -3, -8, -2, 28, 8, -40, 5, 9, -3, -4, -64, -6, 21, 2, 4, 30, -19, 51, -1, 0, 9, -8, -23, 24, 9, -4, -7, -19, -6, 21, 7, -3, 8, -2, -41, 6, -7, 6, 0, -6, 1, -11, -3, -11, -8, 4, -10, 23, -11, -8, -9, 1, -12, -9, -7, 29, 11, -6, 13, -9, -15, -6, 20, 0, -72, -2, 12, -1, -3, 50, -14, -12, -7, -3, -5, 3, 9, -14, 2, -4, -2, 0, -18, -31, -6, -4, 19, 4, 0, -35, 12, 4, 8, 27, -20, -8, -46, 2, -7, 7, 10, -8, 7, -4, -15, -75, -41, -4, -10, 4, 5, 33, -36, -9, 2, -7, -20, 11, -15, 2, -17, -6, 28, 9, 8, -2, -4, -4, -5, -1, 7, -8, 20, -19, -1, -54, 4, 8, 6, 6, 3, -3, -58, 12, -10, -6, -13, -11, 2, 25, 9, -24, -4, -26, -21, 3, 2, -2, 2, -7, -8, 1, -9, -7, 2, 12, 6, 24, -3, -1, 0, -7, 0, -5, -3, -6, 10, -5, 5, -28, 6, -12, -2, 4, 0, 38, 12, -17, -5, -9, -10, 31, 21, 11, 4, -41, -8, 27, 2, 2, -16, -4, 2, -7, -32, -9, 7, 3, -3, -31, 6, -31, -9, 9, 25, 58, 4, 35, -10, 9, 4, -39, 13, -5, 2, 26, -1, -1, 5, 2, 7, 7, -24, 33, -5, 3, 10, 18, 4, -6, 54, 11, -5, -14, -11, -44, 3, -2, 9, -2, 6, -7, -4, -31, 2, -11, -7, -6, -16, -25, -2, 5, 3, 11, 16, -11, -14, -2, 1, -21, -2, -1, -6, -19, -7, 7, -6, -5, 30, -2, -69, -10, 2, 2, 38, -26, 1, -19, 29, 0, -6, 59, -24, 3, -9, 0, -3, -8, 37, -5, 12, -7, -8, -5, -10, 10, -35, 0, -4, 8, 8, -5, 3, 12, 0, -77, -28, 0, 19, 3, -2, 0, 0, -8, 14, 2, 0, 39, -4, -4, 34, 8, -6, -18, 1, 18, -6, -35, 33, -22, 7, -8, -31, 1, 11, -32, -5, -38, -13, -19, -10, 16, -13, 0, 8, 4, -25, 3, 3, -10, -18, -11, -5, -17, 9, -39, 4, -6, 0, 14, 15, 1, 4, 0, -38, 9, -10, 6, -16, -6, 2, -10, 3, -3, 2, 1, 0, -52, 0, 6, 15, -21, -13, -3, -50, -43, -29, 57, -18, -28, 7, 0, -1, 26, 47, 20, 1, 5, 2, -36, 27, -5, 42, -9, -1, 9, -45, -55, 20, 24, -4, -6, -3, -4, 23, 25, -32, -17, 0, -3, -6, 6, 6, 4, 20, 22, -4, 12, -52, -6, -6, 5, 2, -32, 3, -6, -2, -4, -4, -11, 5, -9, 1, -52, -2, 8, -34, -6, -6, 6, -51, -2, -31, 4, -9, 0, 13, 3, 2, 1, 14, 6, 36, 6, 5, 4, -23, -31, -6, -28, -44, -23, -3, -3, -13, 32, 7, 40, 1, -14, 17, -3, -12, 42, 25, 29, 24, -1, -15, 12, -7, -8, -1, -47, 19, -9, -7, -4, 3, -22, -8, -7, 7, 1, 0, -26, 3, -16, 4, -3, 1, -10, -3, 53, -36, 7, -5, 10, -18, 11, 1, 4, -14, -6, -38, 25, 0, 1, 1, -47, -12, -6, -7, 7, 1, 8, -30, 4, 8, -8, 2, -6, -7, -30, -2, -16, -4, -1, -9, 4, 21, 5, 6, 7, -37, -1, -2, 16, 53, -9, 3, -6, 11, -4, 13, -2, -23, -1, -2, -2, -7, 14, 10, -37, 0, 6, -6, 5, -7, 19, 5, -3, 2, 2, -41, 15, 7, -5, 17, 13, -6, -29, -41, -2, 8, 10, -18, 0, 46, 3, 9, -3, -23, 3, -8, 41, 0, 17, 0, -3, -4, -14, -8, 47, -32, -5, -4, -45, -20, -1, -26, 2, 20, 7, 24, 8, 0, 1, 13, 4, -55, -9, 7, -13, -11, 7, 26, -9, 48, 3, 7, -4, -3, -22, 17, 11, 1, 6, -11, 10, 22, 23, 7, 8, 20, -13, 9, -9, -44, 6, 7, 0, 4, 5, -3, 3, 3, -3, -7, 7, 7, 5, 5, -3, -22, -6, 1, 2, -5, -5, 28, -19, 2, 26, 3, 0, -10, 41, 0, -13, -6, 14, 8, 17, 14, 8, 4, 16, 23, -6, 2, 6, 53, 2, 5, 1, -36, -8, -18, -3, -1, 27, -44, 9, -7, -22, -10, -2, -18, 27, -17, -2, 2, -11, 22, -3, -10, 17, 11, -6, -4, -8, 6, 47, -8, 6, 19, -9, -10, 0, 6, -4, 48, -4, 1, -10, -71, 48, -2, -15, 5, -7, -3, -2, 0, -25, 3, -23, -15, 19, -34, 34, -3, -7, -1, 34, 19, -19, -10, -16, 0, 5, 8, -3, 4, -6, -25, 2, -2, 10, -14, -22, 6, -11, -2, 6, 7, -4, -11, 8, 4, -3, -8, -52, 17, 9, -7, -8, -30, 12, 19, 3, 18, -4, -20, 1, -4, -5, 20, -4, 0, 15, 11, -7, 7, 50, -8, 15, -4, -18, -3, -4, 1, -1, 3, 4, 12, -4, 3, 29, 1, -2, 19, 8, -36, -24, 11, -60, -19, -22, 27, 15, 13, 4, 1, 23, 5, -3, -23, -4, 41, -10, -20, -13, 3, -7, 0, 1, -8, -5, 2, -16, -9, -23, 32, 2, 3, 6, 8, 0, 34, -36, 7, -25, -25, 1, -13, 5, -13, -10, 8, 6, -40, 47, -6, -15, 12, 2, -6, -20, 9, 22, 14, 21, -19, -1, 5, 6, -16, 4, -13, -11, 4, -15, 5, -60, 39, -3, -7, 9, 24, 30, -23, -2, 3, 1, 30, 0, -34, 13, -47, -20, -2, -49, -6, -1, 68, -23, -20, -6, 8, -1, 0, 27, 5, -5, 16, 27, -12, 1, 0, 0, 0, 5, 2, -9, 2, -4, 2, -4, 0, 29, 1, 0, -20, -26, -1, -2, 5, 0, -12, 0, -63, -7, -25, -27, -45, -3, -3, -25, -9, 15, 22, -9, -17, 6, 0, -5, 42, 18, -3, 22, -37, -32, -35, -27, -6, -17, -5, -5, -1, -23, -6, 20, -20, -20, 14, 33, -12, -5, -45, 19, -4, 11, -3, -36, 40, -2, -21, -29, -6, -8, 10, -24, -8, -8, -2, 13, -3, -23, 6, -17, -5, 7, -16, 0, -29, -4, 2, -6, 21, 64, 8, -7, 5, -8, -10, 10, 4, 3, 0, -36, 11, 3, -3, 5, 1, -3, -27, -5, 0, 3, 0, 0, 3, -30, -5, -37, 35, 7, 6, 15, 36, 1, 3, -13, -1, 3, 4, 19, 12, -41, 32, 0, -46, 1, 22, -1, -61, 5, -29, -10, -5, 7, -1, -11, -7, -10, 7, -8, 3, 15, -7, -3, -8, -10, -20, -42, 6, -1, -40,
    -- layer=3 filter=0 channel=7
    -9, 4, -16, 24, -1, 0, 49, -37, 12, -12, -1, -5, 0, 11, -22, -5, -36, 19, 0, 6, 0, -3, 10, 32, -11, 49, 4, -4, -16, -15, -14, -32, 4, -18, -19, -10, 0, -11, 8, 6, -9, -17, 11, 3, -5, 0, -9, -3, 20, 3, -5, -27, -4, -7, -3, 15, 54, 0, -2, 22, -40, 11, -12, -2, -7, 27, 14, -11, 4, -16, 9, -3, -1, -7, 1, 4, 7, 18, 27, 5, -7, 6, -13, 9, 5, -23, -20, 5, -4, -1, -3, -16, -2, 0, 36, 0, 6, 2, 8, -5, 21, 1, -4, -17, 27, 13, -17, 12, -3, 14, 13, -2, 3, 31, -2, -9, 5, 23, 0, 5, 3, -9, -40, 24, 15, 6, 11, -13, 4, 6, -16, -8, -11, -7, -17, -9, -6, 0, 6, -1, 6, 0, 2, 0, 3, 0, 20, -34, 2, -20, 6, 2, -6, -10, 0, 0, -3, -5, -9, 2, -25, -1, 18, 21, 2, 0, -2, -7, 51, 30, -16, -26, -13, -5, -10, -8, 62, -21, 17, 0, 16, 12, -21, 2, -1, 6, 21, 19, 12, -3, -4, -1, 12, 12, 15, 7, 1, 24, 7, -2, -1, -48, 4, 5, 27, -20, -10, -2, -8, 7, 26, 11, 4, -3, 2, -33, -2, -34, -4, -7, -15, 0, 23, 22, -6, 0, 3, -4, -39, -10, -21, -48, 0, 2, -6, -12, 0, -49, -28, -8, 33, 6, -1, -16, -8, 23, 33, -8, 59, -3, -12, 8, -18, -18, -1, 0, -26, -10, 30, -35, -1, -43, 10, -6, 12, 4, 6, -6, -6, 8, 0, -6, -9, -16, 29, 43, 6, 11, -41, -2, 2, 18, -17, 1, 12, 8, -5, 1, 9, -6, 4, 26, 7, -21, 5, 1, -25, 16, -5, 2, -11, -1, 28, -49, 9, -5, 10, -30, 6, -19, 24, -46, 23, 0, -3, -2, 30, 23, -18, 4, 3, 28, -30, -11, -6, -24, -6, -22, -2, -16, -17, -7, -37, 0, 10, -3, 4, 51, 8, -19, -34, 3, 1, 0, -5, -2, -2, -7, 0, -7, 29, -4, -14, 0, 3, 0, -13, 7, 1, 0, 1, -3, 2, -9, -7, -11, 3, -4, -9, -36, 2, 0, 1, -4, -2, -5, -31, -59, -1, -10, 16, 6, -34, -14, -7, 23, 23, 6, -9, -10, -25, 1, -4, 56, 5, -19, 25, -2, -59, -5, -7, 0, -5, -4, 13, -1, 11, 6, -12, 0, -3, -17, -12, -5, 19, 7, -42, -15, 13, 18, -23, -7, -11, 0, -9, -6, 2, 4, -4, -8, -12, 0, 1, -13, -3, -3, -26, 10, -3, -1, 6, -21, 12, 0, -3, 5, -3, -63, -40, 2, 0, 0, 16, -10, -23, -4, -7, -4, 0, -19, 3, 2, 1, -2, -7, -2, 29, -6, -18, 0, 9, -1, 15, -6, -7, -5, -44, -9, 9, -4, 0, -22, -46, -19, 5, -8, -6, -6, -1, -8, -12, 35, -4, 7, -1, 2, 11, -11, 4, -5, 6, 5, -21, -1, 4, -10, 0, 26, -43, 3, 4, 12, -4, 5, -10, 18, -5, 0, 16, 0, -8, -23, -7, -5, -1, -1, -23, 4, 59, -35, -5, 36, -1, 4, -27, -24, -12, 45, -11, -3, -36, -14, -31, -25, 4, -38, 4, 19, -3, 2, 0, 20, -5, -3, -21, -8, 6, -22, 11, 32, 3, -50, -3, 46, 4, 1, -28, -18, 0, -5, 0, -52, 4, 17, -32, -3, -1, 2, 3, -39, -5, -27, 2, -2, -12, 3, -5, 5, 5, -61, 0, -3, -2, -8, 13, -12, 0, -27, 4, 1, 5, 0, -31, -12, -32, -7, 14, -1, -3, 0, 8, -11, 22, -9, 0, -15, -18, -17, -8, 13, -5, 17, 4, -10, -2, 13, -4, 5, -1, -48, -4, 5, -7, 1, -12, 0, -6, 8, 0, -26, -51, -29, -27, -29, 2, -7, 2, -6, -6, -9, 36, -21, -4, 0, 2, 3, -17, -38, -36, 17, 5, -8, 6, -3, -4, 25, 20, 6, -7, 13, -9, -2, 17, -8, -55, 18, -2, 0, 20, 3, -10, 2, -14, 2, 7, -9, 5, -1, 0, -23, -23, 26, -5, -11, -35, 4, -9, -4, -9, -25, -20, 7, -3, -31, 0, 34, -1, 2, 4, 36, -24, -27, 8, 21, 7, 0, 4, -1, 0, -1, 0, -59, -6, 21, -23, 13, -3, -12, 8, -8, -3, -39, 4, 0, -11, 26, 1, -10, 15, 13, -21, -2, 27, 33, 11, 3, -6, -2, 3, -23, 10, 0, -38, -3, 8, 18, -2, 11, 18, 41, 48, -4, -33, 1, 17, -12, 3, 7, -15, -3, -30, -24, -25, -17, 25, -3, -20, 20, 3, 2, 1, -46, 5, 7, -5, -14, -40, 24, 3, 41, 16, -2, -7, -11, -7, 8, -33, -26, 0, -12, 20, 0, -5, -44, -3, 1, -20, -1, 4, 9, 4, 4, -35, -1, -37, 4, 32, -18, 0, 0, -41, 15, -27, -47, -6, -32, 5, 4, 16, 5, -2, -3, 12, 30, 0, 19, -1, 11, -4, -30, 0, 22, -18, 12, 34, -7, -19, 17, 0, -1, -4, 9, -14, -10, -2, 4, 4, -3, 0, -13, -1, 2, -20, -33, 7, 0, 6, -7, 11, -9, -4, -6, -4, -5, -64, 10, -1, 25, -10, 5, 17, -23, -3, 0, 1, 8, 1, 18, -16, -24, -2, -22, 41, -6, -8, -4, -1, 30, 24, 0, 0, 14, -7, -4, 23, -10, -11, 6, -15, -1, -21, -5, 41, 6, -6, 8, 15, -2, 23, 28, -4, -17, 7, -3, 11, -2, 9, 2, -13, 41, 13, -9, -55, -9, 18, -23, -3, 20, 0, 3, -17, -7, -9, -3, 0, -10, -7, 25, 16, 61, -4, -4, -44, 7, 14, 0, 1, -6, -4, -24, -28, -2, -14, 0, -44, 21, -10, 6, -8, -2, -18, -29, -3, -3, -7, -7, 3, 4, -7, -10, -16, -11, -1, -4, 31, 46, 2, -1, -14, -4, -8, 0, 11, 26, -28, -5, 0, -26, 1, 25, -14, -55, -8, 39, -16, 6, -13, -21, 20, -3, 6, -4, -2, 3, 39, -5, -3, -7, -8, 10, 1, 1, -3, 37, 1, -1, -5, -26, -4, 7, -5, 41, -23, -48, 6, 2, 3, 0, 7, 6, 17, 5, 19, -36, 0, 1, -17, 28, -20, 60, -7, 0, -7, 10, 0, 17, 9, 49, -39, 33, 0, -10, 0, -14, 4, 17, 1, 2, -12, -21, 25, -9, -22, 8, 0, -20, -1, -5, 10, 4, 13, 5, -6, 52, -16, -28, 0, 1, -25, -37, -11, -52, -2, 34, -3, -3, -9, -5, 6, -1, -7, 11, 33, 4, 6, 5, 13, -2, -6, -17, -12, -6, -10, -10, 18, -2, -5, -27, 14, 4, -7, 1, 7, -33, 16, 1, -4, 21, 2, 4, -11, 14, -30, 47, -24, 4, 3, -24, 8, -5, -9, -6, -4, -37, 0, 6, -17, 33, -8, -6, -71, 19, 7, 0, -47, -48, -11, -59, -1, -11, -4, 2, -22, 12, 1, 5, -2, 7, 6, 25, 28, -32, 4, -2, 11, -5, 4, 0, -17, -9, -3, 26, -29, 0, 0, -3, -9, -12, -4, -8, 0, 0, 16, 6, -21, 5, -4, -9, 5, 4, 25, -10, 14, 16, 40, 3, -7, -9, -7, 2, -14, 6, -24, 4, -5, 7, 1, -33, 11, 4, -1, 16, 25, 12, -10, -26, -1, 5, 21, 9, -8, -1, 0, 30, -6, 9, 7, 55, -3, 19, 5, 5, -5, 8, 2, 6, -6, -38, -5, -19, 23, -55, -27, 5, -8, 21, 0, 0, 2, 10, -2, -40, -2, -8, 13, -4, -5, 15, -10, -30, -24, -23, 33, 2, -18, -30, -11, 33, -8, -4, -1, 5, -21, -14, 15, 15, -10, -25, 40, -6, 4, -5, 4, 6, -10, -7, -4, -35, -4, 28, 17, 12, 25, 3, -6, 18, 19, 0, 45, 23, 7, -10, 36, 2, 2, -11, -3, -23, 15, -1, 41, 10, 2, 3, 30, -4, -42, 49, -4, 16, -5, -14, -33, -14, 24, 4, 8, -28, 10, 0, 6, -1, 24, 1, -43, -30, -3, -5, -6, -11, 0, -60, -8, 3, 17, -14, -4, 0, -11, 4, 6, 13, 5, -4, -31, -8, -13, 3, -11, 6, 8, 5, -29, 2, 9, 1, -1, 8, 0, -3, 0, 1, -4, 10, 4, 0, -24, 0, 0, -1, 25, 0, 4, 13, 0, 2, 3, 10, 8, 0, -32, -41, -1, -33, 16, 1, -47, 1, 0, -10, 3, 3, 7, -24, -48, -5, 0, -14, -19, -36, 10, 0, -36, 2, -39, -6, 14, 12, 68, 0, 11, 1, -30, 3, -4, 36, 6, -5, 23, -5, -17, 36, -6, 3, -20, -2, 24, 8, 21, 1, -1, 0, 7, -8, -36, -8, 1, 14, 4, -3, -4, -22, -6, 5, 23, 4, -12, 0, 0, 0, -7, -41, 19, -3, 5, -6, -6, -13, -44, -7, 0, 4, 13, 2, -6, -3, 2, -7, -4, -5, 10, 1, 5, -13, -5, -6, -12, -32, 4, -3, 49, -8, 8, 1, -21, -49, -46, 10, 3, -18, -5, 0, 2, -28, 10, -15, -18, -4, 2, -11, -8, 0, -4, -6, 0, -7, -16, -4, 5, -6, -4, 16, 23, 0, 2, 12, -7, -3, -28, -31, 5, 0, -35, -4, -32, 4, 4, 8, 5, 9, 19, 0, -42, -62, 0, 3, 2, 0, 25, 12, -28, 28, -1, 5, 9, -14, -37, -23, 4, 42, -27, 15, -5, 2, -3, 9, 7, -18, -16, -7, -12, -8, -2, 21, -34, -31, 6, -38, 1, 3, -13, 37, -6, 9, -8, 9, -8, 37, 19, -2, -17, -20, 31, 6, -7, -9, -6, -1, -5, 3, 3, 7, -5, -20, 14, -11, 35, 3, -22, -7, 10, -43, -13, 4, 3, -8, 38, -4, -77, -11, 21, -8, 0, 8, 15, 10, -54, -7, 31, -29, 20, -27, -7, -4, 5, -41, 18, -6, -5, -6, -8, 2, -1, 15, -7, 28, -3, -8, 14, -10, -26, 0, -16, -4, -5, -1, -35, -6, 0, 13, -24, 0, -1, 8, 37, -11, -10, 12, 5, 6, 6, 2, 0, -3, -5, 3, -2, -5, -6, -36, 8, -2, 1, 31, 22, 0, -28, 11, -39, 14, 2, 0, 10, 6, 21, -3, 38, 48, -34, -9, -7, 1, -8, -20, -3, 0, -11, 8, -7, -8, -15, -3, -6, 31, 0, -5, 9, -14, -4, -11, -10, -1, -1, 1, 60, -15, -11, 7, -5, -3, 4, -12, -24, -5, 0, 9, -16, 49, -42, -28, -14, 29, -7, -23, 6, 37, -15, -5, -16, 35, -2, 3, -5, 18, -4, 19, -24, 9, -7, -4, -9, -7, -6, 0, -3, 2, 7, 1, 7, 2, -3, -19, 35, 32, -5, 6, -18, -5, -46, -5, -4, 43, 2, -6, -4, 10, -83, -22, -4, 16, 29, 9, 13, 0, 0, 26, 1, -3, 6, 34, -16, 48, 8, 1, 16, 0, -2, 6, -7, 18, 10, 43, 6, 19, 8, 12, 4, 5, -7, -3, 20, 4, 27, 19, -2, 26, -7, 2, 4, -9, 26, 17, -6, 19, -56, 0, -27, 6, -11, -41, 0, 2, -18, 0, 16, -7, 19, 13, -7, 9, -19, 15, -7, 28, 6, -2, -18, 5, 0, -4, -19, 11, -3, 11, 29, -1, 9, 7, -3, 6, 0, 2, 0, -1, 11, 6, 30, 22, 7, -3, 3, 4, -36, 1, -3, 2, -1, -1, 25, 0, 6, -3, 1, -5, 4, 9, -8, 1, 3, -63, -1, -38, -16, -51, -7, -4, 18, -1, -6, 1, -6, 6, 17, -7, -1, -10, 49, 7, 0, 33, -50, -3, -38, 3, -1, 2, 22, 4, 9, -3, 5, 2, -10, 8, 27, 8, 0, 11, -22, 6, -34, 5, -59, 10, 17, -2, 4, -2, -7, -19, -40, 12, -1, 5, 34, -2, 1, 5, -24, 54, -7, 5, 24, -18, 3, 10, -53, -20, -11, -2, 0, -1, 0, 20, 29, 0, 1, -5, -9, 20, 29, 5, 5, 4, -3, -11, 3, 0, -7, -5, -2, -10, 18, -4, -23, -8, 0, 4, -35, 3, -3, -1, -15, 4, -4, -1, -56, 12, 0, 17, 14, -13, -1, 18, -2, -9, 2, -58, -16, 10, -52, -11, -13, -5, 8, 3, 0, 7, 39, 10, 0, -9, -8, 53, -7, -9, 0, 0, -103, -10, 12, 9, -1, -3, 64, -8, 7, -30, 0, -6, -6, 21, 30, 0, -63, 42, 54, -43, 0, -9, 19, -1, -28, -11, 4, 8, -40, 30, 32, 55, -5, -25, 24, 5, -5, 0, -4, -56, 0, 12, -7, 0, -18, -7, 31, -48, 19, 1, 8, 15, 0, -3, 21, 58, -30, 0, -3, 39, -8, -46, -3, -7, 0, 41, -25, -54, 4, 15, 1, -8, 0, -13, -9, 3, 5, 5, 17, -4, -46, 1, -13, 1, -10, -9, 0, 10, -14, -6, -21, 13, -37, 17, 12, 2, 0, 3, 24, 33, -55, -4, -27, -7, 11, -40, 33, -3, -48, -87, 4, -13, 0, 8, 1, -3, -5, -44, 0, -48, 0, -6, -13, 39, -50, 6, 14, -12, -17, 26, -39, -24, -7, -63, -1, 8, 4, 1, -3, 30, 7, 2, -14, -3, -36, -30, -1, -7, 4, -6, -2, -6, -2, 20, 3, -5, -17, -1, 6, -10, -11, -6, -35, -54, -9, 0, -19, -5, -31, 5, 0, -23, -32, -9, -2, 0, -32, -48, -13, 0, -48, 9, -14, -5, 4, 6, -8, 2, 28, -3, -7, -14, -12, -15, 2, 1, -7, 44, 7, 43, 6, 9, -3, -1, 45, -14, -11, -7, -9, 2, -15, -64, -14, 9, -34, -1, 5, 31, -1, 1, -18, 5, -4, 25, 0, 7, -73, -6, 29, -1, 11, -38, 7, -7, -7, -2, -9, 32, -39, 9, -6, 6, -8, -6, -9, -74, 3, -53, -16, -57, -40, 22, -37, 35, 4, 46, -75, -2, -34, -2, -16, -2, 10, -14, -11, -19, -9, -5, -10, -40, -6, -7, -37, -7, -41, -75, 9, -24, 10, 1, -3, 17, -72, 1, -21, -25, 4, -5, -11, -16, 6, -32, 5, 50, -19, 3, 93, 2, 0, 16, 35, -4, -13, 18, -2, -17, 3, 11, 4, 41, 1, -29, -97, 9, -5, 3, -45, -20, -15, -9, 33, 30, -33, -1, -17, 28, -6, -14, -18, -17, 13, 36, 19, 0, -40, 7, 0, 11, -28, -7, -34, -2, -13, 2, -40, -1, 1, -17, 26, -1, 7, -11, 6, 5, 5, 2, -42, 2, -1, 12, -2, 7, 4, 2, 0, -21, -22, 6, -7, 34, 5, 2, 7, 20, -4, -17, -28, -32, -8, -16, -28, 6, 29, -19, 7, -24, 21, 4, 7, 24, 6, -2, 12, -10, -16, -15, -48, -3, -20, -6, 14, -1, -42, 1, -38, 14, 15, 45, -13, 20, -2, -23, -26, -9, 3, 5, -9, 25, -1, -29, -30, -4, 26, 34, -43, -1, -2, -1, 43, 0, -10, -4, -38, -12, -2, 2, -4, -5, -8, 0, -44, 20, -28, -1, 7, -1, 3, -32, -34, 1, 8, 10, -40, 22, 10, 0, -3, -10, 7, -19, 5, -4, -1, -5, 3, 1, -15, -9, -61, 19, -4, 3, 1, -14, -9, -7, -29, 22, -8, 0, -15, -46, 17, -17, -3, -35, 6, 10, 2, -4, -1, 14, -3, -3, -61, 14, 12, 8, -6, 6, -7, -11, -22, -5, -1, -1, 0, -40, -40, 3, 8, 17, -43, 2, 26, -17, -3, -2, 11, 13, 28, -11, 0, 1, 8, -23, 23, -1, -24, -38, 16, -86, 0, 7, -15, 10, -37, -2, 2, 0, -56, 35, 34, -19, -1, 7, -4, 4, -1, -6, -6, -10, -1, 39, 52, 3, 3, 13, 16, -47, -6, 4, 6, 34, 2, -4, 28, 30, 4, -6, 8, -14, -33, -24, -16, 5, -18, 48, 7, -15, -5, 44, -4, 3, -17, -10, 0, -3, 6, -56, 17, 4, -18, -1, 10, 0, -4, -5, 9, -2, -1, 0, -26, 36, -6, -16, -28, -10, 0, 4, 35, -8, -42, 0, -9, 11, 26, 12, 13, 4, -40, 15, 18, -4, 4, -10, -1, 5, -4, -32, 5, -59, -1, -9, 6, -5, -37, 3, 7, -1, 4, 38, -15, -50, -10, -22, 3, 0, 4, 0, 0, -3, -1, -4, 4, 4, -26, -21, -17, 14, -3, 6, 0, -5, 0, -13, 0, -4, -5, -22, -39, 4, -15, 0, -10, 17, -9, 2, 32, 8, -20, 12, -1, -30, 1, 1, 2, -6, 28, 8, -21, 3, -4, 2, -9, 0, -4, 2, 0, -10, -2, -8, 6, 30, -24, -37, 9, -4, 4, 13, -8, -58, -1, 18, 0, -7, -37, -40, -3, -5, -2, -42, 34, -26, 0, 25, -6, 27, 3, 21, -6, 19, 0, 0, -60, 0, 7, 0, -66, -22, -9, -7, -40, -3, 2, 3, 0, 10, 2, 0, 11, 2, 21, -2, 3, -22, -5, -16, -14, 0, 14, 11, 0, 23, 2, 1, -11, -25, -18, 3, -9, -29, 47, -18, 10, -15, 0, 6, 8, -3, -3, -52, 0, -9, 2, -21, -19, -50, 1, -29, 30, -3, -3, -17, -41, 12, -2, 14, -8, -21, 8, 4, 5, 25, 0, 8, 3, 0, 33, 7, -7, -47, 8, -7, -19, 2, 29, 0, -2, -46, 18, 0, -4, -11, -24, 4, -7, -6, 14, -33, 20, 1, -7, -8, -2, -19, -12, 3, -7, 0, -5, 32, -42, 1, -19, 6, -13, 5, -10, 47, 0, 2, 24, 6, 19, -8, -17, -5, 4, -7, 45, -7, 9, -35, 18, -1, 0, 0, -105, 3, -1, 11, 1, -6, 1, 5, 6, 1, 5, -6, -2, -63, -9, 4, 0, 7, -5, 16, -26, -20, -1, -24, -35, 1, 19, 0, -1, -19, -3, -6, -4, -11, -40, -9, -48, 12, -16, -45, -68, 16, -17, -20, -5, -9, -41, 2, -6, 3, 12, -38, -29, -37, -1, 7, 60, 4, 23, 1, 6, -41, -49, -16, 5, -10, 8, 3, -26, 1, -2, 6, 2, -1, -7, -3, -62, -43, -3, -17, -8, 45, 2, 0, 3, -33, -23, -10, -5, 14, 1, -13, 10, 4, 0, -19, 16, -10, -29, 8, -6, 1, -10, -28, 0, -3, 4, 2, -6, 0, 0, -1, 39, -5, 1, 2, -20, -2, -13, -4, -13, -18, 2, 2, -39, -17, -2, 29, 10, 7, 0, 7, -5, 3, -20, 48, -4, -6, -4, -59, -10, -7, -4, -6, 2, -3, -43, -9, 1, -7, -10, -13, 21, -4, -2, 4, 37, -8, 11, -19, 5, 0, -14, -1, 2, 19, -2, 0, -5, 7, -12, -7, -15, -3, -23, 85, 12, 2, 21, -28, -39, 63, -2, -5, -41, -15, 36, -5, 1, 41, -6, -18, -2, 3, 0, 42, 1, 11, -5, 3, -2, -9, -14, -1, -14, -24, 5, -11, 5, 0, -34, -34, -32, -3, -3, 31, -4, -46, 28, -5, -13, -19, 15, -2, -4, -36, 0, 6, -6, 0, 1, 9, 0, 12, 7, 0, 5, -1, -28, 6, 2, 36, 5, 3, -4, -9, 35, 1, -70, 27, -66, -7, 4, 9, -21, 6, -20, -3, 17, -40, 6, -30, 30, -2, 17, 0, 7, -8, -6, 14, -5, -5, -4, -15, -5, 23, 9, -6, 44, 30, -31, 6, 20, 0, 59, -41, -20, -13, 4, 17, -21, 7, 3, 0, 20, -28, -6, 0, 5, -8, -5, 20, -29, 20, 3, -38, 0, -4, 3, 30, 22, 4, -3, 0, 26, -5, -66, -6, 29, 0, 4, -2, 24, -3, 0, 16, -14, 28, 27, -13, -7, -4, 5, -5, -42, -40, -7, 4, 2, 8, 1, 0, 19, 31, -8, 0, 0, 36, 1, -22, 0, 1, -18, -52, -4, -17, -14, -13, -7, -16, -8, 35, -12, -9, 8, -1, 85, -15, -9, -10, -6, -17, 0, 23, 2, -1, 10, -3, -18, 32, 2, -7, -15, -50, 25, -19, -52, -18, 5, -11, 1, -7, 6, -9, 42, 4, 24, -3, -1, 15, 5, -11, -2, -2, -31, -14, -10, -6, 35, -42, 7, -19, -19, 4, 25, 22, -22, 5, 15, -4, 10, 5, -11, 1, 4, -15, -1, -5, -58, -15, -9, -10, 7, 22, 52, 7, -1, 7, 30, -16, 13, 44, -6, -24, 29, 30, -10, 39, -4, -16, 2, -7, 31, 0, -3, -7, -18, 0, 8, -46, 14, 10, -2, -3, -6, -26, -20, -20, -5, 43, 3, 7, -46, -12, -13, 0, 18, -14, -13, -30, -1, -58, -8, 42, 9, 17, -23, -48, 1, -1, -23, 15, -5, 14, -23, -15, -14, 4, 17, -2, 10, 7, 0, -4, -16, 1, -13, -3, 4, 2, 7, -1, 33, 6, 1, 2, 2, 5, 18, -5, -1, -21, -6, 9, 10, -26, 2, 7, -2, 5, 4, 57, 5, 17, -1, -17, 17, -7, 26, -14, 5, 0, 9, -7, -4, 28, 14, -9, -7, 14, -35, 9, 2, -5, -27, -21, -47, -1, -27, -1, 24, 14, 33, 7, -9, 20, 6, -92, -65, 3, -20, -9, -14, 20, -16, 2, 30, 3, 55, 40, 40, 0, 3, -4, 27, 0, 6, 1, -19, -25, 7, -24, 12, -20, -6, 3, -57, -9, 1, -2, -4, -13, 0, -5, 32, -1, -9, 1, 19, -12, 21, -1, 1, -9, 2, 0, -2, 5, -6, 7, -6, 11, -8, -4, -3, -5, -8, -5, -6, 49, -12, -2, -20, -9, -5, 5, -40, 6, 0, -1, 1, -8, -2, 8, 2, 12, -2, -24, -13, -8, -52, 9, -6, 7, -1, 2, 3, 5, -6, 4, -9, 0, -7, 38, -21, 3, -5, 20, -9, 0, 29, 20, -5, -2, 17, 25, -32, 6, 3, -8, -12, -54, 3, -7, -45, 28, 23, -8, -5, 5, 7, 17, 14, 30, 4, -8, -82, -7, 13, 14, 2, 2, -28, -22, 1, -1, -9, -11, 3, -9, 34, 2, -13, 9, 20, -26, 0, 4, -9, 0, -9, -8, 18, -20, -3, -7, -6, 44, 16, -25, 2, -6, 1, -64, 5, -5, -18, 20, -7, 14, 4, -3, 4, 0, 2, 33, -15, 8, -54, 1, -17, 0, 1, 0, -13, 0, 3, 8, -29, -24, -44, 31, -44, 0, 3, 3, -50, 13, 0, -7, -9, -1, -37, -27, -7, 10, 7, 19, -20, -1, 3, -45, -1, -8, -4, 5, 2, 5, 3, 0, -13, -98, -28, 0, 17, 2, -34, 7, 19, 56, -7, 3, 4, -15, -3, -2, -3, 23, 3, 3, -6, 0, -38, -13, -9, 21, 0, 43, -13, -12, -13, -41, 27, -1, -14, -9, -40, 1, -23, -3, 32, 28, 4, 7, 24, -1, -9, 39, -3, -16, 28, -2, 3, -5, 17, 11, 10, -24, -10, 6, 9, 4, 5, 1, -5, -3, 0, -9, -7, -4, -20, 3, -18, 3, -21, -13, 39, -34, -9, 6, -7, -3, -12, 27, -15, -4, 2, 5, 38, -4, 24, 28, -3, -3, -2, 24, 0, 21, -6, 7, -43, -6, -8, -8, 9, -20, 5, 42, 16, 9, -4, 0, -1, 1, -8, 40, 28, 3, -41, -3, -5, -31, 6, 7, -44, -33, -30, 25, 18, 22, 7, 44, -5, 5, -25, -4, 7, 19, 11, -4, 6, 4, 13, -7, -5, 3, -6, 19, 5, -4, -6, 34, 30, 12, 6, 17, -17, -5, -8, 25, 8, 0, 19, -2, -3, -13, 45, 13, -10, 42, 1, -3, 24, -7, -26, -5, -5, 9, 1, -5, 11, 11, 21, -5, 2, 0, 42, -7, -33, -19, 22, 47, 0, -6, -14, -32, 12, 4, -14, 11, -1, -8, 7, -38, 5, 18, 6, 16, -39, -22, -1, 7, -14, 3, -3, -17, -17, -32, 57, -5, 8, -5, 22, -7, 8, 2, -12, 1, 12, 36, 9, 4, 13, -2, -25, 4, -7, 1, 5, 3, 24, 1, 2, -13, 34, -2, -6, -39, 1, -3, 10, -24, -3, 31, 11, 37, -5, -10, 2, -6, 0, -36, -2, -32, -31, 6, 1, -36, -28, -8, -87, 7, -24, -20, 36, -1, -10, 2, -55, 6, -41, 3, 30, -18, 6, -26, 27, -10, -10, -22, 1, -8, -8, -4, 18, 12, 2, -36, 23, 1, -1, -3, 7, 2, -1, 4, 22, -9, -18, 6, -4, -31, 0, -3, 15, 19, 2, -3, -79, -58, 41, 0, 6, -3, 3, 18, -2, 2, -4, -2, 16, -39, 6, 4, 1, 1, -13, -22, 8, 0, 0, -6, 7, 11, 1, -8, 22, -29, 0, -4, 33, 40, -19, 1, 7, 6, 1, -1, -54, -5, 3, 31, -6, -5, -4, -1, 7, -25, -8, -15, -29, 7, -42, -48, 3, 0, 2, -6, 7, -2, -21, -10, 2, -4, -7, 6, 2, -3, 0, -4, -44, -5, -11, -34, -7, 4, -17, 9, -23, -1, 3, -8, -1, -45, -12, -8, 17, 16, 18, -25, -12, 0, 10, 4, -47, 33, -6, -3, -55, -25, 45, -58, 5, -21, -31, 0, 0, -3, 6, -5, 9, 54, 35, -8, -9, -10, -27, -42, 9, 2, 3, 9, -3, -1, 34, -36, 0, -6, 3, -4, 10, -46, -7, -7, -17, -3, -8, 0, -7, 32, 0, 7, 0, 5, 3, -1, -3, -30, 2, 3, 49, 7, -16, -2, 6, 30, -9, -3, 0, 3, -10, -24, 9, 20, -30, 1, 6, 3, -10, 30, -57, -10, 6, 4, -8, -59, 0, -1, -26, -6, 0, -7, 5, 7, -2, -2, -5, 0, -4, -28, 5, -6, 11, -26, -49, -6, 11, -13, 24, -10, -10, -42, -13, 32, -46, -10, -1, 1, -11, -6, -11, -9, -1, 0, -14, -12, -9, -11, 9, -16, 23, 1, 0, -30, 18, 0, 11, 16, -17, 3, 4, 6, 29, 21, 2, -3, 27, -1, -5, 21, 11, -57, 16, -6, 6, 6, -3, 14, 16, -53, -5, -3, 43, 0, 0, 1, -7, -6, -6, -4, -11, 39, 15, -26, -26, -9, -3, -29, 9, 14, -12, 57, -1, -4, -7, 30, -6, 8, 0, -17, 27, -22, -24, 11, 0, 7, 3, -6, 0, 17, -2, 0, -9, 25, -5, -4, 25, -49, 5, 34, -44, 9, 0, -2, -8, -9, 1, -9, -4, 8, -17, 5, 4, -64, 3, 6, -32, -2, 36, 23, 25, -35, -48, -46, -3, -1, 12, -6, -11, 16, -11, 17, 11, 5, -8, -16, 0, 7, 2, -7, -3, 5, 16, 21, 45, 2, -2, -24, 7, 7, -4, 15, 9, -13, -4, 5, 1, -10, 0, 17, -2, 27, 0, -15, -19, 2, 4, 5, 2, -2, 16, 2, -15, -34, -21, 13, 2, -18, 8, 29, -43, 15, 1, 22, 0, -1, -2, -31, -12, -9, 16, 9, -1, 9, 2, 25, -4, 19, -6, -23, 9, -31, 41, 0, -11, 11, -8, -53, 0, -43, 31, 4, 0, 2, 13, -8, 2, -13, 0, -3, 13, -19, 0, -4, 2, 3, -45, 6, -1, -3, 2, -4, -12, -5, 3, 16, 21, 0, -30, 4, 4, 12, 5, 8, -2, 36, 0, 28, 5, -16, 39, 3, -31, -44, 8, -10, 20, 3, -5, -34, -10, -7, -27, 39, -10, -13, -21, -5, -14, -9, -99, 9, -25, -2, -17, -24, -22, 8, -3, 38, -9, -21, -53, -1, 0, 0, 26, -10, -8, 12, 50, -7, 38, -7, 38, -5, -1, 0, -11, -2, 12, -8, -47, 16, 4, -30, 58, -8, 3, -6, -51, 8, -24, -7, -6, -19, 3, -3, 17, 0, 13, 11, 42, -39, -19, 8, -9, 0, 3, 6, 7, -6, -5, 0, -10, -1, 18, 2, 0, -11, -4, 0, -70, 22, -19, -7, 0, 5, 3, 7, 3, 46, 13, 3, 7, 39, 1, 23, 8, 29, -17, 20, 0, -5, -31, -4, -24, 6, -1, 3, 5, 7, -42, 5, 2, -4, 2, -11, 2, -8, -4, 42,
    -- layer=3 filter=0 channel=8
    -4, -7, 6, -6, 8, -1, 10, -27, 9, 36, -2, -5, -7, -16, -24, 0, -8, 6, -18, -61, -3, -4, -14, 5, 15, 7, 2, -8, 20, 47, -26, 2, -1, 12, 23, -23, 2, 5, 6, 10, -9, 1, 3, -9, 5, 13, 9, -12, 5, 16, 1, 18, -11, 1, 20, 28, 30, 2, -8, 15, 5, -60, -23, 0, -5, -17, -25, 0, 3, -37, -5, -7, 2, 4, -1, -10, 2, -9, 0, 1, 2, -6, -69, -5, -3, -7, -7, -2, 0, 2, -14, 12, 4, 12, 12, 0, -6, 7, 9, 9, -39, 1, 0, 21, 9, 8, 0, 0, 32, 10, 24, -1, -1, 18, 7, 4, 3, -22, -6, -52, 3, 7, -39, 8, 30, 6, 27, -20, 18, -19, 16, 18, -12, 15, -17, 1, 0, 1, -41, -28, -1, -11, -8, 5, -6, 0, 5, -12, 0, 0, -3, -4, 3, 4, 13, -8, -5, 13, -29, 2, 2, -5, -48, -33, 7, -2, -7, 6, 23, 10, 31, -36, 4, -10, -1, 0, 7, -27, -1, 21, 0, 1, -3, 3, 1, 3, 22, -26, 7, -1, -1, 0, -12, 13, 8, -11, -6, 18, 11, 11, -4, -3, 8, -3, 7, 18, -7, -9, 7, -47, 34, 0, -35, 16, -13, -23, 0, 2, -1, -21, -2, 3, 11, -26, 0, -5, 34, -25, 19, -7, -6, -59, 0, 1, 4, -3, -2, 1, 8, -5, 5, -9, -6, 0, -2, -26, 11, 5, -4, -21, 0, -41, -59, -41, -8, 22, -76, 5, -15, -2, -4, 18, 0, -2, 2, 3, 4, -7, 4, -13, -3, 0, -91, 21, 21, -31, 7, 12, -7, -2, 2, 6, -26, -1, 21, -9, 3, 3, 12, -1, 5, -16, -3, -3, -16, 5, -18, 3, 0, -21, 7, -4, -30, -19, -34, 15, 2, 23, 23, 45, 4, -114, 0, 31, -9, -2, 4, -61, -37, 5, 9, -13, -18, -4, 3, -11, -1, -14, 4, -4, 15, 10, -25, 1, 4, -1, -2, 22, 17, 0, -1, -5, 11, -6, -47, 5, -2, -2, 15, -4, -12, -46, -2, 5, -7, 5, 22, 3, -5, 0, -3, -4, 22, 1, 2, 16, -2, -6, 8, 12, -6, -9, -1, 11, 7, -19, -10, 17, 4, -6, 13, 3, -4, -20, 2, -36, -17, 0, -7, 5, -16, -4, 10, -21, -16, 15, -2, -12, 45, 0, 20, 6, -31, -2, -12, -8, 12, -14, 8, -17, -3, -39, -20, -7, -5, -2, 14, -70, -10, -3, -40, -1, -7, -11, -28, -3, -5, 0, -28, -6, -46, -10, -2, 9, 0, 16, 0, 5, 0, -3, 27, -27, -3, -6, 5, -12, 4, -26, -6, -1, 3, -3, 0, 4, -7, -8, 2, -8, 3, -14, 4, -5, 1, -3, 6, -2, 0, 0, -3, -27, 5, 7, 18, 1, 1, -3, -30, -17, -7, 6, -2, -3, -14, 20, -3, -18, 7, 0, -1, 4, -14, 29, -16, 6, -31, 14, 4, 5, -3, 6, -9, 1, 22, 5, 6, 7, 4, 20, 0, -3, 4, -26, -36, 7, 7, 13, 3, -4, 14, 14, 12, 33, 1, -2, 2, -24, 15, 0, -29, -32, -8, 3, -10, 3, -9, 1, 43, -28, -7, 2, 15, 11, -70, -14, -6, 29, -28, -3, 4, -7, -5, -35, -1, -8, -24, -3, 0, -9, 29, -36, 9, 4, 0, 26, -5, -3, 0, 4, 0, -2, -6, 29, -14, -43, -42, 2, 0, -25, -38, -5, 7, -27, 2, 3, 16, 4, -8, 4, 0, 23, -8, 3, -23, -6, -33, -8, 1, 9, -19, -6, -3, 11, -31, -35, -15, -26, 5, -9, 0, 9, 0, 52, -6, -6, 2, 18, 4, -2, -28, -5, 23, -1, -3, 6, 2, 15, -7, 5, 1, -41, 5, -22, 0, 0, -70, -4, -1, 4, 5, -4, 0, 0, -1, -20, -16, 14, -19, 10, 2, -8, 5, -2, -6, -1, -6, 1, -6, 26, 27, 17, 5, 18, -5, -3, -13, -19, 6, -4, -1, 1, -11, 6, -15, -3, -25, -22, -2, -4, -15, 5, -46, 9, 6, 30, 8, -8, -7, -6, 17, 8, -27, -7, -16, -4, -9, -6, -6, -6, 0, 2, 18, -3, -4, -13, 20, -6, 8, -10, -7, 5, -33, -6, 0, 5, -8, 0, 11, 33, -13, -4, -8, -10, -30, 13, -11, 7, -7, -54, -6, 24, -10, 30, -3, 9, -12, -56, 0, -10, 18, -42, 11, -4, 7, -59, 7, -1, -4, 6, 5, 3, -15, -10, 2, 0, -2, 15, -7, 0, 3, -27, 0, -43, -25, 2, -34, 5, 4, -8, -34, -6, 5, 28, 32, -22, -5, -9, 1, 4, -1, 0, 4, -1, -5, -5, -1, -6, -12, -7, -6, -16, 16, -2, 3, -30, 18, -14, -27, 11, -8, 17, 5, -6, 0, 36, -3, -20, 39, -10, -26, 4, 6, -50, -14, -6, 22, -18, -39, 9, -1, -5, 16, 38, 14, -9, 12, 51, 2, -4, 5, -47, -27, -4, -7, 11, 4, -4, -13, -31, 1, 5, 1, -7, -1, -6, -18, 3, 5, -1, -6, -12, 18, 1, 2, -7, -1, 10, -41, 3, -4, 1, 7, 8, -44, -5, 16, 7, 1, 6, 24, -6, -6, -4, 3, 2, 0, 4, 0, -15, -27, 2, -1, -23, 4, -20, 6, 5, -5, -55, 0, 24, 3, -9, 26, 7, 0, 11, -9, 39, -8, -6, 4, 0, -3, 1, -30, 6, -18, 45, -2, -11, -35, -1, -17, -10, -23, -14, -37, 5, 14, -6, -49, 4, 8, -12, -8, 2, 0, 3, 27, -25, 6, -18, -46, 6, 18, -10, 14, 0, 2, -7, -1, -5, -44, 0, -1, -21, -1, -21, -8, -33, -3, 2, 20, -8, -17, 5, 3, 13, -3, -10, -56, -5, 4, -6, -10, -32, -15, -6, -6, 4, -2, -11, -5, -4, -1, -1, -6, 0, -28, 0, 14, -5, 0, 1, 6, 6, 1, 6, -30, 4, -2, 4, -2, 16, -32, -34, 4, -8, 4, -1, -12, -2, 9, 26, -7, 5, -20, -28, 20, -9, -4, 7, 0, -6, -31, 3, 2, -2, 3, -31, 13, 7, -9, 0, -28, -2, 20, -25, -4, -9, -15, -12, 22, 16, 0, 0, -13, 12, 9, 9, -16, 31, -14, 1, 3, -2, -27, 13, 7, -32, 8, 5, 7, 24, -27, 22, 1, 0, -4, 7, 6, -1, 1, -16, 0, 10, -37, 3, 11, -12, -9, -16, 10, 3, -6, 22, -11, -2, -5, 2, -11, 5, -2, 4, -8, -15, -24, 3, -11, -11, -15, -4, 0, -44, 6, -9, 6, -2, 4, -8, 7, 17, -24, 1, 18, -7, -36, -3, -10, 11, -10, 5, -8, -4, -11, -66, 36, 4, -3, -4, -6, 7, -24, -2, -30, -7, 15, 14, 45, -10, -2, -12, 20, -4, -32, 2, 3, 22, 1, 0, 3, 14, 5, -5, 1, 4, 7, 0, -10, 0, 22, -13, 14, -12, -15, 5, 0, 1, -22, 2, -8, -5, -6, -8, -4, -5, 3, 3, 0, 0, -15, -10, -1, -1, 10, -8, 2, -1, -24, -5, 0, 30, 6, 4, 5, -2, -21, -19, 0, 0, -45, -8, -33, -1, 2, -10, 0, 0, 1, 1, 13, -29, -42, 5, 2, -13, -1, 8, -17, -6, 22, -9, 4, 0, -4, -8, 9, 16, 18, -4, -11, -13, -6, -5, -11, 16, -1, 2, -13, 15, -15, -2, -19, 1, 9, -41, -44, 6, 1, 8, 3, 45, -4, -32, -7, 0, -5, 0, 5, 3, -14, 13, 8, 23, 20, 24, 2, -6, -6, -2, 4, -1, -38, -4, 10, 2, -5, 15, 8, -30, 6, -5, 24, 34, -42, -7, -52, -19, 6, 29, -10, 2, -6, 13, -18, -33, 15, -5, -25, 17, -5, -8, 4, 5, 1, -3, -15, -8, 11, 12, -9, 3, 19, 6, -10, -31, -8, -25, 0, -13, -1, 7, -57, 5, -4, -27, -10, -9, 9, -6, 17, 8, 0, -8, 12, -6, 8, 14, -32, 1, 1, -5, 21, 30, -2, -25, -8, 7, -3, -9, -22, 5, -27, -6, 33, 6, -11, -3, -1, -3, 3, 1, 1, -4, 3, 22, -33, -6, 13, -8, -5, 38, 14, 0, 5, -11, -6, 2, -53, 6, 2, 15, 23, -5, -27, -36, 6, -2, -3, -5, 16, 3, -4, 4, 2, -3, -8, -10, -9, 13, -6, 4, -1, 13, -5, -14, 5, -6, -7, 15, 0, 17, -10, -7, -24, -9, 6, -70, -7, -61, 4, -1, 5, 15, -11, -5, 5, 16, -16, 33, -3, -12, 40, -7, -10, -5, 17, -9, -33, 0, 6, 3, -6, 1, 5, 9, -16, -5, 7, -6, 4, -4, -16, -7, 3, 7, 26, 20, -8, -19, -11, 8, -19, 2, -39, -9, -1, 11, -6, 9, -40, 32, -1, 6, -17, -14, -55, 7, -3, -1, -2, 11, 22, -6, 13, -14, -7, 0, 3, -1, -5, 4, -11, 3, 4, -2, 0, 5, 9, 0, -20, -5, -26, -32, -2, 6, 0, -22, 3, 0, -21, -2, 4, -9, 32, 22, -12, -40, 0, 40, 5, -31, -5, -3, -10, 32, -14, -2, -40, 14, 13, -5, 3, 4, -8, 2, 52, 5, -8, -1, -7, 17, -11, -9, 3, 41, 12, 0, -23, 22, -2, -8, -33, -9, -14, 18, 1, 0, -8, -9, 33, -4, -5, 3, -13, -2, 4, 4, -12, -10, 27, -35, 0, -8, 30, 44, -29, -15, -1, -2, 3, -90, 2, 4, -6, 16, 0, 16, 0, -1, -4, 11, 19, -20, -4, -32, 0, 32, -9, 0, 7, -18, 10, -2, -10, 7, 49, -45, -71, -3, 7, -13, -7, -9, 8, -29, -3, -1, -7, 4, 2, 5, 2, 4, -1, 0, 2, 2, -2, 0, -9, 10, 2, 3, 0, -7, -17, -51, 52, 18, 13, -1, 0, 7, 27, 33, -18, 7, 26, -1, -31, 25, 22, -9, 3, 47, 25, -12, 6, -30, -7, 1, -4, 0, -7, -2, -2, 6, -29, 16, 40, 0, -7, 0, 31, 2, -5, -14, 7, 15, -20, -1, 5, -3, -6, -8, -5, 0, -5, -2, 2, 4, 42, -6, 1, -8, -7, 2, 0, 23, 11, 2, 2, -40, -5, -7, -27, -5, 17, 5, 0, 0, -1, 2, -16, -71, -2, 16, -9, -5, -9, 0, 24, -27, -28, 36, 18, 5, -20, -1, 1, -1, 2, -31, -3, -4, 0, 15, -18, -23, -17, -6, 2, 7, -8, -6, -2, 4, -7, -3, 8, 24, -1, 3, -15, 15, -38, 0, 2, -21, -3, -35, 5, -52, -6, -23, 1, 13, -22, -21, -3, -3, 31, -26, -13, -20, -4, -6, 0, 1, 7, -9, 3, 22, -26, -8, -5, 5, 1, 0, 2, 22, 13, -39, 24, -14, -14, 5, -31, -26, -2, -1, -16, 5, 0, -2, -12, -27, 3, -10, -8, 1, -6, -4, 7, 6, 0, 1, -46, -23, -43, 27, 0, -12, -27, -5, -8, -33, -6, -25, 29, 14, -3, 22, 5, 7, -7, -26, 4, -1, -50, -5, -49, 0, 7, -16, 24, -2, -21, -9, -13, 39, -2, 42, -6, -40, 9, -5, 14, 12, -9, 6, 9, -22, -58, -1, 35, -32, -13, 8, 9, -8, -3, 17, -4, -23, 4, 27, -39, -4, -13, -3, 10, 26, 30, 23, -39, 9, -1, -6, -25, 0, -8, -2, -1, 8, -32, -7, -23, -6, 5, -2, 38, 5, -4, 0, 5, 9, -28, -2, -4, 32, -24, -2, -7, 18, 9, -4, -3, 35, 3, -21, -20, -7, 3, -10, 27, -4, -2, 9, 1, -22, 16, -8, 2, 11, -7, 0, -12, -5, 1, 35, -3, -6, -48, -1, -17, -7, -17, 0, 1, 8, 42, 9, -23, 23, 3, 8, 16, -2, 7, 0, 30, -8, 37, -36, -43, 0, -14, 9, -26, 13, 4, -4, 33, 8, -41, -7, -26, 0, -5, -5, -8, -23, -7, -1, -1, -14, -67, -7, -2, -13, 6, 31, -3, -3, 4, 11, 35, -2, 30, 2, -8, 2, -8, -1, 6, 0, -3, -3, 2, -3, -6, -10, -3, 12, 4, 7, 26, -21, -12, 7, -9, 2, 7, -5, -1, 8, -1, -7, -5, -3, 1, 26, -7, 2, 4, -54, -3, 2, 8, 6, 16, -7, -9, -7, -2, -4, 4, -8, 4, 6, -6, -4, 35, -4, -4, -20, 23, 0, 30, 2, 9, 0, -14, 16, -28, 32, 1, 0, 0, -25, -2, -5, -12, -28, 22, 12, -9, 2, -6, -2, 10, -1, -4, 5, -2, 12, 26, 11, -5, 3, -9, -56, 0, -10, 7, 21, -9, -17, -63, -9, 3, 10, -24, 12, -1, 25, 0, 31, -9, 1, -13, -8, 0, -6, -12, -15, 19, -38, -16, 5, -25, -32, 15, -17, -1, -64, -8, 3, 5, -3, 6, 7, 1, -52, 19, 1, 17, 4, 26, 2, 2, 32, -6, -9, 5, 2, 17, -44, 38, 53, -4, 5, 7, 4, 8, 61, 16, -1, 29, -15, -1, -28, -49, -15, 38, -11, 19, -12, 3, -2, -5, 5, 0, 3, 0, 14, -5, -5, -28, 7, 13, -5, 11, 0, 30, -13, 3, 12, -13, 24, 9, 0, -1, 1, -30, 3, -7, -2, 4, -6, 3, 39, 46, 28, -5, -5, -10, -5, -2, -19, 52, 6, 0, -36, 44, -1, 15, 3, -26, 41, -3, -1, -32, -6, -6, 23, 28, 3, -2, -10, -8, -7, 16, -21, -32, 21, -5, -8, -38, 5, -11, 7, -14, -37, 21, -5, 3, 5, 8, -11, 10, -4, 5, 24, -17, 19, 11, -5, -7, -4, 8, 34, 0, -2, 1, -18, -31, -3, -46, 6, 3, -17, 3, -22, 0, -7, -1, 6, -24, -18, 8, -1, 20, -7, 10, -17, 26, -34, 11, 0, -5, 7, -3, 3, 12, -10, 21, 0, -9, 0, 2, 11, -31, -49, 7, 4, 16, -13, -22, -23, -10, 2, -6, 4, 24, 39, 17, -10, 8, -5, 10, 5, 0, -8, -3, -23, 0, -9, 5, -1, 20, 33, -16, -1, 6, -1, -8, 25, 32, 11, 13, 3, 4, -61, -32, -5, -2, 8, -3, 12, 12, -1, -72, 8, 0, 31, 4, 0, -32, -37, -24, 11, -3, -19, -6, -16, 3, 13, -5, 19, -5, 0, -9, -4, -27, 4, 22, 8, 24, 17, -1, 9, -4, -28, 7, -5, 6, -4, 0, 1, -6, 6, -6, 15, 12, 45, -23, 3, -6, -4, -23, 1, -3, -11, -8, -3, -37, -23, 0, -6, -10, -10, -10, 3, 0, 3, -3, -2, -40, 0, -1, -19, -39, 4, 13, 40, 1, -2, -3, 4, -9, -4, 19, -56, -6, -9, 35, 6, 5, -32, 5, -43, 49, -9, -3, 1, -4, 2, 23, 2, 7, 69, 62, -7, 32, 1, -12, 5, 0, -8, -31, -7, -41, -43, 17, -20, -3, -8, 12, -7, -10, 10, 44, 21, 29, -4, -2, 0, -11, 18, 25, -9, -6, -5, -15, -5, 9, 1, 44, -24, 5, 4, -32, 19, -2, -5, 10, -14, 12, 5, -2, -3, 1, -1, 10, -4, -2, -15, 44, 23, -35, 3, 2, 8, -14, -12, 5, 2, 0, -3, -3, -5, -39, 4, 43, -7, -1, 0, 6, 19, 1, 8, -27, -23, -3, 6, -48, 36, -20, -13, 1, 4, -1, -7, -6, 12, 19, -7, -3, 6, 21, 9, 28, -1, 3, -3, 5, -6, 29, 3, 3, -5, 3, 16, 41, -8, 2, 2, -17, -2, -18, -14, -6, -6, 14, 4, 10, 33, 6, -5, -2, 32, -15, -1, 25, 25, -10, 30, -5, -2, 2, 31, 24, -28, -7, 5, -16, 28, -6, 8, 2, -22, 10, -8, -3, 0, -6, 29, -1, 45, -102, -8, 1, -3, -37, -23, -19, 16, 5, 19, 2, -3, 19, 12, -10, -8, -3, 27, 26, -45, 1, 4, -21, -3, 6, 24, -4, -54, -6, 1, -1, -5, 6, -8, 0, -62, 4, -2, 18, -8, 19, -3, 4, 41, 8, -4, 1, 2, -21, -65, 46, 2, -20, -9, 7, 0, -16, -3, 3, -3, 50, -14, -5, 2, -68, -15, 26, 3, 10, 1, -3, 14, -10, 3, 0, -38, -7, 18, -2, 2, -36, 2, 9, 0, 24, -12, 44, -1, -18, 23, 0, 21, 4, -6, 1, 1, 1, -8, 3, -1, -5, 6, -4, -7, 10, 17, -6, -49, -2, -12, -2, -22, -11, -1, -1, 24, 3, 4, 13, -5, 3, 56, -3, 0, -43, 6, -6, -3, -1, 6, -15, 4, -10, 3, 45, 5, -30, 20, 17, -10, -24, 4, 5, 1, -5, -18, -19, -5, 2, 7, 39, 24, 8, -9, -6, 0, -30, 30, 18, 1, 4, -4, 18, 59, -10, -2, 5, 8, -46, -23, -55, -3, 1, -26, -8, 10, -5, 39, -3, 9, -69, 25, 1, -17, -5, -7, 50, 8, 18, -20, -3, -10, 5, 6, 3, -18, 1, 2, 12, 0, 3, 26, 1, 0, 10, -21, 38, 46, 17, -32, 11, 0, -4, 22, -17, 6, 7, -36, 41, 19, -4, -7, -24, -18, -7, 0, 3, 32, -1, -5, -31, 4, 2, 33, 4, 22, -14, 5, -5, 18, 0, 43, -26, 16, -5, -23, -32, -2, -3, -8, 3, -12, -2, 5, -43, 0, 7, 6, 24, -3, 14, 4, -52, -15, 0, -18, -12, -7, 17, -44, 16, -11, 3, -6, 18, -9, -6, -3, 2, -23, 12, 20, -1, -19, -10, -8, 0, 40, 17, -15, -2, -4, 21, 4, -2, 16, -11, 22, 51, 2, 6, -4, -52, -4, -6, 6, -27, -3, -15, 7, 6, -6, -6, 3, -4, -8, -2, -9, -8, -5, 1, 7, 0, -6, -13, -8, -3, -13, 0, -8, -3, 0, -3, -44, -6, -18, -4, -8, -29, -2, 14, -11, 0, -20, -26, 6, 3, 13, -9, -2, 3, -14, -3, 37, 33, -1, 27, 7, 4, 0, 41, -3, 24, 0, -21, -23, 23, 0, 0, -32, -37, 2, -21, -6, 56, -49, 22, 50, 15, -1, -9, 32, 13, 2, 1, 2, -35, 5, -18, -5, 41, -8, 2, -8, -9, 11, -7, -8, -34, -53, -24, 0, -6, 1, -2, -21, 24, 7, 0, -1, -24, 8, 30, 6, -6, 0, -2, -41, 4, 3, 5, 2, -7, -14, 28, 6, -9, -14, 7, -4, -21, -30, 6, 0, 33, -16, -8, -1, 0, 9, -36, -52, -1, 16, 0, -62, -12, -13, 30, 5, -7, 6, -15, 9, 0, -5, -5, 3, -1, 8, 23, 7, -9, 0, -3, 37, -39, 9, -2, 35, 30, 7, -29, 20, 3, -5, -6, 16, -11, -62, -7, -2, -12, -16, 9, -1, -15, -31, 15, 0, -9, -6, 21, 3, 15, -87, -8, -10, 49, -16, -62, -30, -4, -29, -51, -29, -7, -11, 0, 5, 3, 2, -31, -2, -9, -9, 2, 55, 1, -40, -6, 23, 4, 0, -5, 4, 33, -1, -7, -56, -27, 17, -47, -10, 9, 3, -56, -33, -8, 44, -2, 0, 7, -7, 4, -4, 1, -27, 11, 5, 17, 7, 18, -7, 6, -43, -7, -12, 6, 8, 25, -8, 67, 14, -15, 1, 8, -12, -18, -4, -31, 1, -12, -60, -47, -18, -16, -7, 9, -49, 10, -3, 0, -19, 2, 0, -10, -4, 4, 17, 1, -2, -17, 9, -26, 0, -28, 7, -22, 8, 7, -7, -14, -67, 2, 0, 5, -14, -24, -36, 4, -13, -8, 4, 41, -65, 22, -14, -2, -3, 8, -2, 4, 21, -39, -3, 2, 27, 4, -5, 18, 0, -3, 75, -6, -3, 30, 0, -51, -31, -21, 1, -42, -11, 8, -4, -38, -37, -34, 11, -28, -8, -50, -4, 1, 9, -7, -13, -36, -3, 1, -54, 23, -9, -37, -5, 0, -19, -30, 13, 22, -77, -8, 3, 3, -53, -10, -7, -14, 31, -48, -13, -32, -38, 15, -52, -2, -19, 7, -32, 6, 15, -1, -36, -6, 3, -35, 0, -6, 7, 26, -7, -6, -2, 0, -2, 7, 6, -42, 1, 7, 7, 1, 4, -7, 25, -19, -9, -23, 5, 25, 0, 9, -50, 0, 0, 13, -12, -1, 66, 3, -33, -12, 2, 21, 45, -11, 6, -2, -63, 4, 4, 17, -78, -32, -32, 0, -17, -34, 3, -7, 3, 15, -8, -18, -7, -9, -11, -42, 10, -4, -40, -9, -22, -5, 6, 20, 8, 4, -20, 18, 6, -4, -24, 0, -2, 0, 7, 24, 4, -28, 37, 4, -39, 8, -3, 50, 0, 4, 5, 12, -35, -24, -40, -8, -1, -4, -17, 7, -40, -43, 25, 1, 1, 4, 0, -3, 54, 30, 3, -29, 9, 1, -2, 32, 11, 1, -6, -2, -5, 0, 44, -11, -7, -12, 6, 13, -6, -1, 2, -8, -4, -42, 0, 6, -41, 19, -1, -28, 33, -7, -10, -8, -27, 0, 3, -3, 5, -3, -4, -24, 1, -32, 31, -12, -43, 2, -1, 1, -32, 10, 0, 0, 14, -9, 44, -7, 4, -48, -5, 3, 5, 9, -2, -44, -9, -16, 17, -3, 44, 2, 9, 35, -1, -15, 2, -24, -29, 38, -31, 28, 1, -26, 0, -16, 12, -6, 0, 21, 2, -30, -1, 13, 29, 1, 13, -1, -16, -1, 5, -33, -9, -22, 3, 7, -2, -3, -13, -29, 9, 17, -7, -33, 37, 1, 0, 3, 3, 11, 9, 2, 5, -9, 4, 6, -8, -29, 2, 8, -18, -5, 4, -5, -45, -3, 2, 35, 3, 4, -3, -30, 25, 9, -15, -5, -1, 5, -11, 4, -14, 19, -18, 0, 0, 19, -31, -31, -10, -5, 6, -2, 7, 28, -1, 6, -7, -6, 4, 29, -7, 1, 15, 2, -6, -6, 34, -3, 0, 18, -11, 28, 0, -6, -5, -1, 36, 7, 3, -19, 16, -10, 22, 4, 0, -74, 13, 8, -7, -6, -10, 1, -11, -2, -5, -7, -2, -11, -29, 4, 0, -5, -48, 3, -7, -5, -1, -8, 4, 20, 15, -2, 4, -2, -36, -7, 0, 15, -28, -48, -2, -3, 0, 21, 9, 15, -9, -4, -3, -28, 22, 2, 54, 6, 4, -5, -5, 0, 6, 0, -1, 24, -2, 46, 2, 24, 8, 5, 5, -1, -7, -2, -3, -5, 1, 56, 2, 0, -10, 5, -12, -12, -55, 28, -2, -18, -13, 12, -4, 14, -3, 16, 13, -92, -3, 4, 7, -9, -6, -1, 23, 1, 40, 6, 3, 18, 53, -18, 1, -10, -31, -4, 31, 29, 55, 0, -41, -11, -14, -6, 3, -40, 17, 4, 9, -8, 5, 34, -60, -35, -5, -7, 9, -3, 2, 2, 10, -68, 3, -7, -11, 2, 6, 15, 9, 14, 35, -8, 5, 7, -2, 23, -6, -11, -6, -5, -1, -8, 5, -41, -5, -38, -1, -5, -1, -3, 0, 0, -1, -12, -36, -1, 8, -1, 3, 47, -19, 0, 0, -6, 2, -11, 32, 10, -12, 1, -8, 7, 19, 1, -1, -24, 60, -86, -6, -19, -4, -6, -24, -7, -44, 1, -18, -8, 0, 21, -51, 0, -1, 21, 14, -4, 30, 4, -34, 5, 5, 0, 0, -2, 15, -82, -9, 7, 6, 0, 4, -6, 23, -9, -13, 31, -38, 18, 30, 13, -5, 4, 2, 25, -8, -24, -48, 5, 7, 2, -12, 19, -10, -6, -4, 3, -42, -1, -8, 10, -21, -3, -11, -7, 29, -52, 6, 7, 6, 15, -43, 24, 11, 2, -26, -16, 2, -7, -9, -4, 13, 17, 3, -29, 14, 4, -16, -20, 8, -6, 32, -59, -16, 6, 41, 4, -37, 0, 65, -8, -44, -4, 4, 29, 63, -46, 7, -17, -22, 0, -2, -25, -57, -11, -26, 9, -16, 1, 7, -5, -6, 25, 7, 8, -8, -22, 22, -58, -6, 8, 0, -13, -3, -2, 12, -31, 3, -11, 9, 8, 1, -5, -2, 24, 1, 1, -11, -5, -3, -3, -5, 4, 18, -2, -9, -1, 35, -5, 7, 3, -23, 1, 1, 15, -9, -9, -29, 2, -6, 4, 23, -10, -23, -12, 7, -2, 28, 48, 1, 26, -27, -7, 29, 17, -4, -22, 6, 16, -1, -7, 1, -19, -6, -25, 32, -11, 5, -6, -26, 23, 0, 22, 6, -21, -5, 15, -41, 17, -4, -30, 45, -7, 0, 5, -3, 4, 11, 31, 2, 21, 17, -6, -55, -62, -12, 0, 0, -3, -32, 39, -6, 4, -10, -2, -23, -10, -5, -3, -7, 35, -14, -16, 0, -6, 0, -1, -35, -1, -8, -3, 6, 6, -1, 4, -5, 11, -9, -8, 2, -19, -3, -16, -2, 31, -24, 0, -1, -27, -35, 35, -2, 1, 11, 0, -44, -4, 10, 14, -35, -8, -2, 44, 22, 28, -8, 0, 7, -4, -1, 2, -8, 5, 1, 3, 15, 5, 1, 6, 16, -4, 1, -17, 7, -4, 4, 7, 11, -24, -24, 1, 6, -7, 43, -20, 3, 6, -7, 2, 17, 2, 2, -32, 33, 0, 27, -3, -7, -27, 1, -36, -8, -8, -37, 58, 31, -9, -10, -2, -26, 6, 3, -38, 3, -11, 24, -19, -6, 24, 3, 7, -31, -8, 5, -7, -67, -37, 0, -10, 10, -24, -35, 40, -5, -8, -4, -9, -40, -2, -56, 1, -9, 0, 0, -4, -5, -3, -7, 1, 1, -70, -1, 20, -4, -6, -18, -5, -7, -2, -7, 0, 2, 5, 2, -14, -2, 7, -8, 4, -53, 32, 3, -15, 2, 18, 14, -6, 0, -10, -65, 0, -12, 1, 18, -4, -3, 6, -11, 7, 8, 7, 2, -18, 46, -2, -10, -41, -16, 16, 5, 13, 19, -1, -6, 30, -8, 4, -7, -13, -6, -2, 15, -6, 1, 5, -37, -33, -14, 0, -17, -5, 8, -4, 11, 16, 1, 2, 7, -15, 4, 11, -1, -11, 13, -9, -8, 16, 1, -14, -58, -37, 18, -56, -5, -3, 4, -18, -25, -46, 19, 9, -21, -14, 10, 5, -3, -10, -25, 27, -5, 9, -7, 22, -1, -20, -4, -5, -8, -26, -9, 5, -4, 8, 10, -6, 44, -11, 6, 1, 1, -9, -18, -15, -29, 2, -63, -5, -49, 7, -5, 0, 11, 1, -50, -3, -2, -36, 8, 6, -3, 14, -1, -3, 5, 1, -4, 0, -13, -15, 1, -19, 1, 5, 6, 9, -1, 9, 10, 47, -71, -14, -34, 12, -37, -2, 18, 12, -11, 22, -25, 20, -10, 19, -11, 5, 28, -4, -10, 6, -30, 5, -4, 21, 5, -65, -40, -12, 41, -21, 1, 5, 6, -6, -32, -10, -2, -3, -35, 71, -19, -10, -16, -5, -10, 17, -3, -15, 11, 2, 43, 1, 2, -46, 9, -7, -5, 1, -40, 8, -1, 36, -21, -24, -21, 3, 0, -8, 30, 6, -6, 21, -27, -10, 3, -5, -69, -4, -11, 2, 26, -20, -26, 9, 0, 14, 0, -6, 10, -9, 4, 15, 3, 17, 0, -45, -6, 4, 14, 9, 9, -16, 36, 1, 2, -1, 0, 12, -5, 9, 2, -14, -1, 7, 0, 0, 11, -1, -3, -1, -31, 6, 0, 0, 14, 1, -1, 27, -50, 1, 10, -15, 0, 32, 38, -10, -5, -49, 0, -6, -52, 26, -5, 11, -40, 0, 37, 30, -1, 44, -4, -12, 4, -8, 3, -40, 11, -29, 6, 58, 59, 6, -18, 19, 1, -14, -6, -14, 0, -2, 2, -1, -5, -31, -3, 19, -16, -4, 0, -8, 4, 55, -1, 29, -27, -5, 17, 17, 10, 7, -1, -20, -25, -31, 0, -4, 5, 6, -10, -37, -5, 9, -18, 2, 2, -47, 6, -4, -1, 2, -14, -1, 3, -8, 2, 9, -4, -12, 3, 16, -20, -9, 3, -5, -65, 7, 4, -26, 6, -5, -5, -22, -23, 11, -69, -1, 21, -10, -68, -8, -36, -6, -7, -15, 3, -13, 30, -7, 4, 5, -8, 4, -1, 46, 6, 2, 0, 7, 3, 4, -3, 2, 11,
    -- layer=3 filter=0 channel=9
    -30, -3, 13, 36, 4, -8, -7, 22, -26, -21, 1, 7, -4, 41, 35, 1, 7, -11, 11, -39, 0, 8, -9, 10, -47, 16, -5, 2, 9, -11, 9, 52, 7, 5, 0, -16, 4, 2, -1, 3, -3, 31, 19, 6, -12, 1, 0, -31, -15, 23, 9, -10, 0, 0, 0, 21, 23, 5, -5, 34, -13, -18, -4, -4, 0, 17, 22, -45, 7, 13, -4, 5, -9, -1, -2, 8, -8, 34, 14, 5, -6, -1, 14, -1, 6, 24, -3, -8, -3, 1, 14, -33, 4, 41, 12, 6, -3, 1, -17, -21, -2, 7, -9, -23, 7, 4, -37, 2, -11, 11, -18, -8, 4, 9, 0, 4, 5, 35, -6, -17, -7, -6, -40, 19, -18, 8, -13, 9, -1, 31, -7, -60, 0, -19, -3, -9, 8, -9, -26, 10, 9, -6, 2, 5, -3, -11, 14, -15, -5, 15, -6, 2, -5, -28, 16, 6, 2, 3, -15, 7, 5, 0, 9, -6, -7, 0, 12, -4, -31, -18, -39, -34, -17, -2, 0, -8, -29, -50, -8, 22, 21, 5, -44, -6, -12, -1, -6, 42, 5, -3, 1, -34, 17, 0, 2, 0, -6, -9, -8, 21, 0, -56, 5, 4, -13, -43, 0, 1, -14, 26, -29, 7, -24, -5, -4, -6, -8, -28, -10, 1, 0, 2, -2, 8, 6, -1, -10, 2, 8, 5, 17, -20, 8, -2, 8, 4, 7, 6, -11, 4, -11, 0, -7, 20, 1, -12, 25, 14, 17, -32, -29, -8, -2, 17, 0, 5, 24, 5, -3, 22, -6, -46, 6, -11, 27, 3, -5, -1, 7, 38, -8, 10, -1, 30, -34, -28, -3, -23, -8, 5, -1, -32, 27, -45, -33, 24, -6, 21, 19, -24, 0, -9, 0, -12, -36, 6, 8, 0, 0, 1, 20, 8, -6, 38, 32, 3, 10, -61, -46, -3, -8, 14, 16, 5, -18, 4, 17, 26, 25, 3, 9, -54, 25, 30, 16, 12, 5, -30, 3, 14, 15, 8, -15, -9, 25, -3, 0, -33, 17, -3, -48, 6, -4, 2, 20, -7, 0, -1, 1, -1, -18, -43, 5, -6, 4, -1, 10, -7, -7, -1, -7, 6, 39, 3, 6, 13, 0, 8, 1, -25, 3, -2, -3, 18, 2, -7, 37, -14, -2, 3, 37, -2, 41, -12, -7, 10, 24, 1, -9, 33, 40, -9, -24, -6, -11, 4, -16, 3, 26, 0, -2, 6, 32, -1, 35, -32, -15, -60, 24, -6, -1, 1, 18, -1, -3, -2, 26, -14, -39, 15, 25, 3, 21, 26, -5, -4, -4, 1, 40, 7, -23, 5, -9, -17, 0, 20, 0, -57, 9, 6, 6, -8, -82, -4, 6, -14, 5, 31, -2, 7, 10, -6, -9, -10, -3, -3, -1, -1, 3, 14, 4, 4, 6, -11, -16, -1, 6, 3, 10, 20, 3, 0, -3, -11, -2, 4, -8, -8, 2, 7, 5, -2, -63, -23, 3, 12, -6, 29, 5, 32, 4, -44, 14, 0, 0, 0, -4, 2, 1, 0, 3, 0, -11, 1, 8, 3, -4, 0, 59, 5, -6, -3, -13, 4, -27, 20, 0, 6, -6, 11, -4, -11, -8, 5, -11, 10, 16, -4, -37, -3, -31, 0, -11, 0, -2, 14, -8, 14, 5, -5, 14, -29, 21, 41, 5, 6, -7, 22, -8, -5, -5, -17, 5, 24, -9, 1, -4, 10, -18, 19, -19, 18, 11, 33, 0, 3, 25, -16, 6, -1, 2, 11, -3, -32, 0, -6, -11, -10, 18, 3, -11, -37, -6, 3, -1, 1, -1, 1, -1, -11, -43, -6, -3, -9, -6, -7, -3, -29, -7, -1, 6, -3, 19, -39, 7, 16, 9, 7, -4, 7, -23, -9, -3, -2, 5, 0, -16, -11, 8, -7, -9, 1, 9, -1, -1, 4, 8, -8, -1, 6, 6, -7, -1, -3, -13, -4, 11, -5, -19, 5, 13, 37, 28, -8, -6, -39, -3, -1, 8, -6, -17, -23, 10, -11, -5, -1, -15, -10, 29, 0, -1, -33, 11, 5, -5, -19, -20, 0, 2, -6, -13, 5, -12, 5, 26, -3, -9, -2, 31, 0, 26, -24, -14, -7, -27, -3, -9, -2, -11, -7, 19, 30, -1, -7, -55, -3, 1, 1, 20, 13, -3, -3, -2, 5, -14, -17, -4, -6, -3, 3, 14, -13, -17, -25, -1, -4, -19, -31, -2, -4, 3, -8, 17, 1, -96, 14, -9, -4, -4, 5, -7, -34, -16, 9, 24, 34, 0, 1, -48, -5, 31, 39, -4, 28, -5, 0, 4, 3, 10, 15, 18, -5, -4, -6, -5, 18, -3, 15, 2, -3, -13, -26, -53, 7, 1, -16, -5, 3, -23, 15, 6, 11, -7, 13, -18, -16, 15, 21, -9, -7, -2, -31, -8, 6, 7, 19, 15, -48, 2, 16, 0, 5, 3, -13, 1, 3, 9, 5, 5, 11, 13, -1, -2, 25, 8, 1, 21, -3, -31, -2, 6, 29, 7, -7, 2, 43, -1, 10, 0, 0, -20, 34, -14, -31, -31, -22, 0, 2, 7, 3, -2, -2, 21, 14, -16, -41, 1, -13, 2, -19, 0, 2, 4, 4, -9, 1, -4, 4, 8, 7, -18, 6, 7, -4, -8, -6, -6, -3, 2, 3, -25, 4, 4, 23, -8, 0, 3, -1, -33, 1, 0, 0, -1, 6, 1, -7, -2, 1, 21, 4, 16, -2, -5, -10, -7, 16, 6, 50, 4, 3, 3, 0, 0, 1, 6, -11, -1, -69, -27, -7, 0, -1, 35, 3, -20, -7, -26, 19, 0, 0, 29, -17, -40, -7, -25, 5, -13, 1, -21, -7, 4, 0, -7, 14, 40, 4, 49, 0, -13, 12, -26, -25, 44, 0, 3, -14, -22, 0, -3, 7, 0, 0, 21, -4, 9, -8, 2, -10, 40, -8, 0, -2, -14, -7, 24, -3, -1, -11, -2, 10, -34, -1, 1, -25, -3, -13, -20, -1, -3, 2, -6, 3, 4, 2, -5, 0, 0, -2, 22, -6, 24, -9, 6, 10, -16, -14, 0, 7, 3, -37, -4, 3, -25, 11, -37, 20, 0, 3, -5, -18, -1, 29, -22, -50, 11, -2, -13, 6, -25, -3, -7, 3, -2, 4, 12, 6, -5, -3, -3, -26, 26, -12, -4, -6, -11, -2, -19, 5, -7, 7, 0, 15, -6, -36, -6, 5, -7, 9, 22, -6, -7, -36, -27, 4, 6, 2, 26, 32, -12, -6, 9, 6, -6, -5, -14, 37, 5, 28, -7, -14, -5, 2, 4, 5, 2, 22, -45, -8, 1, 9, 9, 18, -9, -12, 4, 29, -2, -3, 12, 12, 23, 3, -4, -4, -33, -2, 43, -7, -21, 5, 12, 9, -1, 13, -9, 1, -3, 7, -5, -8, 2, -24, 10, -6, -7, -5, -7, 3, -1, -11, -5, 0, -2, -4, -36, -25, 7, 63, -1, -9, -5, 0, -16, 30, -41, 3, -21, 2, 4, 4, -69, -6, -25, -39, 28, -15, 1, 9, 10, -6, -4, 47, 8, 20, 6, 4, -43, 25, -15, -7, -22, -12, 3, 23, 22, 2, 3, -12, -2, -16, 2, -4, -2, 15, 0, 3, 7, -5, 36, -9, -10, 13, -3, -3, 11, -6, -5, 33, 6, 0, -4, -21, -37, -2, 20, 3, -27, 0, -9, 8, 17, 1, 7, 6, -11, 0, -40, 0, 9, -8, -43, -41, 40, -11, 25, 16, -64, 4, 14, -4, 13, 26, -5, 2, 4, 15, 45, -9, 27, -6, 8, 11, -27, 5, 0, -10, 0, 9, 17, -21, 6, -2, -7, -26, 8, 9, -34, -10, -10, -31, 0, -8, -6, 2, -2, 8, -34, 5, -2, 3, -16, -21, -2, -2, -7, -48, -5, -1, 7, -7, -7, 14, 3, 0, -9, -3, -14, 18, -9, 28, -8, 22, -9, -50, -19, -22, -6, -61, -8, 19, -26, -1, -7, 14, 9, 41, 2, -2, 26, 32, 1, -1, 1, -10, -5, -7, -50, 3, -10, -94, -17, 33, 4, 0, -10, 30, -2, -27, -14, 7, 8, -45, -41, -11, -2, -16, 7, 48, 5, -6, 13, -10, 9, -31, 19, 2, -22, -16, 13, -15, 4, 5, -1, 1, 1, 18, -12, -11, -5, -2, 0, 40, 33, 5, -15, -17, -4, -19, 8, -36, -5, -13, 3, 26, 15, 15, 0, 7, -5, 13, -6, -35, 26, 8, -22, 8, -22, 0, 21, 2, -1, 9, -5, 0, -14, 13, -10, -9, 5, 2, -34, 5, -5, 0, 3, -1, -22, 7, -4, 36, -5, 0, -2, -29, 9, -14, -3, 31, 7, 15, 5, -15, -3, 0, -33, -4, -10, -5, -11, -11, -51, 7, -8, 19, -13, -9, -1, -5, 13, 9, 6, 18, 39, -6, 8, 5, -7, -13, -32, 2, -22, -64, -6, 32, -4, -45, 3, -2, 6, 4, 10, -33, -53, 20, -8, -9, 19, 2, -2, -2, 2, 2, 24, 3, 0, -10, 39, -28, 0, 5, 29, -1, 9, 3, 30, -25, -12, -3, -4, -7, 0, 14, -53, -4, -4, -7, -28, -10, 0, 0, -4, 0, 5, -34, -6, 5, -5, 6, 7, -2, 42, -6, -10, 3, -5, -3, 19, -5, 6, 1, -4, 0, 2, 2, 18, -2, -52, -29, -4, 0, -8, -15, 1, -20, -17, -36, -1, 5, -5, 0, -6, -7, 7, 3, 2, 0, 10, -1, -4, -2, -7, -66, -7, 5, 3, 20, -6, -6, -29, 0, -7, 1, -33, 12, -5, -5, 0, 5, -2, 1, 9, -7, 41, -17, 19, -4, 1, 6, -28, 5, 14, -7, 8, 4, -15, -11, -43, 22, 5, -23, 25, -26, 5, -1, 8, -6, -6, 34, -55, 5, -10, 18, -24, -18, -2, 16, -10, 3, 4, -3, -4, -28, -3, -6, 2, 19, 9, -28, -28, -3, -4, 41, -24, -7, 3, -52, 0, 0, 1, -5, 3, 3, -1, -14, -19, 2, -19, -5, 2, -5, 2, 14, 4, 0, 0, 1, -7, -13, -37, 1, 32, 5, 0, -7, -6, -66, 10, 0, 0, -60, -15, -12, -12, -7, 14, -2, 0, -3, -8, -8, 0, -3, -1, -34, 2, -18, -7, -9, -2, -5, 53, -6, 36, -2, -10, -28, 4, -45, -14, 2, 4, -9, 8, -2, 28, 6, -6, -5, 5, 6, 28, -63, 39, 6, -6, -18, 16, -4, -10, -24, 21, 5, 0, 17, -13, -1, 14, -2, -48, -29, 4, -5, 21, -4, 2, 2, -5, -40, 27, -8, -2, -7, 20, 34, -10, -21, 21, 2, 47, 3, -5, -2, 18, -14, 6, 0, -4, 11, 5, -41, -2, -3, -2, 14, -22, -8, 18, 0, -2, -5, -50, -7, -11, 5, -6, -24, 38, 22, -37, 7, -6, -25, 4, -9, -4, 0, -4, -4, -12, 16, -4, 4, -32, -17, -14, -19, 4, -17, 0, 0, 0, 0, -2, -2, -27, 0, -13, 5, -7, 12, -2, -47, 8, 54, 12, 2, 0, 0, 25, 34, 10, -1, -68, 0, 19, -27, 9, 41, 17, -3, 12, -27, 5, -5, -3, -12, -5, 5, -22, -20, -18, -9, 9, -26, -3, -10, -2, -2, -2, -18, -13, 6, -3, -3, -6, -32, 2, 14, -7, 21, -4, 3, 26, -8, -7, 1, 9, 7, -44, 16, -7, 28, -8, 30, -39, 16, -33, -78, -11, 42, 0, -9, -26, -17, 6, -3, 25, 0, 4, 5, -5, 11, 0, -30, 0, -17, 46, -14, -20, -6, -5, -4, 4, 0, -52, 0, -25, 5, -13, -3, -19, -5, -1, 8, -5, -8, -46, -2, -19, 3, 3, -1, 0, -7, -3, -1, 7, 3, 23, -4, 6, -7, -14, -3, 5, -29, 0, -7, 5, -14, -4, 28, 0, 18, 3, -7, -62, 10, 11, -37, -3, 32, -1, 6, 0, -19, -14, 5, -34, 0, 17, -28, -20, 17, 18, 8, -9, -4, 10, -4, 12, -25, 17, -9, 9, -46, 1, -9, 6, -9, -24, 0, 14, -3, -17, 17, -26, -9, -15, 4, 9, -5, -6, 3, -14, 0, -3, 3, 0, -13, 0, 13, -4, -50, 0, -6, -16, -42, 35, -1, -6, -14, 5, -53, -9, 1, 6, 3, -52, -2, -31, 9, 3, -9, -3, -25, 6, 1, -1, -5, 3, 5, -33, 8, 38, -31, -6, 1, -18, 16, 12, 8, -15, -8, 3, -8, 3, -36, -8, -40, 0, 0, -4, -20, 0, 8, -8, 22, 0, 10, -34, 0, 0, -4, -2, -5, -6, -8, -3, -9, -8, 0, -5, 37, -19, 6, 9, 36, 5, -2, 37, 18, -2, 4, 13, 3, 42, -9, 8, 4, -5, 4, -17, -2, -48, 3, 25, -22, -6, -3, 4, -4, -93, 42, 10, -5, 14, -17, 34, 16, -8, 43, 5, 13, -1, -1, 0, -44, -9, 52, 32, -6, 15, 3, 5, 28, -13, -30, -5, -16, -2, -3, 43, -11, 2, -10, -3, -51, -28, -50, 19, -3, -7, 38, 14, 24, 4, -1, 0, -3, 2, -6, 8, -10, 1, -42, -23, 1, -12, 3, 2, -3, -5, 15, -8, 0, 1, 0, 1, -31, 29, 42, 10, -7, -1, -1, -22, -9, -14, 12, 3, 13, -10, 18, 11, -8, 1, 38, 48, 0, -2, 63, 5, 0, -6, -19, 5, -15, -3, 6, -15, 9, -26, 5, 68, -17, -18, 1, 33, 1, -8, -45, -4, -5, -5, -4, -30, -15, 0, 10, 7, -3, 26, -45, -48, 26, -7, -5, -11, 0, -4, 51, -10, -5, 1, 32, 7, -4, -28, -10, 0, -33, 5, 7, 13, 7, 36, 14, 20, -7, -8, -2, -6, -8, 10, 6, -6, 5, 1, 7, -1, 7, -7, -10, 5, -39, -10, 0, -6, 2, -24, -33, -11, -4, -1, 8, 12, 10, -9, 33, 8, -9, 30, -8, -20, -7, -2, -15, -9, 47, -12, -11, 16, 22, -3, 31, 5, 8, 11, 4, -2, -11, -7, -5, 0, 0, 6, 2, -4, 32, 2, -10, 2, -3, -5, 59, -3, -3, -19, -10, -7, 2, 1, 16, 17, 33, -20, 29, 1, 38, 31, 22, -2, 21, -1, -1, 20, -13, -4, 1, 10, -10, -17, 29, -8, 1, 5, 15, -4, -5, -48, 35, 61, -18, -5, 19, 45, 0, 1, 18, -35, 18, -15, -22, -4, -23, -22, -9, -7, 5, 1, 0, 31, 0, -2, 4, -1, -16, 0, -2, 23, -35, -4, -15, -5, 55, 8, 5, 12, -26, 55, 37, -5, 6, -36, -3, 3, -6, 16, -29, -1, -27, 4, -27, 5, 43, 0, -16, 18, -6, -12, -5, -6, 3, -8, 14, -65, -10, 32, -4, -20, 0, 19, 7, 5, -2, -30, 1, 13, -7, -7, -1, 1, -9, -15, -6, 0, 4, 13, -1, -14, 0, -6, -20, -36, 0, 0, -30, -1, -3, 5, 8, -5, 25, 57, 15, -3, -7, -11, 7, 10, 1, -1, -11, -22, 0, -9, -32, -35, -7, -48, 9, -26, 4, 5, 6, -2, 1, 42, -7, -67, 0, -21, 1, -31, 18, 20, 3, 0, -3, -6, 6, 6, -1, -3, -26, -1, -50, 77, 0, 58, 0, 62, -5, -2, -8, 3, -8, -7, 5, 11, 0, -9, 12, 32, -38, 0, 2, 29, -6, 26, 2, -8, 8, -7, -47, 5, -6, 20, -9, 3, -6, -68, 6, 9, -4, 1, -5, 0, -8, -4, 4, -18, -9, -43, -6, 13, -14, -11, -4, 8, 14, 16, -2, -17, -8, 0, 0, 63, -55, -10, 23, -8, -6, 3, 16, -7, 22, 7, -36, 8, -6, -43, -29, 29, 2, -5, -8, -5, 6, -10, 5, 5, 0, 0, -25, 17, 7, 6, 49, -15, 0, 13, 22, 5, -6, -3, 7, 0, -34, 6, 1, -2, -21, 7, 9, 30, -11, -23, -4, -8, 0, 14, 21, -6, 10, 2, 0, 45, 13, 3, 14, 3, 50, 14, -8, 5, 6, -6, 23, -3, 0, 49, -2, -5, 14, 24, -3, -1, -24, 3, -48, -7, 2, 20, 1, -5, 0, 3, -28, -3, -19, -35, 0, -10, -7, -40, -30, 0, -3, 1, -6, 0, 0, 10, -1, -4, -15, -1, -8, -12, -8, 17, -4, -6, 14, -9, -10, 0, -5, -16, 26, -11, 49, -18, 5, -2, -1, 30, 7, 3, 2, 13, -15, -12, -36, 1, -12, -3, -14, 1, -11, 0, 3, -4, 4, -4, -34, -2, -16, -4, -7, 28, 18, -46, -6, 10, 15, 16, -45, -23, -23, -13, -5, 32, -7, -7, 0, -17, 0, -10, -5, 0, 7, 12, -38, -33, 5, 7, 26, 0, -5, 1, 27, -23, 3, 7, -3, 16, -7, -5, -2, 45, -17, 0, -2, 29, 0, 3, 28, -25, -15, -19, -1, -5, 3, 30, -32, 30, 31, 3, -9, -3, -10, -6, -6, 0, -22, 11, 6, -2, -8, -30, -53, -32, -6, -3, 15, -1, 4, -5, -21, -4, 3, 19, 23, -5, -9, 3, 12, 40, -4, 42, -11, 18, -7, -4, 0, 1, 27, -9, -6, 17, -7, -4, -13, 13, 8, -25, -32, 0, 18, 6, 4, -9, -10, -4, 16, -17, -2, 3, 6, 9, 2, 4, 50, 9, -38, 0, -15, -17, 8, 29, -30, -5, -12, -7, 0, 27, 0, -27, 22, -14, -2, 25, 25, 4, -3, 0, 17, 2, 10, -35, -2, -2, -45, -6, 8, -19, -2, 4, -3, 13, -14, 2, 8, 0, 42, 1, -14, -4, 17, 1, 39, -14, 4, -5, -4, 3, -38, -4, -8, -11, -6, -4, 4, 0, -12, 10, -61, 35, 1, 28, 11, -9, 2, 0, 31, -32, -3, -11, -8, -29, -9, 2, -2, -1, 1, -1, -10, 5, 4, 21, 0, -40, -6, 6, 37, 8, -14, -7, -8, -27, 3, -7, -5, -7, 12, -32, -3, -13, 4, -5, -3, 4, 5, 21, -7, 8, -7, 5, -4, -37, -5, -5, -7, -6, -4, 9, -11, -3, -22, 0, -4, -4, 6, 57, -19, -4, 19, -9, 3, -16, -54, -3, -11, 18, 8, -6, -5, -42, 5, -5, 31, 25, 7, 14, 8, 11, 3, 41, -6, 8, -2, -37, -13, 16, -32, -17, 2, 5, -19, 6, -5, 6, 6, -48, -13, 0, -28, 0, -2, 3, 28, -6, -7, -8, -4, -1, 4, -4, 7, 0, -32, 3, -8, 9, 4, 5, -9, -61, 1, 6, 2, 3, 5, -4, -16, -16, 0, 9, -10, -19, 44, 21, -2, 6, -8, -14, -15, -7, -10, 3, -4, 0, 5, 13, -3, -5, 0, -5, -8, -46, 7, 4, -3, 9, 0, 1, 5, 13, 1, 18, -4, 9, -9, 0, 5, 5, 10, -5, -11, -2, -3, -45, -8, 15, 1, 5, 6, -5, 3, -20, -5, 6, 8, -9, -52, -9, 10, -5, 1, -9, 6, -45, -4, -10, 1, -18, 17, -35, -32, -8, -5, -4, -14, -18, -9, 18, 21, -44, 3, 1, 2, -37, -30, 3, -15, -1, -5, 15, 28, -20, 33, 2, -59, 59, 31, -4, -10, 7, 26, -4, 4, 10, -7, 6, 5, -13, -37, -44, 5, 5, -42, 5, -7, -48, -25, -55, -15, -5, 27, 61, -32, -3, -9, -8, -5, -27, -57, -4, 25, -8, 0, -1, 0, -1, 2, 6, -5, 3, -7, 28, -3, 35, -1, -3, -43, 5, 8, 4, -4, 10, 18, -42, -7, -52, -1, -3, -2, -2, -61, 24, -7, 6, -7, 12, -17, 35, 5, 13, -30, 2, -2, -9, -31, -7, -3, 5, 10, 6, 0, 6, 2, 28, -13, 27, 3, -14, -12, 23, -50, -48, -42, 3, 41, -7, -5, 10, 1, -35, -5, -6, 6, -7, -2, -19, 8, -1, -76, 1, -10, -21, 8, -12, -59, 24, 5, -7, 11, 23, 3, -22, 5, -20, -29, -4, -1, -39, 0, -26, 16, -45, 25, 27, -8, -2, 0, -14, -5, 45, 3, 44, 19, 31, -5, -1, -3, 3, 11, 17, 2, -13, 15, 43, 8, -34, 0, 10, 2, -16, -6, 5, 9, -2, -1, -37, 19, -5, 11, -18, -24, 15, 5, 18, -10, 3, 6, -6, -8, 6, -52, 7, 4, -58, 5, 2, 3, -43, -16, -11, -39, 7, -11, -1, 5, 0, -8, -3, -59, -3, -6, 13, -10, -3, 7, 3, -78, -15, 39, -29, -6, 1, -25, 39, 28, 0, -49, -44, 10, -52, -50, 16, -9, -13, -8, -3, -70, -1, -2, -10, -37, -1, -4, -53, 6, -29, -37, 0, -22, 3, -2, 4, -23, -19, 0, 0, 9, -9, -19, -14, -11, 10, 9, 6, 41, -38, -4, -4, 7, -4, 22, 20, 4, -38, 4, -32, -5, -10, -1, 7, 1, -29, -25, -40, -70, -5, 6, 13, -13, -8, 2, -8, 27, -8, -1, -1, 29, 1, -11, -7, 5, 9, 3, 22, 2, -31, 0, 5, 27, -21, 0, -25, -5, -15, 11, -79, 6, 6, -7, -1, 3, -41, -33, -9, 7, -6, -7, 30, 1, -9, -10, 1, -9, -24, 0, -3, 3, 31, -6, -10, -26, 0, -10, -3, -2, 2, 26, -55, 5, -12, -21, -40, -4, 18, -4, -4, 44, 37, 7, 6, -81, -47, -4, 14, 12, 11, 0, -21, 0, 29, 8, -31, 4, 13, 0, 23, -27, 28, 3, -1, -46, -6, -3, 12, -7, -76, -9, -9, 11, -41, 47, -46, -3, -23, -3, -25, -19, 5, 0, -77, 5, 27, -6, -53, 36, 1, 36, -24, -20, -5, 1, -22, 3, 20, -3, 5, 0, -6, 25, 28, 6, 2, 2, -25, -24, -54, 6, -5, -6, -7, -13, 7, -5, 2, 0, 15, 4, 22, -5, -4, 34, 3, 9, -27, -45, 0, -5, 22, 8, -7, -4, -12, -13, -23, -74, 4, -11, -6, -28, 6, -1, -14, 24, 11, -3, -67, 30, -8, 1, -4, 0, 5, -7, 1, -5, -1, 3, 1, -13, -11, -10, -9, 8, 48, -3, -21, 1, 1, -7, 0, 16, 63, 33, -10, -6, 4, -36, -37, -8, -3, -1, -42, -15, 6, -4, 14, 12, -12, -20, -5, 0, 0, -17, -14, 6, 0, -37, 23, 5, 5, 1, -7, -20, -6, -5, 49, -9, 3, 2, 58, 5, -66, 25, -4, -19, 5, 3, -36, 27, 19, -10, 5, 5, 24, 44, 9, 0, -1, -31, 17, -15, -8, 13, 4, 0, -8, -4, 5, -7, -1, -5, -22, -5, 0, -1, 3, 9, -6, 1, -8, 6, 1, 3, -2, -21, 3, -17, 5, -9, -5, -7, 11, -30, 0, -9, -3, -1, 3, -9, 12, 4, 16, -8, 0, 0, 2, -27, 1, 0, -7, 5, -9, 19, -5, 1, 2, -9, 6, -5, 18, -19, -8, -14, 20, -22, 3, 19, -15, -9, 1, -8, 34, 15, -9, 4, -2, -2, -6, 7, -4, -50, 7, -17, 12, 11, 7, -4, -29, -8, 2, 20, 22, -2, -50, -8, 8, -12, 2, -5, -28, 0, -11, -35, -34, 10, -13, 7, 1, -6, 22, 35, 28, 29, -12, -3, 24, -4, -12, 4, -9, -17, -7, 1, -3, -11, -18, -15, 28, 4, 6, -20, -38, 3, -13, -10, -6, -2, 14, 31, 15, -7, -15, -33, 30, 3, -2, -7, -4, 12, -4, 20, 6, -51, -1, -5, 13, 4, -8, 1, -27, 27, -8, 6, 2, 21, 7, -2, 5, 8, -9, -64, -16, 3, -18, 5, -2, 0, -4, -52, 20, 22, -49, 12, 16, -9, 22, -3, 2, 0, 10, -3, -10, -33, 29, 28, 4, -12, 16, -7, -9, 1, 6, 24, -6, -1, -8, -32, 37, -79, 3, -6, 6, -7, -13, 4, 15, -45, -17, 1, -2, 39, -13, -11, -4, -9, -3, 9, -50, -3, -34, 1, -3, -27, 9, -5, -20, -61, 10, 5, -2, 26, 67, -27, 13, 0, 7, -42, 0, 10, 29, 12, -33, 1, 7, 12, 9, 17, 7, 20, 0, 14, -2, -30, 0, 2, 19, -6, 20, 7, 0, 38, -20, 25, -11, -2, -19, -2, 8, 0, -2, -2, -35, 0, 0, 33, 3, 2, -2, -2, 10, 10, -3, -3, 0, 6, 20, -9, 9, 4, 4, 4, 2, 17, 0, -9, 3, 9, -9, -11, 12, 33, 8, -7, -14, -2, 11, 0, -8, -29, 10, -6, 6, 16, -23, 0, 5, 5, 1, -14, 18, 13, 2, -2, 12, 0, 19, 6, -19, 0, -21, -10, -33, -13, 3, 1, -20, -7, -48, 0, -10, 12, -39, 32, 2, -5, -21, -14, 2, -2, 6, 6, 5, 6, -27, 0, 29, 16, 3, 53, -39, -35, -5, -5, 10, 8, -19, -3, 0, -18, -5, -43, -6, 2, 3, -9, -5, 26, 0, 6, 0, 0, -4, -1, 8, -5, 2, 0, -11, -8, -22, -4, -8, 17, -11, 4, 2, -64, 10, 7, 39, 22, 0, 3, 33, 0, -12, 9, 4, -27, 0, 0, 3, 22, -6, 29, 4, -3, -6, 21, 1, -7, -6, -6, -4, 0, 27, -3, 3, -2, 4, -7, 21, 3, -7, -13, 20, -1, -20, 8, -8, 3, -54, -10, -9, 7, 2, -8, 5, 14, -52, 0, 25, -60, -30, -4, 0, 3, -15, 0, -25, -26, -2, -2, 48, 25, 31, 10, -2, -7, 15, -11, -10, -10, -1, 4, 7, -25, 18, 1, 3, -4, 17, 14, -51, -29, -2, -29, 9, 7, 18, 2, -12, -2, 0, 14, 26, -81, -76, -4, -11, 22, -4, -32, 8, 13, -1, 7, 2, 5, -3, -2, -6, -2, 0, -2, -16, 4, 2, 10, -4, 24, -12, 4, -5, 7, 22, 36, 12, 24, -22, -1, -2, -3, 8, -18, 17, -3, 25, -7, 23, -60, 26, 8, 9, -43, -2, -6, -7, -53, -3, 2, -4, 4, 2, -24, 2, -4, 24, -2, 13, -4, 1, -18, 7, -11, -31, -19, -20, 19, 0, 0, 6, -8, 8, 8, 2, 3, -3, 8, 24, -32, -4, -77, 7, 12, -10, -12, -10, -5, -6, 5, 4, 32, 33, -8, -40, 4, -27, -42, -3, 0, -60, -3, 36, 0, -28, 6, 5, -2, 0, 0, 18, -1, 34, 5, 19, 8, 11, 0, 0, 3, 6, 14, 3, 2, -3, 10, -9, -19, -1, 0, 1, -3, 32, -5, -2, -13, -9, -6, 9, -3, 3, 1, -11, -29, -32, 5, -32, -19, -40, 9, -5, -60, 0, -43, -20, -10, 39, 24, -4, -8, -61, -1, -22, -13, 26, 14, 17, -5, 9, -10, 0, -47, -35, -9, -69, 8, 5, 37, 6, 14, 22, 2, 9, -34, -7, 5, 23, 2, -8, -11, 21, -5, -57, -16, -36, -9, 5, -13, 39, -34, -2, -5, 5, 5, 3, 1, 46, -21, -17, -14, -9, -19, -8, 0, 2, -39, 11, 11, 26, 1, 6, 31, -3, -24, 1, 8, 0, 26, 7, -3, -37, 7, 2, -3, -44, 0, -58, -67, -3, -14, 4, 0, 18, 6, -37, -12, -4, -28, -10, 5, 0, -62, -50, 7, -25, 24, -10, 5, 4, 29, 7, -60, -8, -31, 34, 35, -7, -9, -33, -7, 0, 32, 2, 8, 39, 0, -8, 1, -7, -2, 6, -1, -45, -4, 0, -17, -6, -7, 13, 3, 18, -1, -2, 1, -11, -1, -29, 3, -7, -19, -7, 2, -13, 34, -5, -6, -8, 3, 7, 2, -66, 33, 7, 18, 9, 8, 9, -5, -7, -8, 38, -4, 6, -20, -56, 1, -13, -1, -27, 5, 7, 4, -46, -7, 8, 3, 25, -8, -17, -25, 35, -15, -12, -41, -6, -29, 1, 6, -55, 1, -3, -26, -25, 15, -36, -2, -38, 8, -31, -14, 0, 2, -26, 2, -35, 5, -4, -39, 5, 46, 9, 16, 5, 7, 12, 0, -5, 2, 7, -8, 5, 19, -26, 4, -5, -9, -1, 26, -49, 4, -5, -10, -16, -9, 8, 3, -1, 0, -7, -4, 3, 3, -10, 35, -8, 0, 36, -61, 0, -6, -26, -11, 3, -3, -24, 9, 0, -1, 5, -43, 7, 4, 3, 5, -24, 12, 8, 5, -4, -15, 0, 6, -5, 2, 2, 6, 27, -1, 6, -1, 0, 56, -26, 2, 0, -46,

    others => 0);
end iwght_package;
