library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 0, 0, 13, 36, 23, 20, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 18, 22, 16, 43, 28, 27, 11, 0, 
    35, 7, 0, 0, 0, 26, 37, 29, 27, 6, 19, 26, 11, 10, 0, 
    71, 48, 8, 34, 51, 60, 46, 17, 18, 0, 64, 40, 13, 17, 7, 
    63, 71, 3, 0, 9, 30, 45, 44, 22, 21, 58, 29, 20, 15, 20, 
    75, 51, 19, 0, 0, 30, 80, 50, 26, 28, 57, 32, 17, 31, 11, 
    84, 66, 75, 24, 28, 45, 25, 19, 2, 23, 15, 40, 18, 3, 0, 
    78, 75, 66, 33, 27, 34, 17, 26, 35, 32, 36, 3, 0, 0, 0, 
    52, 67, 67, 17, 68, 20, 58, 77, 56, 23, 4, 19, 33, 20, 20, 
    66, 79, 52, 60, 131, 90, 66, 63, 56, 48, 55, 61, 65, 70, 69, 
    80, 69, 60, 101, 89, 59, 61, 58, 55, 55, 59, 62, 74, 74, 67, 
    82, 68, 66, 107, 65, 59, 63, 57, 60, 64, 75, 77, 78, 70, 106, 
    90, 76, 84, 52, 61, 63, 67, 63, 61, 66, 71, 66, 60, 86, 80, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 31, 0, 0, 0, 10, 1, 
    0, 61, 0, 1, 0, 4, 0, 0, 0, 48, 0, 0, 0, 0, 38, 
    0, 46, 0, 61, 0, 12, 0, 0, 0, 65, 0, 0, 0, 0, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 125, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 29, 26, 0, 0, 0, 87, 0, 0, 0, 10, 0, 
    0, 0, 7, 0, 44, 42, 0, 0, 0, 52, 0, 0, 14, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 0, 26, 0, 0, 0, 0, 15, 16, 
    0, 0, 0, 38, 0, 0, 21, 0, 1, 0, 0, 0, 32, 28, 0, 
    13, 0, 0, 117, 0, 17, 25, 0, 0, 0, 14, 19, 20, 0, 0, 
    28, 0, 0, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 29, 45, 0, 0, 0, 0, 0, 0, 0, 3, 7, 0, 0, 9, 
    0, 0, 82, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 33, 0, 0, 
    
    -- channel=2
    92, 96, 96, 97, 97, 90, 100, 113, 104, 77, 61, 67, 74, 80, 84, 
    94, 105, 99, 100, 97, 80, 77, 85, 57, 24, 0, 2, 29, 59, 77, 
    60, 74, 106, 107, 105, 84, 55, 27, 1, 0, 0, 0, 0, 6, 58, 
    0, 10, 88, 104, 87, 53, 5, 0, 0, 0, 0, 0, 0, 0, 26, 
    0, 0, 59, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 54, 78, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 31, 86, 13, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 28, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 15, 5, 0, 0, 12, 50, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 67, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    186, 193, 189, 194, 191, 188, 198, 194, 187, 181, 165, 159, 167, 170, 158, 
    181, 189, 194, 201, 191, 227, 227, 193, 172, 134, 161, 143, 126, 139, 163, 
    182, 136, 192, 195, 194, 234, 191, 126, 97, 162, 222, 174, 167, 105, 142, 
    200, 104, 200, 191, 208, 158, 213, 163, 146, 160, 239, 173, 142, 98, 94, 
    259, 237, 242, 176, 324, 303, 277, 181, 138, 98, 247, 206, 140, 125, 86, 
    286, 280, 259, 219, 240, 277, 299, 210, 168, 122, 326, 199, 144, 151, 112, 
    275, 325, 192, 198, 172, 237, 336, 259, 204, 190, 295, 186, 140, 150, 167, 
    313, 313, 222, 208, 172, 292, 326, 222, 176, 205, 262, 192, 133, 184, 160, 
    354, 326, 276, 196, 226, 204, 198, 189, 153, 236, 168, 158, 97, 132, 183, 
    329, 329, 298, 202, 245, 168, 179, 279, 213, 182, 155, 67, 97, 178, 200, 
    265, 326, 302, 212, 397, 265, 271, 311, 233, 145, 88, 111, 145, 173, 170, 
    204, 270, 296, 377, 456, 199, 163, 156, 137, 131, 138, 147, 154, 171, 166, 
    178, 181, 229, 448, 255, 149, 151, 140, 135, 133, 143, 161, 180, 170, 176, 
    174, 149, 187, 362, 172, 154, 159, 143, 139, 150, 162, 163, 158, 158, 219, 
    193, 149, 163, 174, 139, 124, 143, 146, 157, 173, 170, 144, 167, 243, 175, 
    
    -- channel=4
    118, 126, 120, 123, 119, 116, 130, 133, 123, 112, 98, 98, 98, 106, 103, 
    117, 125, 126, 128, 119, 111, 121, 121, 95, 52, 38, 46, 63, 91, 101, 
    110, 99, 125, 129, 125, 132, 98, 55, 31, 22, 50, 33, 37, 47, 89, 
    64, 28, 124, 124, 119, 66, 69, 33, 24, 38, 65, 48, 35, 29, 58, 
    50, 52, 116, 80, 98, 49, 79, 46, 33, 0, 64, 49, 29, 27, 21, 
    39, 78, 119, 78, 111, 86, 93, 57, 39, 3, 81, 54, 34, 25, 13, 
    31, 84, 105, 117, 61, 64, 114, 57, 64, 19, 79, 41, 19, 26, 41, 
    45, 73, 44, 87, 46, 96, 80, 67, 60, 49, 73, 51, 27, 47, 66, 
    60, 64, 45, 61, 48, 57, 69, 50, 40, 54, 85, 49, 17, 60, 95, 
    75, 63, 70, 12, 84, 21, 28, 66, 36, 80, 41, 10, 23, 78, 108, 
    57, 64, 70, 14, 62, 36, 33, 76, 51, 1, 0, 0, 0, 15, 20, 
    11, 40, 60, 59, 115, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 110, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    0, 2, 0, 5, 5, 0, 0, 4, 8, 5, 3, 0, 0, 6, 12, 
    1, 0, 0, 6, 0, 0, 26, 9, 10, 0, 11, 8, 0, 0, 6, 
    26, 0, 0, 6, 0, 0, 43, 18, 0, 0, 23, 17, 31, 0, 0, 
    90, 0, 0, 0, 24, 0, 14, 22, 7, 0, 53, 2, 34, 22, 0, 
    72, 0, 30, 0, 5, 6, 52, 48, 27, 0, 13, 51, 4, 39, 0, 
    50, 0, 44, 5, 0, 6, 50, 36, 66, 0, 60, 64, 0, 24, 20, 
    49, 30, 0, 58, 0, 0, 12, 39, 66, 0, 69, 45, 0, 0, 25, 
    35, 34, 18, 21, 0, 0, 84, 11, 39, 0, 41, 54, 0, 0, 18, 
    45, 0, 93, 0, 22, 0, 24, 16, 0, 18, 0, 64, 0, 0, 0, 
    14, 0, 101, 0, 40, 6, 0, 21, 15, 13, 51, 0, 0, 0, 11, 
    0, 0, 90, 0, 86, 19, 0, 14, 62, 34, 0, 0, 0, 0, 0, 
    0, 0, 19, 0, 97, 57, 0, 0, 12, 0, 0, 0, 0, 0, 5, 
    11, 0, 0, 12, 127, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 0, 0, 81, 33, 0, 11, 0, 0, 0, 0, 0, 1, 0, 8, 
    32, 0, 0, 1, 11, 0, 0, 0, 0, 0, 10, 0, 0, 18, 44, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 0, 4, 4, 30, 8, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 20, 0, 0, 0, 52, 3, 7, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 5, 0, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 6, 
    25, 0, 0, 0, 0, 63, 42, 49, 28, 2, 0, 0, 0, 0, 0, 
    0, 14, 0, 0, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 3, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 63, 9, 17, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=7
    0, 2, 4, 0, 0, 7, 0, 0, 2, 0, 3, 11, 7, 0, 0, 
    2, 3, 4, 0, 7, 31, 0, 1, 0, 31, 0, 0, 11, 15, 0, 
    0, 38, 1, 0, 2, 7, 0, 0, 11, 42, 0, 0, 0, 4, 21, 
    0, 57, 0, 10, 0, 28, 0, 0, 0, 44, 0, 0, 0, 0, 46, 
    0, 15, 0, 58, 0, 0, 0, 0, 0, 75, 0, 0, 1, 0, 9, 
    0, 12, 0, 0, 73, 0, 0, 0, 0, 129, 0, 0, 8, 0, 0, 
    0, 0, 0, 0, 58, 47, 0, 0, 0, 96, 0, 0, 3, 12, 0, 
    0, 0, 0, 0, 27, 43, 0, 0, 0, 50, 0, 0, 17, 0, 0, 
    0, 0, 0, 35, 0, 1, 0, 0, 24, 0, 11, 0, 17, 17, 0, 
    0, 0, 0, 44, 0, 0, 36, 0, 0, 0, 0, 4, 34, 20, 0, 
    58, 0, 0, 114, 0, 0, 26, 0, 0, 0, 7, 13, 16, 13, 0, 
    31, 33, 0, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 26, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 22, 0, 0, 
    
    -- channel=8
    63, 69, 68, 70, 67, 65, 71, 75, 67, 52, 42, 45, 53, 61, 59, 
    67, 72, 73, 72, 68, 69, 65, 56, 34, 17, 14, 14, 21, 39, 56, 
    43, 37, 68, 73, 71, 49, 32, 14, 13, 13, 21, 17, 15, 16, 41, 
    28, 25, 60, 67, 58, 30, 35, 21, 11, 12, 25, 17, 10, 12, 25, 
    22, 34, 58, 46, 59, 44, 32, 21, 10, 4, 29, 26, 15, 15, 14, 
    9, 22, 60, 42, 17, 30, 38, 29, 20, 11, 27, 15, 13, 12, 16, 
    14, 17, 35, 54, 27, 27, 31, 23, 24, 7, 20, 16, 8, 11, 25, 
    17, 17, 22, 35, 28, 31, 22, 13, 24, 23, 23, 15, 8, 20, 39, 
    15, 10, 12, 15, 23, 9, 21, 18, 17, 20, 18, 8, 8, 32, 58, 
    15, 14, 17, 0, 23, 15, 12, 27, 21, 18, 4, 0, 20, 45, 53, 
    0, 12, 14, 12, 35, 25, 5, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 16, 21, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 3, 2, 0, 0, 
    7, 0, 0, 0, 0, 2, 4, 4, 6, 10, 9, 5, 0, 0, 0, 
    6, 9, 0, 0, 0, 0, 3, 6, 7, 6, 3, 0, 3, 3, 0, 
    5, 10, 0, 0, 0, 0, 0, 2, 3, 0, 2, 4, 0, 0, 12, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 37, 0, 0, 0, 0, 28, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 10, 3, 11, 10, 0, 0, 
    37, 26, 0, 0, 0, 0, 30, 10, 0, 0, 0, 0, 0, 0, 0, 
    45, 56, 0, 0, 95, 54, 1, 7, 0, 0, 30, 22, 10, 19, 0, 
    0, 0, 0, 0, 0, 0, 25, 24, 29, 13, 0, 0, 0, 9, 34, 
    14, 0, 0, 0, 0, 2, 0, 6, 9, 0, 0, 9, 0, 12, 16, 
    9, 19, 24, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 2, 0, 0, 0, 0, 7, 6, 0, 0, 0, 0, 0, 3, 
    0, 0, 10, 2, 2, 0, 2, 53, 0, 0, 0, 0, 14, 0, 0, 
    0, 0, 0, 46, 128, 92, 0, 0, 0, 13, 41, 52, 19, 0, 0, 
    0, 0, 17, 11, 0, 0, 0, 0, 0, 0, 1, 0, 10, 5, 4, 
    10, 0, 0, 0, 0, 5, 2, 1, 5, 12, 19, 25, 0, 0, 35, 
    7, 3, 0, 0, 0, 6, 17, 6, 1, 7, 0, 0, 0, 21, 0, 
    9, 3, 0, 0, 0, 0, 0, 0, 20, 27, 10, 6, 44, 35, 14, 
    
    -- channel=12
    51, 50, 52, 52, 55, 48, 53, 57, 54, 44, 37, 40, 41, 45, 47, 
    55, 52, 56, 52, 55, 52, 41, 42, 32, 31, 19, 23, 33, 43, 45, 
    30, 53, 54, 55, 57, 56, 22, 26, 19, 33, 1, 10, 15, 33, 45, 
    0, 61, 50, 58, 43, 40, 19, 6, 15, 35, 0, 12, 4, 14, 55, 
    0, 37, 33, 62, 15, 10, 0, 0, 9, 43, 11, 0, 17, 9, 37, 
    0, 14, 18, 29, 24, 0, 0, 7, 3, 59, 0, 0, 20, 9, 12, 
    0, 4, 25, 24, 52, 23, 4, 0, 0, 57, 0, 0, 19, 17, 7, 
    0, 0, 13, 21, 45, 23, 0, 10, 0, 49, 0, 0, 20, 12, 25, 
    0, 0, 0, 25, 3, 19, 10, 15, 27, 32, 14, 0, 20, 38, 48, 
    0, 0, 0, 33, 0, 8, 25, 5, 5, 4, 2, 14, 32, 51, 41, 
    17, 0, 0, 40, 0, 0, 7, 0, 0, 4, 7, 4, 11, 21, 9, 
    10, 0, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 3, 15, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 8, 0, 7, 8, 7, 6, 0, 
    13, 0, 0, 0, 0, 0, 5, 0, 18, 0, 0, 2, 0, 5, 0, 
    32, 19, 0, 0, 14, 0, 0, 0, 12, 0, 24, 12, 2, 5, 0, 
    9, 55, 0, 0, 0, 0, 21, 0, 15, 0, 23, 5, 2, 0, 0, 
    17, 24, 3, 0, 0, 4, 37, 21, 0, 0, 14, 12, 4, 8, 0, 
    35, 35, 34, 0, 0, 17, 0, 0, 0, 0, 0, 23, 1, 0, 0, 
    25, 33, 41, 16, 17, 0, 0, 2, 13, 7, 32, 7, 0, 0, 0, 
    28, 22, 44, 0, 15, 11, 41, 60, 47, 24, 17, 31, 52, 49, 42, 
    103, 50, 17, 16, 113, 80, 77, 72, 70, 69, 79, 83, 81, 87, 84, 
    111, 89, 10, 69, 77, 72, 79, 73, 73, 74, 82, 83, 97, 96, 84, 
    111, 98, 68, 102, 65, 74, 75, 75, 77, 82, 97, 103, 101, 93, 138, 
    111, 103, 99, 90, 81, 83, 86, 75, 72, 78, 91, 84, 69, 109, 113, 
    
    -- channel=14
    56, 57, 57, 54, 52, 54, 62, 63, 52, 45, 44, 48, 47, 48, 44, 
    54, 59, 59, 57, 54, 28, 41, 51, 43, 11, 0, 3, 29, 48, 45, 
    39, 67, 60, 59, 60, 40, 22, 9, 8, 0, 0, 0, 0, 28, 46, 
    0, 28, 54, 55, 38, 24, 0, 0, 0, 15, 0, 0, 0, 0, 46, 
    0, 0, 33, 41, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 23, 
    0, 0, 31, 41, 29, 10, 0, 0, 0, 20, 0, 0, 0, 0, 0, 
    0, 0, 42, 25, 23, 7, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 15, 12, 0, 0, 0, 8, 0, 0, 0, 3, 13, 
    0, 0, 0, 0, 2, 7, 0, 0, 1, 0, 17, 0, 8, 18, 39, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 9, 28, 31, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    74, 68, 75, 75, 72, 66, 78, 81, 71, 55, 46, 51, 57, 64, 63, 
    73, 72, 77, 75, 78, 30, 76, 52, 38, 21, 7, 12, 24, 53, 61, 
    26, 53, 78, 76, 78, 25, 36, 24, 35, 0, 16, 16, 2, 34, 42, 
    6, 20, 76, 72, 45, 46, 18, 31, 8, 25, 9, 18, 10, 15, 32, 
    31, 0, 79, 89, 17, 44, 16, 18, 0, 31, 21, 26, 6, 7, 25, 
    51, 0, 86, 51, 0, 57, 4, 26, 0, 14, 20, 26, 12, 11, 18, 
    71, 0, 65, 49, 0, 27, 3, 23, 8, 0, 23, 18, 7, 14, 27, 
    49, 0, 47, 32, 45, 12, 14, 9, 28, 2, 15, 14, 13, 17, 53, 
    17, 0, 28, 1, 44, 17, 27, 0, 30, 0, 25, 10, 10, 34, 60, 
    4, 7, 2, 0, 37, 34, 26, 0, 27, 28, 0, 9, 8, 35, 57, 
    0, 13, 0, 14, 3, 31, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 28, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=16
    93, 92, 92, 92, 92, 92, 92, 92, 92, 93, 94, 92, 91, 92, 92, 
    94, 92, 92, 93, 92, 92, 92, 92, 92, 108, 91, 87, 92, 92, 92, 
    95, 94, 93, 92, 92, 94, 93, 103, 100, 86, 82, 92, 94, 93, 93, 
    88, 93, 92, 92, 95, 103, 86, 89, 76, 72, 66, 69, 94, 93, 93, 
    102, 90, 86, 93, 94, 83, 80, 86, 91, 100, 115, 117, 108, 85, 94, 
    56, 64, 84, 94, 98, 110, 114, 111, 105, 97, 67, 58, 65, 63, 91, 
    107, 98, 83, 72, 86, 74, 41, 31, 49, 98, 112, 117, 100, 112, 96, 
    29, 45, 64, 68, 71, 53, 53, 101, 100, 83, 64, 44, 42, 42, 65, 
    0, 61, 53, 64, 91, 105, 101, 89, 77, 91, 93, 100, 104, 105, 89, 
    87, 111, 111, 112, 111, 100, 96, 83, 82, 81, 80, 72, 59, 61, 63, 
    45, 50, 64, 71, 75, 83, 94, 95, 90, 83, 70, 61, 52, 45, 51, 
    11, 0, 18, 8, 0, 0, 4, 16, 16, 17, 15, 24, 61, 52, 37, 
    0, 2, 5, 3, 0, 0, 6, 71, 60, 65, 72, 44, 18, 32, 44, 
    13, 0, 0, 0, 0, 0, 0, 20, 27, 3, 0, 13, 32, 38, 54, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 29, 31, 42, 57, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 10, 43, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 8, 0, 
    15, 26, 1, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 59, 0, 
    0, 0, 0, 1, 0, 0, 12, 46, 71, 0, 0, 0, 0, 0, 0, 
    38, 36, 0, 27, 0, 3, 46, 0, 0, 0, 0, 3, 20, 22, 25, 
    162, 0, 14, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 13, 15, 
    0, 40, 0, 0, 0, 14, 51, 25, 28, 32, 48, 47, 6, 0, 25, 
    0, 6, 0, 0, 0, 1, 94, 0, 0, 0, 0, 0, 16, 18, 26, 
    0, 2, 5, 0, 2, 2, 66, 5, 0, 0, 35, 30, 0, 14, 15, 
    0, 1, 6, 5, 7, 10, 35, 11, 34, 50, 4, 0, 7, 11, 14, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 12, 2, 1, 2, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 15, 108, 95, 51, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 34, 9, 0, 0, 0, 0, 0, 0, 
    
    -- channel=19
    441, 438, 438, 438, 438, 439, 439, 440, 436, 439, 435, 438, 438, 438, 438, 
    442, 439, 439, 439, 438, 438, 438, 439, 438, 431, 370, 412, 440, 438, 439, 
    437, 437, 439, 441, 440, 443, 433, 442, 387, 344, 333, 382, 441, 440, 442, 
    419, 434, 438, 442, 444, 449, 391, 424, 369, 370, 349, 380, 440, 439, 443, 
    285, 285, 366, 435, 439, 432, 420, 432, 428, 432, 415, 373, 341, 324, 435, 
    343, 363, 426, 394, 392, 384, 343, 358, 380, 419, 371, 363, 357, 342, 432, 
    243, 240, 300, 330, 411, 259, 168, 210, 314, 428, 408, 374, 340, 365, 333, 
    76, 231, 258, 280, 345, 336, 355, 415, 333, 296, 265, 237, 254, 281, 328, 
    69, 380, 339, 378, 412, 425, 402, 364, 334, 338, 325, 334, 302, 297, 276, 
    258, 275, 281, 284, 287, 290, 294, 260, 259, 236, 230, 200, 185, 199, 221, 
    69, 58, 88, 74, 82, 98, 126, 137, 150, 138, 120, 124, 144, 189, 216, 
    28, 17, 89, 56, 5, 0, 39, 144, 104, 101, 126, 178, 221, 207, 222, 
    52, 0, 17, 14, 0, 0, 66, 250, 252, 238, 205, 150, 159, 216, 266, 
    114, 0, 0, 0, 0, 0, 7, 128, 117, 71, 98, 180, 217, 232, 293, 
    112, 13, 0, 0, 0, 0, 6, 43, 63, 145, 214, 210, 222, 259, 309, 
    
    -- channel=20
    95, 94, 94, 94, 94, 94, 94, 96, 95, 93, 92, 94, 94, 94, 94, 
    95, 94, 94, 94, 94, 94, 94, 95, 96, 100, 80, 91, 94, 94, 94, 
    95, 95, 94, 95, 94, 98, 91, 99, 85, 77, 61, 74, 96, 94, 95, 
    83, 86, 93, 96, 97, 106, 84, 90, 51, 42, 29, 51, 91, 91, 93, 
    61, 68, 87, 95, 97, 99, 78, 93, 77, 86, 86, 78, 82, 68, 90, 
    29, 28, 70, 96, 98, 109, 94, 94, 78, 78, 54, 40, 37, 33, 84, 
    53, 47, 84, 58, 77, 18, 0, 0, 40, 94, 97, 93, 94, 79, 70, 
    0, 9, 28, 50, 71, 45, 28, 64, 66, 54, 34, 23, 14, 26, 35, 
    0, 67, 44, 55, 69, 86, 92, 84, 43, 51, 50, 56, 51, 48, 48, 
    12, 50, 43, 46, 40, 42, 32, 20, 27, 15, 14, 14, 3, 10, 17, 
    0, 0, 3, 6, 13, 12, 14, 12, 11, 5, 0, 0, 0, 11, 23, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 6, 28, 32, 32, 
    0, 0, 11, 10, 0, 0, 0, 106, 92, 88, 72, 51, 43, 31, 39, 
    26, 0, 0, 0, 0, 0, 5, 133, 121, 63, 36, 31, 40, 37, 46, 
    32, 0, 0, 0, 0, 0, 0, 44, 33, 25, 47, 43, 42, 40, 46, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 30, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 19, 10, 29, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 27, 0, 36, 2, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 19, 0, 3, 0, 12, 11, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 0, 0, 0, 15, 15, 5, 33, 0, 0, 
    0, 0, 0, 0, 28, 98, 0, 0, 0, 0, 7, 10, 0, 0, 0, 
    0, 0, 10, 0, 0, 25, 0, 17, 1, 13, 22, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 33, 0, 0, 0, 9, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 11, 5, 0, 23, 0, 17, 0, 0, 0, 
    12, 0, 8, 0, 0, 0, 0, 0, 1, 7, 0, 0, 0, 0, 0, 
    26, 0, 22, 34, 15, 0, 0, 29, 4, 0, 0, 0, 0, 1, 0, 
    47, 0, 0, 24, 12, 0, 0, 26, 30, 35, 18, 2, 0, 0, 0, 
    96, 4, 0, 7, 3, 1, 0, 0, 26, 0, 0, 0, 0, 0, 0, 
    85, 13, 5, 4, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    64, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 20, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    53, 60, 41, 0, 0, 0, 16, 14, 0, 0, 0, 0, 0, 0, 6, 
    17, 0, 0, 4, 2, 0, 0, 0, 3, 32, 25, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 
    0, 20, 25, 32, 26, 29, 13, 19, 14, 8, 8, 19, 0, 0, 0, 
    63, 62, 65, 72, 73, 71, 61, 50, 39, 37, 35, 17, 6, 0, 0, 
    5, 8, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 36, 32, 15, 5, 13, 0, 0, 0, 0, 31, 8, 0, 0, 
    0, 5, 6, 12, 8, 7, 0, 0, 6, 24, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 1, 0, 9, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=23
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 28, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 14, 0, 0, 0, 
    0, 20, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 
    0, 0, 0, 0, 0, 0, 7, 8, 17, 0, 0, 0, 0, 34, 0, 
    0, 31, 14, 24, 0, 0, 8, 30, 33, 0, 0, 0, 0, 0, 28, 
    56, 23, 0, 40, 2, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 
    149, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 0, 3, 1, 3, 0, 0, 0, 0, 0, 0, 0, 1, 0, 10, 
    0, 21, 0, 0, 6, 15, 13, 8, 2, 0, 3, 7, 18, 0, 8, 
    0, 38, 0, 0, 0, 12, 79, 0, 0, 0, 5, 0, 0, 2, 22, 
    0, 12, 11, 0, 0, 4, 89, 0, 0, 0, 0, 19, 17, 14, 24, 
    0, 2, 8, 2, 4, 5, 52, 35, 22, 41, 32, 14, 1, 15, 19, 
    0, 0, 0, 0, 2, 4, 24, 30, 30, 24, 0, 0, 7, 10, 15, 
    
    -- channel=24
    20, 20, 20, 20, 20, 20, 19, 21, 21, 18, 18, 19, 20, 20, 20, 
    19, 19, 19, 19, 19, 19, 19, 19, 17, 10, 1, 14, 20, 19, 19, 
    19, 19, 19, 20, 20, 20, 16, 13, 0, 0, 0, 4, 19, 19, 19, 
    9, 12, 17, 19, 20, 20, 12, 17, 12, 10, 9, 8, 12, 14, 16, 
    0, 0, 2, 18, 19, 19, 18, 19, 17, 15, 5, 0, 0, 0, 12, 
    22, 23, 17, 11, 9, 1, 0, 0, 0, 6, 12, 18, 19, 12, 11, 
    0, 0, 0, 6, 11, 0, 0, 0, 12, 16, 9, 1, 2, 0, 0, 
    0, 10, 2, 2, 7, 26, 30, 15, 0, 0, 0, 0, 0, 5, 8, 
    0, 16, 19, 20, 10, 4, 0, 4, 4, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 
    1, 0, 12, 12, 4, 0, 0, 5, 0, 0, 9, 24, 20, 10, 13, 
    13, 0, 0, 5, 3, 1, 10, 65, 77, 65, 34, 13, 19, 13, 10, 
    14, 4, 1, 3, 3, 3, 16, 74, 62, 27, 26, 24, 13, 9, 7, 
    11, 11, 7, 5, 6, 5, 0, 13, 30, 32, 26, 11, 12, 10, 8, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 19, 22, 41, 48, 47, 29, 33, 28, 26, 13, 0, 0, 0, 0, 
    38, 35, 16, 28, 44, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 47, 46, 45, 48, 49, 16, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 37, 41, 42, 44, 44, 28, 0, 1, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 28, 50, 65, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    88, 85, 0, 0, 0, 0, 0, 0, 0, 0, 49, 79, 83, 38, 0, 
    0, 0, 0, 0, 2, 5, 8, 57, 42, 0, 0, 0, 0, 0, 0, 
    0, 70, 0, 0, 0, 102, 111, 0, 0, 0, 0, 32, 44, 64, 26, 
    83, 26, 72, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 
    0, 0, 19, 29, 5, 0, 85, 143, 96, 95, 101, 84, 0, 0, 14, 
    27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 10, 7, 
    23, 2, 0, 0, 0, 2, 0, 0, 0, 0, 57, 32, 0, 0, 0, 
    6, 29, 24, 19, 22, 24, 1, 0, 68, 45, 2, 0, 0, 0, 0, 
    
    -- channel=28
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 
    0, 1, 0, 0, 0, 0, 15, 21, 10, 0, 0, 0, 0, 0, 0, 
    21, 10, 3, 20, 0, 0, 1, 0, 0, 0, 0, 0, 8, 1, 0, 
    46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    7, 29, 1, 7, 13, 16, 31, 0, 4, 3, 7, 0, 0, 5, 16, 
    11, 26, 20, 10, 18, 22, 48, 0, 0, 0, 0, 9, 10, 19, 20, 
    0, 24, 24, 20, 23, 24, 37, 0, 0, 12, 23, 26, 17, 18, 17, 
    0, 28, 28, 28, 27, 28, 34, 30, 22, 36, 21, 17, 19, 17, 15, 
    
    -- channel=29
    34, 34, 34, 34, 34, 34, 34, 34, 31, 36, 37, 34, 34, 34, 34, 
    35, 34, 34, 35, 34, 34, 34, 34, 37, 65, 44, 31, 34, 34, 34, 
    36, 35, 33, 34, 33, 36, 37, 54, 65, 60, 56, 41, 34, 34, 35, 
    39, 40, 36, 33, 34, 49, 28, 37, 30, 36, 27, 28, 41, 38, 36, 
    80, 62, 36, 34, 35, 35, 29, 33, 35, 49, 80, 85, 79, 42, 40, 
    23, 21, 52, 48, 47, 87, 85, 77, 61, 50, 25, 19, 29, 17, 44, 
    93, 75, 52, 21, 61, 48, 33, 2, 5, 55, 73, 79, 66, 82, 55, 
    23, 13, 39, 25, 27, 1, 7, 72, 68, 50, 36, 20, 17, 13, 34, 
    0, 48, 18, 30, 53, 65, 68, 61, 53, 78, 73, 87, 89, 88, 64, 
    93, 98, 103, 102, 96, 87, 88, 72, 74, 65, 80, 68, 58, 53, 45, 
    48, 46, 63, 71, 75, 83, 102, 98, 94, 88, 74, 62, 42, 30, 27, 
    12, 5, 13, 12, 8, 5, 0, 14, 21, 14, 0, 6, 37, 20, 3, 
    1, 7, 8, 2, 0, 0, 0, 0, 0, 0, 23, 0, 0, 5, 11, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 8, 22, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 5, 12, 22, 
    
    -- channel=30
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 15, 5, 2, 2, 63, 53, 47, 34, 27, 4, 0, 0, 0, 
    0, 1, 6, 4, 3, 1, 69, 110, 90, 45, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 20, 40, 23, 5, 0, 0, 0, 0, 0, 
    
    -- channel=31
    12, 10, 10, 10, 11, 10, 11, 11, 12, 9, 6, 11, 10, 10, 10, 
    12, 10, 10, 10, 10, 10, 11, 10, 6, 0, 0, 10, 10, 10, 10, 
    11, 11, 10, 10, 11, 8, 10, 0, 0, 0, 0, 0, 12, 11, 10, 
    4, 4, 9, 12, 10, 0, 11, 6, 10, 1, 0, 2, 7, 7, 9, 
    0, 4, 0, 12, 10, 4, 5, 10, 7, 5, 0, 0, 0, 12, 5, 
    12, 6, 0, 16, 0, 15, 0, 0, 1, 0, 12, 13, 0, 1, 4, 
    0, 0, 4, 13, 0, 13, 0, 0, 18, 4, 4, 1, 5, 0, 4, 
    6, 0, 4, 0, 5, 27, 13, 0, 0, 0, 0, 0, 0, 1, 4, 
    14, 0, 10, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 12, 2, 0, 2, 5, 0, 0, 0, 0, 3, 12, 2, 0, 11, 
    13, 3, 0, 8, 8, 3, 15, 57, 50, 34, 6, 5, 23, 7, 5, 
    12, 6, 1, 4, 5, 4, 24, 20, 16, 7, 24, 13, 8, 13, 4, 
    25, 13, 9, 7, 8, 7, 1, 0, 30, 24, 14, 14, 15, 11, 5, 
    
    -- channel=32
    99, 88, 99, 105, 106, 102, 100, 99, 94, 101, 103, 96, 98, 98, 94, 
    96, 84, 93, 100, 97, 98, 98, 95, 93, 113, 80, 92, 100, 98, 97, 
    91, 78, 85, 89, 86, 87, 90, 88, 88, 108, 64, 98, 102, 91, 91, 
    89, 75, 88, 87, 82, 80, 75, 82, 100, 63, 66, 73, 65, 86, 85, 
    71, 72, 62, 66, 71, 74, 75, 73, 61, 60, 57, 26, 48, 66, 57, 
    28, 29, 51, 32, 36, 37, 61, 65, 56, 46, 29, 42, 66, 26, 46, 
    52, 57, 46, 53, 59, 68, 62, 56, 47, 47, 55, 75, 55, 49, 70, 
    54, 48, 44, 63, 77, 84, 86, 95, 89, 93, 65, 56, 60, 53, 3, 
    80, 89, 75, 90, 101, 104, 94, 73, 61, 54, 41, 58, 65, 62, 56, 
    60, 48, 80, 92, 78, 70, 76, 85, 79, 70, 70, 75, 78, 66, 48, 
    78, 80, 83, 86, 88, 83, 86, 61, 42, 69, 82, 64, 48, 33, 37, 
    61, 79, 84, 57, 45, 56, 74, 62, 55, 47, 47, 42, 28, 29, 15, 
    57, 80, 72, 67, 67, 54, 40, 40, 47, 43, 27, 28, 30, 16, 11, 
    42, 36, 30, 27, 32, 34, 33, 29, 12, 33, 23, 22, 16, 12, 14, 
    12, 9, 11, 12, 11, 16, 23, 24, 22, 32, 18, 15, 13, 12, 18, 
    
    -- channel=33
    0, 16, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 4, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 
    0, 8, 5, 0, 0, 0, 0, 0, 0, 0, 47, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 22, 0, 0, 
    14, 25, 0, 13, 8, 11, 0, 0, 0, 0, 49, 32, 0, 6, 0, 
    4, 0, 0, 19, 10, 0, 2, 2, 14, 12, 39, 0, 0, 0, 0, 
    8, 9, 25, 25, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 10, 0, 0, 0, 0, 0, 9, 0, 28, 0, 0, 0, 0, 
    0, 35, 2, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 3, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 
    0, 1, 1, 2, 4, 2, 0, 0, 23, 0, 0, 0, 0, 2, 0, 
    
    -- channel=34
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=35
    363, 313, 381, 408, 420, 420, 436, 444, 427, 449, 446, 446, 449, 454, 439, 
    373, 318, 386, 412, 420, 417, 424, 427, 428, 450, 335, 436, 452, 453, 437, 
    378, 313, 378, 407, 420, 403, 413, 377, 378, 408, 263, 397, 435, 425, 423, 
    358, 290, 363, 369, 400, 382, 389, 362, 315, 212, 196, 205, 243, 371, 360, 
    205, 198, 212, 226, 250, 261, 266, 280, 209, 202, 178, 166, 244, 295, 226, 
    135, 164, 210, 161, 215, 215, 234, 224, 196, 193, 181, 295, 326, 251, 239, 
    183, 179, 168, 172, 230, 254, 253, 241, 244, 251, 271, 342, 324, 278, 190, 
    214, 223, 231, 277, 305, 322, 326, 324, 305, 306, 236, 279, 305, 254, 176, 
    233, 234, 223, 290, 321, 310, 295, 278, 274, 283, 266, 301, 294, 276, 279, 
    202, 204, 275, 286, 259, 279, 299, 301, 261, 289, 300, 301, 266, 214, 162, 
    217, 261, 264, 255, 245, 250, 290, 192, 156, 253, 252, 208, 164, 126, 123, 
    186, 241, 251, 169, 164, 213, 245, 186, 174, 175, 161, 133, 111, 91, 64, 
    166, 206, 188, 160, 158, 145, 131, 139, 140, 124, 102, 98, 96, 58, 55, 
    84, 71, 75, 78, 99, 101, 98, 98, 79, 136, 79, 73, 58, 55, 60, 
    50, 47, 58, 64, 70, 81, 88, 84, 75, 111, 63, 53, 51, 54, 65, 
    
    -- channel=36
    42, 12, 42, 55, 67, 70, 83, 92, 80, 93, 92, 92, 89, 94, 86, 
    56, 28, 58, 73, 83, 82, 94, 95, 85, 104, 68, 93, 95, 103, 88, 
    71, 37, 69, 85, 98, 87, 101, 89, 85, 99, 48, 87, 100, 106, 93, 
    83, 46, 91, 97, 110, 94, 102, 83, 57, 52, 6, 43, 90, 108, 96, 
    57, 39, 59, 66, 83, 79, 68, 68, 25, 13, 2, 15, 22, 74, 61, 
    0, 1, 19, 0, 13, 12, 10, 18, 6, 7, 0, 35, 55, 84, 38, 
    0, 3, 9, 0, 11, 6, 2, 0, 0, 7, 24, 72, 98, 69, 39, 
    0, 0, 0, 0, 12, 18, 25, 29, 39, 56, 46, 71, 69, 37, 18, 
    16, 12, 4, 22, 31, 30, 27, 29, 32, 45, 27, 49, 54, 61, 70, 
    0, 0, 3, 16, 13, 19, 31, 47, 34, 46, 48, 66, 58, 54, 32, 
    0, 3, 16, 27, 25, 21, 40, 17, 0, 49, 48, 44, 30, 14, 18, 
    0, 8, 17, 0, 0, 13, 49, 14, 3, 23, 23, 2, 9, 0, 1, 
    1, 19, 27, 5, 3, 11, 12, 7, 7, 4, 5, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 6, 0, 0, 0, 0, 6, 
    
    -- channel=37
    22, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 3, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 0, 7, 0, 0, 
    26, 0, 0, 3, 0, 0, 15, 0, 0, 99, 0, 0, 13, 0, 0, 
    25, 0, 0, 0, 3, 0, 16, 20, 26, 41, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 25, 20, 9, 0, 0, 0, 30, 0, 
    0, 0, 19, 0, 0, 0, 0, 19, 0, 4, 0, 0, 61, 0, 52, 
    0, 4, 14, 0, 0, 5, 0, 5, 0, 0, 0, 0, 47, 5, 82, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 38, 0, 0, 4, 75, 8, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 32, 0, 0, 1, 15, 0, 
    21, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 16, 14, 30, 2, 
    0, 0, 0, 10, 0, 0, 34, 32, 0, 0, 8, 27, 18, 14, 7, 
    0, 0, 32, 9, 0, 0, 30, 12, 0, 5, 12, 10, 16, 7, 18, 
    0, 0, 18, 0, 0, 0, 5, 0, 1, 5, 14, 0, 23, 4, 5, 
    1, 1, 1, 0, 0, 0, 0, 7, 0, 23, 5, 4, 8, 0, 5, 
    4, 0, 0, 0, 0, 0, 0, 11, 0, 47, 0, 5, 0, 0, 27, 
    
    -- channel=38
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 79, 24, 85, 67, 0, 0, 
    39, 16, 40, 31, 35, 26, 25, 17, 0, 0, 0, 0, 0, 0, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 11, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 21, 
    0, 0, 0, 0, 0, 0, 0, 28, 23, 0, 0, 22, 12, 9, 0, 
    0, 0, 0, 21, 5, 0, 0, 0, 0, 15, 5, 2, 17, 2, 16, 
    0, 0, 7, 0, 3, 33, 25, 0, 0, 12, 17, 0, 3, 7, 0, 
    25, 39, 21, 10, 0, 0, 11, 17, 6, 0, 6, 4, 8, 0, 0, 
    2, 2, 3, 4, 4, 0, 0, 0, 4, 6, 0, 8, 2, 0, 0, 
    
    -- channel=39
    0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 4, 0, 0, 0, 0, 0, 0, 0, 26, 3, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 7, 0, 56, 13, 0, 0, 2, 
    0, 4, 0, 7, 0, 0, 0, 0, 0, 0, 4, 0, 62, 0, 6, 
    3, 5, 1, 15, 7, 11, 9, 0, 0, 0, 0, 10, 4, 0, 6, 
    20, 2, 0, 14, 4, 0, 0, 0, 0, 0, 27, 8, 0, 24, 0, 
    1, 0, 0, 26, 11, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 
    0, 0, 7, 1, 0, 0, 0, 0, 0, 0, 17, 12, 0, 0, 0, 
    0, 0, 24, 8, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 18, 0, 0, 24, 0, 0, 0, 0, 0, 0, 
    30, 0, 0, 0, 1, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 3, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 
    0, 4, 2, 2, 2, 0, 0, 0, 34, 0, 0, 0, 0, 5, 0, 
    
    -- channel=40
    0, 0, 0, 1, 6, 10, 13, 16, 13, 17, 17, 18, 18, 18, 17, 
    0, 0, 4, 11, 13, 15, 16, 15, 15, 11, 0, 17, 20, 19, 18, 
    8, 5, 11, 19, 21, 18, 19, 10, 10, 9, 0, 8, 18, 20, 21, 
    13, 13, 21, 23, 28, 25, 23, 18, 0, 0, 0, 0, 0, 17, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 12, 12, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 27, 19, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 16, 24, 20, 3, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 11, 14, 13, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 13, 10, 7, 14, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=41
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 19, 24, 
    0, 0, 3, 4, 0, 0, 0, 0, 4, 6, 9, 15, 20, 23, 23, 
    22, 22, 19, 16, 15, 15, 11, 9, 0, 6, 20, 23, 24, 22, 23, 
    
    -- channel=42
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=43
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 
    16, 19, 3, 10, 41, 28, 2, 0, 0, 10, 44, 70, 38, 0, 1, 
    0, 0, 0, 0, 0, 21, 36, 58, 75, 56, 20, 0, 0, 0, 0, 
    36, 56, 75, 64, 33, 20, 12, 0, 0, 0, 0, 0, 0, 33, 107, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 34, 38, 0, 0, 0, 0, 
    28, 46, 6, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 7, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=44
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 4, 12, 0, 0, 
    0, 0, 1, 7, 0, 0, 0, 0, 0, 0, 0, 0, 18, 4, 7, 
    11, 4, 0, 12, 7, 0, 0, 0, 0, 0, 11, 11, 0, 24, 0, 
    2, 0, 0, 9, 0, 0, 0, 0, 0, 0, 10, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 7, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 3, 5, 
    10, 0, 0, 0, 0, 4, 0, 0, 5, 1, 0, 7, 2, 7, 7, 
    3, 0, 0, 0, 0, 3, 0, 2, 3, 6, 3, 10, 2, 10, 12, 
    6, 6, 8, 9, 9, 10, 10, 8, 15, 2, 9, 8, 9, 13, 10, 
    13, 17, 17, 16, 14, 12, 12, 8, 24, 0, 11, 9, 12, 14, 7, 
    
    -- channel=45
    77, 55, 64, 64, 59, 50, 46, 48, 42, 44, 44, 36, 39, 43, 33, 
    67, 43, 50, 50, 46, 41, 43, 43, 38, 73, 25, 32, 37, 41, 31, 
    56, 35, 36, 32, 34, 32, 43, 46, 35, 76, 28, 46, 40, 33, 30, 
    50, 20, 34, 22, 24, 21, 30, 40, 79, 55, 56, 54, 32, 41, 24, 
    54, 48, 48, 47, 42, 44, 45, 64, 48, 57, 53, 3, 23, 29, 29, 
    30, 23, 47, 22, 29, 33, 57, 65, 51, 40, 6, 6, 26, 7, 30, 
    56, 45, 47, 44, 48, 51, 53, 44, 36, 35, 21, 29, 19, 30, 30, 
    51, 36, 32, 51, 61, 65, 67, 73, 68, 74, 35, 16, 20, 17, 0, 
    77, 85, 58, 71, 86, 88, 78, 54, 38, 31, 16, 28, 33, 26, 36, 
    55, 44, 74, 80, 60, 53, 57, 70, 57, 45, 40, 47, 58, 51, 33, 
    71, 75, 74, 79, 81, 65, 77, 52, 23, 58, 67, 55, 44, 35, 40, 
    62, 69, 82, 54, 43, 51, 71, 53, 46, 42, 49, 46, 31, 34, 22, 
    61, 78, 75, 66, 63, 52, 37, 41, 53, 45, 29, 33, 37, 24, 22, 
    44, 38, 36, 33, 39, 40, 38, 33, 13, 42, 30, 27, 24, 21, 20, 
    18, 15, 19, 19, 20, 24, 32, 32, 20, 37, 26, 21, 22, 21, 29, 
    
    -- channel=46
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 
    0, 0, 0, 4, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=47
    0, 6, 0, 0, 0, 7, 3, 0, 2, 5, 17, 10, 16, 0, 18, 
    0, 17, 0, 9, 0, 12, 0, 0, 9, 0, 29, 9, 19, 0, 18, 
    0, 32, 9, 18, 3, 13, 0, 5, 18, 0, 16, 9, 12, 6, 15, 
    1, 38, 10, 19, 16, 18, 12, 0, 0, 0, 0, 4, 13, 3, 33, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 9, 0, 9, 
    0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 20, 6, 0, 0, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 8, 14, 21, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 12, 15, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 3, 1, 3, 18, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    
    -- channel=48
    63, 85, 85, 73, 73, 79, 75, 69, 73, 72, 74, 73, 67, 77, 85, 
    73, 95, 92, 93, 75, 91, 91, 89, 92, 89, 94, 85, 89, 92, 93, 
    75, 94, 93, 77, 53, 41, 49, 37, 46, 48, 46, 60, 92, 94, 96, 
    76, 91, 95, 61, 60, 64, 57, 66, 74, 74, 65, 67, 65, 94, 95, 
    83, 91, 85, 88, 79, 80, 77, 76, 83, 78, 74, 66, 90, 92, 97, 
    80, 93, 100, 83, 76, 77, 78, 81, 82, 78, 76, 92, 94, 91, 93, 
    79, 90, 73, 72, 93, 101, 96, 97, 95, 96, 95, 96, 96, 98, 98, 
    80, 96, 66, 55, 51, 71, 96, 100, 97, 94, 91, 93, 93, 93, 95, 
    81, 94, 95, 79, 75, 30, 57, 76, 97, 104, 95, 94, 95, 95, 97, 
    79, 92, 93, 102, 84, 16, 17, 23, 38, 58, 73, 94, 99, 99, 97, 
    77, 94, 94, 85, 17, 26, 0, 0, 23, 6, 6, 5, 7, 64, 83, 
    89, 113, 111, 110, 112, 91, 83, 99, 101, 93, 91, 87, 99, 101, 101, 
    42, 51, 48, 45, 44, 43, 47, 60, 71, 70, 74, 76, 80, 84, 84, 
    35, 40, 38, 29, 23, 21, 22, 22, 16, 15, 11, 11, 11, 7, 0, 
    15, 13, 10, 9, 8, 4, 7, 3, 4, 2, 4, 6, 0, 0, 48, 
    
    -- channel=49
    10, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    8, 0, 0, 0, 0, 12, 0, 17, 8, 3, 2, 2, 8, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 2, 0, 0, 2, 0, 26, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 34, 94, 15, 13, 31, 23, 81, 18, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 33, 
    0, 0, 0, 0, 0, 6, 2, 9, 0, 4, 0, 0, 14, 27, 0, 
    
    -- channel=50
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=51
    300, 355, 353, 324, 321, 344, 345, 332, 342, 341, 347, 345, 344, 379, 386, 
    303, 354, 367, 348, 302, 326, 330, 320, 340, 340, 338, 326, 372, 387, 393, 
    298, 347, 372, 322, 312, 288, 298, 290, 313, 326, 317, 328, 360, 388, 393, 
    307, 341, 360, 285, 293, 295, 297, 295, 306, 311, 294, 315, 308, 377, 384, 
    332, 342, 352, 357, 309, 310, 307, 319, 326, 318, 314, 321, 374, 381, 381, 
    351, 363, 343, 333, 358, 351, 358, 368, 363, 360, 359, 371, 376, 379, 381, 
    359, 360, 305, 245, 259, 347, 378, 389, 388, 387, 378, 381, 380, 382, 381, 
    364, 392, 375, 336, 236, 208, 304, 381, 392, 381, 375, 377, 378, 377, 376, 
    370, 401, 407, 394, 313, 137, 175, 219, 277, 336, 354, 386, 383, 378, 377, 
    370, 400, 404, 410, 285, 96, 105, 134, 160, 166, 157, 229, 282, 339, 372, 
    360, 395, 398, 389, 272, 259, 150, 159, 286, 223, 204, 201, 211, 330, 352, 
    298, 325, 316, 305, 298, 274, 257, 283, 305, 283, 296, 289, 312, 304, 305, 
    201, 204, 202, 192, 185, 175, 173, 185, 192, 177, 178, 174, 179, 183, 169, 
    137, 127, 122, 113, 117, 103, 100, 102, 105, 97, 88, 94, 93, 87, 94, 
    111, 99, 96, 97, 95, 93, 109, 105, 115, 107, 105, 95, 84, 137, 198, 
    
    -- channel=52
    39, 49, 47, 57, 51, 57, 60, 56, 54, 55, 60, 60, 58, 69, 70, 
    32, 43, 58, 79, 91, 95, 97, 93, 100, 99, 97, 79, 68, 72, 70, 
    34, 38, 61, 99, 96, 90, 93, 89, 89, 95, 88, 78, 74, 68, 67, 
    33, 37, 72, 76, 73, 68, 75, 71, 70, 85, 82, 83, 59, 64, 61, 
    42, 38, 52, 62, 52, 51, 49, 54, 60, 58, 55, 56, 59, 61, 58, 
    56, 58, 55, 51, 45, 44, 46, 52, 51, 49, 49, 46, 61, 60, 57, 
    58, 42, 40, 62, 68, 52, 58, 62, 63, 64, 62, 63, 61, 64, 63, 
    60, 62, 77, 47, 23, 53, 67, 66, 69, 68, 63, 62, 60, 58, 55, 
    67, 72, 74, 83, 70, 23, 27, 77, 86, 72, 56, 62, 63, 61, 56, 
    72, 75, 75, 95, 82, 23, 25, 27, 21, 36, 51, 91, 79, 65, 58, 
    65, 72, 74, 76, 41, 0, 0, 4, 23, 3, 0, 0, 12, 31, 59, 
    77, 89, 90, 90, 87, 94, 60, 46, 69, 61, 52, 56, 40, 53, 59, 
    27, 31, 31, 31, 32, 28, 22, 23, 37, 36, 35, 36, 39, 42, 39, 
    27, 30, 33, 27, 30, 21, 21, 21, 26, 18, 17, 18, 16, 10, 0, 
    22, 16, 18, 16, 17, 7, 15, 13, 14, 13, 17, 19, 0, 11, 18, 
    
    -- channel=53
    0, 0, 26, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 44, 0, 3, 22, 0, 12, 9, 4, 0, 0, 0, 0, 
    0, 0, 5, 13, 13, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 28, 7, 0, 0, 4, 0, 3, 20, 0, 2, 0, 0, 0, 
    0, 0, 0, 17, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 34, 48, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 22, 75, 18, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 149, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 26, 156, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 44, 42, 77, 0, 0, 13, 43, 0, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 25, 0, 0, 1, 2, 0, 0, 0, 0, 0, 
    0, 2, 9, 5, 3, 7, 0, 0, 8, 0, 0, 0, 0, 3, 0, 
    16, 0, 6, 0, 7, 2, 0, 0, 4, 6, 0, 0, 0, 0, 0, 
    22, 3, 2, 0, 3, 0, 4, 0, 7, 5, 5, 5, 0, 0, 8, 
    
    -- channel=54
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 52, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 66, 15, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 20, 7, 0, 0, 48, 89, 59, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 7, 16, 0, 0, 9, 0, 0, 0, 0, 8, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 1, 15, 
    21, 32, 34, 26, 21, 20, 18, 13, 12, 2, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=55
    31, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    26, 0, 0, 0, 6, 0, 0, 2, 0, 0, 0, 5, 14, 0, 0, 
    25, 0, 0, 0, 0, 18, 0, 21, 5, 0, 5, 3, 18, 0, 0, 
    16, 1, 0, 0, 10, 3, 0, 8, 6, 0, 14, 4, 28, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 
    4, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 43, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 43, 42, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 7, 16, 25, 27, 10, 11, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 17, 9, 0, 0, 30, 23, 31, 15, 0, 
    24, 0, 0, 0, 0, 0, 0, 50, 0, 0, 0, 0, 48, 0, 0, 
    19, 0, 0, 0, 0, 0, 2, 20, 0, 0, 1, 2, 0, 0, 3, 
    3, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 31, 
    0, 0, 0, 1, 0, 8, 0, 2, 0, 0, 0, 0, 21, 11, 0, 
    
    -- channel=56
    1, 0, 3, 8, 5, 4, 7, 7, 8, 7, 8, 8, 9, 13, 10, 
    0, 0, 3, 26, 46, 44, 41, 39, 42, 42, 36, 24, 17, 11, 11, 
    0, 0, 6, 31, 34, 37, 39, 36, 30, 33, 37, 33, 16, 9, 8, 
    2, 0, 5, 38, 29, 26, 25, 31, 30, 30, 29, 31, 22, 8, 3, 
    6, 0, 0, 3, 1, 0, 0, 2, 3, 1, 3, 0, 10, 4, 4, 
    9, 5, 0, 0, 8, 7, 9, 10, 11, 9, 9, 5, 3, 4, 6, 
    8, 4, 4, 0, 0, 0, 6, 7, 9, 9, 7, 7, 4, 4, 3, 
    9, 7, 17, 28, 12, 0, 0, 7, 8, 7, 7, 7, 6, 4, 2, 
    13, 11, 11, 16, 25, 6, 0, 0, 0, 5, 3, 8, 7, 5, 3, 
    14, 12, 10, 16, 13, 4, 6, 12, 3, 0, 0, 0, 0, 3, 5, 
    10, 9, 11, 12, 29, 29, 9, 19, 30, 22, 22, 15, 13, 11, 7, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 7, 9, 10, 12, 10, 8, 3, 2, 2, 0, 0, 0, 0, 0, 
    4, 0, 2, 3, 4, 2, 3, 5, 7, 6, 6, 8, 6, 2, 1, 
    14, 7, 7, 7, 8, 9, 13, 12, 13, 13, 13, 10, 2, 7, 0, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=58
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=59
    0, 0, 9, 0, 0, 0, 1, 2, 7, 3, 1, 0, 7, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 25, 7, 17, 29, 27, 24, 10, 0, 0, 0, 
    0, 0, 0, 23, 0, 6, 13, 4, 0, 0, 0, 0, 2, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 35, 30, 28, 25, 28, 24, 21, 2, 0, 0, 0, 
    0, 23, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 32, 109, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 136, 167, 110, 119, 137, 132, 143, 122, 81, 32, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 
    0, 0, 0, 0, 0, 13, 19, 16, 18, 21, 7, 0, 19, 44, 0, 
    
    -- channel=60
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 19, 2, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 16, 15, 13, 17, 8, 6, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 21, 27, 4, 0, 14, 14, 25, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 7, 7, 14, 14, 13, 12, 15, 16, 17, 19, 20, 20, 25, 32, 
    10, 18, 17, 19, 18, 20, 17, 23, 21, 20, 19, 22, 34, 23, 21, 
    
    -- channel=61
    41, 54, 51, 33, 39, 37, 36, 31, 31, 32, 34, 33, 25, 35, 40, 
    49, 67, 59, 20, 0, 19, 18, 9, 19, 22, 22, 14, 46, 46, 41, 
    49, 65, 67, 11, 17, 0, 0, 0, 12, 13, 11, 14, 40, 49, 45, 
    50, 62, 63, 0, 0, 0, 5, 0, 0, 0, 0, 5, 0, 47, 53, 
    52, 62, 58, 65, 48, 51, 44, 46, 50, 49, 41, 40, 45, 55, 54, 
    48, 66, 73, 49, 47, 43, 43, 45, 43, 45, 43, 52, 56, 51, 48, 
    43, 50, 37, 53, 57, 58, 51, 53, 50, 53, 52, 55, 56, 56, 55, 
    43, 53, 32, 15, 35, 47, 54, 50, 52, 51, 48, 50, 52, 53, 54, 
    42, 47, 47, 38, 43, 13, 33, 51, 58, 60, 49, 49, 52, 54, 54, 
    40, 43, 46, 58, 58, 16, 4, 2, 19, 45, 55, 66, 61, 56, 51, 
    40, 45, 46, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 39, 
    70, 82, 82, 82, 84, 72, 68, 73, 80, 68, 74, 66, 81, 80, 74, 
    25, 29, 29, 28, 25, 27, 32, 44, 51, 52, 55, 56, 59, 63, 56, 
    20, 24, 22, 13, 12, 12, 12, 9, 7, 6, 2, 3, 4, 1, 0, 
    0, 4, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 
    
    -- channel=62
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 18, 15, 8, 16, 16, 15, 8, 0, 0, 0, 0, 
    0, 0, 0, 9, 9, 22, 27, 27, 16, 18, 15, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 15, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 3, 0, 0, 0, 18, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=63
    0, 0, 0, 6, 0, 0, 0, 2, 0, 0, 0, 0, 7, 2, 3, 
    0, 0, 0, 22, 23, 24, 24, 31, 29, 22, 23, 35, 0, 0, 3, 
    0, 0, 0, 50, 0, 4, 23, 11, 5, 5, 3, 14, 0, 0, 0, 
    0, 0, 0, 20, 4, 6, 1, 0, 4, 0, 2, 0, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 1, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 20, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 9, 7, 8, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 32, 0, 0, 25, 0, 24, 0, 4, 6, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 1, 2, 5, 7, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 7, 8, 4, 5, 7, 7, 8, 10, 9, 8, 6, 10, 
    21, 8, 7, 8, 11, 7, 11, 14, 13, 15, 17, 13, 6, 11, 0, 
    
    -- channel=64
    0, 0, 0, 3, 6, 0, 0, 0, 7, 10, 13, 0, 22, 0, 0, 
    8, 0, 3, 8, 5, 0, 0, 0, 2, 4, 8, 0, 7, 0, 16, 
    31, 23, 7, 16, 6, 0, 0, 9, 10, 20, 0, 0, 26, 13, 9, 
    1, 0, 9, 18, 0, 0, 8, 7, 0, 7, 0, 11, 34, 24, 40, 
    11, 2, 28, 0, 1, 4, 7, 0, 0, 0, 14, 4, 24, 30, 36, 
    22, 9, 24, 14, 0, 13, 4, 14, 14, 14, 3, 1, 29, 33, 26, 
    11, 5, 24, 30, 23, 15, 12, 20, 20, 20, 20, 25, 19, 21, 16, 
    21, 8, 27, 29, 27, 12, 18, 12, 20, 10, 21, 28, 42, 27, 34, 
    5, 15, 32, 26, 24, 46, 19, 27, 34, 33, 20, 42, 34, 39, 21, 
    28, 37, 29, 22, 34, 11, 42, 39, 29, 44, 32, 30, 35, 12, 0, 
    42, 6, 11, 0, 8, 36, 8, 48, 51, 38, 41, 26, 22, 8, 28, 
    0, 3, 6, 8, 26, 4, 40, 41, 43, 38, 30, 30, 20, 25, 23, 
    48, 36, 27, 9, 19, 17, 33, 52, 38, 38, 33, 34, 23, 11, 22, 
    21, 16, 23, 15, 6, 11, 11, 3, 3, 42, 39, 35, 37, 4, 2, 
    11, 0, 0, 21, 24, 12, 2, 10, 21, 31, 50, 26, 0, 0, 0, 
    
    -- channel=65
    0, 0, 15, 0, 0, 47, 0, 17, 0, 0, 0, 56, 0, 17, 3, 
    0, 5, 0, 0, 0, 22, 0, 32, 0, 6, 0, 70, 0, 49, 0, 
    0, 0, 0, 0, 0, 44, 26, 0, 0, 0, 4, 72, 0, 0, 0, 
    0, 51, 0, 0, 19, 37, 0, 0, 47, 0, 44, 39, 0, 0, 0, 
    0, 54, 0, 0, 32, 0, 0, 58, 4, 24, 0, 10, 0, 0, 0, 
    0, 48, 0, 0, 35, 1, 0, 15, 0, 0, 0, 53, 0, 0, 0, 
    0, 34, 19, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 9, 0, 
    0, 20, 7, 0, 0, 0, 5, 4, 0, 8, 5, 14, 0, 0, 0, 
    9, 14, 0, 0, 13, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 29, 0, 2, 0, 0, 0, 0, 0, 0, 36, 
    0, 18, 0, 17, 13, 0, 53, 0, 0, 0, 0, 0, 0, 9, 2, 
    25, 29, 0, 18, 0, 25, 4, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 4, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 6, 14, 0, 0, 0, 0, 0, 46, 0, 0, 0, 0, 19, 0, 
    0, 0, 55, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 76, 
    
    -- channel=66
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 13, 5, 9, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 16, 14, 7, 9, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 2, 9, 17, 11, 6, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 1, 2, 5, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 9, 11, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 7, 10, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 9, 1, 0, 10, 7, 0, 0, 
    0, 0, 12, 0, 0, 0, 0, 0, 0, 6, 4, 11, 4, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 2, 10, 3, 7, 0, 0, 0, 
    
    -- channel=67
    126, 83, 94, 104, 98, 16, 116, 87, 157, 141, 160, 100, 229, 66, 99, 
    164, 134, 144, 124, 92, 41, 77, 77, 146, 136, 155, 110, 238, 111, 180, 
    158, 115, 128, 129, 74, 28, 108, 149, 118, 150, 91, 147, 289, 193, 202, 
    116, 92, 173, 121, 48, 136, 185, 93, 74, 119, 150, 191, 280, 230, 248, 
    140, 151, 235, 134, 93, 207, 189, 49, 178, 165, 219, 191, 268, 241, 217, 
    149, 140, 234, 199, 174, 197, 178, 210, 239, 228, 216, 178, 278, 222, 211, 
    147, 149, 209, 263, 240, 213, 198, 229, 209, 211, 214, 248, 250, 226, 204, 
    158, 152, 206, 246, 246, 216, 206, 237, 247, 241, 242, 244, 288, 229, 186, 
    163, 209, 215, 210, 233, 246, 241, 259, 276, 268, 254, 265, 255, 210, 150, 
    216, 201, 167, 156, 194, 201, 253, 281, 286, 305, 256, 265, 229, 145, 126, 
    219, 132, 174, 150, 187, 195, 217, 322, 306, 281, 255, 250, 226, 168, 226, 
    181, 283, 260, 186, 214, 188, 265, 300, 295, 277, 263, 263, 231, 190, 217, 
    223, 238, 321, 282, 224, 198, 262, 269, 196, 271, 289, 264, 228, 134, 206, 
    172, 116, 184, 293, 306, 232, 213, 186, 186, 267, 267, 265, 191, 90, 158, 
    171, 73, 94, 213, 311, 324, 279, 244, 215, 208, 232, 190, 155, 150, 204, 
    
    -- channel=68
    23, 3, 3, 0, 16, 0, 15, 4, 34, 28, 41, 0, 79, 3, 12, 
    16, 15, 16, 5, 14, 0, 11, 0, 30, 15, 39, 0, 76, 2, 26, 
    41, 29, 14, 14, 6, 0, 3, 26, 6, 29, 29, 0, 84, 24, 50, 
    23, 0, 29, 14, 0, 18, 46, 9, 4, 16, 25, 22, 86, 40, 71, 
    16, 13, 47, 35, 5, 35, 39, 0, 27, 28, 59, 30, 68, 43, 70, 
    25, 19, 47, 16, 24, 46, 64, 31, 47, 47, 59, 26, 70, 41, 70, 
    23, 11, 31, 58, 71, 66, 65, 57, 75, 70, 62, 52, 72, 36, 59, 
    28, 17, 24, 64, 68, 59, 68, 91, 73, 62, 67, 79, 74, 54, 42, 
    22, 22, 39, 43, 62, 71, 68, 81, 78, 88, 99, 64, 108, 51, 30, 
    37, 38, 32, 38, 41, 78, 63, 76, 91, 92, 79, 88, 74, 32, 15, 
    47, 32, 33, 16, 23, 25, 67, 87, 91, 97, 78, 88, 74, 26, 35, 
    24, 46, 56, 18, 47, 33, 64, 104, 86, 89, 78, 95, 88, 40, 39, 
    58, 87, 93, 64, 39, 53, 70, 108, 69, 84, 93, 85, 90, 22, 40, 
    49, 31, 73, 87, 74, 43, 61, 51, 25, 86, 88, 97, 75, 23, 4, 
    58, 10, 23, 69, 97, 64, 63, 47, 71, 81, 90, 65, 30, 7, 36, 
    
    -- channel=69
    4, 20, 0, 0, 59, 0, 3, 0, 0, 0, 40, 0, 110, 0, 0, 
    0, 11, 9, 0, 64, 0, 0, 0, 4, 0, 39, 0, 98, 0, 13, 
    11, 0, 5, 5, 52, 0, 0, 7, 0, 37, 0, 0, 50, 0, 18, 
    34, 0, 22, 27, 0, 0, 23, 41, 0, 35, 0, 0, 19, 0, 73, 
    32, 0, 58, 23, 0, 0, 79, 0, 0, 0, 2, 0, 11, 0, 125, 
    56, 0, 0, 68, 0, 0, 32, 0, 8, 0, 19, 0, 33, 0, 131, 
    44, 0, 0, 13, 24, 0, 8, 0, 12, 0, 0, 0, 19, 0, 103, 
    28, 0, 0, 0, 0, 24, 0, 0, 4, 0, 8, 0, 47, 0, 90, 
    0, 0, 0, 0, 0, 44, 0, 0, 0, 0, 10, 0, 39, 18, 63, 
    0, 8, 22, 0, 0, 0, 3, 0, 0, 13, 3, 15, 47, 10, 0, 
    57, 0, 40, 0, 0, 9, 0, 4, 7, 18, 2, 11, 28, 0, 0, 
    0, 0, 54, 0, 11, 0, 0, 0, 4, 32, 0, 9, 33, 0, 0, 
    0, 0, 20, 30, 26, 0, 0, 29, 0, 4, 0, 35, 37, 0, 0, 
    38, 0, 0, 0, 43, 3, 0, 21, 0, 0, 0, 35, 73, 0, 0, 
    55, 23, 0, 0, 0, 28, 18, 0, 11, 0, 0, 15, 42, 0, 0, 
    
    -- channel=70
    0, 0, 0, 0, 0, 2, 0, 0, 0, 2, 0, 0, 0, 9, 8, 
    0, 0, 0, 0, 0, 0, 12, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 1, 0, 0, 0, 0, 1, 22, 0, 0, 0, 0, 
    3, 0, 0, 0, 10, 0, 0, 17, 12, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 
    0, 0, 0, 2, 0, 28, 0, 0, 0, 0, 0, 0, 0, 2, 17, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 25, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 20, 0, 
    0, 33, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 
    0, 0, 22, 3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    
    -- channel=71
    0, 0, 6, 0, 0, 47, 0, 12, 0, 6, 0, 57, 0, 30, 4, 
    0, 0, 0, 0, 0, 24, 2, 24, 0, 0, 0, 69, 0, 21, 0, 
    0, 9, 0, 0, 0, 39, 1, 0, 16, 0, 33, 53, 0, 0, 0, 
    0, 50, 0, 0, 1, 17, 0, 0, 42, 0, 21, 24, 0, 0, 0, 
    0, 63, 0, 0, 50, 0, 0, 44, 0, 6, 0, 10, 0, 0, 0, 
    0, 64, 0, 0, 1, 0, 0, 15, 0, 0, 0, 39, 0, 0, 0, 
    0, 29, 12, 0, 0, 0, 0, 0, 0, 4, 8, 0, 0, 1, 0, 
    0, 24, 3, 0, 0, 0, 24, 2, 0, 0, 0, 26, 0, 1, 0, 
    2, 0, 0, 0, 3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 1, 11, 10, 5, 0, 0, 0, 0, 0, 0, 28, 
    0, 31, 0, 17, 0, 0, 46, 0, 0, 0, 0, 0, 0, 2, 0, 
    10, 0, 0, 0, 0, 10, 12, 0, 0, 0, 8, 0, 0, 19, 0, 
    0, 48, 0, 0, 0, 13, 0, 0, 41, 0, 0, 0, 0, 18, 0, 
    0, 13, 73, 0, 0, 0, 0, 0, 9, 4, 6, 0, 0, 43, 18, 
    0, 0, 38, 63, 0, 0, 0, 0, 0, 13, 0, 2, 0, 0, 40, 
    
    -- channel=72
    10, 9, 7, 0, 0, 4, 5, 2, 6, 0, 5, 4, 20, 0, 4, 
    4, 13, 3, 0, 2, 1, 0, 4, 6, 6, 4, 5, 20, 14, 9, 
    2, 0, 0, 0, 1, 5, 11, 8, 0, 2, 0, 7, 21, 6, 12, 
    0, 2, 11, 8, 7, 12, 5, 0, 2, 12, 19, 6, 13, 9, 9, 
    4, 0, 10, 12, 12, 14, 9, 10, 12, 10, 17, 3, 14, 5, 6, 
    8, 0, 1, 13, 13, 18, 37, 26, 21, 19, 18, 18, 11, 2, 14, 
    12, 3, 0, 15, 32, 31, 40, 33, 32, 30, 36, 34, 18, 5, 11, 
    3, 0, 4, 7, 27, 32, 26, 40, 40, 42, 37, 30, 38, 13, 1, 
    9, 8, 1, 0, 11, 34, 35, 36, 36, 32, 38, 31, 31, 16, 7, 
    9, 0, 1, 1, 0, 15, 28, 34, 38, 35, 34, 33, 25, 12, 1, 
    5, 10, 10, 2, 7, 4, 21, 33, 33, 34, 32, 35, 34, 13, 10, 
    17, 39, 29, 9, 5, 7, 22, 36, 32, 34, 36, 40, 35, 16, 0, 
    0, 5, 30, 26, 12, 11, 17, 27, 15, 34, 37, 37, 35, 8, 0, 
    10, 0, 0, 25, 27, 13, 9, 15, 17, 29, 34, 36, 18, 8, 0, 
    11, 6, 4, 0, 27, 25, 20, 9, 19, 21, 20, 15, 21, 11, 14, 
    
    -- channel=73
    0, 5, 0, 0, 7, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=74
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=75
    15, 27, 26, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    12, 33, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 33, 51, 8, 
    0, 0, 0, 0, 0, 45, 49, 0, 0, 0, 0, 0, 15, 6, 3, 
    0, 37, 10, 0, 32, 27, 0, 0, 0, 17, 38, 0, 0, 0, 0, 
    1, 0, 24, 0, 12, 0, 0, 55, 21, 24, 0, 0, 0, 0, 0, 
    0, 0, 0, 70, 28, 0, 13, 16, 6, 0, 0, 9, 0, 0, 0, 
    28, 0, 0, 0, 0, 0, 18, 0, 0, 0, 3, 3, 0, 0, 6, 
    0, 0, 0, 0, 17, 0, 0, 0, 12, 42, 10, 0, 21, 0, 0, 
    20, 12, 0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 5, 19, 
    0, 0, 3, 2, 5, 0, 0, 0, 0, 0, 0, 0, 2, 14, 9, 
    64, 96, 61, 3, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 32, 0, 0, 21, 17, 0, 0, 0, 0, 0, 0, 
    0, 11, 0, 0, 0, 36, 19, 0, 0, 0, 0, 0, 63, 53, 10, 
    
    -- channel=76
    29, 23, 42, 35, 12, 51, 32, 37, 41, 40, 21, 53, 6, 50, 29, 
    30, 25, 34, 31, 7, 48, 34, 43, 33, 38, 25, 61, 10, 46, 29, 
    17, 29, 27, 22, 9, 53, 48, 32, 42, 17, 45, 62, 15, 35, 24, 
    26, 61, 19, 19, 30, 63, 38, 26, 50, 17, 66, 54, 25, 28, 6, 
    19, 62, 12, 19, 46, 43, 19, 45, 52, 49, 43, 55, 31, 24, 0, 
    6, 59, 28, 11, 55, 33, 5, 42, 30, 40, 28, 50, 26, 31, 0, 
    11, 52, 40, 20, 18, 25, 21, 31, 19, 18, 20, 28, 21, 38, 0, 
    18, 46, 30, 23, 20, 13, 31, 15, 20, 24, 16, 24, 0, 30, 0, 
    31, 34, 25, 30, 30, 0, 24, 15, 19, 18, 11, 16, 2, 15, 10, 
    22, 24, 17, 33, 31, 32, 9, 14, 10, 10, 12, 11, 8, 23, 41, 
    10, 40, 22, 49, 32, 20, 40, 11, 6, 4, 14, 14, 13, 29, 36, 
    31, 45, 27, 49, 26, 37, 28, 14, 9, 0, 19, 11, 15, 32, 38, 
    29, 48, 33, 33, 36, 38, 27, 5, 22, 10, 17, 7, 11, 39, 35, 
    22, 47, 63, 43, 35, 47, 45, 30, 39, 17, 11, 2, 4, 37, 57, 
    17, 37, 70, 64, 42, 39, 47, 48, 24, 20, 15, 18, 18, 56, 69, 
    
    -- channel=77
    0, 0, 0, 9, 27, 0, 4, 0, 8, 2, 14, 0, 23, 0, 0, 
    2, 0, 10, 12, 18, 0, 8, 0, 1, 0, 14, 0, 0, 0, 13, 
    26, 2, 4, 18, 8, 0, 0, 15, 9, 27, 0, 0, 8, 4, 5, 
    14, 0, 6, 2, 0, 0, 14, 10, 0, 0, 0, 0, 18, 5, 51, 
    11, 0, 18, 7, 0, 0, 13, 0, 0, 0, 0, 0, 7, 18, 50, 
    16, 5, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 20, 34, 
    0, 1, 8, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 19, 
    7, 1, 1, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 36, 
    0, 0, 22, 17, 10, 0, 0, 0, 0, 0, 0, 0, 4, 12, 5, 
    15, 22, 15, 6, 20, 7, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    35, 0, 1, 1, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    34, 4, 0, 0, 0, 3, 11, 20, 0, 0, 0, 0, 0, 0, 19, 
    18, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 0, 0, 1, 18, 0, 0, 0, 0, 
    
    -- channel=78
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 2, 0, 1, 11, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 15, 11, 1, 0, 0, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 6, 2, 8, 5, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 0, 0, 2, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 5, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 1, 9, 1, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 11, 24, 0, 4, 0, 3, 0, 0, 
    0, 16, 10, 0, 0, 0, 0, 0, 0, 9, 9, 3, 0, 0, 0, 
    0, 0, 13, 2, 0, 0, 0, 0, 0, 9, 19, 0, 0, 0, 0, 
    
    -- channel=79
    1, 33, 4, 10, 4, 21, 9, 32, 13, 27, 8, 43, 0, 9, 27, 
    19, 47, 11, 9, 23, 9, 7, 34, 13, 24, 5, 33, 4, 23, 2, 
    11, 25, 16, 19, 31, 18, 24, 16, 15, 19, 3, 40, 4, 18, 12, 
    8, 1, 20, 11, 52, 15, 17, 27, 16, 32, 3, 42, 3, 21, 0, 
    26, 0, 3, 28, 34, 29, 13, 46, 12, 29, 19, 58, 16, 9, 0, 
    32, 0, 13, 27, 17, 35, 57, 16, 37, 37, 36, 57, 19, 10, 0, 
    37, 1, 31, 26, 46, 29, 45, 23, 40, 34, 38, 38, 40, 21, 19, 
    28, 10, 25, 14, 16, 55, 23, 44, 31, 33, 34, 30, 26, 18, 22, 
    31, 22, 29, 21, 21, 26, 34, 32, 22, 27, 47, 28, 26, 25, 21, 
    19, 22, 25, 12, 3, 32, 24, 21, 38, 12, 41, 26, 6, 14, 33, 
    8, 28, 28, 5, 29, 12, 23, 18, 18, 27, 23, 30, 29, 32, 6, 
    47, 17, 39, 29, 19, 21, 14, 25, 22, 35, 10, 32, 38, 30, 28, 
    12, 31, 47, 51, 25, 31, 15, 14, 30, 27, 22, 30, 24, 52, 24, 
    2, 28, 23, 48, 46, 33, 27, 20, 32, 15, 30, 35, 13, 29, 19, 
    7, 5, 30, 26, 45, 47, 41, 22, 45, 11, 15, 22, 37, 7, 33, 
    
    -- channel=80
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 7, 
    13, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 3, 
    12, 4, 2, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    19, 4, 3, 2, 0, 2, 3, 0, 6, 0, 6, 12, 0, 3, 5, 
    0, 11, 0, 4, 5, 0, 31, 26, 24, 0, 17, 4, 0, 1, 1, 
    0, 14, 21, 19, 0, 28, 30, 11, 0, 8, 22, 7, 0, 0, 1, 
    9, 0, 27, 15, 20, 18, 17, 24, 34, 31, 26, 14, 0, 0, 2, 
    2, 12, 20, 31, 41, 24, 35, 34, 41, 48, 38, 2, 0, 3, 25, 
    12, 4, 34, 53, 0, 38, 26, 0, 16, 5, 0, 0, 0, 0, 32, 
    17, 17, 43, 19, 6, 13, 16, 20, 17, 9, 5, 0, 0, 7, 35, 
    12, 20, 17, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 17, 15, 
    12, 11, 23, 10, 6, 20, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    17, 11, 20, 24, 16, 0, 5, 15, 0, 2, 0, 0, 0, 0, 3, 
    0, 12, 10, 4, 8, 7, 11, 9, 13, 3, 1, 0, 5, 4, 0, 
    
    -- channel=81
    0, 33, 0, 0, 0, 0, 0, 5, 0, 0, 1, 0, 11, 20, 0, 
    0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 11, 4, 6, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 33, 0, 3, 0, 2, 
    0, 4, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 3, 
    0, 7, 0, 0, 3, 0, 0, 1, 0, 10, 0, 0, 6, 0, 0, 
    61, 0, 18, 0, 0, 25, 0, 0, 0, 14, 0, 0, 14, 0, 6, 
    83, 13, 0, 0, 17, 0, 0, 0, 38, 16, 0, 0, 14, 7, 1, 
    0, 65, 0, 0, 17, 0, 0, 1, 0, 0, 0, 0, 19, 23, 0, 
    0, 52, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 47, 37, 0, 
    0, 63, 0, 0, 48, 0, 0, 26, 0, 0, 2, 0, 38, 63, 0, 
    0, 31, 0, 0, 21, 0, 0, 11, 0, 0, 0, 0, 26, 63, 0, 
    0, 6, 0, 0, 0, 19, 29, 0, 0, 0, 0, 11, 26, 22, 0, 
    7, 0, 0, 9, 0, 0, 9, 0, 0, 4, 2, 22, 30, 3, 20, 
    0, 19, 0, 0, 0, 8, 22, 0, 5, 0, 8, 24, 9, 22, 0, 
    2, 20, 0, 14, 1, 4, 0, 0, 0, 0, 11, 10, 0, 0, 18, 
    
    -- channel=82
    49, 37, 63, 65, 72, 72, 68, 54, 36, 21, 25, 24, 25, 21, 20, 
    51, 62, 71, 68, 73, 78, 81, 75, 63, 25, 25, 27, 29, 31, 28, 
    43, 59, 67, 74, 74, 82, 84, 83, 76, 40, 26, 33, 38, 38, 32, 
    45, 45, 68, 70, 76, 87, 83, 77, 71, 73, 63, 53, 39, 39, 37, 
    30, 50, 65, 75, 81, 77, 58, 54, 55, 71, 63, 43, 35, 33, 35, 
    41, 49, 61, 65, 68, 51, 9, 19, 43, 42, 41, 32, 18, 33, 35, 
    11, 50, 42, 48, 45, 32, 36, 19, 5, 15, 20, 10, 7, 31, 30, 
    33, 30, 39, 36, 31, 30, 46, 31, 11, 12, 14, 5, 4, 19, 17, 
    49, 27, 30, 31, 37, 47, 45, 55, 44, 34, 31, 16, 7, 25, 15, 
    54, 35, 15, 27, 12, 29, 44, 31, 37, 20, 7, 4, 6, 21, 1, 
    51, 38, 22, 23, 12, 25, 40, 59, 45, 19, 9, 13, 16, 19, 8, 
    53, 44, 24, 29, 20, 14, 20, 23, 10, 0, 0, 0, 23, 26, 28, 
    56, 52, 40, 30, 40, 45, 48, 31, 6, 0, 0, 0, 1, 24, 31, 
    50, 50, 44, 42, 31, 43, 44, 51, 33, 17, 20, 17, 18, 24, 17, 
    53, 42, 52, 44, 39, 46, 57, 53, 51, 50, 49, 50, 46, 44, 37, 
    
    -- channel=83
    201, 188, 196, 190, 194, 185, 168, 157, 153, 97, 106, 113, 98, 124, 127, 
    234, 237, 195, 209, 210, 202, 194, 179, 164, 95, 89, 116, 137, 150, 118, 
    257, 207, 218, 221, 226, 227, 214, 183, 192, 170, 141, 148, 137, 132, 141, 
    219, 231, 226, 225, 243, 233, 226, 202, 197, 208, 193, 168, 120, 116, 141, 
    203, 215, 234, 233, 234, 235, 215, 213, 208, 178, 200, 198, 105, 134, 140, 
    63, 245, 230, 252, 238, 219, 294, 230, 191, 170, 200, 135, 89, 113, 126, 
    121, 206, 289, 263, 218, 296, 253, 222, 203, 228, 210, 110, 77, 103, 122, 
    171, 168, 283, 245, 268, 305, 280, 279, 296, 288, 246, 122, 70, 138, 153, 
    183, 198, 279, 248, 262, 240, 291, 228, 227, 226, 166, 52, 46, 162, 192, 
    200, 188, 292, 265, 113, 248, 238, 199, 235, 99, 62, 81, 66, 168, 256, 
    223, 198, 274, 197, 72, 91, 99, 144, 129, 67, 53, 53, 86, 163, 269, 
    200, 211, 214, 201, 170, 114, 138, 143, 45, 15, 17, 18, 42, 133, 183, 
    192, 211, 218, 208, 212, 185, 150, 162, 105, 65, 43, 28, 68, 70, 132, 
    204, 172, 225, 183, 189, 156, 186, 199, 146, 152, 125, 135, 136, 134, 149, 
    174, 207, 201, 194, 196, 212, 197, 180, 179, 153, 165, 182, 191, 178, 139, 
    
    -- channel=84
    92, 72, 104, 107, 109, 104, 103, 75, 80, 45, 52, 47, 45, 53, 59, 
    110, 119, 100, 110, 117, 117, 113, 103, 95, 44, 47, 64, 65, 69, 59, 
    113, 108, 107, 119, 119, 125, 123, 115, 110, 66, 61, 67, 72, 74, 64, 
    92, 103, 115, 118, 126, 130, 131, 115, 111, 113, 92, 90, 67, 63, 71, 
    85, 104, 115, 113, 132, 124, 105, 97, 101, 109, 106, 102, 59, 69, 69, 
    41, 94, 117, 119, 120, 92, 94, 116, 94, 78, 94, 72, 48, 60, 64, 
    40, 95, 120, 113, 89, 103, 110, 71, 64, 67, 81, 46, 33, 53, 62, 
    69, 72, 118, 103, 91, 122, 107, 103, 101, 96, 97, 49, 24, 55, 62, 
    96, 67, 110, 97, 108, 97, 140, 114, 114, 111, 99, 35, 14, 62, 78, 
    97, 77, 106, 112, 84, 86, 121, 95, 91, 50, 29, 33, 25, 57, 92, 
    108, 81, 106, 99, 4, 62, 76, 92, 105, 32, 34, 41, 32, 58, 114, 
    103, 90, 89, 82, 61, 44, 51, 61, 24, 13, 7, 7, 30, 56, 95, 
    96, 100, 84, 108, 101, 81, 80, 75, 32, 8, 2, 0, 22, 32, 63, 
    105, 88, 114, 68, 101, 72, 88, 101, 69, 59, 49, 48, 49, 51, 70, 
    94, 91, 103, 90, 80, 99, 105, 103, 90, 85, 86, 90, 90, 88, 65, 
    
    -- channel=85
    57, 0, 7, 0, 16, 8, 19, 0, 48, 0, 0, 12, 4, 0, 33, 
    5, 22, 6, 7, 2, 11, 22, 3, 49, 24, 0, 0, 0, 15, 8, 
    32, 0, 2, 0, 1, 10, 23, 0, 15, 54, 0, 23, 0, 2, 3, 
    41, 0, 3, 0, 9, 8, 18, 17, 0, 10, 18, 45, 6, 0, 0, 
    0, 0, 3, 3, 3, 8, 9, 4, 27, 0, 4, 72, 0, 0, 0, 
    0, 13, 0, 4, 9, 0, 31, 3, 35, 0, 18, 65, 0, 0, 0, 
    0, 0, 13, 16, 0, 0, 31, 41, 0, 0, 55, 43, 0, 0, 0, 
    30, 0, 20, 0, 0, 19, 14, 0, 6, 11, 76, 47, 0, 0, 41, 
    26, 0, 10, 35, 0, 0, 49, 4, 0, 13, 71, 32, 0, 0, 101, 
    32, 0, 3, 127, 0, 0, 69, 0, 66, 30, 17, 17, 0, 0, 128, 
    31, 0, 13, 122, 0, 0, 0, 0, 55, 24, 1, 0, 0, 0, 100, 
    20, 0, 0, 48, 38, 10, 2, 39, 29, 6, 7, 0, 0, 0, 0, 
    0, 3, 11, 0, 46, 16, 0, 46, 40, 21, 22, 0, 0, 0, 0, 
    18, 0, 35, 0, 30, 0, 0, 39, 15, 21, 20, 0, 21, 0, 13, 
    7, 0, 22, 0, 18, 4, 9, 7, 13, 14, 0, 0, 16, 25, 0, 
    
    -- channel=86
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 4, 33, 26, 0, 0, 0, 
    0, 0, 0, 0, 45, 0, 0, 0, 0, 16, 4, 0, 0, 0, 0, 
    0, 0, 0, 12, 0, 68, 34, 20, 40, 0, 15, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 26, 29, 8, 9, 17, 0, 10, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=87
    0, 2, 0, 11, 0, 0, 0, 7, 0, 5, 10, 0, 9, 15, 0, 
    1, 0, 1, 1, 4, 2, 0, 7, 0, 0, 20, 8, 16, 0, 6, 
    0, 16, 0, 5, 6, 0, 0, 10, 2, 0, 8, 0, 8, 12, 8, 
    0, 0, 0, 11, 0, 1, 0, 2, 12, 4, 0, 0, 4, 18, 10, 
    0, 12, 2, 3, 3, 2, 4, 11, 0, 27, 14, 0, 21, 8, 11, 
    96, 0, 14, 0, 0, 41, 0, 0, 0, 28, 0, 0, 20, 9, 16, 
    55, 44, 0, 0, 16, 0, 0, 0, 9, 0, 0, 0, 12, 10, 8, 
    0, 71, 0, 0, 27, 0, 0, 17, 0, 0, 0, 0, 25, 24, 0, 
    0, 58, 0, 0, 29, 23, 0, 8, 12, 0, 0, 0, 46, 46, 0, 
    0, 62, 2, 0, 77, 18, 0, 43, 0, 0, 1, 0, 39, 72, 0, 
    0, 40, 0, 0, 17, 13, 16, 37, 0, 0, 7, 21, 23, 71, 0, 
    0, 14, 14, 0, 0, 5, 2, 0, 0, 4, 2, 17, 43, 21, 26, 
    14, 9, 0, 23, 0, 0, 23, 0, 0, 0, 0, 9, 14, 14, 24, 
    0, 36, 0, 12, 0, 12, 21, 0, 6, 0, 0, 7, 0, 4, 0, 
    13, 13, 0, 11, 0, 0, 4, 4, 0, 6, 14, 14, 0, 0, 18, 
    
    -- channel=88
    61, 64, 61, 66, 66, 66, 66, 56, 48, 31, 34, 36, 35, 39, 39, 
    59, 60, 61, 67, 70, 72, 74, 71, 62, 36, 29, 40, 45, 46, 41, 
    53, 51, 63, 66, 69, 70, 72, 70, 71, 62, 57, 53, 46, 45, 45, 
    45, 53, 61, 66, 70, 72, 74, 67, 63, 67, 64, 53, 41, 43, 44, 
    41, 55, 63, 64, 69, 64, 52, 57, 56, 57, 59, 47, 35, 41, 41, 
    22, 53, 61, 62, 58, 48, 45, 41, 37, 43, 46, 30, 27, 36, 39, 
    36, 42, 56, 52, 52, 51, 47, 49, 46, 43, 40, 28, 25, 34, 37, 
    48, 41, 54, 48, 47, 59, 65, 53, 46, 44, 48, 29, 22, 39, 41, 
    61, 48, 53, 46, 35, 37, 58, 42, 40, 33, 22, 16, 20, 34, 40, 
    58, 44, 45, 40, 17, 38, 50, 62, 57, 25, 26, 34, 29, 34, 42, 
    63, 47, 40, 37, 17, 6, 19, 32, 33, 21, 13, 23, 35, 31, 41, 
    57, 57, 41, 59, 60, 58, 56, 38, 14, 8, 6, 3, 16, 32, 35, 
    61, 60, 51, 43, 56, 46, 52, 60, 44, 29, 24, 19, 22, 22, 29, 
    54, 47, 60, 46, 44, 48, 55, 61, 54, 54, 53, 56, 54, 51, 44, 
    58, 63, 62, 63, 59, 64, 60, 57, 55, 55, 58, 59, 60, 56, 51, 
    
    -- channel=89
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 17, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 5, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 14, 23, 31, 19, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 25, 32, 29, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=90
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=91
    35, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 11, 0, 0, 
    0, 0, 0, 0, 0, 4, 1, 0, 13, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 54, 41, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 10, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 0, 0, 53, 73, 35, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 6, 0, 0, 0, 17, 0, 0, 28, 9, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 26, 7, 0, 21, 23, 0, 0, 35, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 0, 64, 31, 59, 44, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 10, 41, 48, 48, 43, 37, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 0, 23, 29, 42, 52, 52, 28, 0, 
    2, 12, 0, 14, 22, 6, 0, 0, 0, 0, 2, 1, 7, 4, 12, 
    
    -- channel=92
    12, 36, 26, 25, 26, 28, 22, 27, 12, 21, 20, 19, 21, 22, 6, 
    19, 23, 24, 30, 30, 27, 24, 28, 19, 18, 25, 16, 19, 14, 16, 
    16, 32, 28, 28, 29, 28, 24, 31, 23, 12, 30, 14, 18, 17, 17, 
    10, 34, 26, 30, 25, 26, 20, 23, 27, 22, 24, 10, 20, 22, 17, 
    22, 27, 26, 31, 28, 28, 19, 21, 15, 27, 18, 1, 23, 19, 19, 
    44, 27, 31, 24, 27, 34, 7, 9, 8, 29, 12, 2, 29, 20, 22, 
    51, 26, 18, 18, 27, 23, 9, 12, 30, 21, 0, 4, 26, 25, 21, 
    15, 45, 11, 20, 29, 12, 14, 18, 12, 14, 0, 0, 28, 32, 7, 
    6, 40, 11, 3, 29, 23, 0, 16, 12, 6, 0, 11, 36, 37, 0, 
    9, 38, 10, 0, 47, 19, 0, 29, 2, 11, 14, 15, 35, 47, 0, 
    3, 26, 10, 0, 35, 23, 13, 27, 0, 10, 17, 22, 26, 46, 0, 
    6, 14, 21, 3, 15, 14, 19, 15, 14, 20, 20, 30, 31, 25, 21, 
    11, 15, 13, 25, 0, 13, 16, 3, 10, 19, 19, 30, 34, 22, 30, 
    8, 17, 1, 17, 7, 20, 23, 2, 13, 10, 15, 24, 18, 22, 19, 
    13, 18, 6, 13, 11, 16, 14, 11, 14, 11, 18, 20, 12, 13, 17, 
    
    -- channel=93
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 15, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=94
    16, 35, 49, 58, 50, 56, 53, 45, 21, 31, 32, 25, 25, 36, 22, 
    42, 40, 50, 50, 56, 56, 57, 62, 31, 24, 37, 41, 41, 34, 32, 
    26, 42, 49, 56, 54, 58, 57, 67, 51, 16, 34, 33, 45, 44, 37, 
    19, 38, 50, 56, 56, 64, 62, 59, 65, 55, 42, 33, 40, 43, 40, 
    38, 42, 48, 48, 57, 48, 42, 36, 43, 68, 53, 22, 41, 40, 40, 
    62, 25, 41, 44, 47, 26, 7, 38, 31, 42, 36, 15, 37, 37, 41, 
    52, 49, 28, 30, 30, 26, 21, 0, 4, 8, 9, 11, 26, 31, 37, 
    25, 56, 27, 29, 25, 19, 32, 20, 9, 6, 0, 10, 26, 23, 18, 
    42, 43, 21, 24, 33, 33, 37, 47, 43, 41, 23, 16, 36, 28, 0, 
    41, 48, 15, 0, 56, 39, 30, 47, 20, 25, 17, 17, 40, 30, 0, 
    45, 50, 19, 0, 22, 41, 52, 61, 39, 22, 25, 30, 35, 50, 0, 
    50, 44, 27, 9, 17, 28, 33, 19, 16, 15, 8, 23, 38, 53, 23, 
    59, 43, 35, 45, 34, 41, 48, 24, 6, 0, 0, 3, 28, 30, 37, 
    49, 62, 42, 45, 36, 37, 54, 42, 33, 27, 22, 24, 19, 32, 25, 
    45, 51, 48, 47, 35, 46, 54, 54, 49, 47, 51, 49, 42, 38, 42, 
    
    -- channel=95
    69, 52, 50, 48, 48, 50, 56, 51, 37, 30, 25, 25, 32, 30, 34, 
    58, 47, 64, 50, 52, 60, 59, 53, 45, 36, 23, 35, 28, 26, 38, 
    38, 40, 57, 59, 54, 63, 55, 64, 63, 50, 42, 42, 26, 35, 33, 
    59, 39, 54, 59, 59, 66, 59, 59, 53, 56, 55, 44, 26, 32, 32, 
    49, 47, 53, 55, 63, 49, 39, 36, 45, 46, 57, 30, 28, 29, 27, 
    58, 40, 48, 53, 56, 52, 24, 31, 28, 26, 31, 32, 20, 30, 27, 
    22, 52, 38, 36, 63, 33, 57, 23, 24, 26, 30, 29, 23, 27, 22, 
    27, 37, 39, 51, 40, 52, 61, 29, 34, 27, 27, 26, 30, 22, 32, 
    44, 30, 39, 55, 0, 54, 43, 27, 27, 27, 17, 18, 31, 19, 22, 
    30, 40, 25, 14, 19, 28, 44, 26, 26, 32, 30, 14, 27, 23, 0, 
    35, 44, 16, 27, 2, 17, 20, 6, 37, 22, 11, 17, 27, 31, 3, 
    49, 29, 33, 53, 47, 49, 37, 4, 20, 17, 3, 1, 24, 36, 19, 
    48, 35, 40, 47, 61, 19, 32, 45, 33, 21, 17, 16, 13, 30, 7, 
    24, 45, 42, 43, 37, 31, 31, 39, 43, 41, 44, 36, 41, 38, 19, 
    40, 33, 46, 47, 46, 33, 39, 39, 37, 44, 40, 40, 44, 35, 48, 
    
    -- channel=96
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 24, 65, 66, 40, 44, 0, 0, 0, 
    0, 0, 0, 0, 0, 47, 63, 49, 30, 1, 50, 69, 4, 0, 0, 
    0, 0, 0, 0, 12, 9, 20, 0, 0, 27, 90, 95, 43, 0, 0, 
    0, 0, 8, 13, 36, 13, 0, 50, 105, 103, 121, 54, 0, 0, 32, 
    0, 0, 51, 21, 23, 2, 29, 81, 90, 117, 85, 56, 41, 66, 80, 
    0, 71, 69, 30, 5, 0, 17, 82, 121, 71, 53, 57, 104, 86, 69, 
    6, 31, 28, 22, 0, 17, 44, 87, 82, 14, 0, 27, 64, 66, 0, 
    0, 20, 31, 20, 0, 18, 54, 86, 71, 2, 16, 21, 43, 45, 0, 
    0, 19, 50, 53, 68, 92, 102, 106, 66, 31, 31, 11, 13, 3, 0, 
    0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 38, 8, 0, 0, 0, 
    
    -- channel=97
    29, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 3, 1, 
    0, 0, 0, 0, 0, 0, 2, 0, 3, 0, 17, 0, 0, 41, 4, 
    0, 0, 0, 0, 5, 5, 8, 7, 8, 20, 9, 0, 1, 34, 0, 
    5, 12, 11, 9, 13, 14, 12, 15, 14, 15, 0, 15, 14, 3, 0, 
    14, 13, 11, 8, 17, 16, 10, 12, 33, 3, 0, 37, 0, 0, 4, 
    14, 11, 11, 6, 23, 48, 55, 5, 0, 0, 0, 0, 29, 0, 4, 
    12, 10, 1, 20, 28, 0, 0, 0, 0, 97, 57, 0, 5, 4, 0, 
    11, 8, 34, 11, 0, 17, 0, 41, 115, 106, 0, 0, 0, 28, 51, 
    8, 26, 0, 0, 0, 4, 84, 69, 0, 0, 0, 0, 44, 78, 35, 
    40, 87, 0, 14, 0, 29, 96, 4, 0, 0, 0, 0, 30, 0, 0, 
    67, 0, 0, 0, 0, 46, 123, 0, 0, 0, 1, 52, 0, 0, 0, 
    13, 0, 0, 0, 24, 47, 81, 0, 0, 1, 0, 71, 0, 0, 0, 
    11, 8, 6, 0, 74, 42, 64, 0, 0, 37, 0, 7, 14, 0, 11, 
    10, 9, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 10, 
    8, 0, 9, 3, 12, 10, 7, 1, 0, 35, 0, 0, 4, 6, 16, 
    
    -- channel=98
    191, 208, 220, 226, 218, 199, 189, 178, 155, 123, 118, 87, 26, 30, 72, 
    211, 194, 187, 185, 170, 152, 146, 139, 126, 113, 94, 53, 8, 23, 83, 
    145, 145, 142, 136, 129, 120, 119, 118, 111, 108, 40, 0, 19, 51, 87, 
    110, 110, 111, 111, 115, 117, 115, 114, 110, 92, 9, 0, 58, 91, 98, 
    100, 111, 113, 112, 113, 105, 92, 93, 82, 50, 0, 0, 66, 94, 92, 
    109, 111, 112, 112, 100, 65, 0, 0, 0, 0, 0, 0, 2, 47, 81, 
    113, 112, 109, 98, 54, 7, 0, 0, 0, 0, 0, 0, 0, 0, 42, 
    111, 111, 77, 37, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    109, 88, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    96, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=99
    189, 188, 187, 186, 179, 156, 148, 139, 126, 127, 104, 86, 88, 32, 73, 
    168, 169, 163, 136, 124, 114, 112, 106, 98, 92, 86, 105, 45, 41, 82, 
    138, 124, 102, 99, 93, 96, 99, 98, 98, 96, 125, 97, 70, 88, 105, 
    79, 84, 93, 93, 95, 103, 108, 122, 121, 124, 122, 28, 97, 103, 83, 
    85, 90, 95, 98, 99, 117, 139, 143, 154, 195, 117, 80, 97, 83, 77, 
    91, 95, 97, 95, 94, 120, 205, 266, 293, 266, 265, 230, 28, 110, 75, 
    96, 101, 101, 84, 119, 178, 176, 100, 57, 38, 340, 331, 79, 51, 54, 
    100, 102, 85, 139, 131, 93, 132, 86, 155, 317, 411, 382, 114, 27, 86, 
    100, 90, 130, 96, 138, 57, 60, 328, 432, 418, 441, 221, 80, 132, 267, 
    79, 167, 254, 75, 72, 13, 92, 355, 365, 390, 292, 310, 292, 303, 291, 
    79, 254, 203, 97, 12, 10, 133, 346, 381, 136, 101, 157, 339, 278, 173, 
    81, 86, 160, 108, 7, 104, 187, 373, 332, 57, 58, 72, 210, 228, 14, 
    47, 91, 159, 109, 79, 206, 289, 350, 295, 71, 128, 62, 125, 116, 9, 
    56, 85, 137, 88, 113, 155, 173, 181, 125, 73, 119, 53, 28, 0, 0, 
    73, 74, 47, 55, 25, 29, 33, 26, 14, 31, 83, 18, 0, 0, 0, 
    
    -- channel=100
    190, 202, 217, 217, 210, 189, 184, 171, 144, 139, 114, 97, 57, 43, 79, 
    200, 190, 185, 177, 166, 149, 145, 136, 123, 113, 89, 71, 25, 28, 88, 
    153, 147, 143, 134, 125, 118, 120, 117, 113, 105, 80, 43, 28, 70, 100, 
    106, 109, 110, 112, 112, 117, 113, 118, 115, 99, 54, 5, 77, 101, 102, 
    101, 110, 113, 115, 114, 121, 111, 103, 77, 76, 24, 17, 82, 97, 93, 
    108, 112, 114, 114, 96, 72, 85, 89, 95, 91, 31, 29, 35, 68, 83, 
    112, 114, 115, 96, 86, 54, 58, 36, 29, 0, 52, 79, 0, 46, 58, 
    113, 114, 86, 64, 45, 24, 17, 0, 0, 0, 56, 130, 26, 0, 9, 
    113, 85, 46, 34, 32, 0, 0, 44, 73, 80, 88, 73, 6, 0, 34, 
    87, 54, 38, 0, 12, 0, 0, 55, 59, 102, 85, 47, 20, 41, 71, 
    66, 71, 55, 5, 0, 0, 0, 48, 96, 33, 2, 44, 62, 69, 57, 
    57, 0, 28, 12, 0, 0, 0, 51, 96, 0, 5, 0, 36, 56, 9, 
    38, 4, 13, 0, 0, 0, 4, 50, 81, 0, 7, 0, 26, 38, 2, 
    32, 19, 28, 15, 10, 50, 60, 64, 70, 0, 24, 10, 0, 4, 0, 
    39, 3, 0, 0, 0, 0, 0, 0, 0, 0, 20, 1, 0, 0, 0, 
    
    -- channel=101
    7, 20, 6, 17, 25, 21, 8, 28, 6, 31, 20, 11, 25, 0, 13, 
    9, 22, 21, 18, 16, 17, 7, 18, 12, 17, 0, 27, 43, 0, 15, 
    8, 19, 13, 16, 9, 12, 10, 12, 10, 3, 0, 32, 10, 0, 21, 
    8, 8, 11, 15, 6, 10, 7, 11, 7, 0, 65, 0, 4, 16, 18, 
    4, 10, 12, 14, 1, 1, 0, 0, 0, 39, 62, 0, 3, 10, 10, 
    8, 11, 14, 13, 0, 0, 0, 0, 0, 1, 0, 135, 0, 21, 11, 
    9, 13, 20, 0, 0, 0, 27, 43, 9, 0, 0, 192, 22, 0, 0, 
    10, 15, 0, 0, 34, 0, 22, 0, 0, 0, 0, 133, 85, 0, 0, 
    12, 0, 14, 0, 39, 0, 0, 0, 0, 0, 51, 165, 0, 0, 0, 
    0, 0, 140, 0, 58, 0, 0, 0, 0, 24, 0, 58, 0, 0, 33, 
    0, 0, 106, 22, 32, 0, 0, 0, 72, 92, 0, 0, 32, 42, 93, 
    0, 9, 0, 68, 0, 0, 0, 0, 181, 0, 25, 0, 0, 110, 16, 
    0, 0, 0, 61, 0, 0, 0, 0, 178, 0, 51, 0, 0, 111, 0, 
    0, 0, 0, 19, 0, 0, 0, 0, 86, 0, 30, 43, 0, 28, 0, 
    0, 17, 7, 20, 0, 0, 4, 8, 11, 0, 14, 43, 2, 0, 0, 
    
    -- channel=102
    0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 1, 0, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 22, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 0, 0, 
    0, 0, 0, 0, 0, 0, 49, 80, 64, 40, 0, 0, 0, 22, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 44, 0, 22, 38, 0, 0, 0, 0, 58, 0, 0, 0, 
    0, 0, 0, 6, 13, 16, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 6, 0, 25, 0, 0, 0, 0, 72, 45, 82, 0, 0, 27, 
    0, 13, 0, 0, 2, 0, 0, 0, 0, 0, 17, 2, 8, 0, 27, 
    8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 26, 6, 
    0, 3, 0, 16, 16, 65, 73, 78, 75, 0, 26, 20, 27, 46, 1, 
    0, 0, 20, 0, 0, 0, 0, 0, 8, 20, 0, 19, 4, 3, 1, 
    
    -- channel=103
    15, 15, 26, 25, 22, 24, 29, 17, 23, 18, 10, 17, 0, 22, 4, 
    35, 23, 13, 28, 28, 25, 26, 21, 20, 18, 36, 0, 0, 24, 7, 
    26, 19, 25, 23, 24, 22, 20, 19, 18, 23, 43, 0, 0, 14, 3, 
    22, 23, 21, 19, 21, 23, 27, 21, 17, 19, 0, 16, 5, 11, 11, 
    20, 22, 22, 21, 28, 31, 29, 30, 39, 0, 0, 0, 5, 12, 16, 
    22, 22, 20, 20, 40, 61, 42, 4, 4, 0, 30, 0, 40, 0, 12, 
    23, 20, 16, 36, 47, 9, 0, 0, 8, 106, 42, 0, 0, 21, 8, 
    22, 21, 52, 12, 0, 21, 0, 32, 34, 32, 0, 0, 0, 19, 44, 
    21, 48, 0, 23, 0, 20, 70, 63, 0, 0, 0, 0, 40, 40, 9, 
    52, 106, 0, 13, 0, 34, 108, 12, 0, 0, 33, 0, 0, 0, 0, 
    86, 10, 0, 0, 0, 55, 85, 0, 0, 0, 11, 113, 0, 0, 0, 
    44, 18, 10, 0, 26, 42, 90, 0, 0, 11, 0, 62, 32, 0, 2, 
    36, 24, 22, 0, 56, 8, 30, 0, 0, 37, 0, 0, 56, 0, 14, 
    19, 23, 0, 0, 18, 10, 10, 1, 0, 48, 0, 0, 9, 0, 12, 
    15, 6, 3, 0, 0, 1, 0, 0, 0, 30, 0, 0, 4, 5, 15, 
    
    -- channel=104
    149, 142, 138, 137, 128, 118, 113, 107, 93, 77, 77, 63, 28, 21, 61, 
    125, 118, 114, 109, 102, 94, 92, 88, 82, 81, 68, 50, 24, 38, 71, 
    85, 82, 86, 88, 85, 85, 86, 86, 84, 79, 47, 18, 36, 60, 72, 
    74, 82, 84, 85, 86, 89, 91, 88, 85, 69, 28, 14, 61, 74, 73, 
    79, 86, 87, 87, 85, 84, 71, 71, 62, 56, 26, 20, 51, 66, 69, 
    86, 86, 85, 84, 72, 57, 47, 36, 17, 5, 16, 23, 4, 42, 60, 
    86, 87, 83, 69, 55, 14, 0, 0, 0, 0, 6, 27, 7, 3, 32, 
    85, 83, 66, 44, 18, 15, 11, 6, 29, 28, 6, 20, 16, 5, 18, 
    84, 65, 27, 0, 1, 0, 0, 16, 8, 3, 10, 20, 21, 28, 18, 
    68, 50, 20, 0, 3, 0, 0, 0, 0, 4, 0, 19, 17, 6, 10, 
    55, 2, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    47, 3, 0, 5, 0, 0, 0, 3, 10, 0, 5, 0, 0, 4, 9, 
    34, 3, 0, 0, 0, 3, 0, 0, 12, 0, 10, 0, 0, 0, 7, 
    36, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 3, 
    32, 12, 0, 2, 0, 0, 0, 0, 2, 0, 0, 1, 3, 3, 3, 
    
    -- channel=105
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 1, 6, 
    0, 0, 0, 0, 0, 0, 0, 15, 2, 0, 0, 0, 15, 30, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 6, 0, 
    0, 0, 0, 7, 20, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 32, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 20, 37, 0, 0, 0, 0, 17, 23, 0, 0, 0, 24, 
    11, 3, 0, 18, 13, 0, 0, 0, 0, 9, 18, 22, 0, 3, 28, 
    16, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 14, 30, 40, 
    11, 18, 24, 40, 43, 41, 38, 38, 39, 14, 8, 33, 46, 45, 38, 
    
    -- channel=106
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=107
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 6, 0, 4, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 26, 14, 0, 
    0, 0, 0, 0, 0, 0, 11, 20, 16, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 9, 69, 110, 76, 25, 0, 0, 0, 
    0, 0, 0, 0, 0, 61, 78, 9, 0, 0, 87, 59, 0, 5, 0, 
    0, 0, 0, 0, 11, 0, 0, 0, 0, 7, 4, 95, 27, 0, 0, 
    0, 0, 28, 38, 0, 0, 10, 146, 240, 149, 4, 0, 0, 20, 90, 
    0, 19, 0, 0, 0, 0, 10, 37, 0, 0, 0, 0, 68, 135, 36, 
    19, 120, 50, 0, 0, 0, 0, 0, 0, 0, 0, 94, 91, 11, 0, 
    0, 0, 0, 0, 0, 55, 41, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 8, 31, 6, 0, 0, 0, 5, 13, 0, 0, 0, 0, 
    0, 0, 0, 49, 91, 114, 37, 0, 14, 18, 54, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 16, 44, 68, 38, 41, 32, 21, 16, 0, 0, 0, 8, 9, 12, 
    
    -- channel=108
    41, 39, 44, 42, 35, 32, 35, 28, 28, 25, 23, 25, 9, 20, 18, 
    37, 27, 28, 24, 22, 21, 25, 23, 22, 22, 34, 7, 8, 30, 20, 
    21, 17, 17, 16, 20, 18, 20, 23, 23, 26, 18, 3, 15, 31, 16, 
    18, 17, 18, 17, 19, 19, 23, 23, 23, 22, 2, 22, 18, 21, 18, 
    18, 16, 15, 15, 19, 18, 24, 27, 35, 10, 0, 22, 20, 16, 20, 
    17, 14, 15, 16, 25, 31, 15, 0, 0, 0, 6, 0, 29, 11, 15, 
    15, 13, 12, 22, 14, 13, 0, 0, 11, 44, 26, 0, 6, 25, 15, 
    14, 12, 25, 10, 6, 14, 11, 33, 41, 26, 0, 0, 0, 27, 33, 
    11, 24, 9, 8, 1, 25, 31, 26, 0, 0, 0, 0, 26, 13, 17, 
    25, 30, 0, 13, 0, 23, 39, 5, 0, 0, 0, 0, 0, 0, 0, 
    20, 10, 0, 2, 6, 37, 40, 0, 0, 0, 17, 28, 0, 0, 0, 
    18, 0, 12, 0, 26, 30, 27, 0, 0, 16, 7, 37, 0, 0, 8, 
    16, 13, 19, 0, 36, 16, 23, 0, 0, 27, 0, 8, 27, 0, 25, 
    15, 10, 7, 0, 13, 0, 0, 0, 0, 28, 0, 0, 30, 6, 26, 
    14, 13, 18, 10, 18, 18, 17, 16, 18, 31, 0, 5, 23, 25, 28, 
    
    -- channel=109
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 50, 58, 6, 27, 0, 0, 0, 
    0, 0, 0, 0, 0, 19, 46, 41, 15, 0, 39, 37, 9, 18, 0, 
    0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 55, 99, 13, 0, 0, 
    0, 0, 0, 9, 46, 18, 0, 25, 64, 53, 76, 12, 0, 0, 24, 
    0, 0, 39, 17, 23, 0, 0, 60, 53, 100, 64, 16, 21, 45, 56, 
    0, 75, 56, 32, 3, 0, 0, 57, 105, 50, 44, 42, 79, 71, 69, 
    0, 1, 42, 32, 0, 23, 10, 56, 91, 8, 7, 19, 42, 75, 0, 
    0, 13, 44, 14, 0, 5, 32, 50, 66, 3, 13, 12, 47, 45, 0, 
    0, 4, 60, 48, 73, 91, 96, 97, 66, 22, 35, 17, 30, 3, 0, 
    0, 0, 0, 2, 6, 5, 5, 5, 1, 13, 37, 6, 0, 0, 0, 
    
    -- channel=110
    154, 161, 175, 177, 167, 158, 154, 140, 130, 101, 93, 66, 33, 60, 73, 
    164, 152, 155, 156, 145, 134, 131, 120, 112, 101, 78, 49, 11, 55, 80, 
    134, 128, 131, 125, 119, 114, 113, 108, 101, 93, 48, 14, 29, 70, 83, 
    107, 110, 110, 108, 111, 108, 102, 97, 95, 78, 6, 33, 71, 86, 89, 
    104, 112, 113, 110, 110, 100, 88, 73, 43, 2, 0, 24, 65, 88, 89, 
    109, 112, 110, 107, 94, 46, 24, 26, 32, 1, 0, 0, 37, 49, 83, 
    112, 111, 104, 92, 66, 35, 0, 0, 4, 0, 0, 0, 0, 29, 60, 
    112, 105, 71, 35, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    110, 78, 25, 4, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    86, 21, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    81, 10, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 0, 0, 0, 
    57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 9, 
    46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    38, 8, 0, 0, 7, 9, 12, 10, 0, 0, 0, 0, 1, 0, 6, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 0, 
    
    -- channel=111
    108, 103, 102, 108, 100, 90, 85, 82, 70, 48, 61, 48, 0, 29, 46, 
    93, 92, 82, 77, 70, 65, 63, 62, 59, 59, 39, 34, 25, 30, 44, 
    57, 56, 62, 56, 58, 56, 56, 59, 58, 61, 3, 18, 35, 37, 43, 
    51, 56, 55, 57, 59, 57, 52, 56, 60, 49, 0, 35, 55, 47, 50, 
    50, 56, 56, 56, 56, 49, 36, 40, 34, 13, 17, 27, 20, 47, 45, 
    53, 55, 54, 53, 44, 30, 21, 18, 1, 3, 0, 27, 23, 9, 42, 
    56, 56, 48, 45, 24, 0, 0, 4, 0, 33, 0, 0, 26, 0, 23, 
    57, 52, 39, 15, 0, 22, 0, 0, 19, 5, 0, 0, 11, 15, 0, 
    52, 39, 7, 8, 0, 0, 52, 0, 0, 0, 0, 50, 0, 31, 0, 
    54, 0, 1, 0, 18, 14, 24, 0, 0, 1, 6, 1, 0, 0, 0, 
    57, 0, 0, 0, 19, 0, 18, 0, 0, 12, 0, 0, 0, 0, 0, 
    20, 18, 0, 3, 6, 0, 3, 0, 0, 0, 6, 9, 0, 0, 30, 
    23, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 14, 0, 16, 7, 
    20, 5, 0, 12, 0, 0, 0, 0, 0, 0, 0, 13, 0, 18, 2, 
    15, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 13, 5, 5, 7, 
    
    -- channel=112
    21, 21, 20, 28, 18, 7, 14, 17, 13, 11, 10, 8, 3, 0, 0, 
    21, 19, 19, 13, 5, 0, 0, 0, 6, 4, 0, 0, 0, 0, 1, 
    20, 18, 18, 15, 0, 0, 0, 0, 0, 5, 7, 10, 12, 18, 15, 
    13, 12, 5, 0, 0, 0, 0, 0, 0, 0, 10, 11, 12, 11, 2, 
    0, 5, 27, 3, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 
    41, 50, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 
    52, 51, 36, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 19, 
    39, 37, 44, 19, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    36, 36, 24, 27, 30, 31, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    38, 68, 97, 90, 32, 33, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    96, 104, 97, 31, 21, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    122, 93, 48, 23, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    43, 43, 30, 22, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 17, 23, 24, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=113
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 14, 13, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    29, 32, 0, 0, 4, 11, 0, 0, 0, 0, 0, 0, 0, 1, 2, 
    3, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 3, 0, 0, 0, 46, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    6, 16, 16, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39, 15, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 0, 1, 1, 0, 0, 0, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 19, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 12, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    
    -- channel=114
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 15, 11, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 28, 36, 46, 18, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 18, 31, 38, 46, 52, 26, 3, 9, 0, 0, 0, 
    0, 0, 0, 0, 14, 15, 16, 33, 53, 53, 44, 31, 11, 8, 10, 
    0, 0, 0, 0, 8, 8, 17, 30, 39, 47, 56, 44, 32, 23, 15, 
    0, 0, 0, 0, 0, 9, 21, 32, 27, 28, 45, 44, 39, 22, 5, 
    0, 0, 0, 0, 0, 0, 15, 33, 23, 18, 36, 46, 35, 17, 4, 
    0, 0, 0, 0, 0, 0, 8, 25, 24, 17, 28, 38, 31, 20, 23, 
    0, 0, 0, 0, 0, 4, 9, 29, 23, 15, 23, 33, 33, 32, 30, 
    0, 0, 0, 8, 15, 28, 29, 25, 26, 25, 28, 37, 36, 28, 24, 
    0, 0, 0, 0, 0, 23, 21, 4, 22, 28, 16, 25, 38, 33, 32, 
    0, 0, 0, 0, 0, 0, 10, 18, 7, 12, 2, 18, 41, 42, 32, 
    0, 0, 0, 12, 22, 16, 12, 16, 20, 19, 12, 18, 36, 46, 38, 
    0, 15, 28, 30, 31, 23, 24, 37, 37, 31, 25, 28, 38, 45, 42, 
    
    -- channel=115
    151, 146, 142, 157, 151, 150, 148, 126, 120, 109, 95, 80, 62, 53, 52, 
    147, 143, 139, 118, 142, 132, 140, 129, 109, 103, 97, 94, 97, 107, 109, 
    136, 134, 131, 94, 107, 100, 110, 110, 115, 154, 157, 159, 148, 141, 122, 
    126, 129, 120, 80, 84, 95, 100, 120, 134, 138, 159, 164, 137, 133, 115, 
    170, 210, 254, 115, 91, 110, 157, 148, 127, 127, 132, 147, 151, 156, 150, 
    274, 288, 280, 127, 103, 126, 173, 146, 134, 135, 132, 126, 150, 177, 173, 
    266, 265, 254, 202, 113, 133, 165, 141, 148, 150, 134, 117, 151, 153, 153, 
    243, 257, 280, 228, 219, 121, 171, 143, 167, 176, 141, 122, 127, 126, 127, 
    272, 296, 328, 320, 293, 264, 184, 181, 161, 172, 150, 134, 119, 139, 138, 
    378, 437, 450, 396, 283, 282, 186, 188, 159, 169, 168, 151, 124, 119, 76, 
    468, 469, 354, 221, 189, 172, 151, 141, 160, 168, 166, 142, 122, 117, 106, 
    395, 311, 230, 214, 159, 93, 114, 141, 100, 122, 152, 165, 131, 120, 134, 
    201, 195, 178, 178, 172, 146, 137, 127, 113, 134, 195, 174, 144, 118, 122, 
    150, 161, 173, 153, 115, 121, 120, 132, 119, 131, 147, 151, 141, 106, 112, 
    152, 125, 101, 90, 85, 126, 132, 113, 95, 93, 101, 118, 109, 86, 90, 
    
    -- channel=116
    24, 23, 21, 34, 42, 41, 35, 28, 20, 20, 15, 12, 6, 0, 0, 
    22, 24, 26, 23, 52, 53, 55, 38, 25, 19, 14, 13, 11, 12, 17, 
    23, 24, 35, 26, 49, 48, 56, 57, 35, 32, 35, 41, 38, 38, 37, 
    21, 17, 19, 24, 39, 40, 50, 66, 59, 60, 55, 52, 38, 38, 37, 
    15, 25, 65, 32, 38, 42, 53, 64, 71, 64, 67, 62, 45, 54, 53, 
    51, 63, 83, 31, 28, 35, 61, 67, 62, 69, 70, 56, 60, 70, 67, 
    60, 61, 63, 36, 50, 51, 70, 59, 57, 64, 71, 55, 62, 65, 58, 
    49, 53, 71, 72, 38, 22, 60, 63, 60, 65, 67, 58, 58, 39, 43, 
    51, 49, 60, 61, 83, 76, 75, 68, 57, 63, 63, 62, 48, 51, 62, 
    64, 82, 115, 131, 88, 111, 67, 78, 55, 58, 66, 66, 47, 49, 50, 
    103, 122, 90, 94, 77, 88, 65, 68, 63, 64, 67, 64, 50, 51, 50, 
    111, 94, 80, 57, 48, 43, 38, 34, 50, 50, 55, 60, 59, 59, 62, 
    61, 44, 45, 50, 60, 38, 47, 53, 41, 37, 57, 68, 65, 60, 69, 
    38, 44, 58, 61, 53, 57, 38, 60, 49, 45, 64, 58, 67, 62, 61, 
    52, 54, 55, 53, 46, 60, 59, 61, 55, 51, 45, 58, 62, 58, 60, 
    
    -- channel=117
    0, 4, 0, 0, 0, 0, 11, 7, 8, 5, 9, 12, 9, 0, 10, 
    0, 8, 0, 3, 1, 0, 7, 7, 9, 2, 4, 4, 1, 0, 8, 
    0, 2, 14, 0, 5, 0, 0, 0, 0, 0, 0, 4, 5, 8, 14, 
    0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 17, 5, 13, 9, 
    0, 0, 46, 38, 0, 0, 0, 11, 0, 0, 0, 0, 0, 11, 6, 
    0, 0, 69, 36, 0, 0, 5, 13, 0, 0, 0, 0, 0, 3, 13, 
    0, 0, 17, 89, 0, 0, 14, 0, 0, 7, 7, 0, 0, 0, 18, 
    0, 0, 6, 11, 69, 0, 16, 0, 0, 14, 11, 0, 0, 0, 10, 
    0, 0, 0, 37, 14, 50, 0, 15, 0, 7, 7, 8, 0, 0, 20, 
    0, 0, 1, 79, 0, 50, 0, 32, 0, 0, 2, 18, 0, 27, 11, 
    0, 22, 105, 19, 0, 15, 0, 0, 0, 0, 5, 16, 3, 5, 19, 
    21, 32, 40, 19, 45, 0, 0, 30, 0, 0, 0, 12, 16, 0, 41, 
    12, 0, 4, 1, 28, 18, 0, 21, 0, 0, 0, 8, 23, 0, 0, 
    1, 0, 6, 15, 6, 4, 2, 3, 2, 0, 0, 8, 12, 5, 0, 
    9, 13, 11, 12, 0, 0, 12, 18, 10, 7, 0, 1, 21, 1, 5, 
    
    -- channel=118
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 5, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 64, 16, 21, 0, 11, 0, 0, 0, 0, 0, 0, 0, 
    0, 37, 19, 0, 0, 19, 0, 0, 30, 9, 0, 0, 0, 0, 0, 
    23, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 14, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 
    0, 4, 15, 0, 0, 0, 0, 0, 0, 0, 1, 7, 3, 0, 0, 
    
    -- channel=119
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    8, 4, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 4, 5, 2, 0, 
    0, 0, 0, 0, 0, 20, 0, 0, 2, 0, 0, 5, 0, 10, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    2, 10, 0, 0, 0, 0, 8, 0, 2, 0, 0, 0, 1, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 18, 0, 11, 4, 0, 0, 0, 19, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 15, 0, 0, 0, 2, 12, 
    0, 0, 0, 0, 1, 6, 0, 0, 0, 4, 6, 0, 0, 0, 12, 
    0, 0, 0, 0, 15, 12, 0, 0, 0, 1, 3, 0, 0, 5, 7, 
    
    -- channel=120
    5, 6, 5, 10, 15, 15, 15, 11, 8, 8, 7, 6, 6, 6, 8, 
    5, 6, 6, 10, 21, 19, 23, 21, 14, 11, 14, 18, 20, 21, 21, 
    4, 5, 9, 11, 19, 23, 25, 27, 27, 25, 22, 23, 19, 17, 17, 
    6, 6, 14, 21, 16, 20, 27, 34, 30, 24, 23, 22, 20, 21, 25, 
    19, 25, 31, 24, 18, 19, 27, 32, 35, 33, 32, 27, 29, 37, 38, 
    19, 17, 18, 22, 18, 22, 22, 24, 29, 34, 34, 23, 30, 38, 34, 
    10, 12, 17, 27, 20, 14, 25, 26, 25, 29, 32, 26, 24, 24, 20, 
    13, 19, 24, 28, 35, 29, 33, 31, 26, 26, 30, 27, 20, 19, 27, 
    18, 20, 31, 38, 33, 38, 33, 36, 21, 21, 28, 27, 21, 25, 29, 
    35, 34, 28, 29, 19, 31, 29, 34, 22, 21, 28, 29, 20, 23, 32, 
    21, 24, 11, 7, 13, 17, 18, 22, 26, 24, 26, 26, 24, 32, 40, 
    0, 0, 15, 18, 17, 13, 16, 21, 13, 15, 25, 27, 31, 35, 40, 
    7, 5, 10, 21, 31, 29, 19, 24, 23, 17, 23, 24, 33, 38, 37, 
    13, 21, 23, 23, 24, 32, 30, 28, 28, 16, 13, 17, 24, 36, 37, 
    21, 22, 27, 34, 35, 36, 35, 37, 40, 36, 31, 30, 32, 38, 39, 
    
    -- channel=121
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 11, 15, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=122
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=123
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 18, 35, 41, 39, 29, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 13, 5, 0, 0, 0, 
    0, 0, 35, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    67, 76, 41, 5, 0, 0, 9, 0, 0, 0, 0, 0, 0, 14, 16, 
    4, 0, 0, 13, 15, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 73, 54, 13, 0, 0, 0, 0, 0, 0, 0, 4, 
    5, 29, 89, 75, 20, 24, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    86, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 4, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=124
    17, 16, 20, 14, 28, 33, 22, 22, 19, 19, 19, 18, 20, 23, 21, 
    17, 16, 21, 21, 36, 47, 41, 40, 26, 25, 26, 25, 24, 22, 18, 
    19, 19, 13, 30, 48, 59, 65, 61, 44, 30, 23, 22, 17, 14, 14, 
    22, 24, 16, 38, 62, 66, 67, 67, 58, 46, 37, 29, 18, 16, 21, 
    27, 24, 6, 23, 57, 64, 58, 57, 68, 64, 64, 48, 30, 20, 23, 
    14, 10, 0, 16, 50, 69, 53, 57, 66, 66, 68, 66, 40, 22, 17, 
    9, 7, 8, 0, 37, 51, 48, 64, 64, 57, 63, 70, 44, 28, 12, 
    16, 14, 8, 9, 13, 47, 44, 62, 62, 52, 63, 68, 57, 38, 20, 
    19, 21, 14, 2, 18, 11, 37, 49, 64, 55, 61, 65, 66, 35, 17, 
    10, 1, 0, 0, 33, 14, 47, 43, 64, 59, 59, 62, 63, 29, 20, 
    0, 0, 0, 25, 36, 43, 51, 46, 58, 57, 55, 60, 53, 32, 19, 
    0, 0, 0, 20, 30, 60, 55, 35, 61, 62, 55, 54, 40, 38, 15, 
    5, 14, 16, 17, 17, 30, 47, 36, 60, 66, 48, 50, 39, 35, 30, 
    20, 20, 20, 19, 23, 28, 38, 39, 46, 50, 49, 51, 44, 31, 32, 
    17, 20, 25, 25, 30, 32, 28, 28, 32, 36, 43, 39, 32, 30, 27, 
    
    -- channel=125
    12, 12, 7, 15, 0, 0, 0, 4, 6, 5, 6, 6, 2, 0, 0, 
    12, 11, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 11, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 15, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 18, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 1, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 47, 38, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 50, 48, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    84, 60, 9, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 23, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=126
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 1, 6, 7, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 3, 15, 11, 3, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 1, 11, 10, 8, 0, 3, 7, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 10, 8, 8, 17, 18, 14, 
    0, 0, 0, 0, 9, 14, 0, 0, 0, 0, 3, 10, 10, 16, 9, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 4, 1, 2, 4, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 12, 25, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 11, 30, 
    0, 0, 0, 0, 5, 0, 5, 13, 0, 0, 0, 0, 6, 15, 24, 
    0, 0, 0, 0, 0, 4, 0, 0, 4, 0, 0, 0, 14, 31, 17, 
    0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 10, 32, 27, 
    0, 0, 6, 17, 21, 12, 6, 13, 13, 13, 1, 0, 14, 35, 37, 
    11, 21, 25, 29, 37, 25, 20, 29, 32, 24, 23, 25, 27, 42, 40, 
    
    -- channel=127
    10, 11, 10, 13, 22, 26, 21, 13, 12, 11, 11, 11, 11, 10, 12, 
    10, 9, 6, 35, 28, 40, 37, 31, 21, 14, 19, 21, 22, 17, 17, 
    10, 8, 12, 26, 39, 48, 50, 57, 44, 20, 23, 20, 21, 13, 16, 
    13, 9, 7, 42, 45, 43, 55, 62, 51, 38, 33, 25, 18, 21, 25, 
    21, 22, 0, 53, 48, 37, 42, 61, 59, 59, 54, 40, 25, 35, 34, 
    14, 14, 0, 60, 34, 39, 46, 54, 49, 64, 58, 50, 41, 30, 27, 
    11, 14, 15, 25, 35, 40, 49, 54, 40, 52, 56, 63, 34, 18, 16, 
    16, 19, 15, 44, 14, 48, 43, 58, 43, 47, 58, 56, 33, 27, 31, 
    18, 18, 21, 53, 13, 13, 30, 61, 44, 46, 55, 55, 46, 42, 23, 
    25, 15, 27, 9, 26, 5, 40, 62, 47, 49, 53, 58, 50, 33, 30, 
    9, 4, 33, 15, 41, 38, 39, 56, 49, 50, 47, 56, 54, 29, 33, 
    0, 0, 39, 17, 30, 50, 35, 29, 39, 49, 43, 44, 55, 36, 30, 
    22, 11, 16, 27, 35, 38, 29, 35, 45, 51, 29, 48, 45, 39, 33, 
    22, 26, 24, 26, 34, 27, 41, 43, 50, 40, 33, 46, 41, 42, 36, 
    22, 25, 34, 36, 39, 27, 37, 42, 44, 39, 44, 44, 42, 39, 31, 
    
    -- channel=128
    0, 0, 21, 25, 24, 14, 18, 12, 15, 27, 3, 24, 24, 24, 25, 
    0, 4, 14, 27, 39, 34, 34, 37, 46, 37, 10, 44, 38, 35, 34, 
    0, 6, 0, 28, 56, 69, 44, 41, 51, 23, 39, 50, 52, 45, 43, 
    0, 0, 1, 45, 61, 58, 37, 32, 20, 33, 64, 48, 73, 83, 61, 
    23, 33, 45, 42, 42, 68, 63, 56, 32, 41, 47, 59, 75, 62, 48, 
    48, 51, 54, 39, 48, 70, 70, 37, 33, 40, 57, 54, 73, 57, 35, 
    47, 46, 53, 42, 56, 46, 54, 39, 50, 52, 49, 59, 72, 60, 40, 
    49, 49, 53, 27, 57, 72, 50, 66, 51, 44, 69, 60, 75, 81, 61, 
    53, 39, 33, 49, 62, 58, 61, 54, 28, 52, 40, 44, 37, 62, 50, 
    44, 39, 56, 66, 66, 81, 77, 55, 49, 31, 49, 27, 25, 35, 51, 
    54, 59, 51, 59, 58, 69, 56, 72, 59, 58, 29, 26, 45, 41, 34, 
    58, 56, 49, 71, 75, 61, 50, 59, 62, 42, 23, 43, 44, 43, 33, 
    56, 44, 47, 74, 79, 50, 51, 60, 56, 41, 31, 39, 46, 39, 34, 
    55, 41, 35, 65, 52, 45, 54, 48, 41, 28, 26, 33, 32, 25, 30, 
    51, 34, 30, 66, 66, 58, 50, 36, 34, 18, 27, 28, 24, 25, 35, 
    
    -- channel=129
    0, 94, 8, 0, 0, 0, 0, 3, 0, 0, 72, 13, 0, 0, 0, 
    2, 52, 25, 3, 0, 0, 0, 0, 0, 0, 98, 0, 0, 0, 0, 
    1, 16, 71, 13, 17, 0, 0, 0, 0, 1, 36, 0, 0, 0, 0, 
    0, 87, 82, 0, 16, 0, 0, 0, 6, 52, 0, 27, 0, 0, 0, 
    0, 29, 0, 0, 39, 0, 0, 0, 2, 28, 13, 17, 0, 0, 2, 
    0, 0, 0, 0, 16, 0, 0, 0, 4, 27, 9, 22, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 15, 0, 4, 16, 21, 0, 0, 0, 
    0, 0, 0, 45, 0, 0, 0, 0, 0, 10, 0, 5, 0, 0, 0, 
    0, 0, 0, 33, 0, 0, 0, 0, 40, 0, 0, 0, 29, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 9, 0, 0, 
    0, 0, 4, 0, 0, 0, 8, 0, 0, 0, 0, 9, 0, 0, 0, 
    0, 0, 23, 0, 0, 0, 4, 0, 0, 0, 25, 0, 0, 0, 0, 
    0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 13, 0, 0, 9, 0, 0, 0, 0, 3, 0, 0, 12, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 7, 0, 
    
    -- channel=130
    0, 0, 32, 22, 11, 30, 31, 25, 9, 0, 0, 7, 30, 32, 36, 
    0, 0, 29, 14, 0, 0, 0, 3, 2, 0, 0, 0, 14, 22, 27, 
    0, 0, 10, 17, 0, 0, 0, 6, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 3, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 6, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 1, 1, 0, 0, 1, 0, 
    0, 2, 0, 0, 0, 0, 0, 7, 8, 4, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 1, 8, 7, 6, 0, 0, 0, 0, 0, 
    
    -- channel=131
    22, 46, 245, 271, 260, 252, 273, 267, 272, 215, 127, 313, 317, 316, 313, 
    23, 37, 195, 241, 290, 288, 271, 298, 323, 248, 196, 358, 351, 340, 335, 
    28, 34, 124, 250, 306, 337, 231, 231, 253, 210, 313, 349, 373, 369, 368, 
    162, 67, 254, 305, 287, 338, 283, 243, 194, 223, 345, 346, 421, 419, 360, 
    314, 302, 345, 300, 259, 338, 337, 276, 200, 226, 312, 387, 428, 395, 331, 
    352, 342, 357, 296, 301, 338, 322, 228, 234, 239, 310, 374, 441, 408, 333, 
    360, 339, 341, 290, 309, 275, 311, 238, 305, 276, 297, 379, 438, 432, 384, 
    363, 329, 319, 274, 357, 333, 297, 295, 265, 291, 323, 316, 377, 443, 378, 
    371, 294, 302, 325, 353, 372, 351, 316, 235, 278, 295, 260, 252, 319, 329, 
    377, 328, 347, 351, 354, 368, 356, 345, 312, 263, 303, 245, 246, 289, 284, 
    385, 363, 326, 370, 367, 363, 308, 344, 347, 323, 223, 263, 289, 276, 249, 
    380, 363, 320, 386, 394, 340, 331, 341, 345, 280, 228, 278, 285, 281, 243, 
    374, 347, 319, 377, 379, 241, 315, 329, 313, 250, 233, 253, 264, 240, 248, 
    367, 329, 290, 364, 360, 289, 324, 280, 255, 203, 224, 231, 223, 204, 246, 
    320, 300, 272, 336, 364, 342, 277, 234, 222, 168, 213, 225, 217, 222, 237, 
    
    -- channel=132
    0, 0, 104, 93, 89, 100, 102, 96, 84, 54, 25, 99, 114, 114, 118, 
    0, 0, 92, 72, 68, 75, 92, 88, 98, 83, 23, 103, 112, 116, 119, 
    0, 0, 48, 63, 70, 83, 65, 88, 94, 57, 59, 96, 103, 103, 103, 
    1, 0, 46, 89, 63, 87, 54, 56, 51, 39, 92, 80, 101, 113, 98, 
    93, 49, 92, 85, 50, 82, 94, 75, 52, 41, 84, 85, 114, 117, 89, 
    99, 88, 105, 82, 66, 81, 86, 58, 48, 38, 71, 94, 115, 118, 93, 
    102, 92, 108, 89, 63, 61, 84, 49, 69, 52, 68, 89, 114, 117, 90, 
    108, 93, 107, 81, 89, 68, 78, 60, 77, 67, 85, 112, 106, 126, 100, 
    108, 77, 96, 70, 87, 73, 65, 88, 59, 72, 97, 63, 79, 119, 96, 
    107, 75, 87, 90, 82, 100, 91, 76, 62, 79, 95, 87, 62, 88, 76, 
    103, 92, 81, 87, 91, 90, 78, 87, 105, 98, 74, 74, 79, 87, 83, 
    101, 105, 71, 97, 104, 101, 81, 87, 97, 94, 62, 80, 85, 85, 71, 
    103, 108, 72, 90, 112, 69, 102, 97, 103, 85, 70, 76, 85, 79, 73, 
    105, 104, 67, 89, 103, 71, 99, 92, 93, 65, 68, 69, 73, 57, 78, 
    98, 98, 63, 80, 93, 102, 99, 82, 80, 52, 63, 71, 63, 65, 71, 
    
    -- channel=133
    6, 0, 0, 10, 2, 0, 1, 0, 29, 69, 0, 0, 0, 0, 5, 
    3, 0, 0, 0, 0, 10, 0, 0, 9, 94, 0, 0, 4, 2, 6, 
    3, 0, 0, 0, 0, 74, 2, 0, 8, 0, 0, 0, 0, 0, 1, 
    63, 0, 0, 31, 0, 37, 39, 28, 0, 0, 0, 0, 1, 22, 0, 
    36, 0, 0, 61, 0, 0, 27, 54, 0, 0, 0, 0, 2, 54, 0, 
    6, 0, 8, 37, 0, 0, 41, 29, 0, 0, 0, 0, 1, 52, 0, 
    7, 0, 36, 0, 8, 0, 38, 0, 17, 0, 0, 0, 0, 21, 24, 
    20, 0, 72, 0, 20, 1, 16, 16, 0, 0, 9, 0, 0, 14, 0, 
    45, 0, 11, 0, 3, 0, 19, 58, 0, 20, 0, 35, 0, 4, 0, 
    28, 0, 0, 0, 0, 0, 0, 28, 38, 0, 26, 0, 0, 6, 0, 
    4, 31, 0, 1, 0, 43, 0, 0, 27, 33, 0, 0, 0, 24, 2, 
    0, 42, 0, 0, 13, 22, 0, 0, 17, 61, 0, 1, 0, 23, 24, 
    6, 25, 0, 0, 53, 0, 0, 3, 28, 31, 0, 4, 0, 2, 8, 
    15, 27, 0, 0, 44, 0, 15, 8, 25, 12, 0, 2, 24, 0, 0, 
    13, 13, 0, 0, 16, 25, 33, 0, 35, 0, 0, 0, 14, 0, 0, 
    
    -- channel=134
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 15, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 23, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=135
    3, 81, 30, 0, 0, 11, 0, 8, 0, 0, 81, 0, 0, 0, 0, 
    4, 48, 55, 19, 4, 0, 10, 8, 0, 0, 87, 0, 0, 0, 0, 
    1, 18, 87, 9, 34, 0, 0, 16, 0, 24, 21, 2, 0, 0, 0, 
    0, 40, 34, 0, 50, 0, 0, 0, 4, 46, 0, 30, 0, 0, 6, 
    0, 10, 0, 0, 47, 0, 0, 0, 10, 30, 19, 21, 0, 0, 3, 
    0, 0, 0, 0, 20, 0, 0, 0, 3, 22, 11, 35, 0, 0, 0, 
    0, 0, 0, 23, 0, 6, 0, 17, 0, 7, 10, 28, 0, 0, 0, 
    0, 0, 0, 69, 0, 0, 0, 0, 20, 0, 0, 11, 36, 0, 0, 
    0, 0, 0, 17, 0, 0, 0, 0, 18, 0, 0, 0, 31, 0, 37, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 6, 9, 0, 7, 
    0, 0, 20, 0, 0, 0, 17, 0, 0, 0, 10, 5, 0, 0, 0, 
    0, 0, 28, 0, 0, 0, 6, 0, 0, 0, 26, 0, 8, 0, 0, 
    0, 0, 16, 0, 0, 1, 18, 0, 0, 0, 18, 0, 0, 2, 0, 
    0, 0, 17, 6, 0, 0, 0, 0, 0, 0, 8, 0, 0, 19, 4, 
    0, 0, 0, 25, 0, 0, 0, 2, 0, 22, 0, 2, 0, 3, 2, 
    
    -- channel=136
    5, 8, 41, 39, 34, 39, 45, 41, 38, 31, 16, 47, 54, 54, 55, 
    5, 5, 28, 30, 27, 28, 30, 36, 38, 37, 27, 38, 44, 48, 50, 
    7, 5, 17, 32, 23, 26, 17, 18, 17, 20, 25, 22, 29, 32, 36, 
    36, 26, 39, 29, 15, 27, 33, 27, 21, 18, 26, 24, 35, 33, 24, 
    40, 35, 33, 29, 17, 19, 28, 24, 17, 15, 25, 24, 33, 35, 25, 
    33, 30, 30, 32, 24, 21, 21, 19, 21, 16, 22, 20, 29, 35, 29, 
    32, 32, 35, 29, 19, 15, 24, 20, 25, 16, 23, 25, 30, 34, 32, 
    31, 28, 40, 30, 29, 19, 20, 26, 22, 27, 26, 22, 20, 30, 27, 
    30, 20, 36, 34, 24, 28, 25, 27, 25, 27, 34, 32, 17, 19, 23, 
    31, 27, 27, 30, 19, 18, 20, 27, 34, 31, 32, 33, 36, 37, 23, 
    27, 26, 20, 30, 30, 27, 21, 24, 29, 34, 26, 32, 30, 30, 31, 
    26, 28, 20, 26, 30, 32, 33, 31, 32, 32, 30, 29, 30, 34, 30, 
    28, 29, 19, 23, 27, 25, 33, 30, 31, 30, 26, 27, 26, 24, 30, 
    30, 30, 15, 21, 30, 44, 36, 29, 30, 25, 27, 26, 28, 24, 31, 
    23, 29, 15, 15, 25, 30, 30, 28, 29, 24, 25, 28, 29, 30, 25, 
    
    -- channel=137
    34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=138
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=139
    1, 0, 0, 0, 0, 0, 0, 0, 36, 24, 0, 13, 5, 0, 0, 
    1, 0, 0, 0, 27, 0, 0, 0, 0, 15, 32, 3, 0, 0, 0, 
    1, 0, 0, 0, 0, 6, 0, 0, 0, 1, 15, 0, 0, 3, 10, 
    140, 124, 70, 0, 0, 18, 63, 22, 1, 0, 0, 0, 3, 0, 0, 
    38, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 22, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 3, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 3, 0, 37, 30, 11, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 29, 48, 0, 0, 0, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=140
    17, 51, 31, 15, 16, 24, 21, 25, 12, 0, 40, 25, 18, 20, 18, 
    17, 34, 46, 15, 8, 5, 14, 17, 7, 0, 52, 16, 14, 16, 14, 
    17, 23, 67, 15, 8, 0, 9, 16, 5, 12, 31, 17, 8, 9, 10, 
    15, 43, 52, 0, 18, 0, 0, 5, 15, 25, 10, 21, 0, 0, 17, 
    6, 27, 17, 0, 26, 0, 0, 0, 11, 17, 18, 26, 2, 1, 29, 
    13, 16, 14, 0, 15, 0, 0, 0, 10, 13, 16, 29, 9, 4, 28, 
    17, 16, 2, 16, 8, 6, 0, 4, 1, 13, 12, 28, 11, 7, 15, 
    13, 14, 0, 35, 0, 0, 0, 0, 13, 8, 4, 20, 21, 4, 13, 
    9, 20, 0, 17, 0, 3, 0, 0, 25, 0, 11, 9, 37, 11, 32, 
    13, 13, 7, 3, 9, 0, 0, 0, 0, 12, 6, 16, 14, 13, 25, 
    15, 2, 17, 4, 1, 0, 15, 0, 0, 0, 13, 18, 10, 3, 10, 
    15, 5, 26, 0, 0, 0, 12, 2, 0, 0, 26, 9, 11, 1, 8, 
    15, 16, 28, 1, 0, 0, 13, 4, 0, 1, 22, 8, 9, 10, 11, 
    14, 19, 34, 7, 0, 0, 7, 8, 3, 11, 22, 11, 6, 23, 13, 
    15, 25, 27, 14, 0, 0, 0, 13, 5, 20, 17, 15, 11, 18, 16, 
    
    -- channel=141
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 8, 28, 12, 5, 13, 0, 1, 1, 0, 0, 0, 
    0, 0, 0, 2, 17, 12, 0, 3, 0, 0, 17, 0, 9, 28, 2, 
    0, 0, 0, 0, 2, 20, 18, 22, 2, 0, 2, 1, 8, 7, 0, 
    0, 0, 5, 0, 7, 26, 27, 0, 2, 0, 9, 0, 12, 0, 0, 
    0, 0, 6, 0, 10, 0, 22, 0, 19, 14, 1, 0, 9, 2, 0, 
    0, 0, 0, 0, 15, 25, 15, 18, 2, 3, 20, 21, 8, 24, 0, 
    4, 0, 0, 0, 7, 10, 13, 23, 0, 0, 0, 0, 0, 14, 0, 
    0, 0, 10, 6, 17, 31, 23, 8, 0, 0, 13, 0, 0, 0, 0, 
    2, 10, 4, 2, 2, 22, 10, 14, 14, 18, 0, 0, 0, 0, 0, 
    5, 8, 2, 17, 20, 9, 0, 1, 12, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 20, 35, 0, 0, 5, 9, 0, 0, 0, 11, 0, 0, 
    4, 0, 0, 16, 11, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 20, 15, 14, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=142
    0, 45, 28, 8, 12, 24, 18, 13, 0, 0, 23, 6, 15, 17, 19, 
    0, 31, 38, 8, 0, 0, 12, 4, 0, 0, 11, 0, 0, 6, 11, 
    0, 12, 32, 4, 0, 0, 3, 20, 11, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 22, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 7, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 3, 0, 0, 1, 8, 1, 5, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 4, 5, 6, 2, 0, 9, 1, 
    0, 0, 0, 0, 0, 0, 5, 12, 3, 13, 4, 3, 0, 7, 4, 
    
    -- channel=143
    1, 38, 24, 29, 24, 40, 38, 37, 22, 25, 41, 26, 43, 45, 45, 
    4, 26, 1, 40, 6, 30, 29, 30, 24, 33, 21, 28, 35, 42, 42, 
    7, 8, 0, 39, 2, 10, 18, 16, 10, 32, 0, 27, 25, 26, 29, 
    14, 44, 9, 34, 0, 16, 24, 9, 13, 28, 2, 29, 27, 17, 33, 
    39, 29, 22, 40, 0, 11, 15, 13, 11, 23, 19, 12, 28, 37, 36, 
    33, 33, 25, 47, 7, 14, 4, 28, 0, 19, 18, 15, 26, 37, 42, 
    35, 40, 41, 9, 5, 23, 4, 34, 0, 6, 27, 15, 32, 30, 50, 
    39, 35, 30, 2, 22, 3, 19, 10, 15, 42, 9, 44, 19, 18, 48, 
    28, 33, 20, 15, 20, 6, 18, 0, 42, 40, 8, 31, 27, 26, 41, 
    34, 42, 10, 19, 16, 13, 14, 20, 25, 27, 15, 25, 38, 22, 23, 
    33, 31, 15, 24, 27, 14, 12, 23, 20, 11, 35, 21, 15, 27, 27, 
    33, 26, 17, 18, 15, 40, 16, 26, 18, 32, 26, 24, 12, 29, 23, 
    34, 36, 28, 10, 0, 59, 10, 27, 22, 32, 18, 29, 14, 24, 21, 
    37, 38, 39, 8, 21, 39, 16, 25, 28, 38, 17, 26, 25, 24, 24, 
    39, 30, 51, 0, 23, 16, 34, 21, 20, 32, 23, 21, 27, 23, 19, 
    
    -- channel=144
    70, 71, 77, 72, 57, 54, 48, 53, 73, 80, 81, 75, 64, 55, 54, 
    90, 88, 89, 93, 82, 88, 91, 99, 98, 90, 70, 75, 82, 75, 56, 
    97, 97, 93, 92, 58, 71, 74, 78, 73, 74, 50, 74, 83, 70, 46, 
    97, 101, 92, 94, 69, 97, 122, 110, 103, 84, 98, 70, 72, 53, 60, 
    97, 96, 111, 96, 80, 111, 108, 105, 106, 111, 102, 63, 84, 72, 39, 
    90, 101, 88, 94, 70, 88, 92, 102, 102, 100, 102, 100, 78, 98, 97, 
    86, 94, 80, 63, 60, 89, 100, 79, 74, 91, 81, 72, 91, 94, 100, 
    89, 81, 38, 83, 94, 80, 59, 70, 75, 72, 62, 74, 75, 87, 75, 
    67, 63, 58, 65, 57, 59, 71, 44, 0, 7, 29, 0, 26, 78, 82, 
    84, 80, 48, 46, 51, 58, 60, 61, 100, 83, 94, 85, 83, 81, 64, 
    84, 70, 34, 40, 35, 30, 34, 66, 52, 65, 61, 50, 56, 54, 66, 
    97, 94, 23, 33, 36, 32, 58, 51, 29, 67, 57, 75, 81, 54, 53, 
    97, 58, 34, 65, 45, 18, 11, 14, 14, 16, 69, 74, 41, 17, 49, 
    88, 98, 84, 61, 52, 35, 3, 6, 24, 66, 76, 80, 24, 19, 60, 
    98, 90, 75, 55, 48, 32, 14, 17, 26, 41, 65, 56, 24, 21, 48, 
    
    -- channel=145
    0, 0, 0, 0, 0, 3, 8, 20, 5, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 19, 17, 16, 1, 3, 8, 40, 0, 0, 0, 13, 
    0, 0, 0, 0, 59, 10, 0, 0, 0, 18, 0, 14, 0, 0, 0, 
    0, 0, 0, 0, 24, 3, 0, 0, 0, 0, 0, 50, 1, 0, 17, 
    0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 7, 38, 0, 0, 
    0, 0, 0, 0, 17, 2, 0, 0, 12, 0, 0, 15, 2, 0, 0, 
    0, 0, 34, 0, 0, 0, 4, 0, 0, 0, 0, 0, 6, 13, 52, 
    0, 0, 25, 0, 14, 15, 0, 0, 54, 67, 0, 43, 64, 11, 66, 
    0, 0, 0, 0, 14, 0, 1, 39, 0, 0, 0, 0, 0, 0, 93, 
    0, 0, 2, 0, 0, 19, 35, 0, 23, 0, 0, 29, 0, 12, 84, 
    0, 0, 21, 5, 0, 0, 10, 0, 70, 0, 0, 1, 0, 0, 93, 
    0, 0, 35, 0, 0, 0, 0, 7, 30, 96, 0, 0, 0, 23, 101, 
    1, 0, 0, 0, 0, 0, 9, 19, 24, 15, 0, 0, 0, 43, 78, 
    0, 0, 0, 0, 0, 0, 4, 7, 11, 10, 9, 0, 0, 28, 97, 
    
    -- channel=146
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=147
    410, 409, 410, 362, 312, 319, 340, 370, 418, 427, 421, 407, 402, 387, 360, 
    453, 452, 453, 357, 275, 266, 274, 302, 325, 345, 368, 396, 418, 405, 360, 
    458, 457, 444, 334, 175, 238, 238, 250, 239, 247, 280, 410, 422, 368, 324, 
    456, 460, 406, 348, 209, 320, 355, 283, 281, 275, 337, 335, 393, 383, 333, 
    450, 456, 399, 259, 217, 267, 270, 258, 276, 283, 310, 323, 417, 431, 370, 
    405, 449, 330, 272, 147, 204, 227, 214, 216, 222, 249, 278, 359, 459, 457, 
    375, 377, 296, 222, 209, 230, 226, 190, 189, 236, 211, 214, 305, 353, 429, 
    369, 286, 195, 320, 187, 170, 143, 145, 111, 102, 111, 109, 134, 223, 332, 
    362, 265, 238, 212, 138, 198, 206, 203, 171, 196, 250, 186, 213, 264, 304, 
    382, 281, 175, 131, 125, 142, 136, 147, 273, 226, 244, 226, 248, 206, 198, 
    373, 283, 157, 124, 90, 75, 129, 195, 111, 201, 163, 173, 205, 163, 224, 
    366, 270, 102, 179, 146, 72, 97, 98, 98, 198, 221, 259, 168, 138, 127, 
    323, 266, 207, 232, 153, 95, 39, 43, 55, 164, 338, 310, 118, 63, 160, 
    319, 326, 259, 221, 157, 122, 47, 55, 93, 196, 227, 273, 71, 71, 165, 
    309, 288, 269, 187, 139, 112, 81, 84, 95, 122, 163, 184, 95, 72, 163, 
    
    -- channel=148
    90, 79, 95, 89, 77, 66, 62, 61, 73, 98, 97, 95, 90, 83, 76, 
    96, 95, 110, 84, 51, 53, 52, 72, 88, 92, 94, 92, 103, 112, 89, 
    99, 99, 106, 54, 0, 0, 0, 0, 0, 19, 58, 92, 107, 109, 83, 
    99, 103, 85, 74, 5, 27, 20, 10, 6, 7, 29, 89, 96, 104, 73, 
    99, 107, 85, 45, 0, 10, 24, 0, 12, 3, 33, 52, 82, 97, 68, 
    96, 115, 59, 27, 0, 0, 1, 2, 2, 1, 27, 26, 77, 99, 99, 
    82, 104, 69, 39, 0, 0, 11, 0, 0, 20, 12, 19, 61, 89, 93, 
    100, 76, 47, 65, 0, 0, 0, 11, 8, 0, 12, 12, 0, 16, 71, 
    88, 55, 40, 52, 1, 30, 4, 0, 0, 0, 6, 0, 0, 26, 32, 
    87, 63, 50, 12, 0, 7, 0, 19, 29, 28, 38, 31, 53, 20, 1, 
    84, 65, 11, 10, 0, 0, 0, 13, 0, 13, 5, 0, 24, 9, 0, 
    69, 63, 22, 7, 7, 0, 9, 34, 3, 35, 25, 55, 26, 17, 0, 
    48, 37, 0, 41, 16, 4, 0, 0, 0, 17, 41, 65, 7, 0, 0, 
    45, 52, 41, 45, 14, 16, 0, 0, 0, 10, 42, 78, 6, 0, 0, 
    37, 34, 40, 24, 10, 13, 0, 0, 0, 0, 10, 52, 0, 0, 0, 
    
    -- channel=149
    1, 0, 11, 36, 0, 0, 0, 0, 0, 0, 2, 0, 27, 0, 26, 
    0, 0, 25, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 
    0, 0, 29, 144, 0, 0, 0, 15, 1, 0, 0, 0, 17, 38, 0, 
    0, 8, 15, 134, 0, 0, 40, 0, 0, 0, 0, 0, 14, 36, 0, 
    0, 19, 42, 96, 0, 0, 26, 0, 0, 0, 12, 0, 0, 34, 1, 
    0, 32, 54, 104, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 49, 11, 74, 0, 0, 19, 10, 0, 0, 14, 0, 0, 0, 0, 
    8, 74, 0, 53, 10, 23, 5, 23, 0, 0, 13, 0, 0, 0, 0, 
    25, 89, 0, 85, 0, 0, 2, 32, 0, 0, 39, 5, 0, 0, 0, 
    30, 123, 0, 63, 0, 23, 0, 0, 21, 0, 12, 0, 0, 46, 0, 
    7, 137, 6, 28, 11, 0, 0, 48, 0, 28, 8, 0, 38, 0, 0, 
    10, 147, 0, 10, 64, 0, 0, 66, 0, 10, 0, 0, 94, 0, 0, 
    0, 101, 0, 11, 51, 41, 1, 0, 0, 0, 5, 89, 48, 0, 0, 
    0, 23, 55, 14, 10, 63, 1, 0, 0, 0, 0, 102, 41, 0, 0, 
    8, 10, 46, 37, 4, 29, 5, 0, 0, 0, 0, 48, 40, 0, 0, 
    
    -- channel=150
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 19, 27, 15, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 8, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 
    0, 0, 0, 14, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 20, 0, 0, 0, 1, 3, 11, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 6, 18, 0, 
    0, 7, 7, 0, 0, 12, 39, 22, 20, 25, 29, 12, 19, 14, 4, 
    0, 0, 0, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 10, 20, 39, 0, 40, 31, 32, 23, 21, 0, 
    0, 0, 0, 0, 3, 22, 0, 0, 26, 6, 15, 0, 20, 0, 0, 
    0, 0, 23, 0, 0, 0, 35, 44, 0, 0, 0, 0, 2, 23, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 4, 14, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 
    
    -- channel=151
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 19, 10, 4, 19, 16, 0, 7, 0, 0, 12, 
    0, 0, 0, 0, 38, 3, 0, 0, 0, 10, 55, 0, 0, 0, 23, 
    0, 0, 0, 0, 64, 13, 0, 0, 0, 3, 0, 42, 0, 0, 0, 
    0, 0, 0, 0, 39, 8, 0, 1, 2, 7, 0, 33, 9, 0, 0, 
    17, 0, 0, 0, 28, 13, 0, 0, 0, 13, 0, 19, 49, 0, 0, 
    7, 0, 0, 0, 5, 0, 0, 0, 16, 0, 0, 30, 33, 27, 14, 
    0, 0, 57, 0, 1, 0, 0, 0, 0, 5, 0, 8, 49, 33, 77, 
    0, 0, 35, 0, 43, 3, 7, 0, 7, 12, 0, 0, 19, 0, 70, 
    0, 0, 24, 0, 25, 0, 12, 51, 0, 11, 0, 5, 9, 0, 104, 
    0, 0, 0, 0, 0, 24, 33, 0, 60, 0, 0, 34, 0, 36, 59, 
    0, 0, 44, 6, 0, 1, 29, 0, 64, 8, 4, 0, 0, 8, 111, 
    0, 0, 0, 0, 0, 0, 3, 12, 25, 102, 0, 0, 0, 34, 93, 
    0, 0, 0, 0, 0, 0, 3, 14, 26, 34, 29, 0, 0, 45, 81, 
    0, 0, 0, 0, 0, 0, 0, 5, 9, 14, 20, 0, 0, 36, 102, 
    
    -- channel=152
    25, 22, 25, 23, 16, 25, 29, 31, 24, 24, 24, 22, 30, 30, 26, 
    23, 22, 24, 14, 0, 0, 0, 0, 0, 1, 14, 20, 23, 28, 23, 
    20, 19, 21, 8, 0, 0, 0, 0, 0, 0, 0, 25, 27, 25, 14, 
    20, 19, 15, 11, 0, 3, 0, 0, 0, 0, 2, 4, 23, 35, 24, 
    20, 21, 7, 0, 0, 0, 0, 0, 0, 0, 0, 2, 19, 27, 32, 
    18, 21, 15, 10, 0, 0, 0, 0, 0, 0, 0, 0, 6, 20, 20, 
    19, 19, 12, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    28, 15, 11, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 25, 12, 0, 0, 8, 2, 11, 24, 24, 28, 26, 16, 11, 1, 
    22, 18, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 21, 7, 1, 0, 0, 0, 5, 0, 1, 0, 0, 5, 2, 0, 
    5, 8, 0, 11, 9, 0, 0, 0, 0, 0, 6, 5, 0, 0, 0, 
    1, 17, 11, 2, 4, 7, 1, 0, 0, 14, 25, 22, 5, 0, 0, 
    1, 2, 6, 0, 0, 7, 4, 3, 3, 0, 0, 5, 2, 0, 0, 
    0, 0, 2, 0, 0, 3, 2, 1, 0, 0, 0, 4, 5, 0, 0, 
    
    -- channel=153
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 18, 12, 6, 20, 2, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 17, 3, 6, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 20, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 4, 29, 31, 27, 18, 0, 0, 0, 14, 15, 0, 
    0, 0, 0, 0, 0, 17, 32, 28, 13, 0, 0, 0, 20, 14, 0, 
    0, 0, 0, 0, 0, 9, 23, 20, 13, 0, 0, 0, 25, 13, 0, 
    
    -- channel=154
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=155
    11, 9, 3, 0, 0, 16, 33, 54, 9, 0, 0, 0, 26, 13, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 20, 58, 64, 67, 29, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 14, 36, 0, 0, 0, 20, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 30, 85, 
    0, 0, 6, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 57, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 17, 0, 0, 0, 0, 9, 80, 165, 158, 154, 174, 121, 17, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 19, 16, 1, 0, 0, 53, 9, 0, 12, 3, 42, 0, 25, 0, 
    0, 0, 0, 64, 37, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 105, 75, 0, 27, 27, 0, 0, 2, 52, 55, 38, 0, 0, 0, 
    0, 0, 1, 0, 0, 19, 20, 17, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 5, 20, 17, 5, 0, 0, 0, 18, 0, 11, 
    
    -- channel=156
    0, 1, 0, 0, 0, 0, 3, 5, 6, 0, 0, 3, 0, 11, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 5, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 9, 0, 0, 29, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 15, 
    0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 0, 20, 
    0, 0, 10, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 1, 0, 0, 4, 1, 0, 11, 0, 0, 3, 0, 0, 11, 
    0, 0, 13, 0, 0, 4, 5, 0, 20, 0, 0, 0, 0, 7, 17, 
    0, 0, 0, 0, 0, 0, 9, 11, 11, 26, 0, 0, 0, 11, 20, 
    0, 0, 0, 0, 0, 0, 12, 11, 8, 19, 0, 0, 0, 15, 10, 
    0, 0, 0, 0, 0, 0, 5, 5, 3, 0, 0, 0, 0, 15, 17, 
    
    -- channel=157
    16, 14, 23, 24, 17, 8, 7, 4, 23, 26, 23, 17, 6, 5, 1, 
    30, 29, 40, 61, 73, 75, 72, 82, 76, 46, 22, 19, 24, 18, 0, 
    36, 36, 44, 56, 50, 58, 57, 62, 68, 58, 10, 22, 27, 18, 1, 
    36, 43, 34, 80, 57, 71, 96, 96, 85, 71, 72, 22, 16, 9, 13, 
    35, 41, 77, 78, 76, 90, 91, 94, 90, 87, 84, 32, 25, 19, 0, 
    28, 53, 28, 83, 64, 74, 82, 90, 91, 79, 84, 61, 21, 37, 36, 
    29, 49, 33, 25, 58, 82, 94, 75, 70, 92, 68, 57, 68, 51, 36, 
    37, 44, 0, 55, 77, 60, 53, 61, 68, 62, 55, 66, 62, 59, 30, 
    20, 25, 21, 52, 39, 42, 44, 28, 0, 0, 11, 0, 4, 58, 41, 
    31, 49, 41, 17, 52, 46, 54, 36, 82, 64, 76, 68, 73, 59, 18, 
    32, 39, 23, 28, 28, 25, 15, 56, 29, 43, 40, 18, 47, 25, 27, 
    58, 66, 18, 18, 30, 26, 49, 40, 26, 42, 42, 65, 46, 61, 4, 
    60, 21, 22, 56, 31, 20, 15, 15, 7, 0, 39, 62, 34, 11, 18, 
    56, 70, 56, 59, 42, 28, 5, 7, 16, 62, 51, 76, 14, 15, 28, 
    72, 64, 60, 50, 41, 26, 12, 15, 21, 33, 49, 53, 18, 16, 15, 
    
    -- channel=158
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 0, 21, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=159
    18, 18, 6, 30, 11, 16, 23, 21, 7, 17, 21, 21, 28, 30, 34, 
    14, 14, 4, 22, 0, 0, 0, 0, 0, 10, 22, 9, 18, 33, 29, 
    11, 10, 9, 2, 0, 0, 0, 0, 0, 0, 25, 3, 17, 25, 34, 
    12, 1, 21, 0, 0, 0, 0, 0, 0, 0, 0, 8, 19, 24, 26, 
    11, 3, 8, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 10, 30, 
    11, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 11, 10, 
    1, 8, 12, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 
    1, 20, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 37, 0, 24, 0, 4, 0, 0, 4, 16, 0, 0, 0, 0, 0, 
    7, 23, 0, 27, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 12, 
    5, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 23, 
    0, 17, 0, 0, 5, 0, 0, 2, 0, 0, 0, 0, 19, 0, 30, 
    0, 2, 0, 0, 0, 3, 0, 0, 8, 0, 0, 0, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 18, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 
    
    
    others => 0);
end gold_package;
