library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=2
    0, 0, 39, 
    0, 0, 291, 
    0, 0, 0, 
    
    -- channel=3
    459, 98, 382, 
    258, 0, 0, 
    0, 0, 29, 
    
    -- channel=4
    177, 0, 403, 
    0, 0, 183, 
    0, 3, 39, 
    
    -- channel=5
    489, 0, 17, 
    0, 374, 0, 
    0, 0, 0, 
    
    -- channel=6
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=7
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=8
    313, 0, 249, 
    160, 168, 239, 
    0, 0, 0, 
    
    -- channel=9
    0, 0, 0, 
    0, 282, 90, 
    181, 287, 269, 
    
    -- channel=10
    67, 0, 80, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=11
    0, 0, 0, 
    0, 0, 16, 
    312, 0, 0, 
    
    -- channel=12
    355, 0, 281, 
    6, 207, 0, 
    178, 187, 458, 
    
    -- channel=13
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=14
    0, 0, 130, 
    0, 117, 0, 
    0, 0, 0, 
    
    -- channel=15
    370, 303, 152, 
    237, 0, 136, 
    0, 0, 0, 
    
    -- channel=16
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=17
    0, 0, 78, 
    0, 203, 257, 
    0, 172, 0, 
    
    -- channel=18
    66, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=19
    18, 0, 0, 
    0, 0, 5, 
    0, 0, 0, 
    
    -- channel=20
    435, 54, 586, 
    206, 250, 199, 
    197, 0, 0, 
    
    -- channel=21
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=22
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=23
    254, 330, 203, 
    279, 124, 11, 
    0, 0, 0, 
    
    -- channel=24
    157, 0, 54, 
    177, 79, 0, 
    0, 0, 0, 
    
    -- channel=25
    85, 31, 0, 
    0, 0, 0, 
    0, 319, 309, 
    
    -- channel=26
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=27
    0, 0, 0, 
    0, 0, 0, 
    0, 555, 494, 
    
    -- channel=28
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=29
    0, 0, 0, 
    0, 0, 0, 
    0, 350, 0, 
    
    -- channel=30
    0, 0, 0, 
    0, 0, 0, 
    155, 0, 0, 
    
    -- channel=31
    0, 0, 0, 
    0, 0, 0, 
    0, 304, 549, 
    
    -- channel=32
    0, 0, 80, 
    124, 23, 145, 
    0, 0, 0, 
    
    -- channel=33
    0, 68, 227, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=34
    589, 188, 347, 
    235, 0, 52, 
    80, 0, 0, 
    
    -- channel=35
    82, 97, 365, 
    471, 0, 0, 
    0, 0, 0, 
    
    -- channel=36
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=37
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=38
    0, 0, 0, 
    0, 0, 0, 
    0, 171, 55, 
    
    -- channel=39
    0, 260, 2, 
    0, 140, 0, 
    59, 0, 0, 
    
    -- channel=40
    0, 0, 0, 
    287, 106, 159, 
    0, 0, 0, 
    
    -- channel=41
    347, 128, 196, 
    368, 249, 0, 
    0, 62, 168, 
    
    -- channel=42
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=43
    0, 0, 0, 
    0, 111, 0, 
    0, 50, 0, 
    
    -- channel=44
    0, 0, 128, 
    85, 0, 0, 
    0, 0, 0, 
    
    -- channel=45
    0, 0, 11, 
    0, 162, 160, 
    0, 0, 0, 
    
    -- channel=46
    0, 0, 67, 
    0, 125, 105, 
    0, 68, 0, 
    
    -- channel=47
    0, 0, 134, 
    0, 258, 0, 
    0, 0, 0, 
    
    -- channel=48
    0, 244, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=49
    0, 0, 0, 
    0, 11, 167, 
    0, 0, 0, 
    
    -- channel=50
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=51
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=52
    0, 112, 66, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=53
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=54
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=55
    89, 0, 25, 
    186, 0, 0, 
    0, 258, 477, 
    
    -- channel=56
    72, 0, 0, 
    0, 14, 0, 
    0, 0, 0, 
    
    -- channel=57
    0, 0, 0, 
    0, 148, 101, 
    0, 0, 28, 
    
    -- channel=58
    20, 0, 0, 
    150, 0, 0, 
    0, 0, 0, 
    
    -- channel=59
    55, 103, 109, 
    172, 511, 273, 
    314, 0, 0, 
    
    -- channel=60
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 79, 
    
    -- channel=61
    0, 0, 0, 
    0, 0, 0, 
    0, 33, 0, 
    
    -- channel=62
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=63
    0, 0, 0, 
    0, 0, 0, 
    0, 6, 70, 
    
    -- channel=64
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=65
    206, 211, 137, 
    335, 0, 0, 
    0, 0, 0, 
    
    -- channel=66
    0, 0, 0, 
    9, 69, 0, 
    0, 0, 0, 
    
    -- channel=67
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=68
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=69
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=70
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=71
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=72
    86, 131, 0, 
    236, 138, 259, 
    118, 0, 0, 
    
    -- channel=73
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=74
    0, 0, 0, 
    271, 263, 242, 
    448, 0, 0, 
    
    -- channel=75
    76, 0, 67, 
    0, 0, 0, 
    201, 0, 0, 
    
    -- channel=76
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=77
    0, 0, 0, 
    329, 0, 54, 
    0, 251, 255, 
    
    -- channel=78
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 494, 
    
    -- channel=79
    0, 0, 0, 
    0, 0, 0, 
    0, 156, 210, 
    
    -- channel=80
    172, 141, 249, 
    93, 200, 0, 
    182, 109, 223, 
    
    -- channel=81
    0, 148, 235, 
    55, 0, 20, 
    94, 158, 258, 
    
    -- channel=82
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=83
    81, 17, 16, 
    0, 0, 74, 
    0, 0, 0, 
    
    -- channel=84
    0, 0, 0, 
    22, 0, 200, 
    59, 269, 135, 
    
    -- channel=85
    26, 0, 0, 
    0, 0, 102, 
    456, 270, 0, 
    
    -- channel=86
    0, 0, 1, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=87
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=88
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=89
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=90
    380, 35, 198, 
    156, 331, 132, 
    0, 0, 0, 
    
    -- channel=91
    0, 60, 217, 
    395, 295, 151, 
    0, 49, 27, 
    
    -- channel=92
    0, 0, 0, 
    0, 0, 0, 
    0, 11, 0, 
    
    -- channel=93
    30, 0, 148, 
    261, 43, 118, 
    16, 0, 0, 
    
    -- channel=94
    0, 0, 0, 
    155, 146, 67, 
    517, 0, 0, 
    
    -- channel=95
    316, 345, 154, 
    406, 44, 0, 
    411, 59, 319, 
    
    -- channel=96
    0, 65, 0, 
    0, 173, 0, 
    0, 44, 0, 
    
    -- channel=97
    0, 215, 0, 
    0, 0, 46, 
    0, 55, 110, 
    
    -- channel=98
    0, 0, 0, 
    42, 0, 0, 
    0, 181, 0, 
    
    -- channel=99
    321, 0, 214, 
    0, 0, 0, 
    0, 0, 51, 
    
    -- channel=100
    0, 0, 203, 
    82, 332, 0, 
    0, 0, 0, 
    
    -- channel=101
    254, 410, 483, 
    429, 436, 126, 
    0, 0, 0, 
    
    -- channel=102
    313, 312, 149, 
    326, 0, 0, 
    0, 0, 0, 
    
    -- channel=103
    0, 223, 0, 
    206, 98, 32, 
    0, 0, 0, 
    
    -- channel=104
    137, 127, 349, 
    589, 98, 0, 
    402, 0, 0, 
    
    -- channel=105
    0, 151, 27, 
    164, 178, 0, 
    0, 0, 0, 
    
    -- channel=106
    0, 0, 0, 
    0, 0, 0, 
    503, 0, 0, 
    
    -- channel=107
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=108
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=109
    94, 57, 0, 
    246, 0, 0, 
    0, 116, 115, 
    
    -- channel=110
    0, 0, 0, 
    0, 0, 0, 
    159, 0, 0, 
    
    -- channel=111
    0, 0, 130, 
    65, 55, 0, 
    0, 0, 11, 
    
    -- channel=112
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=113
    40, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=114
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=115
    0, 0, 0, 
    0, 0, 278, 
    88, 60, 0, 
    
    -- channel=116
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=117
    369, 310, 0, 
    0, 0, 97, 
    0, 0, 0, 
    
    -- channel=118
    0, 0, 0, 
    0, 0, 15, 
    0, 0, 0, 
    
    -- channel=119
    0, 0, 0, 
    0, 0, 0, 
    0, 111, 0, 
    
    -- channel=120
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=121
    24, 92, 91, 
    451, 324, 191, 
    304, 0, 0, 
    
    -- channel=122
    0, 0, 0, 
    0, 0, 43, 
    0, 0, 0, 
    
    -- channel=123
    31, 0, 10, 
    0, 80, 68, 
    0, 0, 0, 
    
    -- channel=124
    0, 0, 276, 
    265, 0, 223, 
    122, 262, 148, 
    
    -- channel=125
    0, 262, 5, 
    0, 0, 129, 
    27, 132, 423, 
    
    -- channel=126
    60, 0, 6, 
    0, 0, 96, 
    0, 196, 484, 
    
    -- channel=127
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    
    others => 0);
end gold_package;
